
module Fetch_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n2, n4, n7, n9, n11, n12, n13, n14, n17, n18, n19,
         n22, n23, n24, n30, n38, n39, n42, n45, n47, n49, n50, n54, n55, n56,
         n57, n58, n59, n61, n62, n63, n64, n65, n69, n70, n71, n73, n76, n77,
         n79, n82, n85, n86, n87, n89, n94, n95, n96, n97, n101, n102, n103,
         n104, n109, n110, n114, n115, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n132, n133, n134,
         n135, n136, n137, n138, n139;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2_X1 U13 ( .A(n7), .B(A[9]), .Z(SUM[9]) );
  XOR2_X1 U20 ( .A(n12), .B(A[8]), .Z(SUM[8]) );
  XOR2_X1 U23 ( .A(n13), .B(A[7]), .Z(SUM[7]) );
  XOR2_X1 U24 ( .A(A[12]), .B(n14), .Z(SUM[12]) );
  XOR2_X1 U40 ( .A(n54), .B(A[31]), .Z(SUM[31]) );
  NAND3_X1 U86 ( .A1(A[4]), .A2(A[2]), .A3(A[9]), .ZN(n56) );
  XOR2_X1 U105 ( .A(n64), .B(A[18]), .Z(SUM[18]) );
  XOR2_X1 U106 ( .A(n58), .B(A[16]), .Z(SUM[16]) );
  XOR2_X1 U107 ( .A(n77), .B(A[6]), .Z(SUM[6]) );
  XOR2_X1 U108 ( .A(A[2]), .B(A[3]), .Z(SUM[3]) );
  XOR2_X1 U109 ( .A(n18), .B(A[4]), .Z(SUM[4]) );
  XOR2_X1 U110 ( .A(n70), .B(A[10]), .Z(SUM[10]) );
  XOR2_X1 U111 ( .A(n89), .B(A[24]), .Z(SUM[24]) );
  NAND3_X1 U143 ( .A1(n49), .A2(n42), .A3(A[29]), .ZN(n82) );
  NAND3_X1 U144 ( .A1(A[8]), .A2(A[11]), .A3(A[12]), .ZN(n104) );
  NOR2_X1 U2 ( .A1(n19), .A2(n137), .ZN(n23) );
  AND2_X1 U3 ( .A1(n59), .A2(A[14]), .ZN(n2) );
  AND2_X1 U4 ( .A1(n4), .A2(A[26]), .ZN(n39) );
  OR2_X1 U5 ( .A1(n87), .A2(n138), .ZN(n86) );
  NOR2_X1 U6 ( .A1(n76), .A2(n132), .ZN(n12) );
  NAND2_X1 U7 ( .A1(n58), .A2(n85), .ZN(n71) );
  INV_X1 U8 ( .A(n58), .ZN(n134) );
  AND2_X1 U9 ( .A1(n45), .A2(n85), .ZN(n89) );
  AND2_X1 U10 ( .A1(n45), .A2(n85), .ZN(n61) );
  AND2_X1 U11 ( .A1(n101), .A2(n102), .ZN(n58) );
  NAND2_X1 U12 ( .A1(n114), .A2(n115), .ZN(n76) );
  AND2_X1 U14 ( .A1(n101), .A2(n102), .ZN(n45) );
  INV_X1 U15 ( .A(n79), .ZN(n132) );
  AND2_X1 U16 ( .A1(n63), .A2(n94), .ZN(n85) );
  NAND2_X1 U17 ( .A1(n114), .A2(n115), .ZN(n30) );
  XNOR2_X1 U18 ( .A(n38), .B(n138), .ZN(SUM[28]) );
  NOR2_X1 U19 ( .A1(n71), .A2(n87), .ZN(n38) );
  XNOR2_X1 U21 ( .A(n135), .B(n69), .ZN(SUM[5]) );
  NAND4_X1 U22 ( .A1(A[24]), .A2(A[25]), .A3(A[26]), .A4(A[27]), .ZN(n87) );
  NAND4_X1 U25 ( .A1(A[8]), .A2(A[11]), .A3(A[10]), .A4(A[9]), .ZN(n19) );
  AND2_X1 U26 ( .A1(n63), .A2(n94), .ZN(n49) );
  NOR2_X1 U27 ( .A1(n87), .A2(n138), .ZN(n42) );
  NOR2_X1 U28 ( .A1(n55), .A2(n56), .ZN(n102) );
  NAND4_X1 U29 ( .A1(A[3]), .A2(A[5]), .A3(A[6]), .A4(A[7]), .ZN(n55) );
  NOR2_X1 U30 ( .A1(n24), .A2(n96), .ZN(n94) );
  NAND2_X1 U31 ( .A1(A[16]), .A2(A[17]), .ZN(n24) );
  NOR2_X1 U32 ( .A1(n110), .A2(n137), .ZN(n109) );
  NAND4_X1 U33 ( .A1(A[8]), .A2(A[11]), .A3(A[10]), .A4(A[9]), .ZN(n110) );
  NOR2_X1 U34 ( .A1(n76), .A2(n17), .ZN(n59) );
  NAND2_X1 U35 ( .A1(n18), .A2(A[13]), .ZN(n17) );
  NOR2_X1 U36 ( .A1(n103), .A2(n104), .ZN(n101) );
  NAND4_X1 U37 ( .A1(A[14]), .A2(A[15]), .A3(A[13]), .A4(A[10]), .ZN(n103) );
  NOR2_X1 U38 ( .A1(n96), .A2(n97), .ZN(n57) );
  NAND2_X1 U39 ( .A1(A[16]), .A2(A[17]), .ZN(n97) );
  AND2_X1 U41 ( .A1(n79), .A2(A[4]), .ZN(n69) );
  INV_X1 U42 ( .A(A[5]), .ZN(n135) );
  INV_X1 U43 ( .A(A[28]), .ZN(n138) );
  NOR2_X1 U44 ( .A1(n76), .A2(n22), .ZN(n7) );
  NAND2_X1 U45 ( .A1(n18), .A2(A[8]), .ZN(n22) );
  NOR2_X1 U46 ( .A1(n133), .A2(n135), .ZN(n77) );
  INV_X1 U47 ( .A(n69), .ZN(n133) );
  XNOR2_X1 U48 ( .A(n117), .B(A[22]), .ZN(SUM[22]) );
  NAND3_X1 U49 ( .A1(n45), .A2(n9), .A3(A[21]), .ZN(n117) );
  XNOR2_X1 U50 ( .A(n118), .B(A[20]), .ZN(SUM[20]) );
  NAND2_X1 U51 ( .A1(n57), .A2(n58), .ZN(n118) );
  XNOR2_X1 U52 ( .A(n119), .B(A[21]), .ZN(SUM[21]) );
  NAND2_X1 U53 ( .A1(n58), .A2(n9), .ZN(n119) );
  AND2_X1 U54 ( .A1(n69), .A2(n11), .ZN(n13) );
  NOR2_X1 U55 ( .A1(n135), .A2(n136), .ZN(n11) );
  INV_X1 U56 ( .A(A[6]), .ZN(n136) );
  XNOR2_X1 U57 ( .A(n120), .B(A[14]), .ZN(SUM[14]) );
  NAND2_X1 U58 ( .A1(n109), .A2(n59), .ZN(n120) );
  XNOR2_X1 U59 ( .A(n121), .B(A[25]), .ZN(SUM[25]) );
  NAND2_X1 U60 ( .A1(A[24]), .A2(n89), .ZN(n121) );
  NOR2_X1 U61 ( .A1(n62), .A2(n19), .ZN(n14) );
  OR2_X1 U62 ( .A1(n30), .A2(n132), .ZN(n62) );
  XNOR2_X1 U63 ( .A(A[17]), .B(n122), .ZN(SUM[17]) );
  NAND2_X1 U64 ( .A1(n58), .A2(A[16]), .ZN(n122) );
  NOR3_X1 U65 ( .A1(n134), .A2(n82), .A3(n139), .ZN(n54) );
  INV_X1 U66 ( .A(A[30]), .ZN(n139) );
  AND2_X1 U67 ( .A1(A[3]), .A2(A[2]), .ZN(n18) );
  NAND2_X1 U68 ( .A1(A[19]), .A2(A[18]), .ZN(n96) );
  AND2_X1 U69 ( .A1(A[7]), .A2(A[6]), .ZN(n115) );
  AND2_X1 U70 ( .A1(A[5]), .A2(A[4]), .ZN(n114) );
  XOR2_X1 U71 ( .A(n123), .B(A[30]), .Z(SUM[30]) );
  NOR2_X1 U72 ( .A1(n134), .A2(n82), .ZN(n123) );
  XNOR2_X1 U73 ( .A(n95), .B(A[23]), .ZN(SUM[23]) );
  NAND2_X1 U74 ( .A1(n65), .A2(A[22]), .ZN(n95) );
  AND3_X1 U75 ( .A1(n9), .A2(n45), .A3(A[21]), .ZN(n65) );
  XNOR2_X1 U76 ( .A(n124), .B(A[13]), .ZN(SUM[13]) );
  NAND2_X1 U77 ( .A1(n23), .A2(n12), .ZN(n124) );
  XNOR2_X1 U78 ( .A(n125), .B(A[15]), .ZN(SUM[15]) );
  NAND2_X1 U79 ( .A1(n2), .A2(n109), .ZN(n125) );
  XNOR2_X1 U80 ( .A(n126), .B(A[26]), .ZN(SUM[26]) );
  NAND2_X1 U81 ( .A1(n61), .A2(n4), .ZN(n126) );
  XNOR2_X1 U82 ( .A(n127), .B(A[11]), .ZN(SUM[11]) );
  NAND2_X1 U83 ( .A1(n70), .A2(A[10]), .ZN(n127) );
  XNOR2_X1 U84 ( .A(n128), .B(A[19]), .ZN(SUM[19]) );
  NAND2_X1 U85 ( .A1(n64), .A2(A[18]), .ZN(n128) );
  XNOR2_X1 U87 ( .A(n129), .B(A[27]), .ZN(SUM[27]) );
  NAND2_X1 U88 ( .A1(n61), .A2(n39), .ZN(n129) );
  AND3_X1 U89 ( .A1(n73), .A2(A[9]), .A3(A[8]), .ZN(n70) );
  NOR2_X1 U90 ( .A1(n30), .A2(n132), .ZN(n73) );
  XNOR2_X1 U91 ( .A(n130), .B(A[29]), .ZN(SUM[29]) );
  OR2_X1 U92 ( .A1(n71), .A2(n86), .ZN(n130) );
  AND2_X1 U93 ( .A1(n57), .A2(A[20]), .ZN(n9) );
  INV_X1 U94 ( .A(A[12]), .ZN(n137) );
  AND2_X1 U95 ( .A1(A[2]), .A2(A[3]), .ZN(n79) );
  AND2_X1 U96 ( .A1(n45), .A2(n50), .ZN(n64) );
  AND2_X1 U97 ( .A1(A[16]), .A2(A[17]), .ZN(n50) );
  AND2_X1 U98 ( .A1(A[24]), .A2(A[25]), .ZN(n4) );
  AND2_X1 U99 ( .A1(n47), .A2(A[20]), .ZN(n63) );
  AND3_X1 U100 ( .A1(A[22]), .A2(A[21]), .A3(A[23]), .ZN(n47) );
  INV_X1 U101 ( .A(A[2]), .ZN(SUM[2]) );
endmodule


module Fetch ( CLK, RST, ZERO_FLAG, PC_EXT, INS_IN, Bubble_in, HDU_INS_IN, 
        HDU_PC_IN, HDU_NPC_IN, PC_OUT, ADDR_OUT, NPC_OUT, INS_OUT );
  input [31:0] PC_EXT;
  input [31:0] INS_IN;
  input [31:0] HDU_INS_IN;
  input [31:0] HDU_PC_IN;
  input [31:0] HDU_NPC_IN;
  output [31:0] PC_OUT;
  output [31:0] ADDR_OUT;
  output [31:0] NPC_OUT;
  output [31:0] INS_OUT;
  input CLK, RST, ZERO_FLAG, Bubble_in;
  wire   n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, sig_RST, \sig_NPC[9] ,
         \sig_NPC[8] , \sig_NPC[7] , \sig_NPC[6] , \sig_NPC[5] , \sig_NPC[4] ,
         \sig_NPC[3] , \sig_NPC[31] , \sig_NPC[30] , \sig_NPC[2] ,
         \sig_NPC[29] , \sig_NPC[28] , \sig_NPC[27] , \sig_NPC[26] ,
         \sig_NPC[25] , \sig_NPC[24] , \sig_NPC[23] , \sig_NPC[22] ,
         \sig_NPC[21] , \sig_NPC[20] , \sig_NPC[1] , \sig_NPC[19] ,
         \sig_NPC[18] , \sig_NPC[17] , \sig_NPC[16] , \sig_NPC[15] ,
         \sig_NPC[14] , \sig_NPC[13] , \sig_NPC[12] , \sig_NPC[11] ,
         \sig_NPC[10] , \sig_NPC[0] , \sig_INS[9] , \sig_INS[8] , \sig_INS[7] ,
         \sig_INS[6] , \sig_INS[5] , \sig_INS[4] , \sig_INS[3] , \sig_INS[31] ,
         \sig_INS[30] , \sig_INS[2] , \sig_INS[29] , \sig_INS[28] ,
         \sig_INS[27] , \sig_INS[26] , \sig_INS[25] , \sig_INS[24] ,
         \sig_INS[23] , \sig_INS[22] , \sig_INS[21] , \sig_INS[20] ,
         \sig_INS[1] , \sig_INS[19] , \sig_INS[18] , \sig_INS[17] ,
         \sig_INS[16] , \sig_INS[15] , \sig_INS[14] , \sig_INS[13] ,
         \sig_INS[12] , \sig_INS[11] , \sig_INS[10] , \sig_INS[0] ,
         \PC_MUX_OUT[9] , \PC_MUX_OUT[8] , \PC_MUX_OUT[7] , \PC_MUX_OUT[6] ,
         \PC_MUX_OUT[5] , \PC_MUX_OUT[4] , \PC_MUX_OUT[3] , \PC_MUX_OUT[31] ,
         \PC_MUX_OUT[30] , \PC_MUX_OUT[2] , \PC_MUX_OUT[29] , \PC_MUX_OUT[28] ,
         \PC_MUX_OUT[27] , \PC_MUX_OUT[26] , \PC_MUX_OUT[25] ,
         \PC_MUX_OUT[24] , \PC_MUX_OUT[23] , \PC_MUX_OUT[22] ,
         \PC_MUX_OUT[21] , \PC_MUX_OUT[20] , \PC_MUX_OUT[1] , \PC_MUX_OUT[19] ,
         \PC_MUX_OUT[18] , \PC_MUX_OUT[17] , \PC_MUX_OUT[16] ,
         \PC_MUX_OUT[15] , \PC_MUX_OUT[14] , \PC_MUX_OUT[13] ,
         \PC_MUX_OUT[12] , \PC_MUX_OUT[11] , \PC_MUX_OUT[10] , \PC_MUX_OUT[0] ,
         n49;
  assign ADDR_OUT[27] = n27;
  assign ADDR_OUT[26] = n28;
  assign ADDR_OUT[23] = n29;
  assign ADDR_OUT[22] = n30;
  assign ADDR_OUT[21] = n31;
  assign ADDR_OUT[19] = n32;
  assign ADDR_OUT[18] = n33;
  assign ADDR_OUT[17] = n34;
  assign ADDR_OUT[16] = n35;
  assign ADDR_OUT[15] = n36;
  assign ADDR_OUT[14] = n37;
  assign ADDR_OUT[13] = n38;
  assign ADDR_OUT[11] = n39;
  assign ADDR_OUT[10] = n40;
  assign ADDR_OUT[9] = n41;
  assign ADDR_OUT[8] = n42;
  assign ADDR_OUT[7] = n43;
  assign ADDR_OUT[6] = n44;
  assign ADDR_OUT[5] = n45;
  assign ADDR_OUT[4] = n46;
  assign ADDR_OUT[3] = n47;
  assign ADDR_OUT[2] = n48;

  mux21_NBIT32_0 NPC_or_NPC_HDU ( .A(PC_EXT), .B(HDU_NPC_IN), .S(Bubble_in), 
        .Z({\sig_NPC[31] , \sig_NPC[30] , \sig_NPC[29] , \sig_NPC[28] , 
        \sig_NPC[27] , \sig_NPC[26] , \sig_NPC[25] , \sig_NPC[24] , 
        \sig_NPC[23] , \sig_NPC[22] , \sig_NPC[21] , \sig_NPC[20] , 
        \sig_NPC[19] , \sig_NPC[18] , \sig_NPC[17] , \sig_NPC[16] , 
        \sig_NPC[15] , \sig_NPC[14] , \sig_NPC[13] , \sig_NPC[12] , 
        \sig_NPC[11] , \sig_NPC[10] , \sig_NPC[9] , \sig_NPC[8] , \sig_NPC[7] , 
        \sig_NPC[6] , \sig_NPC[5] , \sig_NPC[4] , \sig_NPC[3] , \sig_NPC[2] , 
        \sig_NPC[1] , \sig_NPC[0] }) );
  mux21_NBIT32_5 PC_or_PC_HDU ( .A({ADDR_OUT[31:28], n27, n28, ADDR_OUT[25:24], 
        n29, n30, n31, ADDR_OUT[20], n32, n33, n34, n35, n36, n37, n38, 
        ADDR_OUT[12], n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
        ADDR_OUT[1:0]}), .B(HDU_PC_IN), .S(Bubble_in), .Z({\PC_MUX_OUT[31] , 
        \PC_MUX_OUT[30] , \PC_MUX_OUT[29] , \PC_MUX_OUT[28] , \PC_MUX_OUT[27] , 
        \PC_MUX_OUT[26] , \PC_MUX_OUT[25] , \PC_MUX_OUT[24] , \PC_MUX_OUT[23] , 
        \PC_MUX_OUT[22] , \PC_MUX_OUT[21] , \PC_MUX_OUT[20] , \PC_MUX_OUT[19] , 
        \PC_MUX_OUT[18] , \PC_MUX_OUT[17] , \PC_MUX_OUT[16] , \PC_MUX_OUT[15] , 
        \PC_MUX_OUT[14] , \PC_MUX_OUT[13] , \PC_MUX_OUT[12] , \PC_MUX_OUT[11] , 
        \PC_MUX_OUT[10] , \PC_MUX_OUT[9] , \PC_MUX_OUT[8] , \PC_MUX_OUT[7] , 
        \PC_MUX_OUT[6] , \PC_MUX_OUT[5] , \PC_MUX_OUT[4] , \PC_MUX_OUT[3] , 
        \PC_MUX_OUT[2] , \PC_MUX_OUT[1] , \PC_MUX_OUT[0] }) );
  mux21_NBIT32_4 INS_or_HDU_INS ( .A(INS_IN), .B(HDU_INS_IN), .S(Bubble_in), 
        .Z({\sig_INS[31] , \sig_INS[30] , \sig_INS[29] , \sig_INS[28] , 
        \sig_INS[27] , \sig_INS[26] , \sig_INS[25] , \sig_INS[24] , 
        \sig_INS[23] , \sig_INS[22] , \sig_INS[21] , \sig_INS[20] , 
        \sig_INS[19] , \sig_INS[18] , \sig_INS[17] , \sig_INS[16] , 
        \sig_INS[15] , \sig_INS[14] , \sig_INS[13] , \sig_INS[12] , 
        \sig_INS[11] , \sig_INS[10] , \sig_INS[9] , \sig_INS[8] , \sig_INS[7] , 
        \sig_INS[6] , \sig_INS[5] , \sig_INS[4] , \sig_INS[3] , \sig_INS[2] , 
        \sig_INS[1] , \sig_INS[0] }) );
  regn_N32_0 PC ( .DIN({\sig_NPC[31] , \sig_NPC[30] , \sig_NPC[29] , 
        \sig_NPC[28] , \sig_NPC[27] , \sig_NPC[26] , \sig_NPC[25] , 
        \sig_NPC[24] , \sig_NPC[23] , \sig_NPC[22] , \sig_NPC[21] , 
        \sig_NPC[20] , \sig_NPC[19] , \sig_NPC[18] , \sig_NPC[17] , 
        \sig_NPC[16] , \sig_NPC[15] , \sig_NPC[14] , \sig_NPC[13] , 
        \sig_NPC[12] , \sig_NPC[11] , \sig_NPC[10] , \sig_NPC[9] , 
        \sig_NPC[8] , \sig_NPC[7] , \sig_NPC[6] , \sig_NPC[5] , \sig_NPC[4] , 
        \sig_NPC[3] , \sig_NPC[2] , \sig_NPC[1] , \sig_NPC[0] }), .CLK(CLK), 
        .EN(1'b1), .RST(RST), .DOUT({ADDR_OUT[31:28], n27, n28, 
        ADDR_OUT[25:24], n29, n30, n31, ADDR_OUT[20], n32, n33, n34, n35, n36, 
        n37, n38, ADDR_OUT[12], n39, n40, n41, n42, n43, n44, n45, n46, n47, 
        n48, ADDR_OUT[1:0]}) );
  regn_N32_10 PC_reg ( .DIN({\PC_MUX_OUT[31] , \PC_MUX_OUT[30] , 
        \PC_MUX_OUT[29] , \PC_MUX_OUT[28] , \PC_MUX_OUT[27] , \PC_MUX_OUT[26] , 
        \PC_MUX_OUT[25] , \PC_MUX_OUT[24] , \PC_MUX_OUT[23] , \PC_MUX_OUT[22] , 
        \PC_MUX_OUT[21] , \PC_MUX_OUT[20] , \PC_MUX_OUT[19] , \PC_MUX_OUT[18] , 
        \PC_MUX_OUT[17] , \PC_MUX_OUT[16] , \PC_MUX_OUT[15] , \PC_MUX_OUT[14] , 
        \PC_MUX_OUT[13] , \PC_MUX_OUT[12] , \PC_MUX_OUT[11] , \PC_MUX_OUT[10] , 
        \PC_MUX_OUT[9] , \PC_MUX_OUT[8] , \PC_MUX_OUT[7] , \PC_MUX_OUT[6] , 
        \PC_MUX_OUT[5] , \PC_MUX_OUT[4] , \PC_MUX_OUT[3] , \PC_MUX_OUT[2] , 
        \PC_MUX_OUT[1] , \PC_MUX_OUT[0] }), .CLK(CLK), .EN(1'b1), .RST(sig_RST), .DOUT(PC_OUT) );
  regn_N32_9 IR ( .DIN({\sig_INS[31] , \sig_INS[30] , \sig_INS[29] , 
        \sig_INS[28] , \sig_INS[27] , \sig_INS[26] , \sig_INS[25] , 
        \sig_INS[24] , \sig_INS[23] , \sig_INS[22] , \sig_INS[21] , 
        \sig_INS[20] , \sig_INS[19] , \sig_INS[18] , \sig_INS[17] , 
        \sig_INS[16] , \sig_INS[15] , \sig_INS[14] , \sig_INS[13] , 
        \sig_INS[12] , \sig_INS[11] , \sig_INS[10] , \sig_INS[9] , 
        \sig_INS[8] , \sig_INS[7] , \sig_INS[6] , \sig_INS[5] , \sig_INS[4] , 
        \sig_INS[3] , \sig_INS[2] , \sig_INS[1] , \sig_INS[0] }), .CLK(CLK), 
        .EN(1'b1), .RST(sig_RST), .DOUT(INS_OUT) );
  Fetch_DW01_add_3 add_54 ( .A({ADDR_OUT[31:28], n27, n28, ADDR_OUT[25:24], 
        n29, n30, n31, ADDR_OUT[20], n32, n33, n34, n35, n36, n37, n38, 
        ADDR_OUT[12], n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
        ADDR_OUT[1:0]}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(NPC_OUT) );
  NOR2_X1 U3 ( .A1(ZERO_FLAG), .A2(n49), .ZN(sig_RST) );
  INV_X1 U4 ( .A(RST), .ZN(n49) );
endmodule


module instruction_type ( INST_IN, Rtype, Itype, Jtype );
  input [31:0] INST_IN;
  output Rtype, Itype, Jtype;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  NAND3_X1 U15 ( .A1(INST_IN[26]), .A2(n14), .A3(INST_IN[30]), .ZN(n12) );
  NOR2_X1 U1 ( .A1(n4), .A2(n14), .ZN(Jtype) );
  NOR3_X1 U2 ( .A1(n4), .A2(INST_IN[27]), .A3(INST_IN[26]), .ZN(Rtype) );
  OAI21_X1 U3 ( .B1(INST_IN[31]), .B2(n5), .A(n6), .ZN(Itype) );
  NAND4_X1 U4 ( .A1(INST_IN[31]), .A2(INST_IN[26]), .A3(n7), .A4(INST_IN[27]), 
        .ZN(n6) );
  AOI21_X1 U5 ( .B1(INST_IN[29]), .B2(n8), .A(n13), .ZN(n5) );
  NOR2_X1 U6 ( .A1(INST_IN[30]), .A2(INST_IN[28]), .ZN(n7) );
  OAI21_X1 U7 ( .B1(INST_IN[30]), .B2(INST_IN[26]), .A(n12), .ZN(n8) );
  OR4_X1 U8 ( .A1(INST_IN[28]), .A2(INST_IN[29]), .A3(INST_IN[30]), .A4(
        INST_IN[31]), .ZN(n4) );
  INV_X1 U9 ( .A(INST_IN[27]), .ZN(n14) );
  INV_X1 U10 ( .A(n9), .ZN(n13) );
  OAI21_X1 U11 ( .B1(n10), .B2(n11), .A(INST_IN[28]), .ZN(n9) );
  AOI21_X1 U12 ( .B1(INST_IN[26]), .B2(INST_IN[30]), .A(INST_IN[27]), .ZN(n10)
         );
  NOR3_X1 U13 ( .A1(INST_IN[26]), .A2(INST_IN[29]), .A3(n15), .ZN(n11) );
  INV_X1 U14 ( .A(INST_IN[30]), .ZN(n15) );
endmodule


module instruction_decomposition ( INST_IN, Rtype, Itype, Jtype, ADD_RS1, 
        ADD_RS2, ADD_WR, IMM );
  input [31:0] INST_IN;
  output [4:0] ADD_RS1;
  output [4:0] ADD_RS2;
  output [4:0] ADD_WR;
  output [31:0] IMM;
  input Rtype, Itype, Jtype;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, \IMM[31] , n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45;
  assign IMM[25] = \IMM[31] ;
  assign IMM[26] = \IMM[31] ;
  assign IMM[27] = \IMM[31] ;
  assign IMM[28] = \IMM[31] ;
  assign IMM[29] = \IMM[31] ;
  assign IMM[30] = \IMM[31] ;
  assign IMM[31] = \IMM[31] ;

  NAND3_X1 U68 ( .A1(INST_IN[29]), .A2(INST_IN[27]), .A3(INST_IN[31]), .ZN(n26) );
  NAND3_X1 U69 ( .A1(INST_IN[26]), .A2(Itype), .A3(n27), .ZN(n25) );
  NOR2_X1 U2 ( .A1(n43), .A2(n37), .ZN(ADD_RS2[4]) );
  NOR2_X1 U3 ( .A1(n23), .A2(n42), .ZN(ADD_RS1[4]) );
  NAND2_X1 U4 ( .A1(Jtype), .A2(n23), .ZN(n19) );
  INV_X1 U5 ( .A(n22), .ZN(n44) );
  NOR2_X1 U6 ( .A1(n23), .A2(n41), .ZN(ADD_RS1[3]) );
  NOR2_X1 U7 ( .A1(n43), .A2(n36), .ZN(ADD_RS2[3]) );
  NOR2_X1 U8 ( .A1(n23), .A2(n38), .ZN(ADD_RS1[0]) );
  NOR2_X1 U9 ( .A1(n43), .A2(n33), .ZN(ADD_RS2[0]) );
  OAI21_X1 U10 ( .B1(Jtype), .B2(Itype), .A(n45), .ZN(n22) );
  NOR2_X1 U11 ( .A1(Itype), .A2(Rtype), .ZN(n23) );
  NOR2_X1 U12 ( .A1(n23), .A2(n39), .ZN(ADD_RS1[1]) );
  NOR2_X1 U13 ( .A1(n43), .A2(n34), .ZN(ADD_RS2[1]) );
  NOR2_X1 U14 ( .A1(n23), .A2(n40), .ZN(ADD_RS1[2]) );
  NOR2_X1 U15 ( .A1(n43), .A2(n35), .ZN(ADD_RS2[2]) );
  OR2_X1 U16 ( .A1(n32), .A2(n21), .ZN(n20) );
  INV_X1 U17 ( .A(Rtype), .ZN(n45) );
  NAND2_X1 U18 ( .A1(Itype), .A2(n45), .ZN(n21) );
  OAI221_X1 U19 ( .B1(n21), .B2(n33), .C1(n28), .C2(n45), .A(n19), .ZN(
        ADD_WR[0]) );
  OAI221_X1 U20 ( .B1(n21), .B2(n34), .C1(n29), .C2(n45), .A(n19), .ZN(
        ADD_WR[1]) );
  OAI221_X1 U21 ( .B1(n21), .B2(n35), .C1(n30), .C2(n45), .A(n19), .ZN(
        ADD_WR[2]) );
  OAI221_X1 U22 ( .B1(n21), .B2(n36), .C1(n31), .C2(n45), .A(n19), .ZN(
        ADD_WR[3]) );
  OAI221_X1 U23 ( .B1(n21), .B2(n37), .C1(n32), .C2(n45), .A(n19), .ZN(
        ADD_WR[4]) );
  OAI21_X1 U24 ( .B1(n19), .B2(n42), .A(n20), .ZN(\IMM[31] ) );
  OAI21_X1 U25 ( .B1(n19), .B2(n33), .A(n20), .ZN(IMM[16]) );
  OAI21_X1 U26 ( .B1(n19), .B2(n34), .A(n20), .ZN(IMM[17]) );
  OAI21_X1 U27 ( .B1(n19), .B2(n35), .A(n20), .ZN(IMM[18]) );
  OAI21_X1 U28 ( .B1(n19), .B2(n36), .A(n20), .ZN(IMM[19]) );
  OAI21_X1 U29 ( .B1(n19), .B2(n37), .A(n20), .ZN(IMM[20]) );
  OAI21_X1 U30 ( .B1(n19), .B2(n38), .A(n20), .ZN(IMM[21]) );
  OAI21_X1 U31 ( .B1(n19), .B2(n39), .A(n20), .ZN(IMM[22]) );
  OAI21_X1 U32 ( .B1(n19), .B2(n40), .A(n20), .ZN(IMM[23]) );
  OAI21_X1 U33 ( .B1(n19), .B2(n41), .A(n20), .ZN(IMM[24]) );
  NOR2_X1 U34 ( .A1(n32), .A2(n22), .ZN(IMM[15]) );
  NOR2_X1 U35 ( .A1(n22), .A2(n28), .ZN(IMM[11]) );
  NOR2_X1 U36 ( .A1(n22), .A2(n29), .ZN(IMM[12]) );
  NOR2_X1 U37 ( .A1(n22), .A2(n30), .ZN(IMM[13]) );
  NOR2_X1 U38 ( .A1(n22), .A2(n31), .ZN(IMM[14]) );
  INV_X1 U39 ( .A(n24), .ZN(n43) );
  OAI21_X1 U40 ( .B1(n25), .B2(n26), .A(n45), .ZN(n24) );
  INV_X1 U41 ( .A(INST_IN[16]), .ZN(n33) );
  INV_X1 U42 ( .A(INST_IN[17]), .ZN(n34) );
  INV_X1 U43 ( .A(INST_IN[18]), .ZN(n35) );
  INV_X1 U44 ( .A(INST_IN[19]), .ZN(n36) );
  INV_X1 U45 ( .A(INST_IN[20]), .ZN(n37) );
  INV_X1 U46 ( .A(INST_IN[15]), .ZN(n32) );
  NOR2_X1 U47 ( .A1(INST_IN[30]), .A2(INST_IN[28]), .ZN(n27) );
  INV_X1 U48 ( .A(INST_IN[21]), .ZN(n38) );
  INV_X1 U49 ( .A(INST_IN[22]), .ZN(n39) );
  INV_X1 U50 ( .A(INST_IN[23]), .ZN(n40) );
  INV_X1 U51 ( .A(INST_IN[24]), .ZN(n41) );
  INV_X1 U52 ( .A(INST_IN[25]), .ZN(n42) );
  INV_X1 U53 ( .A(INST_IN[11]), .ZN(n28) );
  INV_X1 U54 ( .A(INST_IN[12]), .ZN(n29) );
  INV_X1 U55 ( .A(INST_IN[13]), .ZN(n30) );
  INV_X1 U56 ( .A(INST_IN[14]), .ZN(n31) );
  AND2_X1 U57 ( .A1(INST_IN[0]), .A2(n44), .ZN(IMM[0]) );
  AND2_X1 U58 ( .A1(INST_IN[1]), .A2(n44), .ZN(IMM[1]) );
  AND2_X1 U59 ( .A1(INST_IN[2]), .A2(n44), .ZN(IMM[2]) );
  AND2_X1 U60 ( .A1(INST_IN[3]), .A2(n44), .ZN(IMM[3]) );
  AND2_X1 U61 ( .A1(INST_IN[4]), .A2(n44), .ZN(IMM[4]) );
  AND2_X1 U62 ( .A1(INST_IN[5]), .A2(n44), .ZN(IMM[5]) );
  AND2_X1 U63 ( .A1(INST_IN[6]), .A2(n44), .ZN(IMM[6]) );
  AND2_X1 U64 ( .A1(INST_IN[7]), .A2(n44), .ZN(IMM[7]) );
  AND2_X1 U65 ( .A1(INST_IN[8]), .A2(n44), .ZN(IMM[8]) );
  AND2_X1 U66 ( .A1(INST_IN[9]), .A2(n44), .ZN(IMM[9]) );
  AND2_X1 U67 ( .A1(INST_IN[10]), .A2(n44), .ZN(IMM[10]) );
endmodule


module register_file_NBIT_ADD5_NBIT_DATA32 ( CLK, RST, ENABLE, RD1, RD2, WR, 
        ADD_WR, ADD_RS1, ADD_RS2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RST, ENABLE, RD1, RD2, WR;
  wire   n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3174, n3175, n3176, n3177, n3178, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n938, n939, n950, n955, n956, n966, n971,
         n972, n982, n987, n988, n998, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n749,
         n824, n825, n826, n834, n835, n836, n837, n838, n840, n841, n842,
         n843, n844, n845, n847, n848, n849, n871, n872, n873, n876, n877,
         n878, n888, n889, n890, n893, n894, n895, n905, n906, n907, n910,
         n911, n912, n922, n923, n924, n927, n928, n929, n941, n942, n943,
         n946, n947, n948, n961, n962, n963, n967, n968, n969, n981, n983,
         n984, n989, n990, n991, n1002, n1003, n1004, n1007, n1008, n1009,
         n1019, n1020, n1021, n1024, n1025, n1026, n1036, n1037, n1038, n1041,
         n1042, n1043, n1053, n1054, n1055, n1058, n1059, n1060, n1070, n1071,
         n1072, n1075, n1076, n1077, n1087, n1088, n1089, n1092, n1093, n1094,
         n1104, n1105, n1106, n1109, n1110, n1111, n1121, n1122, n1123, n1126,
         n1127, n1128, n1138, n1139, n1140, n1143, n1144, n1145, n1155, n1156,
         n1157, n1160, n1161, n1162, n1172, n1173, n1174, n1177, n1178, n1179,
         n1189, n1190, n1191, n1194, n1195, n1196, n1206, n1207, n1208, n1211,
         n1212, n1213, n1223, n1224, n1225, n1228, n1229, n1230, n1240, n1241,
         n1242, n1245, n1246, n1247, n1257, n1258, n1259, n1262, n1263, n1264,
         n1274, n1275, n1276, n1279, n1280, n1281, n1291, n1292, n1293, n1296,
         n1297, n1298, n1308, n1309, n1310, n1313, n1314, n1315, n1325, n1326,
         n1327, n1330, n1331, n1332, n1342, n1343, n1344, n1347, n1348, n1349,
         n1359, n1360, n1361, n1364, n1365, n1366, n1376, n1377, n1378, n1381,
         n1382, n1383, n1393, n1394, n1397, n1398, n1399, n1400, n1401, n1402,
         n1406, n1412, n1413, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1427, n1437, n1438, n1439, n1447, n1448, n1449, n1450, n1451, n1453,
         n1454, n1455, n1456, n1457, n1458, n1460, n1461, n1462, n1481, n1482,
         n1483, n1486, n1487, n1488, n1498, n1499, n1500, n1503, n1504, n1505,
         n1515, n1516, n1517, n1520, n1521, n1522, n1532, n1533, n1534, n1537,
         n1538, n1539, n1549, n1550, n1551, n1554, n1555, n1556, n1566, n1567,
         n1568, n1571, n1572, n1573, n1583, n1584, n1585, n1588, n1589, n1590,
         n1600, n1601, n1602, n1605, n1606, n1607, n1617, n1618, n1619, n1622,
         n1623, n1624, n1634, n1635, n1636, n1639, n1640, n1641, n1651, n1652,
         n1653, n1656, n1657, n1658, n1668, n1669, n1670, n1673, n1674, n1675,
         n1685, n1686, n1687, n1690, n1691, n1692, n1702, n1703, n1704, n1707,
         n1708, n1709, n1719, n1720, n1721, n1724, n1725, n1726, n1736, n1737,
         n1738, n1741, n1742, n1743, n1753, n1754, n1755, n1758, n1759, n1760,
         n1770, n1771, n1772, n1775, n1776, n1777, n1787, n1788, n1789, n1792,
         n1793, n1794, n1804, n1805, n1806, n1809, n1810, n1811, n1821, n1822,
         n1823, n1826, n1827, n1828, n1838, n1839, n1840, n1843, n1844, n1845,
         n1855, n1856, n1857, n1860, n1861, n1862, n1872, n1873, n1874, n1877,
         n1878, n1879, n1889, n1890, n1891, n1894, n1895, n1896, n1906, n1907,
         n1908, n1911, n1912, n1913, n1923, n1924, n1925, n1928, n1929, n1930,
         n1940, n1941, n1942, n1945, n1946, n1947, n1957, n1958, n1959, n1962,
         n1963, n1964, n1974, n1975, n1976, n1979, n1980, n1981, n1993, n1994,
         n1997, n1998, n1999, n2000, n2001, n2002, n2006, n2012, n2013, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902;

  DFFR_X1 \REGISTERS_reg[10][31]  ( .D(n3430), .CK(CLK), .RN(n6444), .Q(n5712), 
        .QN(n2318) );
  DFFR_X1 \REGISTERS_reg[10][30]  ( .D(n3429), .CK(CLK), .RN(n6444), .Q(n5713), 
        .QN(n2322) );
  DFFR_X1 \REGISTERS_reg[10][29]  ( .D(n3428), .CK(CLK), .RN(n6444), .Q(n5714), 
        .QN(n2326) );
  DFFR_X1 \REGISTERS_reg[10][28]  ( .D(n3427), .CK(CLK), .RN(n6444), .Q(n5715), 
        .QN(n2330) );
  DFFR_X1 \REGISTERS_reg[10][27]  ( .D(n3426), .CK(CLK), .RN(n6445), .Q(n5716), 
        .QN(n2334) );
  DFFR_X1 \REGISTERS_reg[10][26]  ( .D(n3425), .CK(CLK), .RN(n6445), .Q(n5717), 
        .QN(n2338) );
  DFFR_X1 \REGISTERS_reg[10][25]  ( .D(n3424), .CK(CLK), .RN(n6445), .Q(n5718), 
        .QN(n2342) );
  DFFR_X1 \REGISTERS_reg[10][24]  ( .D(n3423), .CK(CLK), .RN(n6445), .Q(n5719), 
        .QN(n2346) );
  DFFR_X1 \REGISTERS_reg[10][23]  ( .D(n3422), .CK(CLK), .RN(n6445), .Q(n5720), 
        .QN(n2350) );
  DFFR_X1 \REGISTERS_reg[10][22]  ( .D(n3421), .CK(CLK), .RN(n6445), .Q(n5721), 
        .QN(n2354) );
  DFFR_X1 \REGISTERS_reg[10][21]  ( .D(n3420), .CK(CLK), .RN(n6445), .Q(n5722), 
        .QN(n2358) );
  DFFR_X1 \REGISTERS_reg[10][20]  ( .D(n3419), .CK(CLK), .RN(n6445), .Q(n5723), 
        .QN(n2362) );
  DFFR_X1 \REGISTERS_reg[10][19]  ( .D(n3418), .CK(CLK), .RN(n6443), .Q(n5724), 
        .QN(n2366) );
  DFFR_X1 \REGISTERS_reg[10][18]  ( .D(n3417), .CK(CLK), .RN(n6443), .Q(n5725), 
        .QN(n2370) );
  DFFR_X1 \REGISTERS_reg[10][17]  ( .D(n3416), .CK(CLK), .RN(n6443), .Q(n5726), 
        .QN(n2374) );
  DFFR_X1 \REGISTERS_reg[10][16]  ( .D(n3415), .CK(CLK), .RN(n6443), .Q(n5727), 
        .QN(n2378) );
  DFFR_X1 \REGISTERS_reg[10][15]  ( .D(n3414), .CK(CLK), .RN(n6444), .Q(n5728), 
        .QN(n2382) );
  DFFR_X1 \REGISTERS_reg[10][14]  ( .D(n3413), .CK(CLK), .RN(n6444), .Q(n5729), 
        .QN(n2386) );
  DFFR_X1 \REGISTERS_reg[10][13]  ( .D(n3412), .CK(CLK), .RN(n6444), .Q(n5730), 
        .QN(n2390) );
  DFFR_X1 \REGISTERS_reg[10][12]  ( .D(n3411), .CK(CLK), .RN(n6444), .Q(n5731), 
        .QN(n2394) );
  DFFR_X1 \REGISTERS_reg[10][11]  ( .D(n3410), .CK(CLK), .RN(n6444), .Q(n5732), 
        .QN(n2398) );
  DFFR_X1 \REGISTERS_reg[10][10]  ( .D(n3409), .CK(CLK), .RN(n6444), .Q(n5733), 
        .QN(n2402) );
  DFFR_X1 \REGISTERS_reg[10][9]  ( .D(n3408), .CK(CLK), .RN(n6444), .Q(n5734), 
        .QN(n2406) );
  DFFR_X1 \REGISTERS_reg[10][8]  ( .D(n3407), .CK(CLK), .RN(n6444), .Q(n5735), 
        .QN(n2410) );
  DFFR_X1 \REGISTERS_reg[10][7]  ( .D(n3406), .CK(CLK), .RN(n6443), .Q(n5736), 
        .QN(n2414) );
  DFFR_X1 \REGISTERS_reg[10][6]  ( .D(n3405), .CK(CLK), .RN(n6443), .Q(n5737), 
        .QN(n2418) );
  DFFR_X1 \REGISTERS_reg[10][5]  ( .D(n3404), .CK(CLK), .RN(n6443), .Q(n5738), 
        .QN(n2422) );
  DFFR_X1 \REGISTERS_reg[10][4]  ( .D(n3403), .CK(CLK), .RN(n6443), .Q(n5739), 
        .QN(n2426) );
  DFFR_X1 \REGISTERS_reg[10][3]  ( .D(n3402), .CK(CLK), .RN(n6443), .Q(n5740), 
        .QN(n2430) );
  DFFR_X1 \REGISTERS_reg[10][2]  ( .D(n3401), .CK(CLK), .RN(n6443), .Q(n5741), 
        .QN(n2434) );
  DFFR_X1 \REGISTERS_reg[10][1]  ( .D(n3400), .CK(CLK), .RN(n6443), .Q(n5742), 
        .QN(n2438) );
  DFFR_X1 \REGISTERS_reg[10][0]  ( .D(n3399), .CK(CLK), .RN(n6443), .Q(n5743), 
        .QN(n2442) );
  DFFR_X1 \REGISTERS_reg[11][31]  ( .D(n3398), .CK(CLK), .RN(n6442), .Q(n5548), 
        .QN(n2319) );
  DFFR_X1 \REGISTERS_reg[11][30]  ( .D(n3397), .CK(CLK), .RN(n6442), .Q(n5549), 
        .QN(n2323) );
  DFFR_X1 \REGISTERS_reg[11][29]  ( .D(n3396), .CK(CLK), .RN(n6442), .Q(n5550), 
        .QN(n2327) );
  DFFR_X1 \REGISTERS_reg[11][28]  ( .D(n3395), .CK(CLK), .RN(n6442), .Q(n5551), 
        .QN(n2331) );
  DFFR_X1 \REGISTERS_reg[11][27]  ( .D(n3394), .CK(CLK), .RN(n6441), .Q(n5552), 
        .QN(n2335) );
  DFFR_X1 \REGISTERS_reg[11][26]  ( .D(n3393), .CK(CLK), .RN(n6441), .Q(n5553), 
        .QN(n2339) );
  DFFR_X1 \REGISTERS_reg[11][25]  ( .D(n3392), .CK(CLK), .RN(n6441), .Q(n5554), 
        .QN(n2343) );
  DFFR_X1 \REGISTERS_reg[11][24]  ( .D(n3391), .CK(CLK), .RN(n6441), .Q(n5555), 
        .QN(n2347) );
  DFFR_X1 \REGISTERS_reg[11][23]  ( .D(n3390), .CK(CLK), .RN(n6442), .Q(n5556), 
        .QN(n2351) );
  DFFR_X1 \REGISTERS_reg[11][22]  ( .D(n3389), .CK(CLK), .RN(n6442), .Q(n5557), 
        .QN(n2355) );
  DFFR_X1 \REGISTERS_reg[11][21]  ( .D(n3388), .CK(CLK), .RN(n6442), .Q(n5558), 
        .QN(n2359) );
  DFFR_X1 \REGISTERS_reg[11][20]  ( .D(n3387), .CK(CLK), .RN(n6442), .Q(n5559), 
        .QN(n2363) );
  DFFR_X1 \REGISTERS_reg[11][19]  ( .D(n3386), .CK(CLK), .RN(n6442), .Q(n5560), 
        .QN(n2367) );
  DFFR_X1 \REGISTERS_reg[11][18]  ( .D(n3385), .CK(CLK), .RN(n6442), .Q(n5561), 
        .QN(n2371) );
  DFFR_X1 \REGISTERS_reg[11][17]  ( .D(n3384), .CK(CLK), .RN(n6442), .Q(n5562), 
        .QN(n2375) );
  DFFR_X1 \REGISTERS_reg[11][16]  ( .D(n3383), .CK(CLK), .RN(n6442), .Q(n5563), 
        .QN(n2379) );
  DFFR_X1 \REGISTERS_reg[11][15]  ( .D(n3382), .CK(CLK), .RN(n6440), .Q(n5564), 
        .QN(n2383) );
  DFFR_X1 \REGISTERS_reg[11][14]  ( .D(n3381), .CK(CLK), .RN(n6440), .Q(n5565), 
        .QN(n2387) );
  DFFR_X1 \REGISTERS_reg[11][13]  ( .D(n3380), .CK(CLK), .RN(n6440), .Q(n5566), 
        .QN(n2391) );
  DFFR_X1 \REGISTERS_reg[11][12]  ( .D(n3379), .CK(CLK), .RN(n6440), .Q(n5567), 
        .QN(n2395) );
  DFFR_X1 \REGISTERS_reg[11][11]  ( .D(n3378), .CK(CLK), .RN(n6441), .Q(n5568), 
        .QN(n2399) );
  DFFR_X1 \REGISTERS_reg[11][10]  ( .D(n3377), .CK(CLK), .RN(n6441), .Q(n5569), 
        .QN(n2403) );
  DFFR_X1 \REGISTERS_reg[11][9]  ( .D(n3376), .CK(CLK), .RN(n6441), .Q(n5570), 
        .QN(n2407) );
  DFFR_X1 \REGISTERS_reg[11][8]  ( .D(n3375), .CK(CLK), .RN(n6441), .Q(n5571), 
        .QN(n2411) );
  DFFR_X1 \REGISTERS_reg[11][7]  ( .D(n3374), .CK(CLK), .RN(n6441), .Q(n5572), 
        .QN(n2415) );
  DFFR_X1 \REGISTERS_reg[11][6]  ( .D(n3373), .CK(CLK), .RN(n6441), .Q(n5573), 
        .QN(n2419) );
  DFFR_X1 \REGISTERS_reg[11][5]  ( .D(n3372), .CK(CLK), .RN(n6441), .Q(n5574), 
        .QN(n2423) );
  DFFR_X1 \REGISTERS_reg[11][4]  ( .D(n3371), .CK(CLK), .RN(n6441), .Q(n5575), 
        .QN(n2427) );
  DFFR_X1 \REGISTERS_reg[11][3]  ( .D(n3370), .CK(CLK), .RN(n6452), .Q(n5576), 
        .QN(n2431) );
  DFFR_X1 \REGISTERS_reg[11][2]  ( .D(n3369), .CK(CLK), .RN(n6452), .Q(n5577), 
        .QN(n2435) );
  DFFR_X1 \REGISTERS_reg[11][1]  ( .D(n3368), .CK(CLK), .RN(n6452), .Q(n5578), 
        .QN(n2439) );
  DFFR_X1 \REGISTERS_reg[11][0]  ( .D(n3367), .CK(CLK), .RN(n6452), .Q(n5579), 
        .QN(n2443) );
  DFFR_X1 \REGISTERS_reg[14][31]  ( .D(n3366), .CK(CLK), .RN(n6447), .Q(n5236), 
        .QN(n2316) );
  DFFR_X1 \REGISTERS_reg[14][30]  ( .D(n3365), .CK(CLK), .RN(n6447), .Q(n5238), 
        .QN(n2320) );
  DFFR_X1 \REGISTERS_reg[14][29]  ( .D(n3364), .CK(CLK), .RN(n6447), .Q(n5239), 
        .QN(n2324) );
  DFFR_X1 \REGISTERS_reg[14][28]  ( .D(n3363), .CK(CLK), .RN(n6447), .Q(n5240), 
        .QN(n2328) );
  DFFR_X1 \REGISTERS_reg[14][27]  ( .D(n3362), .CK(CLK), .RN(n6457), .Q(n5241), 
        .QN(n2332) );
  DFFR_X1 \REGISTERS_reg[14][26]  ( .D(n3361), .CK(CLK), .RN(n6457), .Q(n5242), 
        .QN(n2336) );
  DFFR_X1 \REGISTERS_reg[14][25]  ( .D(n3360), .CK(CLK), .RN(n6457), .Q(n5243), 
        .QN(n2340) );
  DFFR_X1 \REGISTERS_reg[14][24]  ( .D(n3359), .CK(CLK), .RN(n6457), .Q(n5244), 
        .QN(n2344) );
  DFFR_X1 \REGISTERS_reg[14][23]  ( .D(n3358), .CK(CLK), .RN(n6458), .Q(n5245), 
        .QN(n2348) );
  DFFR_X1 \REGISTERS_reg[14][22]  ( .D(n3357), .CK(CLK), .RN(n6458), .Q(n5246), 
        .QN(n2352) );
  DFFR_X1 \REGISTERS_reg[14][21]  ( .D(n3356), .CK(CLK), .RN(n6458), .Q(n5247), 
        .QN(n2356) );
  DFFR_X1 \REGISTERS_reg[14][20]  ( .D(n3355), .CK(CLK), .RN(n6458), .Q(n5248), 
        .QN(n2360) );
  DFFR_X1 \REGISTERS_reg[14][19]  ( .D(n3354), .CK(CLK), .RN(n6458), .Q(n5249), 
        .QN(n2364) );
  DFFR_X1 \REGISTERS_reg[14][18]  ( .D(n3353), .CK(CLK), .RN(n6458), .Q(n5250), 
        .QN(n2368) );
  DFFR_X1 \REGISTERS_reg[14][17]  ( .D(n3352), .CK(CLK), .RN(n6458), .Q(n5251), 
        .QN(n2372) );
  DFFR_X1 \REGISTERS_reg[14][16]  ( .D(n3351), .CK(CLK), .RN(n6458), .Q(n5252), 
        .QN(n2376) );
  DFFR_X1 \REGISTERS_reg[14][15]  ( .D(n3350), .CK(CLK), .RN(n6456), .Q(n5253), 
        .QN(n2380) );
  DFFR_X1 \REGISTERS_reg[14][14]  ( .D(n3349), .CK(CLK), .RN(n6456), .Q(n5254), 
        .QN(n2384) );
  DFFR_X1 \REGISTERS_reg[14][13]  ( .D(n3348), .CK(CLK), .RN(n6456), .Q(n5255), 
        .QN(n2388) );
  DFFR_X1 \REGISTERS_reg[14][12]  ( .D(n3347), .CK(CLK), .RN(n6456), .Q(n5256), 
        .QN(n2392) );
  DFFR_X1 \REGISTERS_reg[14][11]  ( .D(n3346), .CK(CLK), .RN(n6457), .Q(n5257), 
        .QN(n2396) );
  DFFR_X1 \REGISTERS_reg[14][10]  ( .D(n3345), .CK(CLK), .RN(n6457), .Q(n5258), 
        .QN(n2400) );
  DFFR_X1 \REGISTERS_reg[14][9]  ( .D(n3344), .CK(CLK), .RN(n6457), .Q(n5259), 
        .QN(n2404) );
  DFFR_X1 \REGISTERS_reg[14][8]  ( .D(n3343), .CK(CLK), .RN(n6457), .Q(n5260), 
        .QN(n2408) );
  DFFR_X1 \REGISTERS_reg[14][7]  ( .D(n3342), .CK(CLK), .RN(n6457), .Q(n5261), 
        .QN(n2412) );
  DFFR_X1 \REGISTERS_reg[14][6]  ( .D(n3341), .CK(CLK), .RN(n6457), .Q(n5262), 
        .QN(n2416) );
  DFFR_X1 \REGISTERS_reg[14][5]  ( .D(n3340), .CK(CLK), .RN(n6457), .Q(n5263), 
        .QN(n2420) );
  DFFR_X1 \REGISTERS_reg[14][4]  ( .D(n3339), .CK(CLK), .RN(n6457), .Q(n5264), 
        .QN(n2424) );
  DFFR_X1 \REGISTERS_reg[14][3]  ( .D(n3338), .CK(CLK), .RN(n6456), .Q(n5265), 
        .QN(n2428) );
  DFFR_X1 \REGISTERS_reg[14][2]  ( .D(n3337), .CK(CLK), .RN(n6456), .Q(n5266), 
        .QN(n2432) );
  DFFR_X1 \REGISTERS_reg[14][1]  ( .D(n3336), .CK(CLK), .RN(n6456), .Q(n5267), 
        .QN(n2436) );
  DFFR_X1 \REGISTERS_reg[14][0]  ( .D(n3335), .CK(CLK), .RN(n6456), .Q(n5237), 
        .QN(n2440) );
  DFFR_X1 \REGISTERS_reg[15][31]  ( .D(n3334), .CK(CLK), .RN(n6455), .Q(n5745), 
        .QN(n2317) );
  DFFR_X1 \REGISTERS_reg[15][30]  ( .D(n3333), .CK(CLK), .RN(n6455), .Q(n5746), 
        .QN(n2321) );
  DFFR_X1 \REGISTERS_reg[15][29]  ( .D(n3332), .CK(CLK), .RN(n6455), .Q(n5747), 
        .QN(n2325) );
  DFFR_X1 \REGISTERS_reg[15][28]  ( .D(n3331), .CK(CLK), .RN(n6455), .Q(n5748), 
        .QN(n2329) );
  DFFR_X1 \REGISTERS_reg[15][27]  ( .D(n3330), .CK(CLK), .RN(n6456), .Q(n5749), 
        .QN(n2333) );
  DFFR_X1 \REGISTERS_reg[15][26]  ( .D(n3329), .CK(CLK), .RN(n6456), .Q(n5750), 
        .QN(n2337) );
  DFFR_X1 \REGISTERS_reg[15][25]  ( .D(n3328), .CK(CLK), .RN(n6456), .Q(n5751), 
        .QN(n2341) );
  DFFR_X1 \REGISTERS_reg[15][24]  ( .D(n3327), .CK(CLK), .RN(n6456), .Q(n5752), 
        .QN(n2345) );
  DFFR_X1 \REGISTERS_reg[15][23]  ( .D(n3326), .CK(CLK), .RN(n6454), .Q(n5753), 
        .QN(n2349) );
  DFFR_X1 \REGISTERS_reg[15][22]  ( .D(n3325), .CK(CLK), .RN(n6454), .Q(n5754), 
        .QN(n2353) );
  DFFR_X1 \REGISTERS_reg[15][21]  ( .D(n3324), .CK(CLK), .RN(n6454), .Q(n5755), 
        .QN(n2357) );
  DFFR_X1 \REGISTERS_reg[15][20]  ( .D(n3323), .CK(CLK), .RN(n6454), .Q(n5756), 
        .QN(n2361) );
  DFFR_X1 \REGISTERS_reg[15][19]  ( .D(n3322), .CK(CLK), .RN(n6455), .Q(n5757), 
        .QN(n2365) );
  DFFR_X1 \REGISTERS_reg[15][18]  ( .D(n3321), .CK(CLK), .RN(n6455), .Q(n5758), 
        .QN(n2369) );
  DFFR_X1 \REGISTERS_reg[15][17]  ( .D(n3320), .CK(CLK), .RN(n6455), .Q(n5759), 
        .QN(n2373) );
  DFFR_X1 \REGISTERS_reg[15][16]  ( .D(n3319), .CK(CLK), .RN(n6455), .Q(n5760), 
        .QN(n2377) );
  DFFR_X1 \REGISTERS_reg[15][15]  ( .D(n3318), .CK(CLK), .RN(n6455), .Q(n5761), 
        .QN(n2381) );
  DFFR_X1 \REGISTERS_reg[15][14]  ( .D(n3317), .CK(CLK), .RN(n6455), .Q(n5762), 
        .QN(n2385) );
  DFFR_X1 \REGISTERS_reg[15][13]  ( .D(n3316), .CK(CLK), .RN(n6455), .Q(n5763), 
        .QN(n2389) );
  DFFR_X1 \REGISTERS_reg[15][12]  ( .D(n3315), .CK(CLK), .RN(n6455), .Q(n5764), 
        .QN(n2393) );
  DFFR_X1 \REGISTERS_reg[15][11]  ( .D(n3314), .CK(CLK), .RN(n6453), .Q(n5765), 
        .QN(n2397) );
  DFFR_X1 \REGISTERS_reg[15][10]  ( .D(n3313), .CK(CLK), .RN(n6453), .Q(n5766), 
        .QN(n2401) );
  DFFR_X1 \REGISTERS_reg[15][9]  ( .D(n3312), .CK(CLK), .RN(n6453), .Q(n5767), 
        .QN(n2405) );
  DFFR_X1 \REGISTERS_reg[15][8]  ( .D(n3311), .CK(CLK), .RN(n6453), .Q(n5768), 
        .QN(n2409) );
  DFFR_X1 \REGISTERS_reg[15][7]  ( .D(n3310), .CK(CLK), .RN(n6454), .Q(n5769), 
        .QN(n2413) );
  DFFR_X1 \REGISTERS_reg[15][6]  ( .D(n3309), .CK(CLK), .RN(n6454), .Q(n5770), 
        .QN(n2417) );
  DFFR_X1 \REGISTERS_reg[15][5]  ( .D(n3308), .CK(CLK), .RN(n6454), .Q(n5771), 
        .QN(n2421) );
  DFFR_X1 \REGISTERS_reg[15][4]  ( .D(n3307), .CK(CLK), .RN(n6454), .Q(n5772), 
        .QN(n2425) );
  DFFR_X1 \REGISTERS_reg[15][3]  ( .D(n3306), .CK(CLK), .RN(n6454), .Q(n5773), 
        .QN(n2429) );
  DFFR_X1 \REGISTERS_reg[15][2]  ( .D(n3305), .CK(CLK), .RN(n6454), .Q(n5774), 
        .QN(n2433) );
  DFFR_X1 \REGISTERS_reg[15][1]  ( .D(n3304), .CK(CLK), .RN(n6454), .Q(n5775), 
        .QN(n2437) );
  DFFR_X1 \REGISTERS_reg[15][0]  ( .D(n3303), .CK(CLK), .RN(n6454), .Q(n5776), 
        .QN(n2441) );
  DFFR_X1 \REGISTERS_reg[18][30]  ( .D(n3301), .CK(CLK), .RN(n6460), .Q(n5453), 
        .QN(n2250) );
  DFFR_X1 \REGISTERS_reg[18][29]  ( .D(n3300), .CK(CLK), .RN(n6460), .Q(n5454), 
        .QN(n2249) );
  DFFR_X1 \REGISTERS_reg[18][28]  ( .D(n3299), .CK(CLK), .RN(n6460), .Q(n5455), 
        .QN(n2248) );
  DFFR_X1 \REGISTERS_reg[18][27]  ( .D(n3298), .CK(CLK), .RN(n6460), .Q(n5456), 
        .QN(n2247) );
  DFFR_X1 \REGISTERS_reg[18][26]  ( .D(n3297), .CK(CLK), .RN(n6460), .Q(n5457), 
        .QN(n2246) );
  DFFR_X1 \REGISTERS_reg[18][25]  ( .D(n3296), .CK(CLK), .RN(n6460), .Q(n5458), 
        .QN(n2245) );
  DFFR_X1 \REGISTERS_reg[18][24]  ( .D(n3295), .CK(CLK), .RN(n6460), .Q(n5459), 
        .QN(n2244) );
  DFFR_X1 \REGISTERS_reg[18][23]  ( .D(n3294), .CK(CLK), .RN(n6458), .Q(n5460), 
        .QN(n2243) );
  DFFR_X1 \REGISTERS_reg[18][22]  ( .D(n3293), .CK(CLK), .RN(n6458), .Q(n5461), 
        .QN(n2242) );
  DFFR_X1 \REGISTERS_reg[18][21]  ( .D(n3292), .CK(CLK), .RN(n6458), .Q(n5462), 
        .QN(n2241) );
  DFFR_X1 \REGISTERS_reg[18][20]  ( .D(n3291), .CK(CLK), .RN(n6458), .Q(n5463), 
        .QN(n2240) );
  DFFR_X1 \REGISTERS_reg[18][19]  ( .D(n3290), .CK(CLK), .RN(n6459), .Q(n5464), 
        .QN(n2239) );
  DFFR_X1 \REGISTERS_reg[18][18]  ( .D(n3289), .CK(CLK), .RN(n6459), .Q(n5465), 
        .QN(n2238) );
  DFFR_X1 \REGISTERS_reg[18][17]  ( .D(n3288), .CK(CLK), .RN(n6459), .Q(n5466), 
        .QN(n2237) );
  DFFR_X1 \REGISTERS_reg[18][16]  ( .D(n3287), .CK(CLK), .RN(n6459), .Q(n5467), 
        .QN(n2236) );
  DFFR_X1 \REGISTERS_reg[18][15]  ( .D(n3286), .CK(CLK), .RN(n6459), .Q(n5468), 
        .QN(n2235) );
  DFFR_X1 \REGISTERS_reg[18][14]  ( .D(n3285), .CK(CLK), .RN(n6459), .Q(n5469), 
        .QN(n2234) );
  DFFR_X1 \REGISTERS_reg[18][13]  ( .D(n3284), .CK(CLK), .RN(n6459), .Q(n5470), 
        .QN(n2233) );
  DFFR_X1 \REGISTERS_reg[18][12]  ( .D(n3283), .CK(CLK), .RN(n6459), .Q(n5471), 
        .QN(n2232) );
  DFFR_X1 \REGISTERS_reg[18][11]  ( .D(n3282), .CK(CLK), .RN(n6387), .Q(n5472), 
        .QN(n2231) );
  DFFR_X1 \REGISTERS_reg[18][10]  ( .D(n3281), .CK(CLK), .RN(n6387), .Q(n5473), 
        .QN(n2230) );
  DFFR_X1 \REGISTERS_reg[18][9]  ( .D(n3280), .CK(CLK), .RN(n6387), .Q(n5474), 
        .QN(n2229) );
  DFFR_X1 \REGISTERS_reg[18][8]  ( .D(n3279), .CK(CLK), .RN(n6387), .Q(n5475), 
        .QN(n2228) );
  DFFR_X1 \REGISTERS_reg[18][7]  ( .D(n3278), .CK(CLK), .RN(n6387), .Q(n5476), 
        .QN(n2227) );
  DFFR_X1 \REGISTERS_reg[18][6]  ( .D(n3277), .CK(CLK), .RN(n6387), .Q(n5477), 
        .QN(n2226) );
  DFFR_X1 \REGISTERS_reg[18][5]  ( .D(n3276), .CK(CLK), .RN(n6387), .Q(n5478), 
        .QN(n2225) );
  DFFR_X1 \REGISTERS_reg[18][4]  ( .D(n3275), .CK(CLK), .RN(n6387), .Q(n5479), 
        .QN(n2224) );
  DFFR_X1 \REGISTERS_reg[18][3]  ( .D(n3274), .CK(CLK), .RN(n6387), .Q(n5480), 
        .QN(n2223) );
  DFFR_X1 \REGISTERS_reg[18][2]  ( .D(n3273), .CK(CLK), .RN(n6387), .Q(n5481), 
        .QN(n2222) );
  DFFR_X1 \REGISTERS_reg[18][1]  ( .D(n3272), .CK(CLK), .RN(n6388), .Q(n5482), 
        .QN(n2221) );
  DFFR_X1 \REGISTERS_reg[18][0]  ( .D(n3271), .CK(CLK), .RN(n6388), .Q(n5486), 
        .QN(n2220) );
  DFFR_X1 \REGISTERS_reg[19][31]  ( .D(n3270), .CK(CLK), .RN(n6386), .Q(n5515), 
        .QN(n2219) );
  DFFR_X1 \REGISTERS_reg[19][30]  ( .D(n3269), .CK(CLK), .RN(n6386), .Q(n5516), 
        .QN(n2218) );
  DFFR_X1 \REGISTERS_reg[19][29]  ( .D(n3268), .CK(CLK), .RN(n6386), .Q(n5517), 
        .QN(n2217) );
  DFFR_X1 \REGISTERS_reg[19][28]  ( .D(n3267), .CK(CLK), .RN(n6386), .Q(n5518), 
        .QN(n2216) );
  DFFR_X1 \REGISTERS_reg[19][27]  ( .D(n3266), .CK(CLK), .RN(n6386), .Q(n5519), 
        .QN(n2215) );
  DFFR_X1 \REGISTERS_reg[19][26]  ( .D(n3265), .CK(CLK), .RN(n6386), .Q(n5520), 
        .QN(n2214) );
  DFFR_X1 \REGISTERS_reg[19][25]  ( .D(n3264), .CK(CLK), .RN(n6386), .Q(n5521), 
        .QN(n2213) );
  DFFR_X1 \REGISTERS_reg[19][24]  ( .D(n3263), .CK(CLK), .RN(n6386), .Q(n5522), 
        .QN(n2212) );
  DFFR_X1 \REGISTERS_reg[19][23]  ( .D(n3262), .CK(CLK), .RN(n6386), .Q(n5523), 
        .QN(n2211) );
  DFFR_X1 \REGISTERS_reg[19][22]  ( .D(n3261), .CK(CLK), .RN(n6386), .Q(n5524), 
        .QN(n2210) );
  DFFR_X1 \REGISTERS_reg[19][21]  ( .D(n3260), .CK(CLK), .RN(n6387), .Q(n5525), 
        .QN(n2209) );
  DFFR_X1 \REGISTERS_reg[19][20]  ( .D(n3259), .CK(CLK), .RN(n6387), .Q(n5526), 
        .QN(n2208) );
  DFFR_X1 \REGISTERS_reg[19][19]  ( .D(n3258), .CK(CLK), .RN(n6385), .Q(n5527), 
        .QN(n2207) );
  DFFR_X1 \REGISTERS_reg[19][18]  ( .D(n3257), .CK(CLK), .RN(n6385), .Q(n5528), 
        .QN(n2206) );
  DFFR_X1 \REGISTERS_reg[19][17]  ( .D(n3256), .CK(CLK), .RN(n6385), .Q(n5529), 
        .QN(n2205) );
  DFFR_X1 \REGISTERS_reg[19][16]  ( .D(n3255), .CK(CLK), .RN(n6385), .Q(n5530), 
        .QN(n2204) );
  DFFR_X1 \REGISTERS_reg[19][15]  ( .D(n3254), .CK(CLK), .RN(n6385), .Q(n5531), 
        .QN(n2203) );
  DFFR_X1 \REGISTERS_reg[19][14]  ( .D(n3253), .CK(CLK), .RN(n6385), .Q(n5532), 
        .QN(n2202) );
  DFFR_X1 \REGISTERS_reg[19][13]  ( .D(n3252), .CK(CLK), .RN(n6385), .Q(n5533), 
        .QN(n2201) );
  DFFR_X1 \REGISTERS_reg[19][12]  ( .D(n3251), .CK(CLK), .RN(n6385), .Q(n5534), 
        .QN(n2200) );
  DFFR_X1 \REGISTERS_reg[19][11]  ( .D(n3250), .CK(CLK), .RN(n6385), .Q(n5535), 
        .QN(n2199) );
  DFFR_X1 \REGISTERS_reg[19][10]  ( .D(n3249), .CK(CLK), .RN(n6385), .Q(n5536), 
        .QN(n2198) );
  DFFR_X1 \REGISTERS_reg[19][9]  ( .D(n3248), .CK(CLK), .RN(n6386), .Q(n5537), 
        .QN(n2197) );
  DFFR_X1 \REGISTERS_reg[19][8]  ( .D(n3247), .CK(CLK), .RN(n6386), .Q(n5538), 
        .QN(n2196) );
  DFFR_X1 \REGISTERS_reg[19][7]  ( .D(n3246), .CK(CLK), .RN(n6385), .Q(n5539), 
        .QN(n2195) );
  DFFR_X1 \REGISTERS_reg[19][6]  ( .D(n3245), .CK(CLK), .RN(n6384), .Q(n5540), 
        .QN(n2194) );
  DFFR_X1 \REGISTERS_reg[19][5]  ( .D(n3244), .CK(CLK), .RN(n6384), .Q(n5541), 
        .QN(n2193) );
  DFFR_X1 \REGISTERS_reg[19][4]  ( .D(n3243), .CK(CLK), .RN(n6384), .Q(n5542), 
        .QN(n2192) );
  DFFR_X1 \REGISTERS_reg[19][3]  ( .D(n3242), .CK(CLK), .RN(n6384), .Q(n5543), 
        .QN(n2191) );
  DFFR_X1 \REGISTERS_reg[19][2]  ( .D(n3241), .CK(CLK), .RN(n6384), .Q(n5544), 
        .QN(n2190) );
  DFFR_X1 \REGISTERS_reg[19][1]  ( .D(n3240), .CK(CLK), .RN(n6384), .Q(n5545), 
        .QN(n2189) );
  DFFR_X1 \REGISTERS_reg[19][0]  ( .D(n3239), .CK(CLK), .RN(n6385), .Q(n5680), 
        .QN(n2188) );
  DFFR_X1 \REGISTERS_reg[25][31]  ( .D(n3142), .CK(CLK), .RN(n6394), .Q(n5137), 
        .QN(n2187) );
  DFFR_X1 \REGISTERS_reg[25][30]  ( .D(n3141), .CK(CLK), .RN(n6394), .Q(n5138), 
        .QN(n2186) );
  DFFR_X1 \REGISTERS_reg[25][29]  ( .D(n3140), .CK(CLK), .RN(n6394), .Q(n5139), 
        .QN(n2185) );
  DFFR_X1 \REGISTERS_reg[25][28]  ( .D(n3139), .CK(CLK), .RN(n6394), .Q(n5140), 
        .QN(n2184) );
  DFFR_X1 \REGISTERS_reg[25][27]  ( .D(n3138), .CK(CLK), .RN(n6394), .Q(n5141), 
        .QN(n2183) );
  DFFR_X1 \REGISTERS_reg[25][26]  ( .D(n3137), .CK(CLK), .RN(n6394), .Q(n5142), 
        .QN(n2182) );
  DFFR_X1 \REGISTERS_reg[25][25]  ( .D(n3136), .CK(CLK), .RN(n6394), .Q(n5143), 
        .QN(n2181) );
  DFFR_X1 \REGISTERS_reg[25][24]  ( .D(n3135), .CK(CLK), .RN(n6394), .Q(n5144), 
        .QN(n2180) );
  DFFR_X1 \REGISTERS_reg[25][23]  ( .D(n3134), .CK(CLK), .RN(n6394), .Q(n5145), 
        .QN(n2179) );
  DFFR_X1 \REGISTERS_reg[25][22]  ( .D(n3133), .CK(CLK), .RN(n6394), .Q(n5146), 
        .QN(n2178) );
  DFFR_X1 \REGISTERS_reg[25][21]  ( .D(n3132), .CK(CLK), .RN(n6395), .Q(n5147), 
        .QN(n2177) );
  DFFR_X1 \REGISTERS_reg[25][20]  ( .D(n3131), .CK(CLK), .RN(n6395), .Q(n5148), 
        .QN(n2176) );
  DFFR_X1 \REGISTERS_reg[25][19]  ( .D(n3130), .CK(CLK), .RN(n6405), .Q(n5149), 
        .QN(n2175) );
  DFFR_X1 \REGISTERS_reg[25][18]  ( .D(n3129), .CK(CLK), .RN(n6405), .Q(n5150), 
        .QN(n2174) );
  DFFR_X1 \REGISTERS_reg[25][17]  ( .D(n3128), .CK(CLK), .RN(n6405), .Q(n5151), 
        .QN(n2173) );
  DFFR_X1 \REGISTERS_reg[25][16]  ( .D(n3127), .CK(CLK), .RN(n6405), .Q(n5152), 
        .QN(n2172) );
  DFFR_X1 \REGISTERS_reg[25][15]  ( .D(n3126), .CK(CLK), .RN(n6405), .Q(n5153), 
        .QN(n2171) );
  DFFR_X1 \REGISTERS_reg[25][14]  ( .D(n3125), .CK(CLK), .RN(n6405), .Q(n5154), 
        .QN(n2170) );
  DFFR_X1 \REGISTERS_reg[25][13]  ( .D(n3124), .CK(CLK), .RN(n6405), .Q(n5155), 
        .QN(n2169) );
  DFFR_X1 \REGISTERS_reg[25][12]  ( .D(n3123), .CK(CLK), .RN(n6405), .Q(n5156), 
        .QN(n2168) );
  DFFR_X1 \REGISTERS_reg[25][11]  ( .D(n3122), .CK(CLK), .RN(n6405), .Q(n5157), 
        .QN(n2167) );
  DFFR_X1 \REGISTERS_reg[25][10]  ( .D(n3121), .CK(CLK), .RN(n6405), .Q(n5158), 
        .QN(n2166) );
  DFFR_X1 \REGISTERS_reg[25][9]  ( .D(n3120), .CK(CLK), .RN(n6405), .Q(n5159), 
        .QN(n2165) );
  DFFR_X1 \REGISTERS_reg[25][8]  ( .D(n3119), .CK(CLK), .RN(n6405), .Q(n5160), 
        .QN(n2164) );
  DFFR_X1 \REGISTERS_reg[25][7]  ( .D(n3118), .CK(CLK), .RN(n6404), .Q(n5161), 
        .QN(n2163) );
  DFFR_X1 \REGISTERS_reg[25][6]  ( .D(n3117), .CK(CLK), .RN(n6404), .Q(n5162), 
        .QN(n2162) );
  DFFR_X1 \REGISTERS_reg[25][5]  ( .D(n3116), .CK(CLK), .RN(n6404), .Q(n5163), 
        .QN(n2161) );
  DFFR_X1 \REGISTERS_reg[25][4]  ( .D(n3115), .CK(CLK), .RN(n6404), .Q(n5164), 
        .QN(n2160) );
  DFFR_X1 \REGISTERS_reg[25][3]  ( .D(n3114), .CK(CLK), .RN(n6404), .Q(n5165), 
        .QN(n2159) );
  DFFR_X1 \REGISTERS_reg[25][2]  ( .D(n3113), .CK(CLK), .RN(n6404), .Q(n5166), 
        .QN(n2158) );
  DFFR_X1 \REGISTERS_reg[25][1]  ( .D(n3112), .CK(CLK), .RN(n6404), .Q(n5167), 
        .QN(n2157) );
  DFFR_X1 \REGISTERS_reg[25][0]  ( .D(n3111), .CK(CLK), .RN(n6404), .Q(n5171), 
        .QN(n2156) );
  DFFR_X1 \REGISTERS_reg[29][31]  ( .D(n3078), .CK(CLK), .RN(n6408), .Q(n5234), 
        .QN(n2059) );
  DFFR_X1 \REGISTERS_reg[29][30]  ( .D(n3077), .CK(CLK), .RN(n6408), .Q(n5268), 
        .QN(n2058) );
  DFFR_X1 \REGISTERS_reg[29][29]  ( .D(n3076), .CK(CLK), .RN(n6408), .Q(n5269), 
        .QN(n2057) );
  DFFR_X1 \REGISTERS_reg[29][28]  ( .D(n3075), .CK(CLK), .RN(n6408), .Q(n5270), 
        .QN(n2056) );
  DFFR_X1 \REGISTERS_reg[29][27]  ( .D(n3074), .CK(CLK), .RN(n6407), .Q(n5271), 
        .QN(n2055) );
  DFFR_X1 \REGISTERS_reg[29][26]  ( .D(n3073), .CK(CLK), .RN(n6407), .Q(n5272), 
        .QN(n2054) );
  DFFR_X1 \REGISTERS_reg[29][25]  ( .D(n3072), .CK(CLK), .RN(n6407), .Q(n5273), 
        .QN(n2053) );
  DFFR_X1 \REGISTERS_reg[29][24]  ( .D(n3071), .CK(CLK), .RN(n6407), .Q(n5274), 
        .QN(n2052) );
  DFFR_X1 \REGISTERS_reg[29][23]  ( .D(n3070), .CK(CLK), .RN(n6407), .Q(n5275), 
        .QN(n2051) );
  DFFR_X1 \REGISTERS_reg[29][22]  ( .D(n3069), .CK(CLK), .RN(n6407), .Q(n5276), 
        .QN(n2050) );
  DFFR_X1 \REGISTERS_reg[29][21]  ( .D(n3068), .CK(CLK), .RN(n6407), .Q(n5277), 
        .QN(n2049) );
  DFFR_X1 \REGISTERS_reg[29][20]  ( .D(n3067), .CK(CLK), .RN(n6407), .Q(n5278), 
        .QN(n2048) );
  DFFR_X1 \REGISTERS_reg[29][19]  ( .D(n3066), .CK(CLK), .RN(n6407), .Q(n5279), 
        .QN(n2047) );
  DFFR_X1 \REGISTERS_reg[29][18]  ( .D(n3065), .CK(CLK), .RN(n6407), .Q(n5280), 
        .QN(n2046) );
  DFFR_X1 \REGISTERS_reg[29][17]  ( .D(n3064), .CK(CLK), .RN(n6407), .Q(n5281), 
        .QN(n2045) );
  DFFR_X1 \REGISTERS_reg[29][16]  ( .D(n3063), .CK(CLK), .RN(n6407), .Q(n5282), 
        .QN(n2044) );
  DFFR_X1 \REGISTERS_reg[29][15]  ( .D(n3062), .CK(CLK), .RN(n6406), .Q(n5283), 
        .QN(n2043) );
  DFFR_X1 \REGISTERS_reg[29][14]  ( .D(n3061), .CK(CLK), .RN(n6406), .Q(n5284), 
        .QN(n2042) );
  DFFR_X1 \REGISTERS_reg[29][13]  ( .D(n3060), .CK(CLK), .RN(n6406), .Q(n5285), 
        .QN(n2041) );
  DFFR_X1 \REGISTERS_reg[29][12]  ( .D(n3059), .CK(CLK), .RN(n6406), .Q(n5286), 
        .QN(n2040) );
  DFFR_X1 \REGISTERS_reg[29][11]  ( .D(n3058), .CK(CLK), .RN(n6406), .Q(n5287), 
        .QN(n2039) );
  DFFR_X1 \REGISTERS_reg[29][10]  ( .D(n3057), .CK(CLK), .RN(n6406), .Q(n5288), 
        .QN(n2038) );
  DFFR_X1 \REGISTERS_reg[29][9]  ( .D(n3056), .CK(CLK), .RN(n6406), .Q(n5289), 
        .QN(n2037) );
  DFFR_X1 \REGISTERS_reg[29][8]  ( .D(n3055), .CK(CLK), .RN(n6406), .Q(n5290), 
        .QN(n2036) );
  DFFR_X1 \REGISTERS_reg[29][7]  ( .D(n3054), .CK(CLK), .RN(n6406), .Q(n5291), 
        .QN(n2035) );
  DFFR_X1 \REGISTERS_reg[29][6]  ( .D(n3053), .CK(CLK), .RN(n6406), .Q(n5292), 
        .QN(n2034) );
  DFFR_X1 \REGISTERS_reg[29][5]  ( .D(n3052), .CK(CLK), .RN(n6406), .Q(n5293), 
        .QN(n2033) );
  DFFR_X1 \REGISTERS_reg[29][4]  ( .D(n3051), .CK(CLK), .RN(n6406), .Q(n5294), 
        .QN(n2032) );
  DFFR_X1 \REGISTERS_reg[29][3]  ( .D(n3050), .CK(CLK), .RN(n6416), .Q(n5295), 
        .QN(n2031) );
  DFFR_X1 \REGISTERS_reg[29][2]  ( .D(n3049), .CK(CLK), .RN(n6416), .Q(n5296), 
        .QN(n2030) );
  DFFR_X1 \REGISTERS_reg[29][1]  ( .D(n3048), .CK(CLK), .RN(n6416), .Q(n5297), 
        .QN(n2029) );
  DFFR_X1 \REGISTERS_reg[29][0]  ( .D(n3047), .CK(CLK), .RN(n6416), .Q(n5235), 
        .QN(n2028) );
  DFF_X1 \OUT2_reg[31]  ( .D(n3015), .CK(CLK), .Q(OUT2[31]), .QN(n7551) );
  DFF_X1 \OUT2_reg[30]  ( .D(n3016), .CK(CLK), .Q(OUT2[30]), .QN(n2655) );
  DFF_X1 \OUT2_reg[29]  ( .D(n3017), .CK(CLK), .Q(OUT2[29]), .QN(n2656) );
  DFF_X1 \OUT2_reg[28]  ( .D(n3018), .CK(CLK), .Q(OUT2[28]), .QN(n2657) );
  DFF_X1 \OUT2_reg[27]  ( .D(n3019), .CK(CLK), .Q(OUT2[27]), .QN(n2658) );
  DFF_X1 \OUT2_reg[26]  ( .D(n3020), .CK(CLK), .Q(OUT2[26]), .QN(n2659) );
  DFF_X1 \OUT2_reg[25]  ( .D(n3021), .CK(CLK), .Q(OUT2[25]), .QN(n2660) );
  DFF_X1 \OUT2_reg[24]  ( .D(n3022), .CK(CLK), .Q(OUT2[24]), .QN(n2661) );
  DFF_X1 \OUT2_reg[23]  ( .D(n3023), .CK(CLK), .Q(OUT2[23]), .QN(n2662) );
  DFF_X1 \OUT2_reg[22]  ( .D(n3024), .CK(CLK), .Q(OUT2[22]), .QN(n2663) );
  DFF_X1 \OUT2_reg[21]  ( .D(n3025), .CK(CLK), .Q(OUT2[21]), .QN(n2664) );
  DFF_X1 \OUT2_reg[20]  ( .D(n3026), .CK(CLK), .Q(OUT2[20]), .QN(n2665) );
  DFF_X1 \OUT2_reg[19]  ( .D(n3027), .CK(CLK), .Q(OUT2[19]), .QN(n2666) );
  DFF_X1 \OUT2_reg[18]  ( .D(n3028), .CK(CLK), .Q(OUT2[18]), .QN(n2667) );
  DFF_X1 \OUT2_reg[17]  ( .D(n3029), .CK(CLK), .Q(OUT2[17]), .QN(n2668) );
  DFF_X1 \OUT2_reg[16]  ( .D(n3030), .CK(CLK), .Q(OUT2[16]), .QN(n2669) );
  DFF_X1 \OUT2_reg[15]  ( .D(n3031), .CK(CLK), .Q(OUT2[15]), .QN(n2670) );
  DFF_X1 \OUT2_reg[14]  ( .D(n3032), .CK(CLK), .Q(OUT2[14]), .QN(n2671) );
  DFF_X1 \OUT2_reg[13]  ( .D(n3033), .CK(CLK), .Q(OUT2[13]), .QN(n2672) );
  DFF_X1 \OUT2_reg[12]  ( .D(n3034), .CK(CLK), .Q(OUT2[12]), .QN(n2673) );
  DFF_X1 \OUT2_reg[11]  ( .D(n3035), .CK(CLK), .Q(OUT2[11]), .QN(n2674) );
  DFF_X1 \OUT2_reg[10]  ( .D(n3036), .CK(CLK), .Q(OUT2[10]), .QN(n2675) );
  DFF_X1 \OUT2_reg[9]  ( .D(n3037), .CK(CLK), .Q(OUT2[9]), .QN(n2676) );
  DFF_X1 \OUT2_reg[8]  ( .D(n3038), .CK(CLK), .Q(OUT2[8]), .QN(n2677) );
  DFF_X1 \OUT2_reg[7]  ( .D(n3039), .CK(CLK), .Q(OUT2[7]), .QN(n2678) );
  DFF_X1 \OUT2_reg[6]  ( .D(n3040), .CK(CLK), .Q(OUT2[6]), .QN(n2679) );
  DFF_X1 \OUT2_reg[5]  ( .D(n3041), .CK(CLK), .Q(OUT2[5]), .QN(n2680) );
  DFF_X1 \OUT2_reg[4]  ( .D(n3042), .CK(CLK), .Q(OUT2[4]), .QN(n2681) );
  DFF_X1 \OUT2_reg[3]  ( .D(n3043), .CK(CLK), .Q(OUT2[3]), .QN(n2682) );
  DFF_X1 \OUT2_reg[2]  ( .D(n3044), .CK(CLK), .Q(OUT2[2]), .QN(n2683) );
  DFF_X1 \OUT2_reg[1]  ( .D(n3045), .CK(CLK), .Q(OUT2[1]), .QN(n2684) );
  DFF_X1 \OUT2_reg[0]  ( .D(n3046), .CK(CLK), .Q(OUT2[0]), .QN(n2685) );
  DFF_X1 \OUT1_reg[31]  ( .D(n3014), .CK(CLK), .Q(OUT1[31]), .QN(n2653) );
  DFF_X1 \OUT1_reg[30]  ( .D(n3013), .CK(CLK), .Q(OUT1[30]), .QN(n2652) );
  DFF_X1 \OUT1_reg[29]  ( .D(n3012), .CK(CLK), .Q(OUT1[29]), .QN(n2651) );
  DFF_X1 \OUT1_reg[28]  ( .D(n3011), .CK(CLK), .Q(OUT1[28]), .QN(n2650) );
  DFF_X1 \OUT1_reg[27]  ( .D(n3010), .CK(CLK), .Q(OUT1[27]), .QN(n2649) );
  DFF_X1 \OUT1_reg[26]  ( .D(n3009), .CK(CLK), .Q(OUT1[26]), .QN(n2648) );
  DFF_X1 \OUT1_reg[25]  ( .D(n3008), .CK(CLK), .Q(OUT1[25]), .QN(n2647) );
  DFF_X1 \OUT1_reg[24]  ( .D(n3007), .CK(CLK), .Q(OUT1[24]), .QN(n2646) );
  DFF_X1 \OUT1_reg[23]  ( .D(n3006), .CK(CLK), .Q(OUT1[23]), .QN(n2645) );
  DFF_X1 \OUT1_reg[22]  ( .D(n3005), .CK(CLK), .Q(OUT1[22]), .QN(n2644) );
  DFF_X1 \OUT1_reg[21]  ( .D(n3004), .CK(CLK), .Q(OUT1[21]), .QN(n2643) );
  DFF_X1 \OUT1_reg[20]  ( .D(n3003), .CK(CLK), .Q(OUT1[20]), .QN(n2642) );
  DFF_X1 \OUT1_reg[19]  ( .D(n3002), .CK(CLK), .Q(OUT1[19]), .QN(n2641) );
  DFF_X1 \OUT1_reg[18]  ( .D(n3001), .CK(CLK), .Q(OUT1[18]), .QN(n2640) );
  DFF_X1 \OUT1_reg[17]  ( .D(n3000), .CK(CLK), .Q(OUT1[17]), .QN(n2639) );
  DFF_X1 \OUT1_reg[16]  ( .D(n2999), .CK(CLK), .Q(OUT1[16]), .QN(n2638) );
  DFF_X1 \OUT1_reg[15]  ( .D(n2998), .CK(CLK), .Q(OUT1[15]), .QN(n2637) );
  DFF_X1 \OUT1_reg[14]  ( .D(n2997), .CK(CLK), .Q(OUT1[14]), .QN(n2636) );
  DFF_X1 \OUT1_reg[13]  ( .D(n2996), .CK(CLK), .Q(OUT1[13]), .QN(n2635) );
  DFF_X1 \OUT1_reg[12]  ( .D(n2995), .CK(CLK), .Q(OUT1[12]), .QN(n2634) );
  DFF_X1 \OUT1_reg[11]  ( .D(n2994), .CK(CLK), .Q(OUT1[11]), .QN(n2633) );
  DFF_X1 \OUT1_reg[10]  ( .D(n2993), .CK(CLK), .Q(OUT1[10]), .QN(n2632) );
  DFF_X1 \OUT1_reg[9]  ( .D(n2992), .CK(CLK), .Q(OUT1[9]), .QN(n2631) );
  DFF_X1 \OUT1_reg[8]  ( .D(n2991), .CK(CLK), .Q(OUT1[8]), .QN(n2630) );
  DFF_X1 \OUT1_reg[7]  ( .D(n2990), .CK(CLK), .Q(OUT1[7]), .QN(n2629) );
  DFF_X1 \OUT1_reg[6]  ( .D(n2989), .CK(CLK), .Q(OUT1[6]), .QN(n2628) );
  DFF_X1 \OUT1_reg[5]  ( .D(n2988), .CK(CLK), .Q(OUT1[5]), .QN(n2627) );
  DFF_X1 \OUT1_reg[4]  ( .D(n2987), .CK(CLK), .Q(OUT1[4]), .QN(n2626) );
  DFF_X1 \OUT1_reg[3]  ( .D(n2986), .CK(CLK), .Q(OUT1[3]), .QN(n2625) );
  DFF_X1 \OUT1_reg[2]  ( .D(n2985), .CK(CLK), .Q(OUT1[2]), .QN(n2624) );
  DFF_X1 \OUT1_reg[1]  ( .D(n2984), .CK(CLK), .Q(OUT1[1]), .QN(n2623) );
  DFF_X1 \OUT1_reg[0]  ( .D(n2983), .CK(CLK), .Q(OUT1[0]), .QN(n6512) );
  DFFR_X1 \REGISTERS_reg[24][31]  ( .D(n3174), .CK(CLK), .RN(n6382), .Q(n2877), 
        .QN(n5880) );
  DFFR_X1 \REGISTERS_reg[24][30]  ( .D(n7656), .CK(CLK), .RN(n6398), .Q(n2876), 
        .QN(n5881) );
  DFFR_X1 \REGISTERS_reg[24][29]  ( .D(n7657), .CK(CLK), .RN(n6397), .Q(n2875), 
        .QN(n5882) );
  DFFR_X1 \REGISTERS_reg[24][28]  ( .D(n7658), .CK(CLK), .RN(n6397), .Q(n2874), 
        .QN(n5883) );
  DFFR_X1 \REGISTERS_reg[24][27]  ( .D(n7659), .CK(CLK), .RN(n6397), .Q(n2873), 
        .QN(n5884) );
  DFFR_X1 \REGISTERS_reg[24][26]  ( .D(n7660), .CK(CLK), .RN(n6397), .Q(n2872), 
        .QN(n5885) );
  DFFR_X1 \REGISTERS_reg[24][25]  ( .D(n7661), .CK(CLK), .RN(n6397), .Q(n2871), 
        .QN(n5886) );
  DFFR_X1 \REGISTERS_reg[24][24]  ( .D(n7662), .CK(CLK), .RN(n6397), .Q(n2870), 
        .QN(n5887) );
  DFFR_X1 \REGISTERS_reg[24][23]  ( .D(n7663), .CK(CLK), .RN(n6397), .Q(n2869), 
        .QN(n5888) );
  DFFR_X1 \REGISTERS_reg[24][22]  ( .D(n7664), .CK(CLK), .RN(n6397), .Q(n2868), 
        .QN(n5889) );
  DFFR_X1 \REGISTERS_reg[24][21]  ( .D(n7665), .CK(CLK), .RN(n6396), .Q(n2867), 
        .QN(n5890) );
  DFFR_X1 \REGISTERS_reg[24][20]  ( .D(n7666), .CK(CLK), .RN(n6396), .Q(n2866), 
        .QN(n5891) );
  DFFR_X1 \REGISTERS_reg[24][19]  ( .D(n7667), .CK(CLK), .RN(n6396), .Q(n2865), 
        .QN(n5892) );
  DFFR_X1 \REGISTERS_reg[24][18]  ( .D(n7668), .CK(CLK), .RN(n6396), .Q(n2864), 
        .QN(n5893) );
  DFFR_X1 \REGISTERS_reg[24][17]  ( .D(n7669), .CK(CLK), .RN(n6396), .Q(n2863), 
        .QN(n5894) );
  DFFR_X1 \REGISTERS_reg[24][16]  ( .D(n7670), .CK(CLK), .RN(n6396), .Q(n2862), 
        .QN(n5895) );
  DFFR_X1 \REGISTERS_reg[24][15]  ( .D(n7671), .CK(CLK), .RN(n6396), .Q(n2861), 
        .QN(n5896) );
  DFFR_X1 \REGISTERS_reg[24][14]  ( .D(n7672), .CK(CLK), .RN(n6396), .Q(n2860), 
        .QN(n5897) );
  DFFR_X1 \REGISTERS_reg[24][13]  ( .D(n7673), .CK(CLK), .RN(n6396), .Q(n2859), 
        .QN(n5898) );
  DFFR_X1 \REGISTERS_reg[24][12]  ( .D(n7674), .CK(CLK), .RN(n6396), .Q(n2858), 
        .QN(n5899) );
  DFFR_X1 \REGISTERS_reg[24][11]  ( .D(n7675), .CK(CLK), .RN(n6396), .Q(n2857), 
        .QN(n5900) );
  DFFR_X1 \REGISTERS_reg[24][10]  ( .D(n7676), .CK(CLK), .RN(n6396), .Q(n2856), 
        .QN(n5901) );
  DFFR_X1 \REGISTERS_reg[24][9]  ( .D(n7677), .CK(CLK), .RN(n6395), .Q(n2855), 
        .QN(n5902) );
  DFFR_X1 \REGISTERS_reg[24][8]  ( .D(n7678), .CK(CLK), .RN(n6395), .Q(n2854), 
        .QN(n5903) );
  DFFR_X1 \REGISTERS_reg[24][7]  ( .D(n7679), .CK(CLK), .RN(n6395), .Q(n2853), 
        .QN(n5904) );
  DFFR_X1 \REGISTERS_reg[24][6]  ( .D(n7680), .CK(CLK), .RN(n6395), .Q(n2852), 
        .QN(n5905) );
  DFFR_X1 \REGISTERS_reg[24][5]  ( .D(n7681), .CK(CLK), .RN(n6395), .Q(n2851), 
        .QN(n5906) );
  DFFR_X1 \REGISTERS_reg[24][4]  ( .D(n7682), .CK(CLK), .RN(n6395), .Q(n2850), 
        .QN(n5907) );
  DFFR_X1 \REGISTERS_reg[24][3]  ( .D(n3146), .CK(CLK), .RN(n6395), .Q(n5483), 
        .QN(n987) );
  DFFR_X1 \REGISTERS_reg[24][2]  ( .D(n3145), .CK(CLK), .RN(n6395), .Q(n5484), 
        .QN(n971) );
  DFFR_X1 \REGISTERS_reg[24][1]  ( .D(n3144), .CK(CLK), .RN(n6395), .Q(n5485), 
        .QN(n955) );
  DFFR_X1 \REGISTERS_reg[24][0]  ( .D(n3143), .CK(CLK), .RN(n6395), .Q(n5583), 
        .QN(n938) );
  DFFR_X1 \REGISTERS_reg[23][3]  ( .D(n3178), .CK(CLK), .RN(n6397), .Q(n5580), 
        .QN(n988) );
  DFFR_X1 \REGISTERS_reg[23][2]  ( .D(n3177), .CK(CLK), .RN(n6397), .Q(n5581), 
        .QN(n972) );
  DFFR_X1 \REGISTERS_reg[23][1]  ( .D(n3176), .CK(CLK), .RN(n6397), .Q(n5582), 
        .QN(n956) );
  DFFR_X1 \REGISTERS_reg[23][0]  ( .D(n3175), .CK(CLK), .RN(n6397), .Q(n5647), 
        .QN(n939) );
  DFFR_X1 \REGISTERS_reg[3][26]  ( .D(n7779), .CK(CLK), .RN(n6428), .Q(n4056), 
        .QN(n5915) );
  DFFR_X1 \REGISTERS_reg[3][25]  ( .D(n7780), .CK(CLK), .RN(n6428), .Q(n4055), 
        .QN(n5916) );
  DFFR_X1 \REGISTERS_reg[3][24]  ( .D(n7781), .CK(CLK), .RN(n6428), .Q(n4054), 
        .QN(n5917) );
  DFFR_X1 \REGISTERS_reg[3][23]  ( .D(n7782), .CK(CLK), .RN(n6427), .Q(n4053), 
        .QN(n5918) );
  DFFR_X1 \REGISTERS_reg[3][22]  ( .D(n7783), .CK(CLK), .RN(n6427), .Q(n4052), 
        .QN(n5919) );
  DFFR_X1 \REGISTERS_reg[3][21]  ( .D(n7784), .CK(CLK), .RN(n6427), .Q(n4051), 
        .QN(n5920) );
  DFFR_X1 \REGISTERS_reg[3][20]  ( .D(n7785), .CK(CLK), .RN(n6427), .Q(n4050), 
        .QN(n5921) );
  DFFR_X1 \REGISTERS_reg[3][19]  ( .D(n7786), .CK(CLK), .RN(n6427), .Q(n4049), 
        .QN(n5922) );
  DFFR_X1 \REGISTERS_reg[3][18]  ( .D(n7787), .CK(CLK), .RN(n6427), .Q(n4048), 
        .QN(n5923) );
  DFFR_X1 \REGISTERS_reg[3][17]  ( .D(n7788), .CK(CLK), .RN(n6427), .Q(n4047), 
        .QN(n5924) );
  DFFR_X1 \REGISTERS_reg[3][16]  ( .D(n7789), .CK(CLK), .RN(n6427), .Q(n4046), 
        .QN(n5925) );
  DFFR_X1 \REGISTERS_reg[3][15]  ( .D(n7790), .CK(CLK), .RN(n6426), .Q(n4045), 
        .QN(n5926) );
  DFFR_X1 \REGISTERS_reg[3][14]  ( .D(n7791), .CK(CLK), .RN(n6426), .Q(n4044), 
        .QN(n5927) );
  DFFR_X1 \REGISTERS_reg[3][13]  ( .D(n7792), .CK(CLK), .RN(n6426), .Q(n4043), 
        .QN(n5928) );
  DFFR_X1 \REGISTERS_reg[3][12]  ( .D(n7793), .CK(CLK), .RN(n6426), .Q(n4042), 
        .QN(n5929) );
  DFFR_X1 \REGISTERS_reg[3][11]  ( .D(n7794), .CK(CLK), .RN(n6426), .Q(n4041), 
        .QN(n5930) );
  DFFR_X1 \REGISTERS_reg[3][10]  ( .D(n7795), .CK(CLK), .RN(n6426), .Q(n4040), 
        .QN(n5931) );
  DFFR_X1 \REGISTERS_reg[3][9]  ( .D(n7796), .CK(CLK), .RN(n6426), .Q(n4039), 
        .QN(n5932) );
  DFFR_X1 \REGISTERS_reg[3][8]  ( .D(n7797), .CK(CLK), .RN(n6426), .Q(n4038), 
        .QN(n5933) );
  DFFR_X1 \REGISTERS_reg[3][7]  ( .D(n7798), .CK(CLK), .RN(n6426), .Q(n4037), 
        .QN(n5934) );
  DFFR_X1 \REGISTERS_reg[3][6]  ( .D(n7799), .CK(CLK), .RN(n6426), .Q(n4036), 
        .QN(n5935) );
  DFFR_X1 \REGISTERS_reg[3][5]  ( .D(n7800), .CK(CLK), .RN(n6426), .Q(n4035), 
        .QN(n5936) );
  DFFR_X1 \REGISTERS_reg[3][4]  ( .D(n7801), .CK(CLK), .RN(n6426), .Q(n4034), 
        .QN(n5937) );
  DFFR_X1 \REGISTERS_reg[3][3]  ( .D(n7802), .CK(CLK), .RN(n6425), .Q(n4033), 
        .QN(n5938) );
  DFFR_X1 \REGISTERS_reg[3][2]  ( .D(n7803), .CK(CLK), .RN(n6425), .Q(n4032), 
        .QN(n5939) );
  DFFR_X1 \REGISTERS_reg[3][1]  ( .D(n7804), .CK(CLK), .RN(n6425), .Q(n4031), 
        .QN(n5940) );
  DFFR_X1 \REGISTERS_reg[3][0]  ( .D(n7805), .CK(CLK), .RN(n6425), .Q(n4030), 
        .QN(n5910) );
  DFFR_X1 \REGISTERS_reg[2][31]  ( .D(n7806), .CK(CLK), .RN(n6420), .Q(n4093), 
        .QN(n5973) );
  DFFR_X1 \REGISTERS_reg[2][30]  ( .D(n7807), .CK(CLK), .RN(n6420), .Q(n4092), 
        .QN(n5975) );
  DFFR_X1 \REGISTERS_reg[2][29]  ( .D(n7808), .CK(CLK), .RN(n6420), .Q(n4091), 
        .QN(n5976) );
  DFFR_X1 \REGISTERS_reg[2][28]  ( .D(n7809), .CK(CLK), .RN(n6420), .Q(n4090), 
        .QN(n5977) );
  DFFR_X1 \REGISTERS_reg[2][27]  ( .D(n7810), .CK(CLK), .RN(n6419), .Q(n4089), 
        .QN(n5978) );
  DFFR_X1 \REGISTERS_reg[2][26]  ( .D(n7811), .CK(CLK), .RN(n6419), .Q(n4088), 
        .QN(n5979) );
  DFFR_X1 \REGISTERS_reg[2][25]  ( .D(n7812), .CK(CLK), .RN(n6419), .Q(n4087), 
        .QN(n5980) );
  DFFR_X1 \REGISTERS_reg[2][24]  ( .D(n7813), .CK(CLK), .RN(n6419), .Q(n4086), 
        .QN(n5981) );
  DFFR_X1 \REGISTERS_reg[2][23]  ( .D(n7814), .CK(CLK), .RN(n6419), .Q(n4085), 
        .QN(n5982) );
  DFFR_X1 \REGISTERS_reg[2][22]  ( .D(n7815), .CK(CLK), .RN(n6419), .Q(n4084), 
        .QN(n5983) );
  DFFR_X1 \REGISTERS_reg[2][21]  ( .D(n7816), .CK(CLK), .RN(n6419), .Q(n4083), 
        .QN(n5984) );
  DFFR_X1 \REGISTERS_reg[2][20]  ( .D(n7817), .CK(CLK), .RN(n6419), .Q(n4082), 
        .QN(n5985) );
  DFFR_X1 \REGISTERS_reg[2][19]  ( .D(n7818), .CK(CLK), .RN(n6418), .Q(n4081), 
        .QN(n5986) );
  DFFR_X1 \REGISTERS_reg[2][18]  ( .D(n7819), .CK(CLK), .RN(n6418), .Q(n4080), 
        .QN(n5987) );
  DFFR_X1 \REGISTERS_reg[2][17]  ( .D(n7820), .CK(CLK), .RN(n6418), .Q(n4079), 
        .QN(n5988) );
  DFFR_X1 \REGISTERS_reg[2][16]  ( .D(n7821), .CK(CLK), .RN(n6418), .Q(n4078), 
        .QN(n5989) );
  DFFR_X1 \REGISTERS_reg[2][15]  ( .D(n7822), .CK(CLK), .RN(n6418), .Q(n4077), 
        .QN(n5990) );
  DFFR_X1 \REGISTERS_reg[2][14]  ( .D(n7823), .CK(CLK), .RN(n6418), .Q(n4076), 
        .QN(n5991) );
  DFFR_X1 \REGISTERS_reg[2][13]  ( .D(n7824), .CK(CLK), .RN(n6418), .Q(n4075), 
        .QN(n5992) );
  DFFR_X1 \REGISTERS_reg[2][12]  ( .D(n7825), .CK(CLK), .RN(n6418), .Q(n4074), 
        .QN(n5993) );
  DFFR_X1 \REGISTERS_reg[2][11]  ( .D(n7826), .CK(CLK), .RN(n6418), .Q(n4073), 
        .QN(n5994) );
  DFFR_X1 \REGISTERS_reg[2][10]  ( .D(n7827), .CK(CLK), .RN(n6418), .Q(n4072), 
        .QN(n5995) );
  DFFR_X1 \REGISTERS_reg[2][9]  ( .D(n7828), .CK(CLK), .RN(n6418), .Q(n4071), 
        .QN(n5996) );
  DFFR_X1 \REGISTERS_reg[2][8]  ( .D(n7829), .CK(CLK), .RN(n6418), .Q(n4070), 
        .QN(n5997) );
  DFFR_X1 \REGISTERS_reg[2][7]  ( .D(n7830), .CK(CLK), .RN(n6417), .Q(n4069), 
        .QN(n5998) );
  DFFR_X1 \REGISTERS_reg[2][6]  ( .D(n7831), .CK(CLK), .RN(n6417), .Q(n4068), 
        .QN(n5999) );
  DFFR_X1 \REGISTERS_reg[2][5]  ( .D(n7832), .CK(CLK), .RN(n6417), .Q(n4067), 
        .QN(n6000) );
  DFFR_X1 \REGISTERS_reg[2][4]  ( .D(n7833), .CK(CLK), .RN(n6417), .Q(n4066), 
        .QN(n6001) );
  DFFR_X1 \REGISTERS_reg[2][3]  ( .D(n7834), .CK(CLK), .RN(n6427), .Q(n4065), 
        .QN(n6002) );
  DFFR_X1 \REGISTERS_reg[2][2]  ( .D(n7835), .CK(CLK), .RN(n6427), .Q(n4064), 
        .QN(n6003) );
  DFFR_X1 \REGISTERS_reg[2][1]  ( .D(n7836), .CK(CLK), .RN(n6427), .Q(n4063), 
        .QN(n6004) );
  DFFR_X1 \REGISTERS_reg[2][0]  ( .D(n7837), .CK(CLK), .RN(n6427), .Q(n4062), 
        .QN(n5974) );
  DFFR_X1 \REGISTERS_reg[28][31]  ( .D(n3110), .CK(CLK), .RN(n6410), .Q(n5681), 
        .QN(n2091) );
  DFFR_X1 \REGISTERS_reg[28][30]  ( .D(n3109), .CK(CLK), .RN(n6410), .Q(n5682), 
        .QN(n2090) );
  DFFR_X1 \REGISTERS_reg[28][29]  ( .D(n3108), .CK(CLK), .RN(n6410), .Q(n5683), 
        .QN(n2089) );
  DFFR_X1 \REGISTERS_reg[28][28]  ( .D(n3107), .CK(CLK), .RN(n6410), .Q(n5684), 
        .QN(n2088) );
  DFFR_X1 \REGISTERS_reg[28][27]  ( .D(n3106), .CK(CLK), .RN(n6410), .Q(n5685), 
        .QN(n2087) );
  DFFR_X1 \REGISTERS_reg[28][26]  ( .D(n3105), .CK(CLK), .RN(n6410), .Q(n5686), 
        .QN(n2086) );
  DFFR_X1 \REGISTERS_reg[28][25]  ( .D(n3104), .CK(CLK), .RN(n6410), .Q(n5687), 
        .QN(n2085) );
  DFFR_X1 \REGISTERS_reg[28][24]  ( .D(n3103), .CK(CLK), .RN(n6410), .Q(n5688), 
        .QN(n2084) );
  DFFR_X1 \REGISTERS_reg[28][23]  ( .D(n3102), .CK(CLK), .RN(n6410), .Q(n5689), 
        .QN(n2083) );
  DFFR_X1 \REGISTERS_reg[28][22]  ( .D(n3101), .CK(CLK), .RN(n6410), .Q(n5690), 
        .QN(n2082) );
  DFFR_X1 \REGISTERS_reg[28][21]  ( .D(n3100), .CK(CLK), .RN(n6410), .Q(n5691), 
        .QN(n2081) );
  DFFR_X1 \REGISTERS_reg[28][20]  ( .D(n3099), .CK(CLK), .RN(n6410), .Q(n5692), 
        .QN(n2080) );
  DFFR_X1 \REGISTERS_reg[28][19]  ( .D(n3098), .CK(CLK), .RN(n6409), .Q(n5693), 
        .QN(n2079) );
  DFFR_X1 \REGISTERS_reg[28][18]  ( .D(n3097), .CK(CLK), .RN(n6409), .Q(n5694), 
        .QN(n2078) );
  DFFR_X1 \REGISTERS_reg[28][17]  ( .D(n3096), .CK(CLK), .RN(n6409), .Q(n5695), 
        .QN(n2077) );
  DFFR_X1 \REGISTERS_reg[28][16]  ( .D(n3095), .CK(CLK), .RN(n6409), .Q(n5696), 
        .QN(n2076) );
  DFFR_X1 \REGISTERS_reg[28][15]  ( .D(n3094), .CK(CLK), .RN(n6409), .Q(n5697), 
        .QN(n2075) );
  DFFR_X1 \REGISTERS_reg[28][14]  ( .D(n3093), .CK(CLK), .RN(n6409), .Q(n5698), 
        .QN(n2074) );
  DFFR_X1 \REGISTERS_reg[28][13]  ( .D(n3092), .CK(CLK), .RN(n6409), .Q(n5699), 
        .QN(n2073) );
  DFFR_X1 \REGISTERS_reg[28][12]  ( .D(n3091), .CK(CLK), .RN(n6409), .Q(n5700), 
        .QN(n2072) );
  DFFR_X1 \REGISTERS_reg[28][11]  ( .D(n3090), .CK(CLK), .RN(n6409), .Q(n5701), 
        .QN(n2071) );
  DFFR_X1 \REGISTERS_reg[28][10]  ( .D(n3089), .CK(CLK), .RN(n6409), .Q(n5702), 
        .QN(n2070) );
  DFFR_X1 \REGISTERS_reg[28][9]  ( .D(n3088), .CK(CLK), .RN(n6409), .Q(n5703), 
        .QN(n2069) );
  DFFR_X1 \REGISTERS_reg[28][8]  ( .D(n3087), .CK(CLK), .RN(n6409), .Q(n5704), 
        .QN(n2068) );
  DFFR_X1 \REGISTERS_reg[28][7]  ( .D(n3086), .CK(CLK), .RN(n6408), .Q(n5705), 
        .QN(n2067) );
  DFFR_X1 \REGISTERS_reg[28][6]  ( .D(n3085), .CK(CLK), .RN(n6408), .Q(n5706), 
        .QN(n2066) );
  DFFR_X1 \REGISTERS_reg[28][5]  ( .D(n3084), .CK(CLK), .RN(n6408), .Q(n5707), 
        .QN(n2065) );
  DFFR_X1 \REGISTERS_reg[28][4]  ( .D(n3083), .CK(CLK), .RN(n6408), .Q(n5708), 
        .QN(n2064) );
  DFFR_X1 \REGISTERS_reg[28][3]  ( .D(n3082), .CK(CLK), .RN(n6408), .Q(n5709), 
        .QN(n2063) );
  DFFR_X1 \REGISTERS_reg[28][2]  ( .D(n3081), .CK(CLK), .RN(n6408), .Q(n5710), 
        .QN(n2062) );
  DFFR_X1 \REGISTERS_reg[28][1]  ( .D(n3080), .CK(CLK), .RN(n6408), .Q(n5711), 
        .QN(n2061) );
  DFFR_X1 \REGISTERS_reg[28][0]  ( .D(n3079), .CK(CLK), .RN(n6408), .Q(n5358), 
        .QN(n2060) );
  DFFR_X1 \REGISTERS_reg[18][31]  ( .D(n3302), .CK(CLK), .RN(n6460), .Q(n5744), 
        .QN(n2251) );
  DFFR_X1 \REGISTERS_reg[27][31]  ( .D(n4541), .CK(CLK), .RN(n6382), .Q(n5391), 
        .QN(n2123) );
  DFFR_X1 \REGISTERS_reg[27][30]  ( .D(n4540), .CK(CLK), .RN(n6401), .Q(n5392), 
        .QN(n2122) );
  DFFR_X1 \REGISTERS_reg[27][29]  ( .D(n4539), .CK(CLK), .RN(n6401), .Q(n5393), 
        .QN(n2121) );
  DFFR_X1 \REGISTERS_reg[27][28]  ( .D(n4538), .CK(CLK), .RN(n6401), .Q(n5394), 
        .QN(n2120) );
  DFFR_X1 \REGISTERS_reg[27][27]  ( .D(n4537), .CK(CLK), .RN(n6401), .Q(n5395), 
        .QN(n2119) );
  DFFR_X1 \REGISTERS_reg[27][26]  ( .D(n4536), .CK(CLK), .RN(n6401), .Q(n5396), 
        .QN(n2118) );
  DFFR_X1 \REGISTERS_reg[27][25]  ( .D(n4535), .CK(CLK), .RN(n6401), .Q(n5397), 
        .QN(n2117) );
  DFFR_X1 \REGISTERS_reg[27][24]  ( .D(n4534), .CK(CLK), .RN(n6401), .Q(n5398), 
        .QN(n2116) );
  DFFR_X1 \REGISTERS_reg[27][23]  ( .D(n4533), .CK(CLK), .RN(n6401), .Q(n5399), 
        .QN(n2115) );
  DFFR_X1 \REGISTERS_reg[27][22]  ( .D(n4532), .CK(CLK), .RN(n6400), .Q(n5400), 
        .QN(n2114) );
  DFFR_X1 \REGISTERS_reg[27][21]  ( .D(n4531), .CK(CLK), .RN(n6400), .Q(n5401), 
        .QN(n2113) );
  DFFR_X1 \REGISTERS_reg[27][20]  ( .D(n4530), .CK(CLK), .RN(n6400), .Q(n5402), 
        .QN(n2112) );
  DFFR_X1 \REGISTERS_reg[27][19]  ( .D(n4529), .CK(CLK), .RN(n6400), .Q(n5403), 
        .QN(n2111) );
  DFFR_X1 \REGISTERS_reg[27][18]  ( .D(n4528), .CK(CLK), .RN(n6400), .Q(n5404), 
        .QN(n2110) );
  DFFR_X1 \REGISTERS_reg[27][17]  ( .D(n4527), .CK(CLK), .RN(n6400), .Q(n5405), 
        .QN(n2109) );
  DFFR_X1 \REGISTERS_reg[27][16]  ( .D(n4526), .CK(CLK), .RN(n6400), .Q(n5406), 
        .QN(n2108) );
  DFFR_X1 \REGISTERS_reg[27][15]  ( .D(n4525), .CK(CLK), .RN(n6400), .Q(n5407), 
        .QN(n2107) );
  DFFR_X1 \REGISTERS_reg[27][14]  ( .D(n4524), .CK(CLK), .RN(n6400), .Q(n5408), 
        .QN(n2106) );
  DFFR_X1 \REGISTERS_reg[27][13]  ( .D(n4523), .CK(CLK), .RN(n6400), .Q(n5409), 
        .QN(n2105) );
  DFFR_X1 \REGISTERS_reg[27][12]  ( .D(n4522), .CK(CLK), .RN(n6400), .Q(n5410), 
        .QN(n2104) );
  DFFR_X1 \REGISTERS_reg[27][11]  ( .D(n4521), .CK(CLK), .RN(n6411), .Q(n5411), 
        .QN(n2103) );
  DFFR_X1 \REGISTERS_reg[27][10]  ( .D(n4520), .CK(CLK), .RN(n6411), .Q(n5412), 
        .QN(n2102) );
  DFFR_X1 \REGISTERS_reg[27][9]  ( .D(n4519), .CK(CLK), .RN(n6411), .Q(n5413), 
        .QN(n2101) );
  DFFR_X1 \REGISTERS_reg[27][8]  ( .D(n4518), .CK(CLK), .RN(n6411), .Q(n5414), 
        .QN(n2100) );
  DFFR_X1 \REGISTERS_reg[27][7]  ( .D(n4517), .CK(CLK), .RN(n6411), .Q(n5415), 
        .QN(n2099) );
  DFFR_X1 \REGISTERS_reg[27][6]  ( .D(n4516), .CK(CLK), .RN(n6411), .Q(n5416), 
        .QN(n2098) );
  DFFR_X1 \REGISTERS_reg[27][5]  ( .D(n4515), .CK(CLK), .RN(n6411), .Q(n5417), 
        .QN(n2097) );
  DFFR_X1 \REGISTERS_reg[27][4]  ( .D(n4514), .CK(CLK), .RN(n6411), .Q(n5418), 
        .QN(n2096) );
  DFFR_X1 \REGISTERS_reg[27][3]  ( .D(n4513), .CK(CLK), .RN(n6411), .Q(n5419), 
        .QN(n2095) );
  DFFR_X1 \REGISTERS_reg[27][2]  ( .D(n4512), .CK(CLK), .RN(n6411), .Q(n5420), 
        .QN(n2094) );
  DFFR_X1 \REGISTERS_reg[27][1]  ( .D(n4511), .CK(CLK), .RN(n6411), .Q(n5421), 
        .QN(n2093) );
  DFFR_X1 \REGISTERS_reg[27][0]  ( .D(n4510), .CK(CLK), .RN(n6411), .Q(n5546), 
        .QN(n2092) );
  DFFR_X1 \REGISTERS_reg[4][31]  ( .D(n4317), .CK(CLK), .RN(n6425), .Q(n5875), 
        .QN(n2315) );
  DFFR_X1 \REGISTERS_reg[4][30]  ( .D(n4316), .CK(CLK), .RN(n6425), .Q(n5298), 
        .QN(n2314) );
  DFFR_X1 \REGISTERS_reg[4][29]  ( .D(n4315), .CK(CLK), .RN(n6425), .Q(n5299), 
        .QN(n2313) );
  DFFR_X1 \REGISTERS_reg[4][28]  ( .D(n4314), .CK(CLK), .RN(n6425), .Q(n5300), 
        .QN(n2312) );
  DFFR_X1 \REGISTERS_reg[4][27]  ( .D(n4313), .CK(CLK), .RN(n6425), .Q(n5301), 
        .QN(n2311) );
  DFFR_X1 \REGISTERS_reg[4][26]  ( .D(n4312), .CK(CLK), .RN(n6425), .Q(n5302), 
        .QN(n2310) );
  DFFR_X1 \REGISTERS_reg[4][25]  ( .D(n4311), .CK(CLK), .RN(n6425), .Q(n5303), 
        .QN(n2309) );
  DFFR_X1 \REGISTERS_reg[4][24]  ( .D(n4310), .CK(CLK), .RN(n6425), .Q(n5304), 
        .QN(n2308) );
  DFFR_X1 \REGISTERS_reg[4][23]  ( .D(n4309), .CK(CLK), .RN(n6424), .Q(n5305), 
        .QN(n2307) );
  DFFR_X1 \REGISTERS_reg[4][22]  ( .D(n4308), .CK(CLK), .RN(n6424), .Q(n5306), 
        .QN(n2306) );
  DFFR_X1 \REGISTERS_reg[4][21]  ( .D(n4307), .CK(CLK), .RN(n6424), .Q(n5307), 
        .QN(n2305) );
  DFFR_X1 \REGISTERS_reg[4][20]  ( .D(n4306), .CK(CLK), .RN(n6424), .Q(n5308), 
        .QN(n2304) );
  DFFR_X1 \REGISTERS_reg[4][19]  ( .D(n4305), .CK(CLK), .RN(n6424), .Q(n5309), 
        .QN(n2303) );
  DFFR_X1 \REGISTERS_reg[4][18]  ( .D(n4304), .CK(CLK), .RN(n6424), .Q(n5310), 
        .QN(n2302) );
  DFFR_X1 \REGISTERS_reg[4][17]  ( .D(n4303), .CK(CLK), .RN(n6424), .Q(n5311), 
        .QN(n2301) );
  DFFR_X1 \REGISTERS_reg[4][16]  ( .D(n4302), .CK(CLK), .RN(n6424), .Q(n5312), 
        .QN(n2300) );
  DFFR_X1 \REGISTERS_reg[4][15]  ( .D(n4301), .CK(CLK), .RN(n6424), .Q(n5313), 
        .QN(n2299) );
  DFFR_X1 \REGISTERS_reg[4][14]  ( .D(n4300), .CK(CLK), .RN(n6424), .Q(n5314), 
        .QN(n2298) );
  DFFR_X1 \REGISTERS_reg[4][13]  ( .D(n4299), .CK(CLK), .RN(n6424), .Q(n5315), 
        .QN(n2297) );
  DFFR_X1 \REGISTERS_reg[4][12]  ( .D(n4298), .CK(CLK), .RN(n6424), .Q(n5316), 
        .QN(n2296) );
  DFFR_X1 \REGISTERS_reg[4][11]  ( .D(n4297), .CK(CLK), .RN(n6423), .Q(n5317), 
        .QN(n2295) );
  DFFR_X1 \REGISTERS_reg[4][10]  ( .D(n4296), .CK(CLK), .RN(n6423), .Q(n5318), 
        .QN(n2294) );
  DFFR_X1 \REGISTERS_reg[4][9]  ( .D(n4295), .CK(CLK), .RN(n6423), .Q(n5319), 
        .QN(n2293) );
  DFFR_X1 \REGISTERS_reg[4][8]  ( .D(n4294), .CK(CLK), .RN(n6423), .Q(n5320), 
        .QN(n2292) );
  DFFR_X1 \REGISTERS_reg[4][7]  ( .D(n4293), .CK(CLK), .RN(n6423), .Q(n5321), 
        .QN(n2291) );
  DFFR_X1 \REGISTERS_reg[4][6]  ( .D(n4292), .CK(CLK), .RN(n6423), .Q(n5322), 
        .QN(n2290) );
  DFFR_X1 \REGISTERS_reg[4][5]  ( .D(n4291), .CK(CLK), .RN(n6423), .Q(n5323), 
        .QN(n2289) );
  DFFR_X1 \REGISTERS_reg[4][4]  ( .D(n4290), .CK(CLK), .RN(n6423), .Q(n5324), 
        .QN(n2288) );
  DFFR_X1 \REGISTERS_reg[4][3]  ( .D(n4289), .CK(CLK), .RN(n6423), .Q(n5325), 
        .QN(n2287) );
  DFFR_X1 \REGISTERS_reg[4][2]  ( .D(n4288), .CK(CLK), .RN(n6423), .Q(n5326), 
        .QN(n2286) );
  DFFR_X1 \REGISTERS_reg[4][1]  ( .D(n4287), .CK(CLK), .RN(n6423), .Q(n5327), 
        .QN(n2285) );
  DFFR_X1 \REGISTERS_reg[4][0]  ( .D(n4286), .CK(CLK), .RN(n6423), .Q(n5876), 
        .QN(n2284) );
  DFFR_X1 \REGISTERS_reg[26][31]  ( .D(n4509), .CK(CLK), .RN(n6404), .Q(n5649), 
        .QN(n2155) );
  DFFR_X1 \REGISTERS_reg[26][30]  ( .D(n4508), .CK(CLK), .RN(n6404), .Q(n5650), 
        .QN(n2154) );
  DFFR_X1 \REGISTERS_reg[26][29]  ( .D(n4507), .CK(CLK), .RN(n6404), .Q(n5651), 
        .QN(n2153) );
  DFFR_X1 \REGISTERS_reg[26][28]  ( .D(n4506), .CK(CLK), .RN(n6404), .Q(n5652), 
        .QN(n2152) );
  DFFR_X1 \REGISTERS_reg[26][27]  ( .D(n4505), .CK(CLK), .RN(n6403), .Q(n5653), 
        .QN(n2151) );
  DFFR_X1 \REGISTERS_reg[26][26]  ( .D(n4504), .CK(CLK), .RN(n6403), .Q(n5654), 
        .QN(n2150) );
  DFFR_X1 \REGISTERS_reg[26][25]  ( .D(n4503), .CK(CLK), .RN(n6403), .Q(n5655), 
        .QN(n2149) );
  DFFR_X1 \REGISTERS_reg[26][24]  ( .D(n4502), .CK(CLK), .RN(n6403), .Q(n5656), 
        .QN(n2148) );
  DFFR_X1 \REGISTERS_reg[26][23]  ( .D(n4501), .CK(CLK), .RN(n6403), .Q(n5657), 
        .QN(n2147) );
  DFFR_X1 \REGISTERS_reg[26][22]  ( .D(n4500), .CK(CLK), .RN(n6403), .Q(n5658), 
        .QN(n2146) );
  DFFR_X1 \REGISTERS_reg[26][21]  ( .D(n4499), .CK(CLK), .RN(n6403), .Q(n5659), 
        .QN(n2145) );
  DFFR_X1 \REGISTERS_reg[26][20]  ( .D(n4498), .CK(CLK), .RN(n6403), .Q(n5660), 
        .QN(n2144) );
  DFFR_X1 \REGISTERS_reg[26][19]  ( .D(n4497), .CK(CLK), .RN(n6403), .Q(n5661), 
        .QN(n2143) );
  DFFR_X1 \REGISTERS_reg[26][18]  ( .D(n4496), .CK(CLK), .RN(n6403), .Q(n5662), 
        .QN(n2142) );
  DFFR_X1 \REGISTERS_reg[26][17]  ( .D(n4495), .CK(CLK), .RN(n6403), .Q(n5663), 
        .QN(n2141) );
  DFFR_X1 \REGISTERS_reg[26][16]  ( .D(n4494), .CK(CLK), .RN(n6403), .Q(n5664), 
        .QN(n2140) );
  DFFR_X1 \REGISTERS_reg[26][15]  ( .D(n4493), .CK(CLK), .RN(n6402), .Q(n5665), 
        .QN(n2139) );
  DFFR_X1 \REGISTERS_reg[26][14]  ( .D(n4492), .CK(CLK), .RN(n6402), .Q(n5666), 
        .QN(n2138) );
  DFFR_X1 \REGISTERS_reg[26][13]  ( .D(n4491), .CK(CLK), .RN(n6402), .Q(n5667), 
        .QN(n2137) );
  DFFR_X1 \REGISTERS_reg[26][12]  ( .D(n4490), .CK(CLK), .RN(n6402), .Q(n5668), 
        .QN(n2136) );
  DFFR_X1 \REGISTERS_reg[26][11]  ( .D(n4489), .CK(CLK), .RN(n6402), .Q(n5669), 
        .QN(n2135) );
  DFFR_X1 \REGISTERS_reg[26][10]  ( .D(n4488), .CK(CLK), .RN(n6402), .Q(n5670), 
        .QN(n2134) );
  DFFR_X1 \REGISTERS_reg[26][9]  ( .D(n4487), .CK(CLK), .RN(n6402), .Q(n5671), 
        .QN(n2133) );
  DFFR_X1 \REGISTERS_reg[26][8]  ( .D(n4486), .CK(CLK), .RN(n6402), .Q(n5672), 
        .QN(n2132) );
  DFFR_X1 \REGISTERS_reg[26][7]  ( .D(n4485), .CK(CLK), .RN(n6402), .Q(n5673), 
        .QN(n2131) );
  DFFR_X1 \REGISTERS_reg[26][6]  ( .D(n4484), .CK(CLK), .RN(n6402), .Q(n5674), 
        .QN(n2130) );
  DFFR_X1 \REGISTERS_reg[26][5]  ( .D(n4483), .CK(CLK), .RN(n6402), .Q(n5675), 
        .QN(n2129) );
  DFFR_X1 \REGISTERS_reg[26][4]  ( .D(n4482), .CK(CLK), .RN(n6402), .Q(n5676), 
        .QN(n2128) );
  DFFR_X1 \REGISTERS_reg[26][3]  ( .D(n4481), .CK(CLK), .RN(n6401), .Q(n5677), 
        .QN(n2127) );
  DFFR_X1 \REGISTERS_reg[26][2]  ( .D(n4480), .CK(CLK), .RN(n6401), .Q(n5678), 
        .QN(n2126) );
  DFFR_X1 \REGISTERS_reg[26][1]  ( .D(n4479), .CK(CLK), .RN(n6401), .Q(n5679), 
        .QN(n2125) );
  DFFR_X1 \REGISTERS_reg[26][0]  ( .D(n4478), .CK(CLK), .RN(n6401), .Q(n5648), 
        .QN(n2124) );
  DFFR_X1 \REGISTERS_reg[17][31]  ( .D(n4413), .CK(CLK), .RN(n6463), .Q(n5168), 
        .QN(n2283) );
  DFFR_X1 \REGISTERS_reg[17][30]  ( .D(n4412), .CK(CLK), .RN(n6463), .Q(n5361), 
        .QN(n2282) );
  DFFR_X1 \REGISTERS_reg[17][29]  ( .D(n4411), .CK(CLK), .RN(n6463), .Q(n5362), 
        .QN(n2281) );
  DFFR_X1 \REGISTERS_reg[17][28]  ( .D(n4410), .CK(CLK), .RN(n6463), .Q(n5363), 
        .QN(n2280) );
  DFFR_X1 \REGISTERS_reg[17][27]  ( .D(n4409), .CK(CLK), .RN(n6462), .Q(n5364), 
        .QN(n2279) );
  DFFR_X1 \REGISTERS_reg[17][26]  ( .D(n4408), .CK(CLK), .RN(n6462), .Q(n5365), 
        .QN(n2278) );
  DFFR_X1 \REGISTERS_reg[17][25]  ( .D(n4407), .CK(CLK), .RN(n6462), .Q(n5366), 
        .QN(n2277) );
  DFFR_X1 \REGISTERS_reg[17][24]  ( .D(n4406), .CK(CLK), .RN(n6462), .Q(n5367), 
        .QN(n2276) );
  DFFR_X1 \REGISTERS_reg[17][23]  ( .D(n4405), .CK(CLK), .RN(n6462), .Q(n5368), 
        .QN(n2275) );
  DFFR_X1 \REGISTERS_reg[17][22]  ( .D(n4404), .CK(CLK), .RN(n6462), .Q(n5369), 
        .QN(n2274) );
  DFFR_X1 \REGISTERS_reg[17][21]  ( .D(n4403), .CK(CLK), .RN(n6462), .Q(n5370), 
        .QN(n2273) );
  DFFR_X1 \REGISTERS_reg[17][20]  ( .D(n4402), .CK(CLK), .RN(n6462), .Q(n5371), 
        .QN(n2272) );
  DFFR_X1 \REGISTERS_reg[17][19]  ( .D(n4401), .CK(CLK), .RN(n6461), .Q(n5372), 
        .QN(n2271) );
  DFFR_X1 \REGISTERS_reg[17][18]  ( .D(n4400), .CK(CLK), .RN(n6461), .Q(n5373), 
        .QN(n2270) );
  DFFR_X1 \REGISTERS_reg[17][17]  ( .D(n4399), .CK(CLK), .RN(n6461), .Q(n5374), 
        .QN(n2269) );
  DFFR_X1 \REGISTERS_reg[17][16]  ( .D(n4398), .CK(CLK), .RN(n6461), .Q(n5375), 
        .QN(n2268) );
  DFFR_X1 \REGISTERS_reg[17][15]  ( .D(n4397), .CK(CLK), .RN(n6461), .Q(n5376), 
        .QN(n2267) );
  DFFR_X1 \REGISTERS_reg[17][14]  ( .D(n4396), .CK(CLK), .RN(n6461), .Q(n5377), 
        .QN(n2266) );
  DFFR_X1 \REGISTERS_reg[17][13]  ( .D(n4395), .CK(CLK), .RN(n6461), .Q(n5378), 
        .QN(n2265) );
  DFFR_X1 \REGISTERS_reg[17][12]  ( .D(n4394), .CK(CLK), .RN(n6461), .Q(n5379), 
        .QN(n2264) );
  DFFR_X1 \REGISTERS_reg[17][11]  ( .D(n4393), .CK(CLK), .RN(n6461), .Q(n5380), 
        .QN(n2263) );
  DFFR_X1 \REGISTERS_reg[17][10]  ( .D(n4392), .CK(CLK), .RN(n6461), .Q(n5381), 
        .QN(n2262) );
  DFFR_X1 \REGISTERS_reg[17][9]  ( .D(n4391), .CK(CLK), .RN(n6461), .Q(n5382), 
        .QN(n2261) );
  DFFR_X1 \REGISTERS_reg[17][8]  ( .D(n4390), .CK(CLK), .RN(n6461), .Q(n5383), 
        .QN(n2260) );
  DFFR_X1 \REGISTERS_reg[17][7]  ( .D(n4389), .CK(CLK), .RN(n6460), .Q(n5384), 
        .QN(n2259) );
  DFFR_X1 \REGISTERS_reg[17][6]  ( .D(n4388), .CK(CLK), .RN(n6460), .Q(n5385), 
        .QN(n2258) );
  DFFR_X1 \REGISTERS_reg[17][5]  ( .D(n4387), .CK(CLK), .RN(n6460), .Q(n5386), 
        .QN(n2257) );
  DFFR_X1 \REGISTERS_reg[17][4]  ( .D(n4386), .CK(CLK), .RN(n6460), .Q(n5387), 
        .QN(n2256) );
  DFFR_X1 \REGISTERS_reg[17][3]  ( .D(n4385), .CK(CLK), .RN(n6459), .Q(n5388), 
        .QN(n2255) );
  DFFR_X1 \REGISTERS_reg[17][2]  ( .D(n4384), .CK(CLK), .RN(n6459), .Q(n5389), 
        .QN(n2254) );
  DFFR_X1 \REGISTERS_reg[17][1]  ( .D(n4383), .CK(CLK), .RN(n6459), .Q(n5390), 
        .QN(n2253) );
  DFFR_X1 \REGISTERS_reg[17][0]  ( .D(n4382), .CK(CLK), .RN(n6459), .Q(n5233), 
        .QN(n2252) );
  DFFR_X1 \REGISTERS_reg[5][31]  ( .D(n4349), .CK(CLK), .RN(n6422), .Q(n5809), 
        .QN(n4029) );
  DFFR_X1 \REGISTERS_reg[5][30]  ( .D(n4348), .CK(CLK), .RN(n6422), .Q(n5810), 
        .QN(n4028) );
  DFFR_X1 \REGISTERS_reg[5][29]  ( .D(n4347), .CK(CLK), .RN(n6422), .Q(n5811), 
        .QN(n4027) );
  DFFR_X1 \REGISTERS_reg[5][28]  ( .D(n4346), .CK(CLK), .RN(n6422), .Q(n5812), 
        .QN(n4026) );
  DFFR_X1 \REGISTERS_reg[5][27]  ( .D(n4345), .CK(CLK), .RN(n6434), .Q(n5813), 
        .QN(n4025) );
  DFFR_X1 \REGISTERS_reg[5][26]  ( .D(n4344), .CK(CLK), .RN(n6434), .Q(n5814), 
        .QN(n4024) );
  DFFR_X1 \REGISTERS_reg[5][25]  ( .D(n4343), .CK(CLK), .RN(n6434), .Q(n5815), 
        .QN(n4023) );
  DFFR_X1 \REGISTERS_reg[5][24]  ( .D(n4342), .CK(CLK), .RN(n6434), .Q(n5816), 
        .QN(n4022) );
  DFFR_X1 \REGISTERS_reg[5][23]  ( .D(n4341), .CK(CLK), .RN(n6434), .Q(n5817), 
        .QN(n4021) );
  DFFR_X1 \REGISTERS_reg[5][22]  ( .D(n4340), .CK(CLK), .RN(n6434), .Q(n5818), 
        .QN(n4020) );
  DFFR_X1 \REGISTERS_reg[5][21]  ( .D(n4339), .CK(CLK), .RN(n6434), .Q(n5819), 
        .QN(n4019) );
  DFFR_X1 \REGISTERS_reg[5][20]  ( .D(n4338), .CK(CLK), .RN(n6434), .Q(n5820), 
        .QN(n4018) );
  DFFR_X1 \REGISTERS_reg[5][19]  ( .D(n4337), .CK(CLK), .RN(n6433), .Q(n5821), 
        .QN(n4017) );
  DFFR_X1 \REGISTERS_reg[5][18]  ( .D(n4336), .CK(CLK), .RN(n6433), .Q(n5822), 
        .QN(n4016) );
  DFFR_X1 \REGISTERS_reg[5][17]  ( .D(n4335), .CK(CLK), .RN(n6433), .Q(n5823), 
        .QN(n4015) );
  DFFR_X1 \REGISTERS_reg[5][16]  ( .D(n4334), .CK(CLK), .RN(n6433), .Q(n5824), 
        .QN(n4014) );
  DFFR_X1 \REGISTERS_reg[5][15]  ( .D(n4333), .CK(CLK), .RN(n6433), .Q(n5825), 
        .QN(n4013) );
  DFFR_X1 \REGISTERS_reg[5][14]  ( .D(n4332), .CK(CLK), .RN(n6433), .Q(n5826), 
        .QN(n4012) );
  DFFR_X1 \REGISTERS_reg[5][13]  ( .D(n4331), .CK(CLK), .RN(n6433), .Q(n5827), 
        .QN(n4011) );
  DFFR_X1 \REGISTERS_reg[5][12]  ( .D(n4330), .CK(CLK), .RN(n6433), .Q(n5828), 
        .QN(n4010) );
  DFFR_X1 \REGISTERS_reg[5][11]  ( .D(n4329), .CK(CLK), .RN(n6433), .Q(n5829), 
        .QN(n4009) );
  DFFR_X1 \REGISTERS_reg[5][10]  ( .D(n4328), .CK(CLK), .RN(n6433), .Q(n5830), 
        .QN(n4008) );
  DFFR_X1 \REGISTERS_reg[5][9]  ( .D(n4327), .CK(CLK), .RN(n6433), .Q(n5831), 
        .QN(n4007) );
  DFFR_X1 \REGISTERS_reg[5][8]  ( .D(n4326), .CK(CLK), .RN(n6433), .Q(n5832), 
        .QN(n4006) );
  DFFR_X1 \REGISTERS_reg[5][7]  ( .D(n4325), .CK(CLK), .RN(n6432), .Q(n5833), 
        .QN(n4005) );
  DFFR_X1 \REGISTERS_reg[5][6]  ( .D(n4324), .CK(CLK), .RN(n6432), .Q(n5834), 
        .QN(n4004) );
  DFFR_X1 \REGISTERS_reg[5][5]  ( .D(n4323), .CK(CLK), .RN(n6432), .Q(n5835), 
        .QN(n4003) );
  DFFR_X1 \REGISTERS_reg[5][4]  ( .D(n4322), .CK(CLK), .RN(n6432), .Q(n5836), 
        .QN(n4002) );
  DFFR_X1 \REGISTERS_reg[5][3]  ( .D(n4321), .CK(CLK), .RN(n6431), .Q(n5837), 
        .QN(n4001) );
  DFFR_X1 \REGISTERS_reg[5][2]  ( .D(n4320), .CK(CLK), .RN(n6431), .Q(n5838), 
        .QN(n4000) );
  DFFR_X1 \REGISTERS_reg[5][1]  ( .D(n4319), .CK(CLK), .RN(n6431), .Q(n5839), 
        .QN(n3999) );
  DFFR_X1 \REGISTERS_reg[5][0]  ( .D(n4318), .CK(CLK), .RN(n6431), .Q(n5840), 
        .QN(n3998) );
  DFFR_X1 \REGISTERS_reg[31][31]  ( .D(n4605), .CK(CLK), .RN(n6413), .Q(n5487), 
        .QN(n2717) );
  DFFR_X1 \REGISTERS_reg[31][30]  ( .D(n4604), .CK(CLK), .RN(n6413), .Q(n5488), 
        .QN(n2716) );
  DFFR_X1 \REGISTERS_reg[31][29]  ( .D(n4603), .CK(CLK), .RN(n6413), .Q(n5489), 
        .QN(n2715) );
  DFFR_X1 \REGISTERS_reg[31][28]  ( .D(n4602), .CK(CLK), .RN(n6413), .Q(n5490), 
        .QN(n2714) );
  DFFR_X1 \REGISTERS_reg[31][27]  ( .D(n4601), .CK(CLK), .RN(n6413), .Q(n5491), 
        .QN(n2713) );
  DFFR_X1 \REGISTERS_reg[31][26]  ( .D(n4600), .CK(CLK), .RN(n6413), .Q(n5492), 
        .QN(n2712) );
  DFFR_X1 \REGISTERS_reg[31][25]  ( .D(n4599), .CK(CLK), .RN(n6413), .Q(n5493), 
        .QN(n2711) );
  DFFR_X1 \REGISTERS_reg[31][24]  ( .D(n4598), .CK(CLK), .RN(n6413), .Q(n5494), 
        .QN(n2710) );
  DFFR_X1 \REGISTERS_reg[31][23]  ( .D(n4597), .CK(CLK), .RN(n6413), .Q(n5495), 
        .QN(n2709) );
  DFFR_X1 \REGISTERS_reg[31][22]  ( .D(n4596), .CK(CLK), .RN(n6413), .Q(n5496), 
        .QN(n2708) );
  DFFR_X1 \REGISTERS_reg[31][21]  ( .D(n4595), .CK(CLK), .RN(n6413), .Q(n5497), 
        .QN(n2707) );
  DFFR_X1 \REGISTERS_reg[31][20]  ( .D(n4594), .CK(CLK), .RN(n6413), .Q(n5498), 
        .QN(n2706) );
  DFFR_X1 \REGISTERS_reg[31][19]  ( .D(n4593), .CK(CLK), .RN(n6412), .Q(n5499), 
        .QN(n2705) );
  DFFR_X1 \REGISTERS_reg[31][18]  ( .D(n4592), .CK(CLK), .RN(n6412), .Q(n5500), 
        .QN(n2704) );
  DFFR_X1 \REGISTERS_reg[31][17]  ( .D(n4591), .CK(CLK), .RN(n6412), .Q(n5501), 
        .QN(n2703) );
  DFFR_X1 \REGISTERS_reg[31][16]  ( .D(n4590), .CK(CLK), .RN(n6412), .Q(n5502), 
        .QN(n2702) );
  DFFR_X1 \REGISTERS_reg[31][15]  ( .D(n4589), .CK(CLK), .RN(n6412), .Q(n5503), 
        .QN(n2701) );
  DFFR_X1 \REGISTERS_reg[31][14]  ( .D(n4588), .CK(CLK), .RN(n6412), .Q(n5504), 
        .QN(n2700) );
  DFFR_X1 \REGISTERS_reg[31][13]  ( .D(n4587), .CK(CLK), .RN(n6412), .Q(n5505), 
        .QN(n2699) );
  DFFR_X1 \REGISTERS_reg[31][12]  ( .D(n4586), .CK(CLK), .RN(n6412), .Q(n5506), 
        .QN(n2698) );
  DFFR_X1 \REGISTERS_reg[31][11]  ( .D(n4585), .CK(CLK), .RN(n6412), .Q(n5507), 
        .QN(n2697) );
  DFFR_X1 \REGISTERS_reg[31][10]  ( .D(n4584), .CK(CLK), .RN(n6412), .Q(n5508), 
        .QN(n2696) );
  DFFR_X1 \REGISTERS_reg[31][9]  ( .D(n4583), .CK(CLK), .RN(n6412), .Q(n5509), 
        .QN(n2695) );
  DFFR_X1 \REGISTERS_reg[31][8]  ( .D(n4582), .CK(CLK), .RN(n6412), .Q(n5510), 
        .QN(n2694) );
  DFFR_X1 \REGISTERS_reg[31][7]  ( .D(n4581), .CK(CLK), .RN(n6417), .Q(n5511), 
        .QN(n2693) );
  DFFR_X1 \REGISTERS_reg[31][6]  ( .D(n4580), .CK(CLK), .RN(n6417), .Q(n5512), 
        .QN(n2692) );
  DFFR_X1 \REGISTERS_reg[31][5]  ( .D(n4579), .CK(CLK), .RN(n6417), .Q(n5513), 
        .QN(n2691) );
  DFFR_X1 \REGISTERS_reg[31][4]  ( .D(n4578), .CK(CLK), .RN(n6417), .Q(n5514), 
        .QN(n2690) );
  DFFR_X1 \REGISTERS_reg[31][3]  ( .D(n4577), .CK(CLK), .RN(n6417), .Q(n998), 
        .QN(n5877) );
  DFFR_X1 \REGISTERS_reg[31][2]  ( .D(n4576), .CK(CLK), .RN(n6417), .Q(n982), 
        .QN(n5878) );
  DFFR_X1 \REGISTERS_reg[31][1]  ( .D(n4575), .CK(CLK), .RN(n6417), .Q(n966), 
        .QN(n5879) );
  DFFR_X1 \REGISTERS_reg[31][0]  ( .D(n4574), .CK(CLK), .RN(n6417), .Q(n950), 
        .QN(n5908) );
  DFFR_X1 \REGISTERS_reg[21][31]  ( .D(n4477), .CK(CLK), .RN(n6394), .Q(n5172), 
        .QN(n2973) );
  DFFR_X1 \REGISTERS_reg[21][30]  ( .D(n4476), .CK(CLK), .RN(n6394), .Q(n5173), 
        .QN(n2972) );
  DFFR_X1 \REGISTERS_reg[21][29]  ( .D(n4475), .CK(CLK), .RN(n6393), .Q(n5174), 
        .QN(n2971) );
  DFFR_X1 \REGISTERS_reg[21][28]  ( .D(n4474), .CK(CLK), .RN(n6393), .Q(n5175), 
        .QN(n2970) );
  DFFR_X1 \REGISTERS_reg[21][27]  ( .D(n4473), .CK(CLK), .RN(n6393), .Q(n5176), 
        .QN(n2969) );
  DFFR_X1 \REGISTERS_reg[21][26]  ( .D(n4472), .CK(CLK), .RN(n6393), .Q(n5177), 
        .QN(n2968) );
  DFFR_X1 \REGISTERS_reg[21][25]  ( .D(n4471), .CK(CLK), .RN(n6393), .Q(n5178), 
        .QN(n2967) );
  DFFR_X1 \REGISTERS_reg[21][24]  ( .D(n4470), .CK(CLK), .RN(n6393), .Q(n5179), 
        .QN(n2966) );
  DFFR_X1 \REGISTERS_reg[21][23]  ( .D(n4469), .CK(CLK), .RN(n6393), .Q(n5180), 
        .QN(n2965) );
  DFFR_X1 \REGISTERS_reg[21][22]  ( .D(n4468), .CK(CLK), .RN(n6393), .Q(n5181), 
        .QN(n2964) );
  DFFR_X1 \REGISTERS_reg[21][21]  ( .D(n4467), .CK(CLK), .RN(n6392), .Q(n5182), 
        .QN(n2963) );
  DFFR_X1 \REGISTERS_reg[21][20]  ( .D(n4466), .CK(CLK), .RN(n6392), .Q(n5183), 
        .QN(n2962) );
  DFFR_X1 \REGISTERS_reg[21][19]  ( .D(n4465), .CK(CLK), .RN(n6392), .Q(n5184), 
        .QN(n2961) );
  DFFR_X1 \REGISTERS_reg[21][18]  ( .D(n4464), .CK(CLK), .RN(n6392), .Q(n5185), 
        .QN(n2960) );
  DFFR_X1 \REGISTERS_reg[21][17]  ( .D(n4463), .CK(CLK), .RN(n6392), .Q(n5186), 
        .QN(n2959) );
  DFFR_X1 \REGISTERS_reg[21][16]  ( .D(n4462), .CK(CLK), .RN(n6392), .Q(n5187), 
        .QN(n2958) );
  DFFR_X1 \REGISTERS_reg[21][15]  ( .D(n4461), .CK(CLK), .RN(n6392), .Q(n5188), 
        .QN(n2957) );
  DFFR_X1 \REGISTERS_reg[21][14]  ( .D(n4460), .CK(CLK), .RN(n6392), .Q(n5189), 
        .QN(n2956) );
  DFFR_X1 \REGISTERS_reg[21][13]  ( .D(n4459), .CK(CLK), .RN(n6392), .Q(n5190), 
        .QN(n2955) );
  DFFR_X1 \REGISTERS_reg[21][12]  ( .D(n4458), .CK(CLK), .RN(n6392), .Q(n5191), 
        .QN(n2954) );
  DFFR_X1 \REGISTERS_reg[21][11]  ( .D(n4457), .CK(CLK), .RN(n6392), .Q(n5192), 
        .QN(n2953) );
  DFFR_X1 \REGISTERS_reg[21][10]  ( .D(n4456), .CK(CLK), .RN(n6392), .Q(n5193), 
        .QN(n2952) );
  DFFR_X1 \REGISTERS_reg[21][9]  ( .D(n4455), .CK(CLK), .RN(n6391), .Q(n5194), 
        .QN(n2951) );
  DFFR_X1 \REGISTERS_reg[21][8]  ( .D(n4454), .CK(CLK), .RN(n6391), .Q(n5195), 
        .QN(n2950) );
  DFFR_X1 \REGISTERS_reg[21][7]  ( .D(n4453), .CK(CLK), .RN(n6391), .Q(n5196), 
        .QN(n2949) );
  DFFR_X1 \REGISTERS_reg[21][6]  ( .D(n4452), .CK(CLK), .RN(n6391), .Q(n5197), 
        .QN(n2948) );
  DFFR_X1 \REGISTERS_reg[21][5]  ( .D(n4451), .CK(CLK), .RN(n6391), .Q(n5198), 
        .QN(n2947) );
  DFFR_X1 \REGISTERS_reg[21][4]  ( .D(n4450), .CK(CLK), .RN(n6391), .Q(n5199), 
        .QN(n2946) );
  DFFR_X1 \REGISTERS_reg[21][3]  ( .D(n4449), .CK(CLK), .RN(n6391), .Q(n5200), 
        .QN(n2945) );
  DFFR_X1 \REGISTERS_reg[21][2]  ( .D(n4448), .CK(CLK), .RN(n6391), .Q(n5201), 
        .QN(n2944) );
  DFFR_X1 \REGISTERS_reg[21][1]  ( .D(n4447), .CK(CLK), .RN(n6391), .Q(n5202), 
        .QN(n2943) );
  DFFR_X1 \REGISTERS_reg[21][0]  ( .D(n4446), .CK(CLK), .RN(n6391), .Q(n5359), 
        .QN(n2942) );
  DFFR_X1 \REGISTERS_reg[12][31]  ( .D(n4221), .CK(CLK), .RN(n6452), .Q(n5615), 
        .QN(n3805) );
  DFFR_X1 \REGISTERS_reg[12][30]  ( .D(n4220), .CK(CLK), .RN(n6452), .Q(n5616), 
        .QN(n3804) );
  DFFR_X1 \REGISTERS_reg[12][29]  ( .D(n4219), .CK(CLK), .RN(n6452), .Q(n5617), 
        .QN(n3803) );
  DFFR_X1 \REGISTERS_reg[12][28]  ( .D(n4218), .CK(CLK), .RN(n6452), .Q(n5618), 
        .QN(n3802) );
  DFFR_X1 \REGISTERS_reg[12][27]  ( .D(n4217), .CK(CLK), .RN(n6451), .Q(n5619), 
        .QN(n3801) );
  DFFR_X1 \REGISTERS_reg[12][26]  ( .D(n4216), .CK(CLK), .RN(n6451), .Q(n5620), 
        .QN(n3800) );
  DFFR_X1 \REGISTERS_reg[12][25]  ( .D(n4215), .CK(CLK), .RN(n6451), .Q(n5621), 
        .QN(n3799) );
  DFFR_X1 \REGISTERS_reg[12][24]  ( .D(n4214), .CK(CLK), .RN(n6451), .Q(n5622), 
        .QN(n3798) );
  DFFR_X1 \REGISTERS_reg[12][23]  ( .D(n4213), .CK(CLK), .RN(n6451), .Q(n5623), 
        .QN(n3797) );
  DFFR_X1 \REGISTERS_reg[12][22]  ( .D(n4212), .CK(CLK), .RN(n6451), .Q(n5624), 
        .QN(n3796) );
  DFFR_X1 \REGISTERS_reg[12][21]  ( .D(n4211), .CK(CLK), .RN(n6451), .Q(n5625), 
        .QN(n3795) );
  DFFR_X1 \REGISTERS_reg[12][20]  ( .D(n4210), .CK(CLK), .RN(n6451), .Q(n5626), 
        .QN(n3794) );
  DFFR_X1 \REGISTERS_reg[12][19]  ( .D(n4209), .CK(CLK), .RN(n6451), .Q(n5627), 
        .QN(n3793) );
  DFFR_X1 \REGISTERS_reg[12][18]  ( .D(n4208), .CK(CLK), .RN(n6451), .Q(n5628), 
        .QN(n3792) );
  DFFR_X1 \REGISTERS_reg[12][17]  ( .D(n4207), .CK(CLK), .RN(n6451), .Q(n5629), 
        .QN(n3791) );
  DFFR_X1 \REGISTERS_reg[12][16]  ( .D(n4206), .CK(CLK), .RN(n6451), .Q(n5630), 
        .QN(n3790) );
  DFFR_X1 \REGISTERS_reg[12][15]  ( .D(n4205), .CK(CLK), .RN(n6450), .Q(n5631), 
        .QN(n3789) );
  DFFR_X1 \REGISTERS_reg[12][14]  ( .D(n4204), .CK(CLK), .RN(n6450), .Q(n5632), 
        .QN(n3788) );
  DFFR_X1 \REGISTERS_reg[12][13]  ( .D(n4203), .CK(CLK), .RN(n6450), .Q(n5633), 
        .QN(n3787) );
  DFFR_X1 \REGISTERS_reg[12][12]  ( .D(n4202), .CK(CLK), .RN(n6450), .Q(n5634), 
        .QN(n3786) );
  DFFR_X1 \REGISTERS_reg[12][11]  ( .D(n4201), .CK(CLK), .RN(n6450), .Q(n5635), 
        .QN(n3785) );
  DFFR_X1 \REGISTERS_reg[12][10]  ( .D(n4200), .CK(CLK), .RN(n6450), .Q(n5636), 
        .QN(n3784) );
  DFFR_X1 \REGISTERS_reg[12][9]  ( .D(n4199), .CK(CLK), .RN(n6450), .Q(n5637), 
        .QN(n3783) );
  DFFR_X1 \REGISTERS_reg[12][8]  ( .D(n4198), .CK(CLK), .RN(n6450), .Q(n5638), 
        .QN(n3782) );
  DFFR_X1 \REGISTERS_reg[12][7]  ( .D(n4197), .CK(CLK), .RN(n6450), .Q(n5639), 
        .QN(n3781) );
  DFFR_X1 \REGISTERS_reg[12][6]  ( .D(n4196), .CK(CLK), .RN(n6450), .Q(n5640), 
        .QN(n3780) );
  DFFR_X1 \REGISTERS_reg[12][5]  ( .D(n4195), .CK(CLK), .RN(n6450), .Q(n5641), 
        .QN(n3779) );
  DFFR_X1 \REGISTERS_reg[12][4]  ( .D(n4194), .CK(CLK), .RN(n6450), .Q(n5642), 
        .QN(n3778) );
  DFFR_X1 \REGISTERS_reg[12][3]  ( .D(n4193), .CK(CLK), .RN(n6449), .Q(n5643), 
        .QN(n3777) );
  DFFR_X1 \REGISTERS_reg[12][2]  ( .D(n4192), .CK(CLK), .RN(n6449), .Q(n5644), 
        .QN(n3776) );
  DFFR_X1 \REGISTERS_reg[12][1]  ( .D(n4191), .CK(CLK), .RN(n6449), .Q(n5645), 
        .QN(n3775) );
  DFFR_X1 \REGISTERS_reg[12][0]  ( .D(n4190), .CK(CLK), .RN(n6449), .Q(n5646), 
        .QN(n3774) );
  DFFR_X1 \REGISTERS_reg[8][31]  ( .D(n4157), .CK(CLK), .RN(n6438), .Q(n5777), 
        .QN(n3933) );
  DFFR_X1 \REGISTERS_reg[8][30]  ( .D(n4156), .CK(CLK), .RN(n6438), .Q(n5778), 
        .QN(n3932) );
  DFFR_X1 \REGISTERS_reg[8][29]  ( .D(n4155), .CK(CLK), .RN(n6438), .Q(n5779), 
        .QN(n3931) );
  DFFR_X1 \REGISTERS_reg[8][28]  ( .D(n4154), .CK(CLK), .RN(n6438), .Q(n5780), 
        .QN(n3930) );
  DFFR_X1 \REGISTERS_reg[8][27]  ( .D(n4153), .CK(CLK), .RN(n6438), .Q(n5781), 
        .QN(n3929) );
  DFFR_X1 \REGISTERS_reg[8][26]  ( .D(n4152), .CK(CLK), .RN(n6438), .Q(n5782), 
        .QN(n3928) );
  DFFR_X1 \REGISTERS_reg[8][25]  ( .D(n4151), .CK(CLK), .RN(n6438), .Q(n5783), 
        .QN(n3927) );
  DFFR_X1 \REGISTERS_reg[8][24]  ( .D(n4150), .CK(CLK), .RN(n6438), .Q(n5784), 
        .QN(n3926) );
  DFFR_X1 \REGISTERS_reg[8][23]  ( .D(n4149), .CK(CLK), .RN(n6438), .Q(n5785), 
        .QN(n3925) );
  DFFR_X1 \REGISTERS_reg[8][22]  ( .D(n4148), .CK(CLK), .RN(n6438), .Q(n5786), 
        .QN(n3924) );
  DFFR_X1 \REGISTERS_reg[8][21]  ( .D(n4147), .CK(CLK), .RN(n6438), .Q(n5787), 
        .QN(n3923) );
  DFFR_X1 \REGISTERS_reg[8][20]  ( .D(n4146), .CK(CLK), .RN(n6438), .Q(n5788), 
        .QN(n3922) );
  DFFR_X1 \REGISTERS_reg[8][19]  ( .D(n4145), .CK(CLK), .RN(n6437), .Q(n5789), 
        .QN(n3921) );
  DFFR_X1 \REGISTERS_reg[8][18]  ( .D(n4144), .CK(CLK), .RN(n6437), .Q(n5790), 
        .QN(n3920) );
  DFFR_X1 \REGISTERS_reg[8][17]  ( .D(n4143), .CK(CLK), .RN(n6437), .Q(n5791), 
        .QN(n3919) );
  DFFR_X1 \REGISTERS_reg[8][16]  ( .D(n4142), .CK(CLK), .RN(n6437), .Q(n5792), 
        .QN(n3918) );
  DFFR_X1 \REGISTERS_reg[8][15]  ( .D(n4141), .CK(CLK), .RN(n6437), .Q(n5793), 
        .QN(n3917) );
  DFFR_X1 \REGISTERS_reg[8][14]  ( .D(n4140), .CK(CLK), .RN(n6437), .Q(n5794), 
        .QN(n3916) );
  DFFR_X1 \REGISTERS_reg[8][13]  ( .D(n4139), .CK(CLK), .RN(n6437), .Q(n5795), 
        .QN(n3915) );
  DFFR_X1 \REGISTERS_reg[8][12]  ( .D(n4138), .CK(CLK), .RN(n6437), .Q(n5796), 
        .QN(n3914) );
  DFFR_X1 \REGISTERS_reg[8][11]  ( .D(n4137), .CK(CLK), .RN(n6437), .Q(n5797), 
        .QN(n3913) );
  DFFR_X1 \REGISTERS_reg[8][10]  ( .D(n4136), .CK(CLK), .RN(n6437), .Q(n5798), 
        .QN(n3912) );
  DFFR_X1 \REGISTERS_reg[8][9]  ( .D(n4135), .CK(CLK), .RN(n6437), .Q(n5799), 
        .QN(n3911) );
  DFFR_X1 \REGISTERS_reg[8][8]  ( .D(n4134), .CK(CLK), .RN(n6437), .Q(n5800), 
        .QN(n3910) );
  DFFR_X1 \REGISTERS_reg[8][7]  ( .D(n4133), .CK(CLK), .RN(n6436), .Q(n5801), 
        .QN(n3909) );
  DFFR_X1 \REGISTERS_reg[8][6]  ( .D(n4132), .CK(CLK), .RN(n6436), .Q(n5802), 
        .QN(n3908) );
  DFFR_X1 \REGISTERS_reg[8][5]  ( .D(n4131), .CK(CLK), .RN(n6436), .Q(n5803), 
        .QN(n3907) );
  DFFR_X1 \REGISTERS_reg[8][4]  ( .D(n4130), .CK(CLK), .RN(n6436), .Q(n5804), 
        .QN(n3906) );
  DFFR_X1 \REGISTERS_reg[8][3]  ( .D(n4129), .CK(CLK), .RN(n6436), .Q(n5805), 
        .QN(n3905) );
  DFFR_X1 \REGISTERS_reg[8][2]  ( .D(n4128), .CK(CLK), .RN(n6436), .Q(n5806), 
        .QN(n3904) );
  DFFR_X1 \REGISTERS_reg[8][1]  ( .D(n4127), .CK(CLK), .RN(n6436), .Q(n5807), 
        .QN(n3903) );
  DFFR_X1 \REGISTERS_reg[8][0]  ( .D(n4126), .CK(CLK), .RN(n6436), .Q(n5808), 
        .QN(n3902) );
  DFFR_X1 \REGISTERS_reg[30][31]  ( .D(n4573), .CK(CLK), .RN(n6416), .Q(n5584), 
        .QN(n2749) );
  DFFR_X1 \REGISTERS_reg[30][30]  ( .D(n4572), .CK(CLK), .RN(n6416), .Q(n5585), 
        .QN(n2748) );
  DFFR_X1 \REGISTERS_reg[30][29]  ( .D(n4571), .CK(CLK), .RN(n6416), .Q(n5586), 
        .QN(n2747) );
  DFFR_X1 \REGISTERS_reg[30][28]  ( .D(n4570), .CK(CLK), .RN(n6416), .Q(n5587), 
        .QN(n2746) );
  DFFR_X1 \REGISTERS_reg[30][27]  ( .D(n4569), .CK(CLK), .RN(n6416), .Q(n5588), 
        .QN(n2745) );
  DFFR_X1 \REGISTERS_reg[30][26]  ( .D(n4568), .CK(CLK), .RN(n6416), .Q(n5589), 
        .QN(n2744) );
  DFFR_X1 \REGISTERS_reg[30][25]  ( .D(n4567), .CK(CLK), .RN(n6416), .Q(n5590), 
        .QN(n2743) );
  DFFR_X1 \REGISTERS_reg[30][24]  ( .D(n4566), .CK(CLK), .RN(n6416), .Q(n5591), 
        .QN(n2742) );
  DFFR_X1 \REGISTERS_reg[30][23]  ( .D(n4565), .CK(CLK), .RN(n6415), .Q(n5592), 
        .QN(n2741) );
  DFFR_X1 \REGISTERS_reg[30][22]  ( .D(n4564), .CK(CLK), .RN(n6415), .Q(n5593), 
        .QN(n2740) );
  DFFR_X1 \REGISTERS_reg[30][21]  ( .D(n4563), .CK(CLK), .RN(n6415), .Q(n5594), 
        .QN(n2739) );
  DFFR_X1 \REGISTERS_reg[30][20]  ( .D(n4562), .CK(CLK), .RN(n6415), .Q(n5595), 
        .QN(n2738) );
  DFFR_X1 \REGISTERS_reg[30][19]  ( .D(n4561), .CK(CLK), .RN(n6415), .Q(n5596), 
        .QN(n2737) );
  DFFR_X1 \REGISTERS_reg[30][18]  ( .D(n4560), .CK(CLK), .RN(n6415), .Q(n5597), 
        .QN(n2736) );
  DFFR_X1 \REGISTERS_reg[30][17]  ( .D(n4559), .CK(CLK), .RN(n6415), .Q(n5598), 
        .QN(n2735) );
  DFFR_X1 \REGISTERS_reg[30][16]  ( .D(n4558), .CK(CLK), .RN(n6415), .Q(n5599), 
        .QN(n2734) );
  DFFR_X1 \REGISTERS_reg[30][15]  ( .D(n4557), .CK(CLK), .RN(n6415), .Q(n5600), 
        .QN(n2733) );
  DFFR_X1 \REGISTERS_reg[30][14]  ( .D(n4556), .CK(CLK), .RN(n6415), .Q(n5601), 
        .QN(n2732) );
  DFFR_X1 \REGISTERS_reg[30][13]  ( .D(n4555), .CK(CLK), .RN(n6415), .Q(n5602), 
        .QN(n2731) );
  DFFR_X1 \REGISTERS_reg[30][12]  ( .D(n4554), .CK(CLK), .RN(n6415), .Q(n5603), 
        .QN(n2730) );
  DFFR_X1 \REGISTERS_reg[30][11]  ( .D(n4553), .CK(CLK), .RN(n6414), .Q(n5604), 
        .QN(n2729) );
  DFFR_X1 \REGISTERS_reg[30][10]  ( .D(n4552), .CK(CLK), .RN(n6414), .Q(n5605), 
        .QN(n2728) );
  DFFR_X1 \REGISTERS_reg[30][9]  ( .D(n4551), .CK(CLK), .RN(n6414), .Q(n5606), 
        .QN(n2727) );
  DFFR_X1 \REGISTERS_reg[30][8]  ( .D(n4550), .CK(CLK), .RN(n6414), .Q(n5607), 
        .QN(n2726) );
  DFFR_X1 \REGISTERS_reg[30][7]  ( .D(n4549), .CK(CLK), .RN(n6414), .Q(n5608), 
        .QN(n2725) );
  DFFR_X1 \REGISTERS_reg[30][6]  ( .D(n4548), .CK(CLK), .RN(n6414), .Q(n5609), 
        .QN(n2724) );
  DFFR_X1 \REGISTERS_reg[30][5]  ( .D(n4547), .CK(CLK), .RN(n6414), .Q(n5610), 
        .QN(n2723) );
  DFFR_X1 \REGISTERS_reg[30][4]  ( .D(n4546), .CK(CLK), .RN(n6414), .Q(n5611), 
        .QN(n2722) );
  DFFR_X1 \REGISTERS_reg[30][3]  ( .D(n4545), .CK(CLK), .RN(n6414), .Q(n5612), 
        .QN(n2721) );
  DFFR_X1 \REGISTERS_reg[30][2]  ( .D(n4544), .CK(CLK), .RN(n6414), .Q(n5613), 
        .QN(n2720) );
  DFFR_X1 \REGISTERS_reg[30][1]  ( .D(n4543), .CK(CLK), .RN(n6414), .Q(n5614), 
        .QN(n2719) );
  DFFR_X1 \REGISTERS_reg[30][0]  ( .D(n4542), .CK(CLK), .RN(n6414), .Q(n5360), 
        .QN(n2718) );
  DFFR_X1 \REGISTERS_reg[20][31]  ( .D(n4445), .CK(CLK), .RN(n6384), .Q(n5105), 
        .QN(n3581) );
  DFFR_X1 \REGISTERS_reg[20][30]  ( .D(n4444), .CK(CLK), .RN(n6384), .Q(n5106), 
        .QN(n3580) );
  DFFR_X1 \REGISTERS_reg[20][29]  ( .D(n4443), .CK(CLK), .RN(n6384), .Q(n5107), 
        .QN(n3579) );
  DFFR_X1 \REGISTERS_reg[20][28]  ( .D(n4442), .CK(CLK), .RN(n6384), .Q(n5108), 
        .QN(n3578) );
  DFFR_X1 \REGISTERS_reg[20][27]  ( .D(n4441), .CK(CLK), .RN(n6384), .Q(n5109), 
        .QN(n3577) );
  DFFR_X1 \REGISTERS_reg[20][26]  ( .D(n4440), .CK(CLK), .RN(n6384), .Q(n5110), 
        .QN(n3576) );
  DFFR_X1 \REGISTERS_reg[20][25]  ( .D(n4439), .CK(CLK), .RN(n6383), .Q(n5111), 
        .QN(n3575) );
  DFFR_X1 \REGISTERS_reg[20][24]  ( .D(n4438), .CK(CLK), .RN(n6383), .Q(n5112), 
        .QN(n3574) );
  DFFR_X1 \REGISTERS_reg[20][23]  ( .D(n4437), .CK(CLK), .RN(n6383), .Q(n5113), 
        .QN(n3573) );
  DFFR_X1 \REGISTERS_reg[20][22]  ( .D(n4436), .CK(CLK), .RN(n6383), .Q(n5114), 
        .QN(n3572) );
  DFFR_X1 \REGISTERS_reg[20][21]  ( .D(n4435), .CK(CLK), .RN(n6383), .Q(n5115), 
        .QN(n3571) );
  DFFR_X1 \REGISTERS_reg[20][20]  ( .D(n4434), .CK(CLK), .RN(n6383), .Q(n5116), 
        .QN(n3570) );
  DFFR_X1 \REGISTERS_reg[20][19]  ( .D(n4433), .CK(CLK), .RN(n6383), .Q(n5117), 
        .QN(n3569) );
  DFFR_X1 \REGISTERS_reg[20][18]  ( .D(n4432), .CK(CLK), .RN(n6383), .Q(n5118), 
        .QN(n3568) );
  DFFR_X1 \REGISTERS_reg[20][17]  ( .D(n4431), .CK(CLK), .RN(n6383), .Q(n5119), 
        .QN(n3567) );
  DFFR_X1 \REGISTERS_reg[20][16]  ( .D(n4430), .CK(CLK), .RN(n6383), .Q(n5120), 
        .QN(n3566) );
  DFFR_X1 \REGISTERS_reg[20][15]  ( .D(n4429), .CK(CLK), .RN(n6383), .Q(n5121), 
        .QN(n3565) );
  DFFR_X1 \REGISTERS_reg[20][14]  ( .D(n4428), .CK(CLK), .RN(n6383), .Q(n5122), 
        .QN(n3564) );
  DFFR_X1 \REGISTERS_reg[20][13]  ( .D(n4427), .CK(CLK), .RN(n6382), .Q(n5123), 
        .QN(n3563) );
  DFFR_X1 \REGISTERS_reg[20][12]  ( .D(n4426), .CK(CLK), .RN(n6382), .Q(n5124), 
        .QN(n3562) );
  DFFR_X1 \REGISTERS_reg[20][11]  ( .D(n4425), .CK(CLK), .RN(n6382), .Q(n5125), 
        .QN(n3561) );
  DFFR_X1 \REGISTERS_reg[20][10]  ( .D(n4424), .CK(CLK), .RN(n6382), .Q(n5126), 
        .QN(n3560) );
  DFFR_X1 \REGISTERS_reg[20][9]  ( .D(n4423), .CK(CLK), .RN(n6382), .Q(n5127), 
        .QN(n3559) );
  DFFR_X1 \REGISTERS_reg[20][8]  ( .D(n4422), .CK(CLK), .RN(n6382), .Q(n5128), 
        .QN(n2982) );
  DFFR_X1 \REGISTERS_reg[20][7]  ( .D(n4421), .CK(CLK), .RN(n6382), .Q(n5129), 
        .QN(n2981) );
  DFFR_X1 \REGISTERS_reg[20][6]  ( .D(n4420), .CK(CLK), .RN(n6382), .Q(n5130), 
        .QN(n2980) );
  DFFR_X1 \REGISTERS_reg[20][5]  ( .D(n4419), .CK(CLK), .RN(n6382), .Q(n5131), 
        .QN(n2979) );
  DFFR_X1 \REGISTERS_reg[20][4]  ( .D(n4418), .CK(CLK), .RN(n6382), .Q(n5132), 
        .QN(n2978) );
  DFFR_X1 \REGISTERS_reg[20][3]  ( .D(n4417), .CK(CLK), .RN(n6393), .Q(n5133), 
        .QN(n2977) );
  DFFR_X1 \REGISTERS_reg[20][2]  ( .D(n4416), .CK(CLK), .RN(n6393), .Q(n5134), 
        .QN(n2976) );
  DFFR_X1 \REGISTERS_reg[20][1]  ( .D(n4415), .CK(CLK), .RN(n6393), .Q(n5135), 
        .QN(n2975) );
  DFFR_X1 \REGISTERS_reg[20][0]  ( .D(n4414), .CK(CLK), .RN(n6393), .Q(n5136), 
        .QN(n2974) );
  DFFR_X1 \REGISTERS_reg[16][31]  ( .D(n4381), .CK(CLK), .RN(n6453), .Q(n5422), 
        .QN(n3677) );
  DFFR_X1 \REGISTERS_reg[16][30]  ( .D(n4380), .CK(CLK), .RN(n6453), .Q(n5423), 
        .QN(n3676) );
  DFFR_X1 \REGISTERS_reg[16][29]  ( .D(n4379), .CK(CLK), .RN(n6453), .Q(n5424), 
        .QN(n3675) );
  DFFR_X1 \REGISTERS_reg[16][28]  ( .D(n4378), .CK(CLK), .RN(n6453), .Q(n5425), 
        .QN(n3674) );
  DFFR_X1 \REGISTERS_reg[16][27]  ( .D(n4377), .CK(CLK), .RN(n6453), .Q(n5426), 
        .QN(n3673) );
  DFFR_X1 \REGISTERS_reg[16][26]  ( .D(n4376), .CK(CLK), .RN(n6453), .Q(n5427), 
        .QN(n3672) );
  DFFR_X1 \REGISTERS_reg[16][25]  ( .D(n4375), .CK(CLK), .RN(n6453), .Q(n5428), 
        .QN(n3671) );
  DFFR_X1 \REGISTERS_reg[16][24]  ( .D(n4374), .CK(CLK), .RN(n6453), .Q(n5429), 
        .QN(n3670) );
  DFFR_X1 \REGISTERS_reg[16][23]  ( .D(n4373), .CK(CLK), .RN(n6452), .Q(n5430), 
        .QN(n3669) );
  DFFR_X1 \REGISTERS_reg[16][22]  ( .D(n4372), .CK(CLK), .RN(n6452), .Q(n5431), 
        .QN(n3668) );
  DFFR_X1 \REGISTERS_reg[16][21]  ( .D(n4371), .CK(CLK), .RN(n6452), .Q(n5432), 
        .QN(n3667) );
  DFFR_X1 \REGISTERS_reg[16][20]  ( .D(n4370), .CK(CLK), .RN(n6452), .Q(n5433), 
        .QN(n3666) );
  DFFR_X1 \REGISTERS_reg[16][19]  ( .D(n4369), .CK(CLK), .RN(n6464), .Q(n5434), 
        .QN(n3665) );
  DFFR_X1 \REGISTERS_reg[16][18]  ( .D(n4368), .CK(CLK), .RN(n6464), .Q(n5435), 
        .QN(n3664) );
  DFFR_X1 \REGISTERS_reg[16][17]  ( .D(n4367), .CK(CLK), .RN(n6464), .Q(n5436), 
        .QN(n3663) );
  DFFR_X1 \REGISTERS_reg[16][16]  ( .D(n4366), .CK(CLK), .RN(n6464), .Q(n5437), 
        .QN(n3662) );
  DFFR_X1 \REGISTERS_reg[16][15]  ( .D(n4365), .CK(CLK), .RN(n6464), .Q(n5438), 
        .QN(n3661) );
  DFFR_X1 \REGISTERS_reg[16][14]  ( .D(n4364), .CK(CLK), .RN(n6464), .Q(n5439), 
        .QN(n3660) );
  DFFR_X1 \REGISTERS_reg[16][13]  ( .D(n4363), .CK(CLK), .RN(n6464), .Q(n5440), 
        .QN(n3659) );
  DFFR_X1 \REGISTERS_reg[16][12]  ( .D(n4362), .CK(CLK), .RN(n6464), .Q(n5441), 
        .QN(n3658) );
  DFFR_X1 \REGISTERS_reg[16][11]  ( .D(n4361), .CK(CLK), .RN(n6463), .Q(n5442), 
        .QN(n3657) );
  DFFR_X1 \REGISTERS_reg[16][10]  ( .D(n4360), .CK(CLK), .RN(n6463), .Q(n5443), 
        .QN(n3656) );
  DFFR_X1 \REGISTERS_reg[16][9]  ( .D(n4359), .CK(CLK), .RN(n6463), .Q(n5444), 
        .QN(n3655) );
  DFFR_X1 \REGISTERS_reg[16][8]  ( .D(n4358), .CK(CLK), .RN(n6463), .Q(n5445), 
        .QN(n3654) );
  DFFR_X1 \REGISTERS_reg[16][7]  ( .D(n4357), .CK(CLK), .RN(n6463), .Q(n5446), 
        .QN(n3653) );
  DFFR_X1 \REGISTERS_reg[16][6]  ( .D(n4356), .CK(CLK), .RN(n6463), .Q(n5447), 
        .QN(n3652) );
  DFFR_X1 \REGISTERS_reg[16][5]  ( .D(n4355), .CK(CLK), .RN(n6463), .Q(n5448), 
        .QN(n3651) );
  DFFR_X1 \REGISTERS_reg[16][4]  ( .D(n4354), .CK(CLK), .RN(n6463), .Q(n5449), 
        .QN(n3650) );
  DFFR_X1 \REGISTERS_reg[16][3]  ( .D(n4353), .CK(CLK), .RN(n6462), .Q(n5450), 
        .QN(n3649) );
  DFFR_X1 \REGISTERS_reg[16][2]  ( .D(n4352), .CK(CLK), .RN(n6462), .Q(n5451), 
        .QN(n3648) );
  DFFR_X1 \REGISTERS_reg[16][1]  ( .D(n4351), .CK(CLK), .RN(n6462), .Q(n5452), 
        .QN(n3647) );
  DFFR_X1 \REGISTERS_reg[16][0]  ( .D(n4350), .CK(CLK), .RN(n6462), .Q(n5547), 
        .QN(n3646) );
  DFFR_X1 \REGISTERS_reg[13][31]  ( .D(n4253), .CK(CLK), .RN(n6449), .Q(n5873), 
        .QN(n3773) );
  DFFR_X1 \REGISTERS_reg[13][30]  ( .D(n4252), .CK(CLK), .RN(n6449), .Q(n5328), 
        .QN(n3772) );
  DFFR_X1 \REGISTERS_reg[13][29]  ( .D(n4251), .CK(CLK), .RN(n6449), .Q(n5329), 
        .QN(n3771) );
  DFFR_X1 \REGISTERS_reg[13][28]  ( .D(n4250), .CK(CLK), .RN(n6449), .Q(n5330), 
        .QN(n3770) );
  DFFR_X1 \REGISTERS_reg[13][27]  ( .D(n4249), .CK(CLK), .RN(n6449), .Q(n5331), 
        .QN(n3769) );
  DFFR_X1 \REGISTERS_reg[13][26]  ( .D(n4248), .CK(CLK), .RN(n6449), .Q(n5332), 
        .QN(n3768) );
  DFFR_X1 \REGISTERS_reg[13][25]  ( .D(n4247), .CK(CLK), .RN(n6449), .Q(n5333), 
        .QN(n3767) );
  DFFR_X1 \REGISTERS_reg[13][24]  ( .D(n4246), .CK(CLK), .RN(n6449), .Q(n5334), 
        .QN(n3766) );
  DFFR_X1 \REGISTERS_reg[13][23]  ( .D(n4245), .CK(CLK), .RN(n6448), .Q(n5335), 
        .QN(n3765) );
  DFFR_X1 \REGISTERS_reg[13][22]  ( .D(n4244), .CK(CLK), .RN(n6448), .Q(n5336), 
        .QN(n3764) );
  DFFR_X1 \REGISTERS_reg[13][21]  ( .D(n4243), .CK(CLK), .RN(n6448), .Q(n5337), 
        .QN(n3763) );
  DFFR_X1 \REGISTERS_reg[13][20]  ( .D(n4242), .CK(CLK), .RN(n6448), .Q(n5338), 
        .QN(n3762) );
  DFFR_X1 \REGISTERS_reg[13][19]  ( .D(n4241), .CK(CLK), .RN(n6448), .Q(n5339), 
        .QN(n3761) );
  DFFR_X1 \REGISTERS_reg[13][18]  ( .D(n4240), .CK(CLK), .RN(n6448), .Q(n5340), 
        .QN(n3760) );
  DFFR_X1 \REGISTERS_reg[13][17]  ( .D(n4239), .CK(CLK), .RN(n6448), .Q(n5341), 
        .QN(n3759) );
  DFFR_X1 \REGISTERS_reg[13][16]  ( .D(n4238), .CK(CLK), .RN(n6448), .Q(n5342), 
        .QN(n3758) );
  DFFR_X1 \REGISTERS_reg[13][15]  ( .D(n4237), .CK(CLK), .RN(n6448), .Q(n5343), 
        .QN(n3757) );
  DFFR_X1 \REGISTERS_reg[13][14]  ( .D(n4236), .CK(CLK), .RN(n6448), .Q(n5344), 
        .QN(n3756) );
  DFFR_X1 \REGISTERS_reg[13][13]  ( .D(n4235), .CK(CLK), .RN(n6448), .Q(n5345), 
        .QN(n3755) );
  DFFR_X1 \REGISTERS_reg[13][12]  ( .D(n4234), .CK(CLK), .RN(n6448), .Q(n5346), 
        .QN(n3754) );
  DFFR_X1 \REGISTERS_reg[13][11]  ( .D(n4233), .CK(CLK), .RN(n6447), .Q(n5347), 
        .QN(n3753) );
  DFFR_X1 \REGISTERS_reg[13][10]  ( .D(n4232), .CK(CLK), .RN(n6447), .Q(n5348), 
        .QN(n3752) );
  DFFR_X1 \REGISTERS_reg[13][9]  ( .D(n4231), .CK(CLK), .RN(n6447), .Q(n5349), 
        .QN(n3751) );
  DFFR_X1 \REGISTERS_reg[13][8]  ( .D(n4230), .CK(CLK), .RN(n6447), .Q(n5350), 
        .QN(n3750) );
  DFFR_X1 \REGISTERS_reg[13][7]  ( .D(n4229), .CK(CLK), .RN(n6447), .Q(n5351), 
        .QN(n3749) );
  DFFR_X1 \REGISTERS_reg[13][6]  ( .D(n4228), .CK(CLK), .RN(n6447), .Q(n5352), 
        .QN(n3748) );
  DFFR_X1 \REGISTERS_reg[13][5]  ( .D(n4227), .CK(CLK), .RN(n6447), .Q(n5353), 
        .QN(n3747) );
  DFFR_X1 \REGISTERS_reg[13][4]  ( .D(n4226), .CK(CLK), .RN(n6447), .Q(n5354), 
        .QN(n3746) );
  DFFR_X1 \REGISTERS_reg[13][3]  ( .D(n4225), .CK(CLK), .RN(n6446), .Q(n5355), 
        .QN(n3745) );
  DFFR_X1 \REGISTERS_reg[13][2]  ( .D(n4224), .CK(CLK), .RN(n6446), .Q(n5356), 
        .QN(n3744) );
  DFFR_X1 \REGISTERS_reg[13][1]  ( .D(n4223), .CK(CLK), .RN(n6446), .Q(n5357), 
        .QN(n3743) );
  DFFR_X1 \REGISTERS_reg[13][0]  ( .D(n4222), .CK(CLK), .RN(n6446), .Q(n5874), 
        .QN(n3742) );
  DFFR_X1 \REGISTERS_reg[9][31]  ( .D(n4189), .CK(CLK), .RN(n6436), .Q(n5841), 
        .QN(n3901) );
  DFFR_X1 \REGISTERS_reg[9][30]  ( .D(n4188), .CK(CLK), .RN(n6436), .Q(n5842), 
        .QN(n3900) );
  DFFR_X1 \REGISTERS_reg[9][29]  ( .D(n4187), .CK(CLK), .RN(n6436), .Q(n5843), 
        .QN(n3899) );
  DFFR_X1 \REGISTERS_reg[9][28]  ( .D(n4186), .CK(CLK), .RN(n6436), .Q(n5844), 
        .QN(n3898) );
  DFFR_X1 \REGISTERS_reg[9][27]  ( .D(n4185), .CK(CLK), .RN(n6435), .Q(n5845), 
        .QN(n3897) );
  DFFR_X1 \REGISTERS_reg[9][26]  ( .D(n4184), .CK(CLK), .RN(n6435), .Q(n5846), 
        .QN(n3896) );
  DFFR_X1 \REGISTERS_reg[9][25]  ( .D(n4183), .CK(CLK), .RN(n6435), .Q(n5847), 
        .QN(n3895) );
  DFFR_X1 \REGISTERS_reg[9][24]  ( .D(n4182), .CK(CLK), .RN(n6435), .Q(n5848), 
        .QN(n3894) );
  DFFR_X1 \REGISTERS_reg[9][23]  ( .D(n4181), .CK(CLK), .RN(n6435), .Q(n5849), 
        .QN(n3893) );
  DFFR_X1 \REGISTERS_reg[9][22]  ( .D(n4180), .CK(CLK), .RN(n6435), .Q(n5850), 
        .QN(n3892) );
  DFFR_X1 \REGISTERS_reg[9][21]  ( .D(n4179), .CK(CLK), .RN(n6435), .Q(n5851), 
        .QN(n3891) );
  DFFR_X1 \REGISTERS_reg[9][20]  ( .D(n4178), .CK(CLK), .RN(n6435), .Q(n5852), 
        .QN(n3890) );
  DFFR_X1 \REGISTERS_reg[9][19]  ( .D(n4177), .CK(CLK), .RN(n6435), .Q(n5853), 
        .QN(n3889) );
  DFFR_X1 \REGISTERS_reg[9][18]  ( .D(n4176), .CK(CLK), .RN(n6435), .Q(n5854), 
        .QN(n3888) );
  DFFR_X1 \REGISTERS_reg[9][17]  ( .D(n4175), .CK(CLK), .RN(n6435), .Q(n5855), 
        .QN(n3887) );
  DFFR_X1 \REGISTERS_reg[9][16]  ( .D(n4174), .CK(CLK), .RN(n6435), .Q(n5856), 
        .QN(n3886) );
  DFFR_X1 \REGISTERS_reg[9][15]  ( .D(n4173), .CK(CLK), .RN(n6434), .Q(n5857), 
        .QN(n3885) );
  DFFR_X1 \REGISTERS_reg[9][14]  ( .D(n4172), .CK(CLK), .RN(n6434), .Q(n5858), 
        .QN(n3884) );
  DFFR_X1 \REGISTERS_reg[9][13]  ( .D(n4171), .CK(CLK), .RN(n6434), .Q(n5859), 
        .QN(n3883) );
  DFFR_X1 \REGISTERS_reg[9][12]  ( .D(n4170), .CK(CLK), .RN(n6434), .Q(n5860), 
        .QN(n3882) );
  DFFR_X1 \REGISTERS_reg[9][11]  ( .D(n4169), .CK(CLK), .RN(n6446), .Q(n5861), 
        .QN(n3881) );
  DFFR_X1 \REGISTERS_reg[9][10]  ( .D(n4168), .CK(CLK), .RN(n6446), .Q(n5862), 
        .QN(n3880) );
  DFFR_X1 \REGISTERS_reg[9][9]  ( .D(n4167), .CK(CLK), .RN(n6446), .Q(n5863), 
        .QN(n3879) );
  DFFR_X1 \REGISTERS_reg[9][8]  ( .D(n4166), .CK(CLK), .RN(n6446), .Q(n5864), 
        .QN(n3878) );
  DFFR_X1 \REGISTERS_reg[9][7]  ( .D(n4165), .CK(CLK), .RN(n6446), .Q(n5865), 
        .QN(n3877) );
  DFFR_X1 \REGISTERS_reg[9][6]  ( .D(n4164), .CK(CLK), .RN(n6446), .Q(n5866), 
        .QN(n3876) );
  DFFR_X1 \REGISTERS_reg[9][5]  ( .D(n4163), .CK(CLK), .RN(n6446), .Q(n5867), 
        .QN(n3875) );
  DFFR_X1 \REGISTERS_reg[9][4]  ( .D(n4162), .CK(CLK), .RN(n6446), .Q(n5868), 
        .QN(n3874) );
  DFFR_X1 \REGISTERS_reg[9][3]  ( .D(n4161), .CK(CLK), .RN(n6445), .Q(n5869), 
        .QN(n3873) );
  DFFR_X1 \REGISTERS_reg[9][2]  ( .D(n4160), .CK(CLK), .RN(n6445), .Q(n5870), 
        .QN(n3872) );
  DFFR_X1 \REGISTERS_reg[9][1]  ( .D(n4159), .CK(CLK), .RN(n6445), .Q(n5871), 
        .QN(n3871) );
  DFFR_X1 \REGISTERS_reg[9][0]  ( .D(n4158), .CK(CLK), .RN(n6445), .Q(n5872), 
        .QN(n3870) );
  DFFR_X1 \REGISTERS_reg[1][31]  ( .D(n4285), .CK(CLK), .RN(n6422), .Q(n5169), 
        .QN(n4094) );
  DFFR_X1 \REGISTERS_reg[1][30]  ( .D(n4284), .CK(CLK), .RN(n6422), .Q(n5203), 
        .QN(n4095) );
  DFFR_X1 \REGISTERS_reg[1][29]  ( .D(n4283), .CK(CLK), .RN(n6422), .Q(n5204), 
        .QN(n4096) );
  DFFR_X1 \REGISTERS_reg[1][28]  ( .D(n4282), .CK(CLK), .RN(n6422), .Q(n5205), 
        .QN(n4097) );
  DFFR_X1 \REGISTERS_reg[1][27]  ( .D(n4281), .CK(CLK), .RN(n6422), .Q(n5206), 
        .QN(n4098) );
  DFFR_X1 \REGISTERS_reg[1][26]  ( .D(n4280), .CK(CLK), .RN(n6422), .Q(n5207), 
        .QN(n4099) );
  DFFR_X1 \REGISTERS_reg[1][25]  ( .D(n4279), .CK(CLK), .RN(n6422), .Q(n5208), 
        .QN(n4100) );
  DFFR_X1 \REGISTERS_reg[1][24]  ( .D(n4278), .CK(CLK), .RN(n6422), .Q(n5209), 
        .QN(n4101) );
  DFFR_X1 \REGISTERS_reg[1][23]  ( .D(n4277), .CK(CLK), .RN(n6421), .Q(n5210), 
        .QN(n4102) );
  DFFR_X1 \REGISTERS_reg[1][22]  ( .D(n4276), .CK(CLK), .RN(n6421), .Q(n5211), 
        .QN(n4103) );
  DFFR_X1 \REGISTERS_reg[1][21]  ( .D(n4275), .CK(CLK), .RN(n6421), .Q(n5212), 
        .QN(n4104) );
  DFFR_X1 \REGISTERS_reg[1][20]  ( .D(n4274), .CK(CLK), .RN(n6421), .Q(n5213), 
        .QN(n4105) );
  DFFR_X1 \REGISTERS_reg[1][19]  ( .D(n4273), .CK(CLK), .RN(n6421), .Q(n5214), 
        .QN(n4106) );
  DFFR_X1 \REGISTERS_reg[1][18]  ( .D(n4272), .CK(CLK), .RN(n6421), .Q(n5215), 
        .QN(n4107) );
  DFFR_X1 \REGISTERS_reg[1][17]  ( .D(n4271), .CK(CLK), .RN(n6421), .Q(n5216), 
        .QN(n4108) );
  DFFR_X1 \REGISTERS_reg[1][16]  ( .D(n4270), .CK(CLK), .RN(n6421), .Q(n5217), 
        .QN(n4109) );
  DFFR_X1 \REGISTERS_reg[1][15]  ( .D(n4269), .CK(CLK), .RN(n6421), .Q(n5218), 
        .QN(n4110) );
  DFFR_X1 \REGISTERS_reg[1][14]  ( .D(n4268), .CK(CLK), .RN(n6421), .Q(n5219), 
        .QN(n4111) );
  DFFR_X1 \REGISTERS_reg[1][13]  ( .D(n4267), .CK(CLK), .RN(n6421), .Q(n5220), 
        .QN(n4112) );
  DFFR_X1 \REGISTERS_reg[1][12]  ( .D(n4266), .CK(CLK), .RN(n6421), .Q(n5221), 
        .QN(n4113) );
  DFFR_X1 \REGISTERS_reg[1][11]  ( .D(n4265), .CK(CLK), .RN(n6420), .Q(n5222), 
        .QN(n4114) );
  DFFR_X1 \REGISTERS_reg[1][10]  ( .D(n4264), .CK(CLK), .RN(n6420), .Q(n5223), 
        .QN(n4115) );
  DFFR_X1 \REGISTERS_reg[1][9]  ( .D(n4263), .CK(CLK), .RN(n6420), .Q(n5224), 
        .QN(n4116) );
  DFFR_X1 \REGISTERS_reg[1][8]  ( .D(n4262), .CK(CLK), .RN(n6420), .Q(n5225), 
        .QN(n4117) );
  DFFR_X1 \REGISTERS_reg[1][7]  ( .D(n4261), .CK(CLK), .RN(n6420), .Q(n5226), 
        .QN(n4118) );
  DFFR_X1 \REGISTERS_reg[1][6]  ( .D(n4260), .CK(CLK), .RN(n6420), .Q(n5227), 
        .QN(n4119) );
  DFFR_X1 \REGISTERS_reg[1][5]  ( .D(n4259), .CK(CLK), .RN(n6420), .Q(n5228), 
        .QN(n4120) );
  DFFR_X1 \REGISTERS_reg[1][4]  ( .D(n4258), .CK(CLK), .RN(n6420), .Q(n5229), 
        .QN(n4121) );
  DFFR_X1 \REGISTERS_reg[1][3]  ( .D(n4257), .CK(CLK), .RN(n6419), .Q(n5230), 
        .QN(n4122) );
  DFFR_X1 \REGISTERS_reg[1][2]  ( .D(n4256), .CK(CLK), .RN(n6419), .Q(n5231), 
        .QN(n4123) );
  DFFR_X1 \REGISTERS_reg[1][1]  ( .D(n4255), .CK(CLK), .RN(n6419), .Q(n5232), 
        .QN(n4124) );
  DFFR_X1 \REGISTERS_reg[1][0]  ( .D(n4254), .CK(CLK), .RN(n6419), .Q(n5170), 
        .QN(n4125) );
  DFFR_X1 \REGISTERS_reg[23][31]  ( .D(n3206), .CK(CLK), .RN(RST), .Q(n4750), 
        .QN(n7521) );
  DFFR_X1 \REGISTERS_reg[23][30]  ( .D(n7683), .CK(CLK), .RN(n6389), .Q(n4748), 
        .QN(n7498) );
  DFFR_X1 \REGISTERS_reg[23][29]  ( .D(n7684), .CK(CLK), .RN(n6388), .Q(n4742), 
        .QN(n7479) );
  DFFR_X1 \REGISTERS_reg[23][28]  ( .D(n7685), .CK(CLK), .RN(n6388), .Q(n4744), 
        .QN(n7460) );
  DFFR_X1 \REGISTERS_reg[23][27]  ( .D(n7686), .CK(CLK), .RN(n6400), .Q(n4746), 
        .QN(n7441) );
  DFFR_X1 \REGISTERS_reg[23][26]  ( .D(n7687), .CK(CLK), .RN(n6399), .Q(n4736), 
        .QN(n7422) );
  DFFR_X1 \REGISTERS_reg[23][25]  ( .D(n7688), .CK(CLK), .RN(n6399), .Q(n4738), 
        .QN(n7403) );
  DFFR_X1 \REGISTERS_reg[23][24]  ( .D(n7689), .CK(CLK), .RN(n6399), .Q(n4740), 
        .QN(n7384) );
  DFFR_X1 \REGISTERS_reg[23][23]  ( .D(n7690), .CK(CLK), .RN(n6399), .Q(n4730), 
        .QN(n7365) );
  DFFR_X1 \REGISTERS_reg[23][22]  ( .D(n7691), .CK(CLK), .RN(n6399), .Q(n4732), 
        .QN(n7346) );
  DFFR_X1 \REGISTERS_reg[23][21]  ( .D(n7692), .CK(CLK), .RN(n6399), .Q(n4734), 
        .QN(n7327) );
  DFFR_X1 \REGISTERS_reg[23][20]  ( .D(n7693), .CK(CLK), .RN(n6399), .Q(n4724), 
        .QN(n7308) );
  DFFR_X1 \REGISTERS_reg[23][19]  ( .D(n7694), .CK(CLK), .RN(n6399), .Q(n4726), 
        .QN(n7289) );
  DFFR_X1 \REGISTERS_reg[23][18]  ( .D(n7695), .CK(CLK), .RN(n6399), .Q(n4728), 
        .QN(n7270) );
  DFFR_X1 \REGISTERS_reg[23][17]  ( .D(n7696), .CK(CLK), .RN(n6399), .Q(n4718), 
        .QN(n7251) );
  DFFR_X1 \REGISTERS_reg[23][16]  ( .D(n7697), .CK(CLK), .RN(n6399), .Q(n4720), 
        .QN(n7232) );
  DFFR_X1 \REGISTERS_reg[23][15]  ( .D(n7698), .CK(CLK), .RN(n6399), .Q(n4722), 
        .QN(n7213) );
  DFFR_X1 \REGISTERS_reg[23][14]  ( .D(n7699), .CK(CLK), .RN(n6398), .Q(n4712), 
        .QN(n7194) );
  DFFR_X1 \REGISTERS_reg[23][13]  ( .D(n7700), .CK(CLK), .RN(n6398), .Q(n4714), 
        .QN(n7175) );
  DFFR_X1 \REGISTERS_reg[23][12]  ( .D(n7701), .CK(CLK), .RN(n6398), .Q(n4716), 
        .QN(n7156) );
  DFFR_X1 \REGISTERS_reg[23][11]  ( .D(n7702), .CK(CLK), .RN(n6398), .Q(n4706), 
        .QN(n7137) );
  DFFR_X1 \REGISTERS_reg[23][10]  ( .D(n7703), .CK(CLK), .RN(n6398), .Q(n4708), 
        .QN(n7118) );
  DFFR_X1 \REGISTERS_reg[23][9]  ( .D(n7704), .CK(CLK), .RN(n6398), .Q(n4710), 
        .QN(n7099) );
  DFFR_X1 \REGISTERS_reg[23][8]  ( .D(n7705), .CK(CLK), .RN(n6398), .Q(n4700), 
        .QN(n7080) );
  DFFR_X1 \REGISTERS_reg[23][7]  ( .D(n7706), .CK(CLK), .RN(n6398), .Q(n4702), 
        .QN(n7061) );
  DFFR_X1 \REGISTERS_reg[23][6]  ( .D(n7707), .CK(CLK), .RN(n6398), .Q(n4704), 
        .QN(n7042) );
  DFFR_X1 \REGISTERS_reg[23][5]  ( .D(n7708), .CK(CLK), .RN(n6398), .Q(n4696), 
        .QN(n7023) );
  DFFR_X1 \REGISTERS_reg[23][4]  ( .D(n7709), .CK(CLK), .RN(n6398), .Q(n4698), 
        .QN(n7004) );
  DFFR_X1 \REGISTERS_reg[22][31]  ( .D(n3238), .CK(CLK), .RN(n6391), .Q(n2941), 
        .QN(n5941) );
  DFFR_X1 \REGISTERS_reg[22][30]  ( .D(n3237), .CK(CLK), .RN(n6391), .Q(n2940), 
        .QN(n5942) );
  DFFR_X1 \REGISTERS_reg[22][29]  ( .D(n3236), .CK(CLK), .RN(n6390), .Q(n2939), 
        .QN(n5943) );
  DFFR_X1 \REGISTERS_reg[22][28]  ( .D(n3235), .CK(CLK), .RN(n6390), .Q(n2938), 
        .QN(n5944) );
  DFFR_X1 \REGISTERS_reg[22][27]  ( .D(n3234), .CK(CLK), .RN(n6390), .Q(n2937), 
        .QN(n5945) );
  DFFR_X1 \REGISTERS_reg[22][26]  ( .D(n3233), .CK(CLK), .RN(n6390), .Q(n2936), 
        .QN(n5946) );
  DFFR_X1 \REGISTERS_reg[22][25]  ( .D(n3232), .CK(CLK), .RN(n6390), .Q(n2935), 
        .QN(n5947) );
  DFFR_X1 \REGISTERS_reg[22][24]  ( .D(n3231), .CK(CLK), .RN(n6390), .Q(n2934), 
        .QN(n5948) );
  DFFR_X1 \REGISTERS_reg[22][23]  ( .D(n3230), .CK(CLK), .RN(n6390), .Q(n2933), 
        .QN(n5949) );
  DFFR_X1 \REGISTERS_reg[22][22]  ( .D(n3229), .CK(CLK), .RN(n6390), .Q(n2932), 
        .QN(n5950) );
  DFFR_X1 \REGISTERS_reg[22][21]  ( .D(n3228), .CK(CLK), .RN(n6390), .Q(n2931), 
        .QN(n5951) );
  DFFR_X1 \REGISTERS_reg[22][20]  ( .D(n3227), .CK(CLK), .RN(n6390), .Q(n2930), 
        .QN(n5952) );
  DFFR_X1 \REGISTERS_reg[22][19]  ( .D(n3226), .CK(CLK), .RN(n6390), .Q(n2929), 
        .QN(n5953) );
  DFFR_X1 \REGISTERS_reg[22][18]  ( .D(n3225), .CK(CLK), .RN(n6390), .Q(n2928), 
        .QN(n5954) );
  DFFR_X1 \REGISTERS_reg[22][17]  ( .D(n3224), .CK(CLK), .RN(n6389), .Q(n2927), 
        .QN(n5955) );
  DFFR_X1 \REGISTERS_reg[22][16]  ( .D(n3223), .CK(CLK), .RN(n6389), .Q(n2926), 
        .QN(n5956) );
  DFFR_X1 \REGISTERS_reg[22][15]  ( .D(n3222), .CK(CLK), .RN(n6389), .Q(n2925), 
        .QN(n5957) );
  DFFR_X1 \REGISTERS_reg[22][14]  ( .D(n3221), .CK(CLK), .RN(n6389), .Q(n2924), 
        .QN(n5958) );
  DFFR_X1 \REGISTERS_reg[22][13]  ( .D(n3220), .CK(CLK), .RN(n6389), .Q(n2923), 
        .QN(n5959) );
  DFFR_X1 \REGISTERS_reg[22][12]  ( .D(n3219), .CK(CLK), .RN(n6389), .Q(n2922), 
        .QN(n5960) );
  DFFR_X1 \REGISTERS_reg[22][11]  ( .D(n3218), .CK(CLK), .RN(n6389), .Q(n2921), 
        .QN(n5961) );
  DFFR_X1 \REGISTERS_reg[22][10]  ( .D(n3217), .CK(CLK), .RN(n6389), .Q(n2920), 
        .QN(n5962) );
  DFFR_X1 \REGISTERS_reg[22][9]  ( .D(n3216), .CK(CLK), .RN(n6389), .Q(n2919), 
        .QN(n5963) );
  DFFR_X1 \REGISTERS_reg[22][8]  ( .D(n3215), .CK(CLK), .RN(n6389), .Q(n2918), 
        .QN(n5964) );
  DFFR_X1 \REGISTERS_reg[22][7]  ( .D(n3214), .CK(CLK), .RN(n6388), .Q(n2917), 
        .QN(n5965) );
  DFFR_X1 \REGISTERS_reg[22][6]  ( .D(n3213), .CK(CLK), .RN(n6388), .Q(n2916), 
        .QN(n5966) );
  DFFR_X1 \REGISTERS_reg[22][5]  ( .D(n3212), .CK(CLK), .RN(n6388), .Q(n2915), 
        .QN(n5967) );
  DFFR_X1 \REGISTERS_reg[22][4]  ( .D(n3211), .CK(CLK), .RN(n6388), .Q(n2914), 
        .QN(n5968) );
  DFFR_X1 \REGISTERS_reg[22][3]  ( .D(n3210), .CK(CLK), .RN(n6388), .Q(n2913), 
        .QN(n5969) );
  DFFR_X1 \REGISTERS_reg[22][2]  ( .D(n3209), .CK(CLK), .RN(n6388), .Q(n2912), 
        .QN(n5970) );
  DFFR_X1 \REGISTERS_reg[22][1]  ( .D(n3208), .CK(CLK), .RN(n6388), .Q(n2911), 
        .QN(n5971) );
  DFFR_X1 \REGISTERS_reg[22][0]  ( .D(n3207), .CK(CLK), .RN(n6388), .Q(n2910), 
        .QN(n5972) );
  DFFR_X1 \REGISTERS_reg[7][31]  ( .D(n7710), .CK(CLK), .RN(n6429), .Q(n4814), 
        .QN(n7535) );
  DFFR_X1 \REGISTERS_reg[7][30]  ( .D(n7711), .CK(CLK), .RN(n6429), .Q(n4780), 
        .QN(n7505) );
  DFFR_X1 \REGISTERS_reg[7][29]  ( .D(n7712), .CK(CLK), .RN(n6429), .Q(n4776), 
        .QN(n7486) );
  DFFR_X1 \REGISTERS_reg[7][28]  ( .D(n7713), .CK(CLK), .RN(n6429), .Q(n4778), 
        .QN(n7467) );
  DFFR_X1 \REGISTERS_reg[7][27]  ( .D(n7714), .CK(CLK), .RN(n6429), .Q(n4754), 
        .QN(n7448) );
  DFFR_X1 \REGISTERS_reg[7][26]  ( .D(n7715), .CK(CLK), .RN(n6429), .Q(n4772), 
        .QN(n7429) );
  DFFR_X1 \REGISTERS_reg[7][25]  ( .D(n7716), .CK(CLK), .RN(n6429), .Q(n4774), 
        .QN(n7410) );
  DFFR_X1 \REGISTERS_reg[7][24]  ( .D(n7717), .CK(CLK), .RN(n6429), .Q(n4766), 
        .QN(n7391) );
  DFFR_X1 \REGISTERS_reg[7][23]  ( .D(n7718), .CK(CLK), .RN(n6428), .Q(n4770), 
        .QN(n7372) );
  DFFR_X1 \REGISTERS_reg[7][22]  ( .D(n7719), .CK(CLK), .RN(n6428), .Q(n4764), 
        .QN(n7353) );
  DFFR_X1 \REGISTERS_reg[7][21]  ( .D(n7720), .CK(CLK), .RN(n6428), .Q(n4760), 
        .QN(n7334) );
  DFFR_X1 \REGISTERS_reg[7][20]  ( .D(n7721), .CK(CLK), .RN(n6428), .Q(n4768), 
        .QN(n7315) );
  DFFR_X1 \REGISTERS_reg[7][19]  ( .D(n7722), .CK(CLK), .RN(n6440), .Q(n4758), 
        .QN(n7296) );
  DFFR_X1 \REGISTERS_reg[7][18]  ( .D(n7723), .CK(CLK), .RN(n6440), .Q(n4756), 
        .QN(n7277) );
  DFFR_X1 \REGISTERS_reg[7][17]  ( .D(n7724), .CK(CLK), .RN(n6440), .Q(n4762), 
        .QN(n7258) );
  DFFR_X1 \REGISTERS_reg[7][16]  ( .D(n7725), .CK(CLK), .RN(n6440), .Q(n4752), 
        .QN(n7239) );
  DFFR_X1 \REGISTERS_reg[7][15]  ( .D(n7726), .CK(CLK), .RN(n6440), .Q(n4782), 
        .QN(n7220) );
  DFFR_X1 \REGISTERS_reg[7][14]  ( .D(n7727), .CK(CLK), .RN(n6440), .Q(n4784), 
        .QN(n7201) );
  DFFR_X1 \REGISTERS_reg[7][13]  ( .D(n7728), .CK(CLK), .RN(n6440), .Q(n4786), 
        .QN(n7182) );
  DFFR_X1 \REGISTERS_reg[7][12]  ( .D(n7729), .CK(CLK), .RN(n6440), .Q(n4788), 
        .QN(n7163) );
  DFFR_X1 \REGISTERS_reg[7][11]  ( .D(n7730), .CK(CLK), .RN(n6439), .Q(n4790), 
        .QN(n7144) );
  DFFR_X1 \REGISTERS_reg[7][10]  ( .D(n7731), .CK(CLK), .RN(n6439), .Q(n4792), 
        .QN(n7125) );
  DFFR_X1 \REGISTERS_reg[7][9]  ( .D(n7732), .CK(CLK), .RN(n6439), .Q(n4794), 
        .QN(n7106) );
  DFFR_X1 \REGISTERS_reg[7][8]  ( .D(n7733), .CK(CLK), .RN(n6439), .Q(n4796), 
        .QN(n7087) );
  DFFR_X1 \REGISTERS_reg[7][7]  ( .D(n7734), .CK(CLK), .RN(n6439), .Q(n4798), 
        .QN(n7068) );
  DFFR_X1 \REGISTERS_reg[7][6]  ( .D(n7735), .CK(CLK), .RN(n6439), .Q(n4800), 
        .QN(n7049) );
  DFFR_X1 \REGISTERS_reg[7][5]  ( .D(n7736), .CK(CLK), .RN(n6439), .Q(n4802), 
        .QN(n7030) );
  DFFR_X1 \REGISTERS_reg[7][4]  ( .D(n7737), .CK(CLK), .RN(n6439), .Q(n4804), 
        .QN(n7011) );
  DFFR_X1 \REGISTERS_reg[7][3]  ( .D(n7738), .CK(CLK), .RN(n6439), .Q(n4806), 
        .QN(n6992) );
  DFFR_X1 \REGISTERS_reg[7][2]  ( .D(n7739), .CK(CLK), .RN(n6439), .Q(n4808), 
        .QN(n6974) );
  DFFR_X1 \REGISTERS_reg[7][1]  ( .D(n7740), .CK(CLK), .RN(n6439), .Q(n4810), 
        .QN(n6956) );
  DFFR_X1 \REGISTERS_reg[7][0]  ( .D(n7741), .CK(CLK), .RN(n6439), .Q(n4812), 
        .QN(n6937) );
  DFFR_X1 \REGISTERS_reg[6][31]  ( .D(n7742), .CK(CLK), .RN(n6432), .QN(n7534)
         );
  DFFR_X1 \REGISTERS_reg[6][30]  ( .D(n7743), .CK(CLK), .RN(n6432), .QN(n7504)
         );
  DFFR_X1 \REGISTERS_reg[6][29]  ( .D(n7744), .CK(CLK), .RN(n6432), .QN(n7485)
         );
  DFFR_X1 \REGISTERS_reg[6][28]  ( .D(n7745), .CK(CLK), .RN(n6432), .QN(n7466)
         );
  DFFR_X1 \REGISTERS_reg[6][27]  ( .D(n7746), .CK(CLK), .RN(n6432), .QN(n7447)
         );
  DFFR_X1 \REGISTERS_reg[6][26]  ( .D(n7747), .CK(CLK), .RN(n6432), .QN(n7428)
         );
  DFFR_X1 \REGISTERS_reg[6][25]  ( .D(n7748), .CK(CLK), .RN(n6432), .QN(n7409)
         );
  DFFR_X1 \REGISTERS_reg[6][24]  ( .D(n7749), .CK(CLK), .RN(n6432), .QN(n7390)
         );
  DFFR_X1 \REGISTERS_reg[6][23]  ( .D(n7750), .CK(CLK), .RN(n6431), .QN(n7371)
         );
  DFFR_X1 \REGISTERS_reg[6][22]  ( .D(n7751), .CK(CLK), .RN(n6431), .QN(n7352)
         );
  DFFR_X1 \REGISTERS_reg[6][21]  ( .D(n7752), .CK(CLK), .RN(n6431), .QN(n7333)
         );
  DFFR_X1 \REGISTERS_reg[6][20]  ( .D(n7753), .CK(CLK), .RN(n6431), .QN(n7314)
         );
  DFFR_X1 \REGISTERS_reg[6][19]  ( .D(n7754), .CK(CLK), .RN(n6431), .QN(n7295)
         );
  DFFR_X1 \REGISTERS_reg[6][18]  ( .D(n7755), .CK(CLK), .RN(n6431), .QN(n7276)
         );
  DFFR_X1 \REGISTERS_reg[6][17]  ( .D(n7756), .CK(CLK), .RN(n6431), .QN(n7257)
         );
  DFFR_X1 \REGISTERS_reg[6][16]  ( .D(n7757), .CK(CLK), .RN(n6431), .QN(n7238)
         );
  DFFR_X1 \REGISTERS_reg[6][15]  ( .D(n7758), .CK(CLK), .RN(n6430), .QN(n7219)
         );
  DFFR_X1 \REGISTERS_reg[6][14]  ( .D(n7759), .CK(CLK), .RN(n6430), .QN(n7200)
         );
  DFFR_X1 \REGISTERS_reg[6][13]  ( .D(n7760), .CK(CLK), .RN(n6430), .QN(n7181)
         );
  DFFR_X1 \REGISTERS_reg[6][12]  ( .D(n7761), .CK(CLK), .RN(n6430), .QN(n7162)
         );
  DFFR_X1 \REGISTERS_reg[6][11]  ( .D(n7762), .CK(CLK), .RN(n6430), .QN(n7143)
         );
  DFFR_X1 \REGISTERS_reg[6][10]  ( .D(n7763), .CK(CLK), .RN(n6430), .QN(n7124)
         );
  DFFR_X1 \REGISTERS_reg[6][9]  ( .D(n7764), .CK(CLK), .RN(n6430), .QN(n7105)
         );
  DFFR_X1 \REGISTERS_reg[6][8]  ( .D(n7765), .CK(CLK), .RN(n6430), .QN(n7086)
         );
  DFFR_X1 \REGISTERS_reg[6][7]  ( .D(n7766), .CK(CLK), .RN(n6430), .QN(n7067)
         );
  DFFR_X1 \REGISTERS_reg[6][6]  ( .D(n7767), .CK(CLK), .RN(n6430), .QN(n7048)
         );
  DFFR_X1 \REGISTERS_reg[6][5]  ( .D(n7768), .CK(CLK), .RN(n6430), .QN(n7029)
         );
  DFFR_X1 \REGISTERS_reg[6][4]  ( .D(n7769), .CK(CLK), .RN(n6430), .QN(n7010)
         );
  DFFR_X1 \REGISTERS_reg[6][3]  ( .D(n7770), .CK(CLK), .RN(n6429), .QN(n6991)
         );
  DFFR_X1 \REGISTERS_reg[6][2]  ( .D(n7771), .CK(CLK), .RN(n6429), .QN(n6973)
         );
  DFFR_X1 \REGISTERS_reg[6][1]  ( .D(n7772), .CK(CLK), .RN(n6429), .QN(n6955)
         );
  DFFR_X1 \REGISTERS_reg[6][0]  ( .D(n7773), .CK(CLK), .RN(n6429), .QN(n6936)
         );
  DFFR_X1 \REGISTERS_reg[3][31]  ( .D(n7774), .CK(CLK), .RN(n6428), .Q(n4061), 
        .QN(n5909) );
  DFFR_X1 \REGISTERS_reg[3][30]  ( .D(n7775), .CK(CLK), .RN(n6428), .Q(n4060), 
        .QN(n5911) );
  DFFR_X1 \REGISTERS_reg[3][29]  ( .D(n7776), .CK(CLK), .RN(n6428), .Q(n4059), 
        .QN(n5912) );
  DFFR_X1 \REGISTERS_reg[3][28]  ( .D(n7777), .CK(CLK), .RN(n6428), .Q(n4058), 
        .QN(n5913) );
  DFFR_X1 \REGISTERS_reg[3][27]  ( .D(n7778), .CK(CLK), .RN(n6428), .Q(n4057), 
        .QN(n5914) );
  AND2_X1 U2 ( .A1(n4662), .A2(ADD_WR[3]), .ZN(n4606) );
  AND2_X1 U3 ( .A1(n4662), .A2(n7590), .ZN(n4607) );
  AND2_X1 U4 ( .A1(n6480), .A2(n7898), .ZN(n4608) );
  AND3_X1 U5 ( .A1(n749), .A2(ADD_WR[3]), .A3(n7589), .ZN(n4609) );
  AND3_X1 U6 ( .A1(ADD_RS1[0]), .A2(ADD_RS1[4]), .A3(n7592), .ZN(n4610) );
  AND2_X1 U7 ( .A1(n4663), .A2(ADD_WR[0]), .ZN(n4611) );
  AND3_X1 U8 ( .A1(ADD_RS1[3]), .A2(ADD_RS1[4]), .A3(n7593), .ZN(n4612) );
  AND2_X1 U9 ( .A1(n6479), .A2(n7900), .ZN(n4613) );
  AND2_X1 U10 ( .A1(n4663), .A2(n6485), .ZN(n4614) );
  AND4_X1 U11 ( .A1(ADD_RS2[3]), .A2(ADD_RS2[4]), .A3(n6237), .A4(n7595), .ZN(
        n4615) );
  AND4_X1 U12 ( .A1(n1999), .A2(n1997), .A3(n6173), .A4(n1998), .ZN(n4616) );
  AND4_X1 U13 ( .A1(ADD_RS2[0]), .A2(ADD_RS2[4]), .A3(n6237), .A4(n7594), .ZN(
        n4617) );
  AND2_X1 U14 ( .A1(n2013), .A2(n6163), .ZN(n4618) );
  AND3_X1 U15 ( .A1(ADD_WR[1]), .A2(n7591), .A3(n6485), .ZN(n4619) );
  AND3_X1 U16 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(n7591), .ZN(n4620) );
  AND2_X1 U17 ( .A1(n6163), .A2(n4613), .ZN(n4621) );
  AND3_X1 U18 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(n6482), .ZN(n4622) );
  AND3_X1 U19 ( .A1(ADD_WR[0]), .A2(n7591), .A3(n6482), .ZN(n4623) );
  AND3_X1 U20 ( .A1(ADD_WR[2]), .A2(n6485), .A3(n6482), .ZN(n4624) );
  AND3_X1 U21 ( .A1(n7591), .A2(n6485), .A3(n6482), .ZN(n4625) );
  AND2_X1 U22 ( .A1(n2012), .A2(n6163), .ZN(n4626) );
  AND3_X1 U23 ( .A1(n1406), .A2(n4608), .A3(n6236), .ZN(n4627) );
  AND3_X1 U24 ( .A1(n1406), .A2(n1413), .A3(n6236), .ZN(n4628) );
  AND3_X1 U25 ( .A1(n1393), .A2(n4608), .A3(n6236), .ZN(n4629) );
  AND2_X1 U26 ( .A1(n1394), .A2(n4617), .ZN(n4630) );
  AND2_X1 U27 ( .A1(n2019), .A2(n4613), .ZN(n4631) );
  AND2_X1 U28 ( .A1(n1419), .A2(n4608), .ZN(n4632) );
  AND2_X1 U29 ( .A1(n2006), .A2(n4621), .ZN(n4633) );
  AND2_X1 U30 ( .A1(n2006), .A2(n4626), .ZN(n4634) );
  AND2_X1 U31 ( .A1(n4609), .A2(n4619), .ZN(n4635) );
  AND2_X1 U32 ( .A1(n4606), .A2(n4614), .ZN(n4636) );
  AND2_X1 U33 ( .A1(n4606), .A2(n4619), .ZN(n4637) );
  AND2_X1 U34 ( .A1(n4606), .A2(n4620), .ZN(n4638) );
  AND2_X1 U35 ( .A1(n4607), .A2(n4620), .ZN(n4639) );
  AND2_X1 U36 ( .A1(n4607), .A2(n4619), .ZN(n4640) );
  AND2_X1 U37 ( .A1(n6489), .A2(n4623), .ZN(n4641) );
  AND2_X1 U38 ( .A1(n6489), .A2(n4622), .ZN(n4642) );
  AND2_X1 U39 ( .A1(n4623), .A2(n4609), .ZN(n4643) );
  AND2_X1 U40 ( .A1(n4622), .A2(n4609), .ZN(n4644) );
  AND2_X1 U41 ( .A1(n4625), .A2(n4609), .ZN(n4645) );
  AND2_X1 U42 ( .A1(n4624), .A2(n4609), .ZN(n4646) );
  AND2_X1 U43 ( .A1(n4611), .A2(n4609), .ZN(n4647) );
  AND2_X1 U44 ( .A1(n4614), .A2(n4609), .ZN(n4648) );
  AND2_X1 U45 ( .A1(n4620), .A2(n4609), .ZN(n4649) );
  AND2_X1 U46 ( .A1(n4625), .A2(n4607), .ZN(n4650) );
  AND2_X1 U47 ( .A1(n4624), .A2(n4607), .ZN(n4651) );
  AND2_X1 U48 ( .A1(n4622), .A2(n4607), .ZN(n4652) );
  AND2_X1 U49 ( .A1(n4623), .A2(n4607), .ZN(n4653) );
  AND2_X1 U50 ( .A1(n4624), .A2(n4606), .ZN(n4654) );
  AND2_X1 U51 ( .A1(n4622), .A2(n4606), .ZN(n4655) );
  AND2_X1 U52 ( .A1(n4623), .A2(n4606), .ZN(n4656) );
  AND2_X1 U53 ( .A1(ENABLE), .A2(n6464), .ZN(n4657) );
  AND2_X1 U54 ( .A1(n4624), .A2(n6489), .ZN(n4658) );
  AND2_X1 U55 ( .A1(n4621), .A2(n4610), .ZN(n4659) );
  AND2_X1 U56 ( .A1(RD1), .A2(n4657), .ZN(n4660) );
  AND2_X1 U57 ( .A1(n1994), .A2(n6163), .ZN(n4661) );
  AND2_X1 U58 ( .A1(n749), .A2(ADD_WR[4]), .ZN(n4662) );
  AND2_X1 U59 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .ZN(n4663) );
  INV_X1 U60 ( .A(n2877), .ZN(n4664) );
  INV_X1 U61 ( .A(n2876), .ZN(n4665) );
  INV_X1 U62 ( .A(n2875), .ZN(n4666) );
  INV_X1 U63 ( .A(n2874), .ZN(n4667) );
  INV_X1 U64 ( .A(n2873), .ZN(n4668) );
  INV_X1 U65 ( .A(n2872), .ZN(n4669) );
  INV_X1 U66 ( .A(n2871), .ZN(n4670) );
  INV_X1 U67 ( .A(n2870), .ZN(n4671) );
  INV_X1 U68 ( .A(n2869), .ZN(n4672) );
  INV_X1 U69 ( .A(n2868), .ZN(n4673) );
  INV_X1 U70 ( .A(n2867), .ZN(n4674) );
  INV_X1 U71 ( .A(n2866), .ZN(n4675) );
  INV_X1 U72 ( .A(n2865), .ZN(n4676) );
  INV_X1 U73 ( .A(n2864), .ZN(n4677) );
  INV_X1 U74 ( .A(n2863), .ZN(n4678) );
  INV_X1 U75 ( .A(n2862), .ZN(n4679) );
  INV_X1 U76 ( .A(n2861), .ZN(n4680) );
  INV_X1 U77 ( .A(n2860), .ZN(n4681) );
  INV_X1 U78 ( .A(n2859), .ZN(n4682) );
  INV_X1 U79 ( .A(n2858), .ZN(n4683) );
  INV_X1 U80 ( .A(n2857), .ZN(n4684) );
  INV_X1 U81 ( .A(n2856), .ZN(n4685) );
  INV_X1 U82 ( .A(n2855), .ZN(n4686) );
  INV_X1 U83 ( .A(n2854), .ZN(n4687) );
  INV_X1 U84 ( .A(n2853), .ZN(n4688) );
  INV_X1 U85 ( .A(n2852), .ZN(n4689) );
  INV_X1 U86 ( .A(n2851), .ZN(n4690) );
  INV_X1 U87 ( .A(n2850), .ZN(n4691) );
  INV_X1 U88 ( .A(n998), .ZN(n4692) );
  INV_X1 U89 ( .A(n982), .ZN(n4693) );
  INV_X1 U90 ( .A(n966), .ZN(n4694) );
  INV_X1 U91 ( .A(n950), .ZN(n4695) );
  INV_X1 U92 ( .A(n4696), .ZN(n4697) );
  INV_X1 U93 ( .A(n4698), .ZN(n4699) );
  INV_X1 U94 ( .A(n4700), .ZN(n4701) );
  INV_X1 U95 ( .A(n4702), .ZN(n4703) );
  INV_X1 U96 ( .A(n4704), .ZN(n4705) );
  INV_X1 U97 ( .A(n4706), .ZN(n4707) );
  INV_X1 U98 ( .A(n4708), .ZN(n4709) );
  INV_X1 U99 ( .A(n4710), .ZN(n4711) );
  INV_X1 U100 ( .A(n4712), .ZN(n4713) );
  INV_X1 U101 ( .A(n4714), .ZN(n4715) );
  INV_X1 U102 ( .A(n4716), .ZN(n4717) );
  INV_X1 U103 ( .A(n4718), .ZN(n4719) );
  INV_X1 U104 ( .A(n4720), .ZN(n4721) );
  INV_X1 U105 ( .A(n4722), .ZN(n4723) );
  INV_X1 U106 ( .A(n4724), .ZN(n4725) );
  INV_X1 U107 ( .A(n4726), .ZN(n4727) );
  INV_X1 U108 ( .A(n4728), .ZN(n4729) );
  INV_X1 U109 ( .A(n4730), .ZN(n4731) );
  INV_X1 U110 ( .A(n4732), .ZN(n4733) );
  INV_X1 U111 ( .A(n4734), .ZN(n4735) );
  INV_X1 U112 ( .A(n4736), .ZN(n4737) );
  INV_X1 U113 ( .A(n4738), .ZN(n4739) );
  INV_X1 U114 ( .A(n4740), .ZN(n4741) );
  INV_X1 U115 ( .A(n4742), .ZN(n4743) );
  INV_X1 U116 ( .A(n4744), .ZN(n4745) );
  INV_X1 U117 ( .A(n4746), .ZN(n4747) );
  INV_X1 U118 ( .A(n4748), .ZN(n4749) );
  INV_X1 U119 ( .A(n4750), .ZN(n4751) );
  INV_X1 U120 ( .A(n4752), .ZN(n4753) );
  INV_X1 U121 ( .A(n4754), .ZN(n4755) );
  INV_X1 U122 ( .A(n4756), .ZN(n4757) );
  INV_X1 U123 ( .A(n4758), .ZN(n4759) );
  INV_X1 U124 ( .A(n4760), .ZN(n4761) );
  INV_X1 U125 ( .A(n4762), .ZN(n4763) );
  INV_X1 U126 ( .A(n4764), .ZN(n4765) );
  INV_X1 U127 ( .A(n4766), .ZN(n4767) );
  INV_X1 U128 ( .A(n4768), .ZN(n4769) );
  INV_X1 U129 ( .A(n4770), .ZN(n4771) );
  INV_X1 U130 ( .A(n4772), .ZN(n4773) );
  INV_X1 U131 ( .A(n4774), .ZN(n4775) );
  INV_X1 U132 ( .A(n4776), .ZN(n4777) );
  INV_X1 U133 ( .A(n4778), .ZN(n4779) );
  INV_X1 U134 ( .A(n4780), .ZN(n4781) );
  INV_X1 U135 ( .A(n4782), .ZN(n4783) );
  INV_X1 U136 ( .A(n4784), .ZN(n4785) );
  INV_X1 U137 ( .A(n4786), .ZN(n4787) );
  INV_X1 U138 ( .A(n4788), .ZN(n4789) );
  INV_X1 U139 ( .A(n4790), .ZN(n4791) );
  INV_X1 U140 ( .A(n4792), .ZN(n4793) );
  INV_X1 U141 ( .A(n4794), .ZN(n4795) );
  INV_X1 U142 ( .A(n4796), .ZN(n4797) );
  INV_X1 U143 ( .A(n4798), .ZN(n4799) );
  INV_X1 U144 ( .A(n4800), .ZN(n4801) );
  INV_X1 U145 ( .A(n4802), .ZN(n4803) );
  INV_X1 U146 ( .A(n4804), .ZN(n4805) );
  INV_X1 U147 ( .A(n4806), .ZN(n4807) );
  INV_X1 U148 ( .A(n4808), .ZN(n4809) );
  INV_X1 U149 ( .A(n4810), .ZN(n4811) );
  INV_X1 U150 ( .A(n4812), .ZN(n4813) );
  INV_X1 U151 ( .A(n4814), .ZN(n4815) );
  BUF_X1 U152 ( .A(n4641), .Z(n6007) );
  NAND2_X1 U153 ( .A1(DATAIN[17]), .A2(n6006), .ZN(n4844) );
  NAND2_X1 U154 ( .A1(DATAIN[24]), .A2(n6007), .ZN(n4826) );
  NAND2_X1 U155 ( .A1(DATAIN[25]), .A2(n6007), .ZN(n4824) );
  NAND2_X1 U156 ( .A1(DATAIN[26]), .A2(n6007), .ZN(n4822) );
  NAND2_X1 U157 ( .A1(DATAIN[27]), .A2(n6007), .ZN(n4820) );
  NAND2_X1 U158 ( .A1(DATAIN[28]), .A2(n6007), .ZN(n4818) );
  NAND2_X1 U159 ( .A1(n5205), .A2(n4816), .ZN(n4817) );
  NAND2_X1 U160 ( .A1(n4817), .A2(n4818), .ZN(n4282) );
  INV_X1 U161 ( .A(n6007), .ZN(n4816) );
  NAND2_X1 U162 ( .A1(n5206), .A2(n4836), .ZN(n4819) );
  NAND2_X1 U163 ( .A1(n4819), .A2(n4820), .ZN(n4281) );
  NAND2_X1 U164 ( .A1(n5207), .A2(n4833), .ZN(n4821) );
  NAND2_X1 U165 ( .A1(n4821), .A2(n4822), .ZN(n4280) );
  NAND2_X1 U166 ( .A1(n5208), .A2(n4830), .ZN(n4823) );
  NAND2_X1 U167 ( .A1(n4823), .A2(n4824), .ZN(n4279) );
  NAND2_X1 U168 ( .A1(n5209), .A2(n4827), .ZN(n4825) );
  NAND2_X1 U169 ( .A1(n4825), .A2(n4826), .ZN(n4278) );
  BUF_X1 U170 ( .A(n4641), .Z(n6006) );
  NAND2_X1 U171 ( .A1(DATAIN[14]), .A2(n6006), .ZN(n4853) );
  NAND2_X1 U172 ( .A1(DATAIN[18]), .A2(n6006), .ZN(n4841) );
  NAND2_X1 U173 ( .A1(DATAIN[19]), .A2(n6006), .ZN(n4838) );
  NAND2_X1 U174 ( .A1(DATAIN[20]), .A2(n6006), .ZN(n4835) );
  NAND2_X1 U175 ( .A1(DATAIN[21]), .A2(n6006), .ZN(n4832) );
  NAND2_X1 U176 ( .A1(DATAIN[22]), .A2(n6006), .ZN(n4829) );
  NAND2_X1 U177 ( .A1(n5211), .A2(n4827), .ZN(n4828) );
  NAND2_X1 U178 ( .A1(n4828), .A2(n4829), .ZN(n4276) );
  INV_X1 U179 ( .A(n6006), .ZN(n4827) );
  NAND2_X1 U180 ( .A1(n5212), .A2(n4830), .ZN(n4831) );
  NAND2_X1 U181 ( .A1(n4831), .A2(n4832), .ZN(n4275) );
  INV_X1 U182 ( .A(n6006), .ZN(n4830) );
  NAND2_X1 U183 ( .A1(n5213), .A2(n4833), .ZN(n4834) );
  NAND2_X1 U184 ( .A1(n4834), .A2(n4835), .ZN(n4274) );
  INV_X1 U185 ( .A(n6006), .ZN(n4833) );
  NAND2_X1 U186 ( .A1(n5214), .A2(n4836), .ZN(n4837) );
  NAND2_X1 U187 ( .A1(n4837), .A2(n4838), .ZN(n4273) );
  INV_X1 U188 ( .A(n6006), .ZN(n4836) );
  NAND2_X1 U189 ( .A1(n5215), .A2(n4839), .ZN(n4840) );
  NAND2_X1 U190 ( .A1(n4840), .A2(n4841), .ZN(n4272) );
  INV_X1 U191 ( .A(n6006), .ZN(n4839) );
  NAND2_X1 U192 ( .A1(n5216), .A2(n4842), .ZN(n4843) );
  NAND2_X1 U193 ( .A1(n4843), .A2(n4844), .ZN(n4271) );
  INV_X1 U194 ( .A(n6006), .ZN(n4842) );
  BUF_X1 U195 ( .A(n4641), .Z(n6005) );
  NAND2_X1 U196 ( .A1(DATAIN[8]), .A2(n6005), .ZN(n4871) );
  NAND2_X1 U197 ( .A1(DATAIN[15]), .A2(n6006), .ZN(n4850) );
  NAND2_X1 U198 ( .A1(DATAIN[16]), .A2(n6006), .ZN(n4847) );
  NAND2_X1 U199 ( .A1(n5217), .A2(n4845), .ZN(n4846) );
  NAND2_X1 U200 ( .A1(n4846), .A2(n4847), .ZN(n4270) );
  INV_X1 U201 ( .A(n6006), .ZN(n4845) );
  NAND2_X1 U202 ( .A1(n5218), .A2(n4848), .ZN(n4849) );
  NAND2_X1 U203 ( .A1(n4849), .A2(n4850), .ZN(n4269) );
  INV_X1 U204 ( .A(n6006), .ZN(n4848) );
  NAND2_X1 U205 ( .A1(n5219), .A2(n4851), .ZN(n4852) );
  NAND2_X1 U206 ( .A1(n4852), .A2(n4853), .ZN(n4268) );
  INV_X1 U207 ( .A(n6006), .ZN(n4851) );
  NAND2_X1 U208 ( .A1(DATAIN[6]), .A2(n6005), .ZN(n4877) );
  NAND2_X1 U209 ( .A1(DATAIN[9]), .A2(n6005), .ZN(n4868) );
  NAND2_X1 U210 ( .A1(DATAIN[10]), .A2(n6005), .ZN(n4865) );
  NAND2_X1 U211 ( .A1(DATAIN[11]), .A2(n6005), .ZN(n4862) );
  NAND2_X1 U212 ( .A1(DATAIN[12]), .A2(n6006), .ZN(n4859) );
  NAND2_X1 U213 ( .A1(DATAIN[13]), .A2(n6006), .ZN(n4856) );
  NAND2_X1 U214 ( .A1(n5220), .A2(n4854), .ZN(n4855) );
  NAND2_X1 U215 ( .A1(n4855), .A2(n4856), .ZN(n4267) );
  INV_X1 U216 ( .A(n6006), .ZN(n4854) );
  NAND2_X1 U217 ( .A1(n5221), .A2(n4857), .ZN(n4858) );
  NAND2_X1 U218 ( .A1(n4858), .A2(n4859), .ZN(n4266) );
  INV_X1 U219 ( .A(n6006), .ZN(n4857) );
  NAND2_X1 U220 ( .A1(n5222), .A2(n4860), .ZN(n4861) );
  NAND2_X1 U221 ( .A1(n4861), .A2(n4862), .ZN(n4265) );
  INV_X1 U222 ( .A(n6005), .ZN(n4860) );
  NAND2_X1 U223 ( .A1(n5223), .A2(n4863), .ZN(n4864) );
  NAND2_X1 U224 ( .A1(n4864), .A2(n4865), .ZN(n4264) );
  INV_X1 U225 ( .A(n6005), .ZN(n4863) );
  NAND2_X1 U226 ( .A1(n5224), .A2(n4866), .ZN(n4867) );
  NAND2_X1 U227 ( .A1(n4867), .A2(n4868), .ZN(n4263) );
  INV_X1 U228 ( .A(n6005), .ZN(n4866) );
  NAND2_X1 U229 ( .A1(n5225), .A2(n4869), .ZN(n4870) );
  NAND2_X1 U230 ( .A1(n4870), .A2(n4871), .ZN(n4262) );
  INV_X1 U231 ( .A(n6005), .ZN(n4869) );
  NAND2_X1 U232 ( .A1(DATAIN[4]), .A2(n6005), .ZN(n4883) );
  NAND2_X1 U233 ( .A1(DATAIN[7]), .A2(n6005), .ZN(n4874) );
  NAND2_X1 U234 ( .A1(n5226), .A2(n4872), .ZN(n4873) );
  NAND2_X1 U235 ( .A1(n4873), .A2(n4874), .ZN(n4261) );
  INV_X1 U236 ( .A(n6005), .ZN(n4872) );
  NAND2_X1 U237 ( .A1(n5227), .A2(n4875), .ZN(n4876) );
  NAND2_X1 U238 ( .A1(n4876), .A2(n4877), .ZN(n4260) );
  INV_X1 U239 ( .A(n6005), .ZN(n4875) );
  NAND2_X1 U240 ( .A1(DATAIN[2]), .A2(n6005), .ZN(n4889) );
  NAND2_X1 U241 ( .A1(DATAIN[5]), .A2(n6005), .ZN(n4880) );
  NAND2_X1 U242 ( .A1(n5228), .A2(n4878), .ZN(n4879) );
  NAND2_X1 U243 ( .A1(n4879), .A2(n4880), .ZN(n4259) );
  INV_X1 U244 ( .A(n6005), .ZN(n4878) );
  NAND2_X1 U245 ( .A1(n5229), .A2(n4881), .ZN(n4882) );
  NAND2_X1 U246 ( .A1(n4882), .A2(n4883), .ZN(n4258) );
  INV_X1 U247 ( .A(n6005), .ZN(n4881) );
  NAND2_X1 U248 ( .A1(DATAIN[0]), .A2(n6005), .ZN(n4895) );
  NAND2_X1 U249 ( .A1(DATAIN[3]), .A2(n6005), .ZN(n4886) );
  NAND2_X1 U250 ( .A1(n5230), .A2(n4884), .ZN(n4885) );
  NAND2_X1 U251 ( .A1(n4885), .A2(n4886), .ZN(n4257) );
  INV_X1 U252 ( .A(n6005), .ZN(n4884) );
  NAND2_X1 U253 ( .A1(n5231), .A2(n4887), .ZN(n4888) );
  NAND2_X1 U254 ( .A1(n4888), .A2(n4889), .ZN(n4256) );
  INV_X1 U255 ( .A(n6005), .ZN(n4887) );
  NAND2_X1 U256 ( .A1(DATAIN[1]), .A2(n6005), .ZN(n4892) );
  NAND2_X1 U257 ( .A1(n5232), .A2(n4890), .ZN(n4891) );
  NAND2_X1 U258 ( .A1(n4891), .A2(n4892), .ZN(n4255) );
  INV_X1 U259 ( .A(n6005), .ZN(n4890) );
  NAND2_X1 U260 ( .A1(n5170), .A2(n4893), .ZN(n4894) );
  NAND2_X1 U261 ( .A1(n4894), .A2(n4895), .ZN(n4254) );
  INV_X1 U262 ( .A(n6005), .ZN(n4893) );
  INV_X1 U263 ( .A(n6075), .ZN(n6074) );
  INV_X1 U264 ( .A(n6075), .ZN(n6073) );
  INV_X1 U265 ( .A(n6093), .ZN(n6091) );
  BUF_X1 U266 ( .A(n6465), .Z(n6464) );
  BUF_X1 U267 ( .A(n7511), .Z(n6180) );
  BUF_X1 U268 ( .A(n7511), .Z(n6179) );
  BUF_X1 U269 ( .A(n6908), .Z(n6127) );
  BUF_X1 U270 ( .A(n6911), .Z(n6138) );
  BUF_X1 U271 ( .A(n6919), .Z(n6167) );
  BUF_X1 U272 ( .A(n6908), .Z(n6128) );
  BUF_X1 U273 ( .A(n6911), .Z(n6139) );
  BUF_X1 U274 ( .A(n6919), .Z(n6168) );
  BUF_X1 U275 ( .A(n7525), .Z(n6202) );
  BUF_X1 U276 ( .A(n7525), .Z(n6203) );
  BUF_X1 U277 ( .A(n4633), .Z(n6124) );
  BUF_X1 U278 ( .A(n4634), .Z(n6135) );
  BUF_X1 U279 ( .A(n6910), .Z(n6130) );
  BUF_X1 U280 ( .A(n6910), .Z(n6131) );
  BUF_X1 U281 ( .A(n4633), .Z(n6125) );
  BUF_X1 U282 ( .A(n4634), .Z(n6136) );
  BUF_X1 U283 ( .A(n7525), .Z(n6204) );
  BUF_X1 U284 ( .A(n6910), .Z(n6132) );
  BUF_X1 U285 ( .A(n4633), .Z(n6126) );
  BUF_X1 U286 ( .A(n4634), .Z(n6137) );
  BUF_X1 U287 ( .A(n6908), .Z(n6129) );
  BUF_X1 U288 ( .A(n6911), .Z(n6140) );
  BUF_X1 U289 ( .A(n6919), .Z(n6169) );
  BUF_X1 U290 ( .A(n7511), .Z(n6181) );
  INV_X1 U291 ( .A(n4902), .ZN(n6288) );
  INV_X1 U292 ( .A(n4902), .ZN(n6289) );
  INV_X1 U293 ( .A(n4901), .ZN(n6326) );
  INV_X1 U294 ( .A(n4901), .ZN(n6325) );
  INV_X1 U295 ( .A(n4900), .ZN(n6271) );
  INV_X1 U296 ( .A(n4900), .ZN(n6272) );
  INV_X1 U297 ( .A(n4899), .ZN(n6309) );
  INV_X1 U298 ( .A(n4899), .ZN(n6308) );
  INV_X1 U299 ( .A(n6102), .ZN(n6100) );
  INV_X1 U300 ( .A(n6111), .ZN(n6109) );
  INV_X1 U301 ( .A(n6102), .ZN(n6101) );
  INV_X1 U302 ( .A(n6111), .ZN(n6110) );
  INV_X1 U303 ( .A(n6057), .ZN(n6056) );
  INV_X1 U304 ( .A(n6057), .ZN(n6055) );
  INV_X1 U305 ( .A(n6066), .ZN(n6065) );
  INV_X1 U306 ( .A(n6066), .ZN(n6064) );
  INV_X1 U307 ( .A(n6084), .ZN(n6082) );
  INV_X1 U308 ( .A(n4897), .ZN(n6119) );
  INV_X1 U309 ( .A(n4897), .ZN(n6120) );
  INV_X1 U310 ( .A(n4898), .ZN(n6133) );
  INV_X1 U311 ( .A(n4898), .ZN(n6134) );
  INV_X1 U312 ( .A(n4896), .ZN(n6182) );
  INV_X1 U313 ( .A(n4896), .ZN(n6183) );
  BUF_X1 U314 ( .A(n1458), .Z(n6274) );
  BUF_X1 U315 ( .A(n1458), .Z(n6273) );
  BUF_X1 U316 ( .A(n845), .Z(n6310) );
  BUF_X1 U317 ( .A(n845), .Z(n6311) );
  BUF_X1 U318 ( .A(n1453), .Z(n6286) );
  BUF_X1 U319 ( .A(n1453), .Z(n6285) );
  BUF_X1 U320 ( .A(n840), .Z(n6322) );
  BUF_X1 U321 ( .A(n840), .Z(n6323) );
  BUF_X1 U322 ( .A(n845), .Z(n6312) );
  BUF_X1 U323 ( .A(n1458), .Z(n6275) );
  BUF_X1 U324 ( .A(n1453), .Z(n6287) );
  BUF_X1 U325 ( .A(n840), .Z(n6324) );
  BUF_X1 U326 ( .A(n4906), .Z(n6149) );
  BUF_X1 U327 ( .A(n4906), .Z(n6150) );
  BUF_X1 U328 ( .A(n4904), .Z(n6223) );
  BUF_X1 U329 ( .A(n4904), .Z(n6224) );
  BUF_X1 U330 ( .A(n4629), .Z(n6208) );
  BUF_X1 U331 ( .A(n4628), .Z(n6196) );
  BUF_X1 U332 ( .A(n4628), .Z(n6197) );
  BUF_X1 U333 ( .A(n4629), .Z(n6209) );
  BUF_X1 U334 ( .A(n4908), .Z(n6229) );
  BUF_X1 U335 ( .A(n4908), .Z(n6230) );
  BUF_X1 U336 ( .A(n4905), .Z(n6146) );
  BUF_X1 U337 ( .A(n4905), .Z(n6147) );
  BUF_X1 U338 ( .A(n4903), .Z(n6220) );
  BUF_X1 U339 ( .A(n4903), .Z(n6221) );
  BUF_X1 U340 ( .A(n7520), .Z(n6187) );
  BUF_X1 U341 ( .A(n7520), .Z(n6188) );
  BUF_X1 U342 ( .A(n7529), .Z(n6214) );
  BUF_X1 U343 ( .A(n7529), .Z(n6215) );
  BUF_X1 U344 ( .A(n4907), .Z(n6155) );
  BUF_X1 U345 ( .A(n4907), .Z(n6156) );
  BUF_X1 U346 ( .A(n4631), .Z(n6159) );
  BUF_X1 U347 ( .A(n4631), .Z(n6158) );
  BUF_X1 U348 ( .A(n4632), .Z(n6217) );
  BUF_X1 U349 ( .A(n4632), .Z(n6218) );
  BUF_X1 U350 ( .A(n7519), .Z(n6185) );
  BUF_X1 U351 ( .A(n7519), .Z(n6184) );
  BUF_X1 U352 ( .A(n6907), .Z(n6121) );
  BUF_X1 U353 ( .A(n6907), .Z(n6122) );
  BUF_X1 U354 ( .A(n4659), .Z(n6164) );
  BUF_X1 U355 ( .A(n6913), .Z(n6141) );
  BUF_X1 U356 ( .A(n6913), .Z(n6142) );
  BUF_X1 U357 ( .A(n7528), .Z(n6211) );
  BUF_X1 U358 ( .A(n7528), .Z(n6212) );
  BUF_X1 U359 ( .A(n7524), .Z(n6199) );
  BUF_X1 U360 ( .A(n7524), .Z(n6200) );
  BUF_X1 U361 ( .A(n4659), .Z(n6165) );
  BUF_X1 U362 ( .A(n4627), .Z(n6193) );
  BUF_X1 U363 ( .A(n4630), .Z(n6205) );
  BUF_X1 U364 ( .A(n4627), .Z(n6194) );
  BUF_X1 U365 ( .A(n4630), .Z(n6206) );
  BUF_X1 U366 ( .A(n7522), .Z(n6190) );
  BUF_X1 U367 ( .A(n4909), .Z(n6152) );
  BUF_X1 U368 ( .A(n4909), .Z(n6153) );
  BUF_X1 U369 ( .A(n7522), .Z(n6191) );
  BUF_X1 U370 ( .A(n6906), .Z(n6116) );
  BUF_X1 U371 ( .A(n6906), .Z(n6117) );
  BUF_X1 U372 ( .A(n4910), .Z(n6226) );
  BUF_X1 U373 ( .A(n4910), .Z(n6227) );
  BUF_X1 U374 ( .A(n6922), .Z(n6170) );
  BUF_X1 U375 ( .A(n6922), .Z(n6171) );
  BUF_X1 U376 ( .A(n6071), .Z(n6075) );
  BUF_X1 U377 ( .A(n6089), .Z(n6093) );
  BUF_X1 U378 ( .A(n835), .Z(n6334) );
  BUF_X1 U379 ( .A(n1448), .Z(n6297) );
  BUF_X1 U380 ( .A(n835), .Z(n6333) );
  BUF_X1 U381 ( .A(n1448), .Z(n6296) );
  BUF_X1 U382 ( .A(n843), .Z(n6317) );
  BUF_X1 U383 ( .A(n843), .Z(n6316) );
  BUF_X1 U384 ( .A(n1456), .Z(n6280) );
  BUF_X1 U385 ( .A(n1456), .Z(n6279) );
  BUF_X1 U386 ( .A(n838), .Z(n6328) );
  BUF_X1 U387 ( .A(n838), .Z(n6327) );
  BUF_X1 U388 ( .A(n1451), .Z(n6291) );
  BUF_X1 U389 ( .A(n1462), .Z(n6266) );
  BUF_X1 U390 ( .A(n849), .Z(n6303) );
  BUF_X1 U391 ( .A(n849), .Z(n6302) );
  BUF_X1 U392 ( .A(n1462), .Z(n6265) );
  BUF_X1 U393 ( .A(n1451), .Z(n6290) );
  BUF_X1 U394 ( .A(n842), .Z(n6320) );
  BUF_X1 U395 ( .A(n842), .Z(n6319) );
  BUF_X1 U396 ( .A(n1455), .Z(n6283) );
  BUF_X1 U397 ( .A(n1455), .Z(n6282) );
  BUF_X1 U398 ( .A(n4904), .Z(n6225) );
  BUF_X1 U399 ( .A(n4906), .Z(n6151) );
  BUF_X1 U400 ( .A(n4629), .Z(n6210) );
  BUF_X1 U401 ( .A(n4628), .Z(n6198) );
  BUF_X1 U402 ( .A(n1461), .Z(n6269) );
  BUF_X1 U403 ( .A(n848), .Z(n6306) );
  BUF_X1 U404 ( .A(n848), .Z(n6305) );
  BUF_X1 U405 ( .A(n1461), .Z(n6268) );
  BUF_X1 U406 ( .A(n837), .Z(n6331) );
  BUF_X1 U407 ( .A(n837), .Z(n6330) );
  BUF_X1 U408 ( .A(n1450), .Z(n6294) );
  BUF_X1 U409 ( .A(n1450), .Z(n6293) );
  BUF_X1 U410 ( .A(n834), .Z(n6337) );
  BUF_X1 U411 ( .A(n1447), .Z(n6300) );
  BUF_X1 U412 ( .A(n834), .Z(n6336) );
  BUF_X1 U413 ( .A(n1447), .Z(n6299) );
  BUF_X1 U414 ( .A(n844), .Z(n6314) );
  BUF_X1 U415 ( .A(n844), .Z(n6313) );
  BUF_X1 U416 ( .A(n1457), .Z(n6277) );
  BUF_X1 U417 ( .A(n1457), .Z(n6276) );
  BUF_X1 U418 ( .A(n4908), .Z(n6231) );
  BUF_X1 U419 ( .A(n835), .Z(n6335) );
  BUF_X1 U420 ( .A(n1448), .Z(n6298) );
  BUF_X1 U421 ( .A(n7520), .Z(n6189) );
  BUF_X1 U422 ( .A(n4903), .Z(n6222) );
  BUF_X1 U423 ( .A(n4905), .Z(n6148) );
  BUF_X1 U424 ( .A(n843), .Z(n6318) );
  BUF_X1 U425 ( .A(n1456), .Z(n6281) );
  BUF_X1 U426 ( .A(n1462), .Z(n6267) );
  BUF_X1 U427 ( .A(n1451), .Z(n6292) );
  BUF_X1 U428 ( .A(n838), .Z(n6329) );
  BUF_X1 U429 ( .A(n849), .Z(n6304) );
  BUF_X1 U430 ( .A(n7529), .Z(n6216) );
  BUF_X1 U431 ( .A(n4907), .Z(n6157) );
  BUF_X1 U432 ( .A(n6907), .Z(n6123) );
  BUF_X1 U433 ( .A(n4632), .Z(n6219) );
  BUF_X1 U434 ( .A(n4631), .Z(n6160) );
  BUF_X1 U435 ( .A(n842), .Z(n6321) );
  BUF_X1 U436 ( .A(n1455), .Z(n6284) );
  BUF_X1 U437 ( .A(n6913), .Z(n6143) );
  BUF_X1 U438 ( .A(n7519), .Z(n6186) );
  BUF_X1 U439 ( .A(n7528), .Z(n6213) );
  BUF_X1 U440 ( .A(n7524), .Z(n6201) );
  BUF_X1 U441 ( .A(n1461), .Z(n6270) );
  BUF_X1 U442 ( .A(n848), .Z(n6307) );
  BUF_X1 U443 ( .A(n1450), .Z(n6295) );
  BUF_X1 U444 ( .A(n837), .Z(n6332) );
  BUF_X1 U445 ( .A(n4627), .Z(n6195) );
  BUF_X1 U446 ( .A(n4630), .Z(n6207) );
  BUF_X1 U447 ( .A(n4659), .Z(n6166) );
  BUF_X1 U448 ( .A(n4909), .Z(n6154) );
  BUF_X1 U449 ( .A(n7522), .Z(n6192) );
  BUF_X1 U450 ( .A(n834), .Z(n6338) );
  BUF_X1 U451 ( .A(n1447), .Z(n6301) );
  BUF_X1 U452 ( .A(n6906), .Z(n6118) );
  BUF_X1 U453 ( .A(n844), .Z(n6315) );
  BUF_X1 U454 ( .A(n1457), .Z(n6278) );
  BUF_X1 U455 ( .A(n4910), .Z(n6228) );
  BUF_X1 U456 ( .A(n6922), .Z(n6172) );
  BUF_X1 U457 ( .A(n6071), .Z(n6076) );
  BUF_X1 U458 ( .A(n6071), .Z(n6077) );
  BUF_X1 U459 ( .A(n6089), .Z(n6094) );
  BUF_X1 U460 ( .A(n6089), .Z(n6095) );
  BUF_X1 U461 ( .A(n6072), .Z(n6078) );
  BUF_X1 U462 ( .A(n6072), .Z(n6079) );
  BUF_X1 U463 ( .A(n6090), .Z(n6096) );
  BUF_X1 U464 ( .A(n6090), .Z(n6097) );
  BUF_X1 U465 ( .A(n6375), .Z(n6465) );
  BUF_X1 U466 ( .A(n6377), .Z(n6472) );
  BUF_X1 U467 ( .A(n6377), .Z(n6471) );
  BUF_X1 U468 ( .A(n6376), .Z(n6470) );
  BUF_X1 U469 ( .A(n6377), .Z(n6473) );
  BUF_X1 U470 ( .A(n6378), .Z(n6475) );
  BUF_X1 U471 ( .A(n6378), .Z(n6474) );
  BUF_X1 U472 ( .A(n6378), .Z(n6476) );
  BUF_X1 U473 ( .A(n6375), .Z(n6466) );
  BUF_X1 U474 ( .A(n6375), .Z(n6467) );
  BUF_X1 U475 ( .A(n6376), .Z(n6469) );
  BUF_X1 U476 ( .A(n6376), .Z(n6468) );
  BUF_X1 U477 ( .A(n6379), .Z(n6477) );
  BUF_X1 U478 ( .A(n6379), .Z(n6478) );
  NOR2_X1 U479 ( .A1(n7898), .A2(n6480), .ZN(n1412) );
  NOR2_X1 U480 ( .A1(n7900), .A2(n6479), .ZN(n2012) );
  NOR3_X1 U481 ( .A1(n7592), .A2(n7593), .A3(n7901), .ZN(n2006) );
  NOR3_X1 U482 ( .A1(n7594), .A2(n7595), .A3(n7899), .ZN(n1406) );
  BUF_X1 U483 ( .A(n6484), .Z(n6033) );
  BUF_X1 U484 ( .A(n6484), .Z(n6032) );
  BUF_X1 U485 ( .A(n4650), .Z(n6014) );
  BUF_X1 U486 ( .A(n4650), .Z(n6015) );
  BUF_X1 U487 ( .A(n6916), .Z(n6161) );
  BUF_X1 U488 ( .A(n6916), .Z(n6162) );
  BUF_X1 U489 ( .A(n7510), .Z(n6176) );
  BUF_X1 U490 ( .A(n7510), .Z(n6177) );
  NAND2_X1 U491 ( .A1(n2023), .A2(n2012), .ZN(n1462) );
  NAND2_X1 U492 ( .A1(n2022), .A2(n2013), .ZN(n1456) );
  NAND2_X1 U493 ( .A1(n2023), .A2(n2013), .ZN(n1455) );
  NAND2_X1 U494 ( .A1(n2022), .A2(n1994), .ZN(n1457) );
  NAND2_X1 U495 ( .A1(n2022), .A2(n4613), .ZN(n1451) );
  NAND2_X1 U496 ( .A1(n2023), .A2(n4613), .ZN(n1450) );
  NAND2_X1 U497 ( .A1(n1422), .A2(n1413), .ZN(n843) );
  NAND2_X1 U498 ( .A1(n1423), .A2(n1413), .ZN(n842) );
  NAND2_X1 U499 ( .A1(n1422), .A2(n1394), .ZN(n844) );
  NAND2_X1 U500 ( .A1(n1423), .A2(n1412), .ZN(n849) );
  NAND2_X1 U501 ( .A1(n1422), .A2(n4608), .ZN(n838) );
  NAND2_X1 U502 ( .A1(n1423), .A2(n4608), .ZN(n837) );
  NAND2_X1 U503 ( .A1(n1394), .A2(n1419), .ZN(n848) );
  BUF_X1 U504 ( .A(n6916), .Z(n6163) );
  NAND2_X1 U505 ( .A1(n1994), .A2(n2019), .ZN(n1461) );
  BUF_X1 U506 ( .A(n4650), .Z(n6016) );
  AND2_X1 U507 ( .A1(n4617), .A2(n4608), .ZN(n4896) );
  BUF_X1 U508 ( .A(n6484), .Z(n6034) );
  BUF_X1 U509 ( .A(n6232), .Z(n6234) );
  BUF_X1 U510 ( .A(n6232), .Z(n6235) );
  BUF_X1 U511 ( .A(n6233), .Z(n6236) );
  BUF_X1 U512 ( .A(n6053), .Z(n6057) );
  BUF_X1 U513 ( .A(n6062), .Z(n6066) );
  BUF_X1 U514 ( .A(n6080), .Z(n6084) );
  BUF_X1 U515 ( .A(n6098), .Z(n6102) );
  BUF_X1 U516 ( .A(n6107), .Z(n6111) );
  AND2_X1 U517 ( .A1(n4612), .A2(n4626), .ZN(n4897) );
  AND2_X1 U518 ( .A1(n4612), .A2(n4661), .ZN(n4898) );
  AND2_X1 U519 ( .A1(n2022), .A2(n2012), .ZN(n1453) );
  AND2_X1 U520 ( .A1(n1422), .A2(n1412), .ZN(n840) );
  NAND2_X1 U521 ( .A1(n1420), .A2(n1394), .ZN(n4899) );
  NAND2_X1 U522 ( .A1(n2020), .A2(n1994), .ZN(n4900) );
  NAND2_X1 U523 ( .A1(n1423), .A2(n1394), .ZN(n4901) );
  NAND2_X1 U524 ( .A1(n2023), .A2(n1994), .ZN(n4902) );
  AND2_X1 U525 ( .A1(n1413), .A2(n1420), .ZN(n835) );
  AND2_X1 U526 ( .A1(n1413), .A2(n1419), .ZN(n834) );
  AND2_X1 U527 ( .A1(n1406), .A2(n1394), .ZN(n845) );
  AND2_X1 U528 ( .A1(n2006), .A2(n1994), .ZN(n1458) );
  AND2_X1 U529 ( .A1(n2013), .A2(n2019), .ZN(n1447) );
  AND2_X1 U530 ( .A1(n2013), .A2(n2020), .ZN(n1448) );
  AND2_X1 U531 ( .A1(n1394), .A2(n1393), .ZN(n4903) );
  AND2_X1 U532 ( .A1(n1412), .A2(n1393), .ZN(n4904) );
  AND2_X1 U533 ( .A1(n1994), .A2(n1993), .ZN(n4905) );
  AND2_X1 U534 ( .A1(n2012), .A2(n1993), .ZN(n4906) );
  BUF_X1 U535 ( .A(n6053), .Z(n6058) );
  BUF_X1 U536 ( .A(n6053), .Z(n6059) );
  BUF_X1 U537 ( .A(n6062), .Z(n6067) );
  BUF_X1 U538 ( .A(n6062), .Z(n6068) );
  BUF_X1 U539 ( .A(n6080), .Z(n6085) );
  BUF_X1 U540 ( .A(n6080), .Z(n6086) );
  BUF_X1 U541 ( .A(n6098), .Z(n6103) );
  BUF_X1 U542 ( .A(n6098), .Z(n6104) );
  BUF_X1 U543 ( .A(n6107), .Z(n6112) );
  BUF_X1 U544 ( .A(n6107), .Z(n6113) );
  BUF_X1 U545 ( .A(n6054), .Z(n6060) );
  BUF_X1 U546 ( .A(n6054), .Z(n6061) );
  BUF_X1 U547 ( .A(n6063), .Z(n6069) );
  BUF_X1 U548 ( .A(n6063), .Z(n6070) );
  BUF_X1 U549 ( .A(n6081), .Z(n6087) );
  BUF_X1 U550 ( .A(n6081), .Z(n6088) );
  BUF_X1 U551 ( .A(n6099), .Z(n6105) );
  BUF_X1 U552 ( .A(n6108), .Z(n6114) );
  NAND2_X1 U553 ( .A1(n2012), .A2(n2019), .ZN(n4907) );
  NAND2_X1 U554 ( .A1(n1412), .A2(n1419), .ZN(n4908) );
  NAND2_X1 U555 ( .A1(n2020), .A2(n2012), .ZN(n4909) );
  NAND2_X1 U556 ( .A1(n1420), .A2(n1412), .ZN(n4910) );
  BUF_X1 U557 ( .A(n7510), .Z(n6178) );
  BUF_X1 U558 ( .A(n6233), .Z(n6237) );
  BUF_X1 U559 ( .A(n6099), .Z(n6106) );
  BUF_X1 U560 ( .A(n6108), .Z(n6115) );
  BUF_X1 U561 ( .A(n6488), .Z(n6071) );
  BUF_X1 U562 ( .A(n6491), .Z(n6089) );
  BUF_X1 U563 ( .A(n6380), .Z(n6377) );
  BUF_X1 U564 ( .A(n6380), .Z(n6378) );
  BUF_X1 U565 ( .A(n6381), .Z(n6375) );
  BUF_X1 U566 ( .A(n6381), .Z(n6376) );
  BUF_X1 U567 ( .A(n6488), .Z(n6072) );
  BUF_X1 U568 ( .A(n6491), .Z(n6090) );
  BUF_X1 U569 ( .A(n6380), .Z(n6379) );
  NOR3_X1 U570 ( .A1(ADD_RS1[0]), .A2(ADD_RS1[4]), .A3(n7592), .ZN(n2022) );
  NOR3_X1 U571 ( .A1(n7593), .A2(ADD_RS1[4]), .A3(n7592), .ZN(n2023) );
  NOR3_X1 U572 ( .A1(ADD_RS2[0]), .A2(ADD_RS2[4]), .A3(n7594), .ZN(n1422) );
  NOR3_X1 U573 ( .A1(n7595), .A2(ADD_RS2[4]), .A3(n7594), .ZN(n1423) );
  NOR2_X1 U574 ( .A1(n7898), .A2(ADD_RS2[1]), .ZN(n1394) );
  NOR3_X1 U575 ( .A1(ADD_RS1[0]), .A2(ADD_RS1[3]), .A3(n7901), .ZN(n1993) );
  NOR3_X1 U576 ( .A1(ADD_RS2[0]), .A2(ADD_RS2[3]), .A3(n7899), .ZN(n1393) );
  NOR2_X1 U577 ( .A1(n6480), .A2(ADD_RS2[2]), .ZN(n1413) );
  NOR2_X1 U578 ( .A1(n7900), .A2(ADD_RS1[1]), .ZN(n1994) );
  NOR3_X1 U579 ( .A1(ADD_RS1[3]), .A2(ADD_RS1[4]), .A3(n7593), .ZN(n2019) );
  NOR3_X1 U580 ( .A1(ADD_RS2[3]), .A2(ADD_RS2[4]), .A3(n7595), .ZN(n1419) );
  NOR2_X1 U581 ( .A1(n6479), .A2(ADD_RS1[2]), .ZN(n2013) );
  NOR3_X1 U582 ( .A1(ADD_RS1[3]), .A2(ADD_RS1[4]), .A3(ADD_RS1[0]), .ZN(n2020)
         );
  NOR3_X1 U583 ( .A1(ADD_RS2[3]), .A2(ADD_RS2[4]), .A3(ADD_RS2[0]), .ZN(n1420)
         );
  INV_X1 U584 ( .A(n4616), .ZN(n6144) );
  INV_X1 U585 ( .A(n4616), .ZN(n6145) );
  BUF_X1 U586 ( .A(n4643), .Z(n6008) );
  BUF_X1 U587 ( .A(n4643), .Z(n6009) );
  BUF_X1 U588 ( .A(n4644), .Z(n6011) );
  BUF_X1 U589 ( .A(n4644), .Z(n6012) );
  BUF_X1 U590 ( .A(n4651), .Z(n6017) );
  BUF_X1 U591 ( .A(n4651), .Z(n6018) );
  BUF_X1 U592 ( .A(n4636), .Z(n6020) );
  BUF_X1 U593 ( .A(n4636), .Z(n6021) );
  BUF_X1 U594 ( .A(n4645), .Z(n6023) );
  BUF_X1 U595 ( .A(n4645), .Z(n6024) );
  BUF_X1 U596 ( .A(n4646), .Z(n6026) );
  BUF_X1 U597 ( .A(n4646), .Z(n6027) );
  BUF_X1 U598 ( .A(n4652), .Z(n6029) );
  BUF_X1 U599 ( .A(n4652), .Z(n6030) );
  BUF_X1 U600 ( .A(n4642), .Z(n6035) );
  BUF_X1 U601 ( .A(n4642), .Z(n6036) );
  BUF_X1 U602 ( .A(n4653), .Z(n6038) );
  BUF_X1 U603 ( .A(n4653), .Z(n6039) );
  BUF_X1 U604 ( .A(n4637), .Z(n6041) );
  BUF_X1 U605 ( .A(n4637), .Z(n6042) );
  BUF_X1 U606 ( .A(n4658), .Z(n6044) );
  BUF_X1 U607 ( .A(n4658), .Z(n6045) );
  BUF_X1 U608 ( .A(n4638), .Z(n6047) );
  BUF_X1 U609 ( .A(n4638), .Z(n6048) );
  BUF_X1 U610 ( .A(n4654), .Z(n6050) );
  BUF_X1 U611 ( .A(n4654), .Z(n6051) );
  BUF_X1 U612 ( .A(n4655), .Z(n6241) );
  BUF_X1 U613 ( .A(n4655), .Z(n6242) );
  BUF_X1 U614 ( .A(n4656), .Z(n6244) );
  BUF_X1 U615 ( .A(n4656), .Z(n6245) );
  BUF_X1 U616 ( .A(n4639), .Z(n6247) );
  BUF_X1 U617 ( .A(n4639), .Z(n6248) );
  BUF_X1 U618 ( .A(n4640), .Z(n6250) );
  BUF_X1 U619 ( .A(n4640), .Z(n6251) );
  BUF_X1 U620 ( .A(n4647), .Z(n6253) );
  BUF_X1 U621 ( .A(n4647), .Z(n6254) );
  BUF_X1 U622 ( .A(n4648), .Z(n6256) );
  BUF_X1 U623 ( .A(n4648), .Z(n6257) );
  BUF_X1 U624 ( .A(n4649), .Z(n6259) );
  BUF_X1 U625 ( .A(n4649), .Z(n6260) );
  BUF_X1 U626 ( .A(n4635), .Z(n6262) );
  BUF_X1 U627 ( .A(n4635), .Z(n6263) );
  BUF_X1 U628 ( .A(n7552), .Z(n6238) );
  BUF_X1 U629 ( .A(n7552), .Z(n6239) );
  BUF_X1 U630 ( .A(n4643), .Z(n6010) );
  BUF_X1 U631 ( .A(n4644), .Z(n6013) );
  BUF_X1 U632 ( .A(n4651), .Z(n6019) );
  BUF_X1 U633 ( .A(n4636), .Z(n6022) );
  BUF_X1 U634 ( .A(n4645), .Z(n6025) );
  BUF_X1 U635 ( .A(n4646), .Z(n6028) );
  BUF_X1 U636 ( .A(n4652), .Z(n6031) );
  BUF_X1 U637 ( .A(n4642), .Z(n6037) );
  BUF_X1 U638 ( .A(n4653), .Z(n6040) );
  BUF_X1 U639 ( .A(n4637), .Z(n6043) );
  BUF_X1 U640 ( .A(n4658), .Z(n6046) );
  BUF_X1 U641 ( .A(n4638), .Z(n6049) );
  BUF_X1 U642 ( .A(n4654), .Z(n6052) );
  BUF_X1 U643 ( .A(n4655), .Z(n6243) );
  BUF_X1 U644 ( .A(n4656), .Z(n6246) );
  BUF_X1 U645 ( .A(n4639), .Z(n6249) );
  BUF_X1 U646 ( .A(n4640), .Z(n6252) );
  BUF_X1 U647 ( .A(n4647), .Z(n6255) );
  BUF_X1 U648 ( .A(n4648), .Z(n6258) );
  BUF_X1 U649 ( .A(n4649), .Z(n6261) );
  BUF_X1 U650 ( .A(n4635), .Z(n6264) );
  BUF_X1 U651 ( .A(n7552), .Z(n6240) );
  INV_X1 U652 ( .A(ADD_RS1[2]), .ZN(n7900) );
  INV_X1 U653 ( .A(ADD_RS2[2]), .ZN(n7898) );
  BUF_X1 U654 ( .A(n7542), .Z(n6232) );
  BUF_X1 U655 ( .A(n7542), .Z(n6233) );
  BUF_X1 U656 ( .A(n6493), .Z(n6107) );
  BUF_X1 U657 ( .A(n6486), .Z(n6053) );
  BUF_X1 U658 ( .A(n6487), .Z(n6062) );
  BUF_X1 U659 ( .A(n6490), .Z(n6080) );
  BUF_X1 U660 ( .A(n6492), .Z(n6098) );
  BUF_X1 U661 ( .A(RST), .Z(n6380) );
  BUF_X1 U662 ( .A(n6493), .Z(n6108) );
  BUF_X1 U663 ( .A(n6486), .Z(n6054) );
  BUF_X1 U664 ( .A(n6487), .Z(n6063) );
  BUF_X1 U665 ( .A(n6490), .Z(n6081) );
  BUF_X1 U666 ( .A(n6492), .Z(n6099) );
  BUF_X1 U667 ( .A(RST), .Z(n6381) );
  NOR4_X1 U668 ( .A1(n7902), .A2(n1400), .A3(n1401), .A4(n1402), .ZN(n1399) );
  XNOR2_X1 U669 ( .A(n7590), .B(ADD_RS1[3]), .ZN(n2001) );
  XNOR2_X1 U670 ( .A(n7589), .B(ADD_RS1[4]), .ZN(n2000) );
  XNOR2_X1 U671 ( .A(ADD_RS2[2]), .B(n7591), .ZN(n1402) );
  XNOR2_X1 U672 ( .A(n7589), .B(ADD_RS2[4]), .ZN(n1400) );
  XNOR2_X1 U673 ( .A(n7590), .B(ADD_RS2[3]), .ZN(n1401) );
  XNOR2_X1 U674 ( .A(ADD_RS1[2]), .B(n7591), .ZN(n2002) );
  BUF_X1 U675 ( .A(n4660), .Z(n6173) );
  BUF_X1 U676 ( .A(n4660), .Z(n6174) );
  AOI21_X1 U677 ( .B1(n6931), .B2(n6930), .A(n6929), .ZN(n7542) );
  AND2_X1 U678 ( .A1(n1397), .A2(n1427), .ZN(n6931) );
  NOR2_X1 U679 ( .A1(n1402), .A2(n6928), .ZN(n6930) );
  NOR3_X1 U680 ( .A1(n1401), .A2(n7902), .A3(n1400), .ZN(n1427) );
  BUF_X1 U681 ( .A(n4660), .Z(n6175) );
  NOR4_X1 U682 ( .A1(n7902), .A2(n2000), .A3(n2001), .A4(n2002), .ZN(n1999) );
  NOR3_X1 U683 ( .A1(n2001), .A2(n7902), .A3(n2000), .ZN(n2027) );
  INV_X1 U684 ( .A(n1398), .ZN(n6928) );
  AOI221_X1 U685 ( .B1(n6275), .B2(n7655), .C1(n6271), .C2(n7867), .A(n1981), 
        .ZN(n1974) );
  AOI221_X1 U686 ( .B1(n6275), .B2(n7654), .C1(n6271), .C2(n7866), .A(n1964), 
        .ZN(n1957) );
  AOI221_X1 U687 ( .B1(n6275), .B2(n7653), .C1(n6271), .C2(n7865), .A(n1947), 
        .ZN(n1940) );
  AOI221_X1 U688 ( .B1(n6275), .B2(n7652), .C1(n6271), .C2(n7864), .A(n1930), 
        .ZN(n1923) );
  AOI221_X1 U689 ( .B1(n6275), .B2(n7651), .C1(n6271), .C2(n7863), .A(n1913), 
        .ZN(n1906) );
  AOI221_X1 U690 ( .B1(n6275), .B2(n7650), .C1(n6271), .C2(n7862), .A(n1896), 
        .ZN(n1889) );
  AOI221_X1 U691 ( .B1(n6275), .B2(n7649), .C1(n6271), .C2(n7861), .A(n1879), 
        .ZN(n1872) );
  AOI221_X1 U692 ( .B1(n6274), .B2(n7648), .C1(n6271), .C2(n7860), .A(n1862), 
        .ZN(n1855) );
  AOI221_X1 U693 ( .B1(n6274), .B2(n7647), .C1(n6271), .C2(n7859), .A(n1845), 
        .ZN(n1838) );
  AOI221_X1 U694 ( .B1(n6274), .B2(n7646), .C1(n6271), .C2(n7858), .A(n1828), 
        .ZN(n1821) );
  AOI221_X1 U695 ( .B1(n6274), .B2(n7645), .C1(n6271), .C2(n7857), .A(n1811), 
        .ZN(n1804) );
  AOI221_X1 U696 ( .B1(n6274), .B2(n7644), .C1(n6271), .C2(n7856), .A(n1794), 
        .ZN(n1787) );
  AOI221_X1 U697 ( .B1(n6274), .B2(n7643), .C1(n6272), .C2(n7855), .A(n1777), 
        .ZN(n1770) );
  AOI221_X1 U698 ( .B1(n6274), .B2(n7642), .C1(n6272), .C2(n7854), .A(n1760), 
        .ZN(n1753) );
  AOI221_X1 U699 ( .B1(n6274), .B2(n7641), .C1(n6272), .C2(n7853), .A(n1743), 
        .ZN(n1736) );
  AOI221_X1 U700 ( .B1(n6274), .B2(n7640), .C1(n6272), .C2(n7852), .A(n1726), 
        .ZN(n1719) );
  AOI221_X1 U701 ( .B1(n6274), .B2(n7639), .C1(n6272), .C2(n7851), .A(n1709), 
        .ZN(n1702) );
  AOI221_X1 U702 ( .B1(n6274), .B2(n7638), .C1(n6272), .C2(n7850), .A(n1692), 
        .ZN(n1685) );
  AOI221_X1 U703 ( .B1(n6274), .B2(n7637), .C1(n6272), .C2(n7849), .A(n1675), 
        .ZN(n1668) );
  AOI221_X1 U704 ( .B1(n6273), .B2(n7636), .C1(n6272), .C2(n7848), .A(n1658), 
        .ZN(n1651) );
  AOI221_X1 U705 ( .B1(n6273), .B2(n7635), .C1(n6272), .C2(n7847), .A(n1641), 
        .ZN(n1634) );
  AOI221_X1 U706 ( .B1(n6273), .B2(n7634), .C1(n6272), .C2(n7846), .A(n1624), 
        .ZN(n1617) );
  AOI221_X1 U707 ( .B1(n6273), .B2(n7633), .C1(n6272), .C2(n7845), .A(n1607), 
        .ZN(n1600) );
  AOI221_X1 U708 ( .B1(n6273), .B2(n7632), .C1(n6272), .C2(n7844), .A(n1590), 
        .ZN(n1583) );
  AOI221_X1 U709 ( .B1(n6273), .B2(n7631), .C1(n6271), .C2(n7843), .A(n1573), 
        .ZN(n1566) );
  AOI221_X1 U710 ( .B1(n6273), .B2(n7630), .C1(n6272), .C2(n7842), .A(n1556), 
        .ZN(n1549) );
  AOI221_X1 U711 ( .B1(n6273), .B2(n7629), .C1(n6271), .C2(n7841), .A(n1539), 
        .ZN(n1532) );
  AOI221_X1 U712 ( .B1(n6273), .B2(n7628), .C1(n6272), .C2(n7840), .A(n1522), 
        .ZN(n1515) );
  AOI221_X1 U713 ( .B1(n6273), .B2(n7627), .C1(n6271), .C2(n7839), .A(n1505), 
        .ZN(n1498) );
  AOI221_X1 U714 ( .B1(n6273), .B2(n7626), .C1(n6272), .C2(n7838), .A(n1488), 
        .ZN(n1481) );
  AOI221_X1 U715 ( .B1(n6273), .B2(n7587), .C1(n6271), .C2(n5103), .A(n1460), 
        .ZN(n1437) );
  AOI221_X1 U716 ( .B1(n6310), .B2(n7588), .C1(n6309), .C2(n5104), .A(n847), 
        .ZN(n824) );
  AOI221_X1 U717 ( .B1(n6310), .B2(n7655), .C1(n6308), .C2(n7867), .A(n878), 
        .ZN(n871) );
  AOI221_X1 U718 ( .B1(n6310), .B2(n7654), .C1(n6309), .C2(n7866), .A(n895), 
        .ZN(n888) );
  AOI221_X1 U719 ( .B1(n6310), .B2(n7653), .C1(n6308), .C2(n7865), .A(n912), 
        .ZN(n905) );
  AOI221_X1 U720 ( .B1(n6310), .B2(n7652), .C1(n6309), .C2(n7864), .A(n929), 
        .ZN(n922) );
  AOI221_X1 U721 ( .B1(n6310), .B2(n7651), .C1(n6308), .C2(n7863), .A(n948), 
        .ZN(n941) );
  AOI221_X1 U722 ( .B1(n6310), .B2(n7650), .C1(n6309), .C2(n7862), .A(n969), 
        .ZN(n961) );
  AOI221_X1 U723 ( .B1(n6310), .B2(n7649), .C1(n6309), .C2(n7861), .A(n991), 
        .ZN(n981) );
  AOI221_X1 U724 ( .B1(n6310), .B2(n7648), .C1(n6309), .C2(n7860), .A(n1009), 
        .ZN(n1002) );
  AOI221_X1 U725 ( .B1(n6310), .B2(n7647), .C1(n6309), .C2(n7859), .A(n1026), 
        .ZN(n1019) );
  AOI221_X1 U726 ( .B1(n6310), .B2(n7646), .C1(n6309), .C2(n7858), .A(n1043), 
        .ZN(n1036) );
  AOI221_X1 U727 ( .B1(n6310), .B2(n7645), .C1(n6309), .C2(n7857), .A(n1060), 
        .ZN(n1053) );
  AOI221_X1 U728 ( .B1(n6311), .B2(n7644), .C1(n6309), .C2(n7856), .A(n1077), 
        .ZN(n1070) );
  AOI221_X1 U729 ( .B1(n6311), .B2(n7643), .C1(n6309), .C2(n7855), .A(n1094), 
        .ZN(n1087) );
  AOI221_X1 U730 ( .B1(n6311), .B2(n7642), .C1(n6309), .C2(n7854), .A(n1111), 
        .ZN(n1104) );
  AOI221_X1 U731 ( .B1(n6311), .B2(n7641), .C1(n6309), .C2(n7853), .A(n1128), 
        .ZN(n1121) );
  AOI221_X1 U732 ( .B1(n6311), .B2(n7640), .C1(n6309), .C2(n7852), .A(n1145), 
        .ZN(n1138) );
  AOI221_X1 U733 ( .B1(n6311), .B2(n7639), .C1(n6309), .C2(n7851), .A(n1162), 
        .ZN(n1155) );
  AOI221_X1 U734 ( .B1(n6311), .B2(n7638), .C1(n6309), .C2(n7850), .A(n1179), 
        .ZN(n1172) );
  AOI221_X1 U735 ( .B1(n6311), .B2(n7637), .C1(n6308), .C2(n7849), .A(n1196), 
        .ZN(n1189) );
  AOI221_X1 U736 ( .B1(n6311), .B2(n7636), .C1(n6308), .C2(n7848), .A(n1213), 
        .ZN(n1206) );
  AOI221_X1 U737 ( .B1(n6311), .B2(n7635), .C1(n6308), .C2(n7847), .A(n1230), 
        .ZN(n1223) );
  AOI221_X1 U738 ( .B1(n6311), .B2(n7634), .C1(n6308), .C2(n7846), .A(n1247), 
        .ZN(n1240) );
  AOI221_X1 U739 ( .B1(n6311), .B2(n7633), .C1(n6308), .C2(n7845), .A(n1264), 
        .ZN(n1257) );
  AOI221_X1 U740 ( .B1(n6312), .B2(n7632), .C1(n6308), .C2(n7844), .A(n1281), 
        .ZN(n1274) );
  AOI221_X1 U741 ( .B1(n6312), .B2(n7631), .C1(n6308), .C2(n7843), .A(n1298), 
        .ZN(n1291) );
  AOI221_X1 U742 ( .B1(n6312), .B2(n7630), .C1(n6308), .C2(n7842), .A(n1315), 
        .ZN(n1308) );
  AOI221_X1 U743 ( .B1(n6312), .B2(n7629), .C1(n6308), .C2(n7841), .A(n1332), 
        .ZN(n1325) );
  AOI221_X1 U744 ( .B1(n6312), .B2(n7628), .C1(n6308), .C2(n7840), .A(n1349), 
        .ZN(n1342) );
  AOI221_X1 U745 ( .B1(n6312), .B2(n7627), .C1(n6308), .C2(n7839), .A(n1366), 
        .ZN(n1359) );
  AOI221_X1 U746 ( .B1(n6312), .B2(n7626), .C1(n6308), .C2(n7838), .A(n1383), 
        .ZN(n1376) );
  AOI221_X1 U747 ( .B1(n6288), .B2(n7897), .C1(n6287), .C2(n7625), .A(n1980), 
        .ZN(n1975) );
  AOI221_X1 U748 ( .B1(n6288), .B2(n7896), .C1(n6287), .C2(n7624), .A(n1963), 
        .ZN(n1958) );
  AOI221_X1 U749 ( .B1(n6288), .B2(n7895), .C1(n6287), .C2(n7623), .A(n1946), 
        .ZN(n1941) );
  AOI221_X1 U750 ( .B1(n6288), .B2(n7894), .C1(n6287), .C2(n7622), .A(n1929), 
        .ZN(n1924) );
  AOI221_X1 U751 ( .B1(n6288), .B2(n7893), .C1(n6287), .C2(n7621), .A(n1912), 
        .ZN(n1907) );
  AOI221_X1 U752 ( .B1(n6288), .B2(n7892), .C1(n6287), .C2(n7620), .A(n1895), 
        .ZN(n1890) );
  AOI221_X1 U753 ( .B1(n6288), .B2(n7891), .C1(n6287), .C2(n7619), .A(n1878), 
        .ZN(n1873) );
  AOI221_X1 U754 ( .B1(n6288), .B2(n7890), .C1(n6286), .C2(n7618), .A(n1861), 
        .ZN(n1856) );
  AOI221_X1 U755 ( .B1(n6288), .B2(n7889), .C1(n6286), .C2(n7617), .A(n1844), 
        .ZN(n1839) );
  AOI221_X1 U756 ( .B1(n6288), .B2(n7888), .C1(n6286), .C2(n7616), .A(n1827), 
        .ZN(n1822) );
  AOI221_X1 U757 ( .B1(n6288), .B2(n7887), .C1(n6286), .C2(n7615), .A(n1810), 
        .ZN(n1805) );
  AOI221_X1 U758 ( .B1(n6288), .B2(n7886), .C1(n6286), .C2(n7614), .A(n1793), 
        .ZN(n1788) );
  AOI221_X1 U759 ( .B1(n6289), .B2(n7885), .C1(n6286), .C2(n7613), .A(n1776), 
        .ZN(n1771) );
  AOI221_X1 U760 ( .B1(n6289), .B2(n7884), .C1(n6286), .C2(n7612), .A(n1759), 
        .ZN(n1754) );
  AOI221_X1 U761 ( .B1(n6289), .B2(n7883), .C1(n6286), .C2(n7611), .A(n1742), 
        .ZN(n1737) );
  AOI221_X1 U762 ( .B1(n6289), .B2(n7882), .C1(n6286), .C2(n7610), .A(n1725), 
        .ZN(n1720) );
  AOI221_X1 U763 ( .B1(n6289), .B2(n7881), .C1(n6286), .C2(n7609), .A(n1708), 
        .ZN(n1703) );
  AOI221_X1 U764 ( .B1(n6289), .B2(n7880), .C1(n6286), .C2(n7608), .A(n1691), 
        .ZN(n1686) );
  AOI221_X1 U765 ( .B1(n6289), .B2(n7879), .C1(n6286), .C2(n7607), .A(n1674), 
        .ZN(n1669) );
  AOI221_X1 U766 ( .B1(n6289), .B2(n7878), .C1(n6285), .C2(n7606), .A(n1657), 
        .ZN(n1652) );
  AOI221_X1 U767 ( .B1(n6289), .B2(n7877), .C1(n6285), .C2(n7605), .A(n1640), 
        .ZN(n1635) );
  AOI221_X1 U768 ( .B1(n6289), .B2(n7876), .C1(n6285), .C2(n7604), .A(n1623), 
        .ZN(n1618) );
  AOI221_X1 U769 ( .B1(n6289), .B2(n7875), .C1(n6285), .C2(n7603), .A(n1606), 
        .ZN(n1601) );
  AOI221_X1 U770 ( .B1(n6289), .B2(n7874), .C1(n6285), .C2(n7602), .A(n1589), 
        .ZN(n1584) );
  AOI221_X1 U771 ( .B1(n6288), .B2(n7873), .C1(n6285), .C2(n7601), .A(n1572), 
        .ZN(n1567) );
  AOI221_X1 U772 ( .B1(n6289), .B2(n7872), .C1(n6285), .C2(n7600), .A(n1555), 
        .ZN(n1550) );
  AOI221_X1 U773 ( .B1(n6288), .B2(n7871), .C1(n6285), .C2(n7599), .A(n1538), 
        .ZN(n1533) );
  AOI221_X1 U774 ( .B1(n6289), .B2(n7870), .C1(n6285), .C2(n7598), .A(n1521), 
        .ZN(n1516) );
  AOI221_X1 U775 ( .B1(n6288), .B2(n7869), .C1(n6285), .C2(n7597), .A(n1504), 
        .ZN(n1499) );
  AOI221_X1 U776 ( .B1(n6289), .B2(n7868), .C1(n6285), .C2(n7596), .A(n1487), 
        .ZN(n1482) );
  AOI221_X1 U777 ( .B1(n6288), .B2(n5101), .C1(n6285), .C2(n7585), .A(n1454), 
        .ZN(n1438) );
  AOI221_X1 U778 ( .B1(n6326), .B2(n5102), .C1(n6322), .C2(n7586), .A(n841), 
        .ZN(n825) );
  AOI221_X1 U779 ( .B1(n6325), .B2(n7897), .C1(n6322), .C2(n7625), .A(n877), 
        .ZN(n872) );
  AOI221_X1 U780 ( .B1(n6326), .B2(n7896), .C1(n6322), .C2(n7624), .A(n894), 
        .ZN(n889) );
  AOI221_X1 U781 ( .B1(n6325), .B2(n7895), .C1(n6322), .C2(n7623), .A(n911), 
        .ZN(n906) );
  AOI221_X1 U782 ( .B1(n6326), .B2(n7894), .C1(n6322), .C2(n7622), .A(n928), 
        .ZN(n923) );
  AOI221_X1 U783 ( .B1(n6325), .B2(n7893), .C1(n6322), .C2(n7621), .A(n947), 
        .ZN(n942) );
  AOI221_X1 U784 ( .B1(n6326), .B2(n7892), .C1(n6322), .C2(n7620), .A(n968), 
        .ZN(n962) );
  AOI221_X1 U785 ( .B1(n6326), .B2(n7891), .C1(n6322), .C2(n7619), .A(n990), 
        .ZN(n983) );
  AOI221_X1 U786 ( .B1(n6326), .B2(n7890), .C1(n6322), .C2(n7618), .A(n1008), 
        .ZN(n1003) );
  AOI221_X1 U787 ( .B1(n6326), .B2(n7889), .C1(n6322), .C2(n7617), .A(n1025), 
        .ZN(n1020) );
  AOI221_X1 U788 ( .B1(n6326), .B2(n7888), .C1(n6322), .C2(n7616), .A(n1042), 
        .ZN(n1037) );
  AOI221_X1 U789 ( .B1(n6326), .B2(n7887), .C1(n6322), .C2(n7615), .A(n1059), 
        .ZN(n1054) );
  AOI221_X1 U790 ( .B1(n6326), .B2(n7886), .C1(n6323), .C2(n7614), .A(n1076), 
        .ZN(n1071) );
  AOI221_X1 U791 ( .B1(n6326), .B2(n7885), .C1(n6323), .C2(n7613), .A(n1093), 
        .ZN(n1088) );
  AOI221_X1 U792 ( .B1(n6326), .B2(n7884), .C1(n6323), .C2(n7612), .A(n1110), 
        .ZN(n1105) );
  AOI221_X1 U793 ( .B1(n6326), .B2(n7883), .C1(n6323), .C2(n7611), .A(n1127), 
        .ZN(n1122) );
  AOI221_X1 U794 ( .B1(n6326), .B2(n7882), .C1(n6323), .C2(n7610), .A(n1144), 
        .ZN(n1139) );
  AOI221_X1 U795 ( .B1(n6326), .B2(n7881), .C1(n6323), .C2(n7609), .A(n1161), 
        .ZN(n1156) );
  AOI221_X1 U796 ( .B1(n6326), .B2(n7880), .C1(n6323), .C2(n7608), .A(n1178), 
        .ZN(n1173) );
  AOI221_X1 U797 ( .B1(n6325), .B2(n7879), .C1(n6323), .C2(n7607), .A(n1195), 
        .ZN(n1190) );
  AOI221_X1 U798 ( .B1(n6325), .B2(n7878), .C1(n6323), .C2(n7606), .A(n1212), 
        .ZN(n1207) );
  AOI221_X1 U799 ( .B1(n6325), .B2(n7877), .C1(n6323), .C2(n7605), .A(n1229), 
        .ZN(n1224) );
  AOI221_X1 U800 ( .B1(n6325), .B2(n7876), .C1(n6323), .C2(n7604), .A(n1246), 
        .ZN(n1241) );
  AOI221_X1 U801 ( .B1(n6325), .B2(n7875), .C1(n6323), .C2(n7603), .A(n1263), 
        .ZN(n1258) );
  AOI221_X1 U802 ( .B1(n6325), .B2(n7874), .C1(n6324), .C2(n7602), .A(n1280), 
        .ZN(n1275) );
  AOI221_X1 U803 ( .B1(n6325), .B2(n7873), .C1(n6324), .C2(n7601), .A(n1297), 
        .ZN(n1292) );
  AOI221_X1 U804 ( .B1(n6325), .B2(n7872), .C1(n6324), .C2(n7600), .A(n1314), 
        .ZN(n1309) );
  AOI221_X1 U805 ( .B1(n6325), .B2(n7871), .C1(n6324), .C2(n7599), .A(n1331), 
        .ZN(n1326) );
  AOI221_X1 U806 ( .B1(n6325), .B2(n7870), .C1(n6324), .C2(n7598), .A(n1348), 
        .ZN(n1343) );
  AOI221_X1 U807 ( .B1(n6325), .B2(n7869), .C1(n6324), .C2(n7597), .A(n1365), 
        .ZN(n1360) );
  AOI221_X1 U808 ( .B1(n6325), .B2(n7868), .C1(n6324), .C2(n7596), .A(n1382), 
        .ZN(n1377) );
  XNOR2_X1 U809 ( .A(ADD_RS2[1]), .B(ADD_WR[1]), .ZN(n1398) );
  XNOR2_X1 U810 ( .A(ADD_RS1[0]), .B(ADD_WR[0]), .ZN(n1997) );
  XNOR2_X1 U811 ( .A(ADD_RS1[1]), .B(ADD_WR[1]), .ZN(n1998) );
  INV_X1 U812 ( .A(WR), .ZN(n7902) );
  XNOR2_X1 U813 ( .A(ADD_RS2[0]), .B(ADD_WR[0]), .ZN(n1397) );
  AOI221_X1 U814 ( .B1(n6299), .B2(n4061), .C1(n6296), .C2(n4093), .A(n1449), 
        .ZN(n1439) );
  AOI221_X1 U815 ( .B1(n6336), .B2(n4030), .C1(n6333), .C2(n4062), .A(n836), 
        .ZN(n826) );
  INV_X1 U816 ( .A(DATAIN[31]), .ZN(n6374) );
  INV_X1 U817 ( .A(DATAIN[4]), .ZN(n6347) );
  INV_X1 U818 ( .A(DATAIN[5]), .ZN(n6348) );
  INV_X1 U819 ( .A(DATAIN[6]), .ZN(n6349) );
  INV_X1 U820 ( .A(DATAIN[7]), .ZN(n6350) );
  INV_X1 U821 ( .A(DATAIN[8]), .ZN(n6351) );
  INV_X1 U822 ( .A(DATAIN[9]), .ZN(n6352) );
  INV_X1 U823 ( .A(DATAIN[10]), .ZN(n6353) );
  INV_X1 U824 ( .A(DATAIN[11]), .ZN(n6354) );
  INV_X1 U825 ( .A(DATAIN[12]), .ZN(n6355) );
  INV_X1 U826 ( .A(DATAIN[13]), .ZN(n6356) );
  INV_X1 U827 ( .A(DATAIN[14]), .ZN(n6357) );
  INV_X1 U828 ( .A(DATAIN[15]), .ZN(n6358) );
  INV_X1 U829 ( .A(DATAIN[16]), .ZN(n6359) );
  INV_X1 U830 ( .A(DATAIN[17]), .ZN(n6360) );
  INV_X1 U831 ( .A(DATAIN[18]), .ZN(n6361) );
  INV_X1 U832 ( .A(DATAIN[19]), .ZN(n6362) );
  INV_X1 U833 ( .A(DATAIN[20]), .ZN(n6363) );
  INV_X1 U834 ( .A(DATAIN[21]), .ZN(n6364) );
  INV_X1 U835 ( .A(DATAIN[22]), .ZN(n6365) );
  INV_X1 U836 ( .A(DATAIN[23]), .ZN(n6366) );
  INV_X1 U837 ( .A(DATAIN[24]), .ZN(n6367) );
  INV_X1 U838 ( .A(DATAIN[25]), .ZN(n6368) );
  INV_X1 U839 ( .A(DATAIN[26]), .ZN(n6369) );
  INV_X1 U840 ( .A(DATAIN[27]), .ZN(n6370) );
  INV_X1 U841 ( .A(DATAIN[28]), .ZN(n6371) );
  INV_X1 U842 ( .A(DATAIN[29]), .ZN(n6372) );
  INV_X1 U843 ( .A(DATAIN[30]), .ZN(n6373) );
  INV_X1 U844 ( .A(n2285), .ZN(n7867) );
  INV_X1 U845 ( .A(n2436), .ZN(n7625) );
  INV_X1 U846 ( .A(n2286), .ZN(n7866) );
  INV_X1 U847 ( .A(n2432), .ZN(n7624) );
  INV_X1 U848 ( .A(n2287), .ZN(n7865) );
  INV_X1 U849 ( .A(n2428), .ZN(n7623) );
  INV_X1 U850 ( .A(n2288), .ZN(n7864) );
  INV_X1 U851 ( .A(n2424), .ZN(n7622) );
  INV_X1 U852 ( .A(n2289), .ZN(n7863) );
  INV_X1 U853 ( .A(n2420), .ZN(n7621) );
  INV_X1 U854 ( .A(n2290), .ZN(n7862) );
  INV_X1 U855 ( .A(n2416), .ZN(n7620) );
  INV_X1 U856 ( .A(n2291), .ZN(n7861) );
  INV_X1 U857 ( .A(n2412), .ZN(n7619) );
  INV_X1 U858 ( .A(n2292), .ZN(n7860) );
  INV_X1 U859 ( .A(n2408), .ZN(n7618) );
  INV_X1 U860 ( .A(n2293), .ZN(n7859) );
  INV_X1 U861 ( .A(n2404), .ZN(n7617) );
  INV_X1 U862 ( .A(n2294), .ZN(n7858) );
  INV_X1 U863 ( .A(n2400), .ZN(n7616) );
  INV_X1 U864 ( .A(n2295), .ZN(n7857) );
  INV_X1 U865 ( .A(n2396), .ZN(n7615) );
  INV_X1 U866 ( .A(n2296), .ZN(n7856) );
  INV_X1 U867 ( .A(n2392), .ZN(n7614) );
  INV_X1 U868 ( .A(n2297), .ZN(n7855) );
  INV_X1 U869 ( .A(n2388), .ZN(n7613) );
  INV_X1 U870 ( .A(n2298), .ZN(n7854) );
  INV_X1 U871 ( .A(n2384), .ZN(n7612) );
  INV_X1 U872 ( .A(n2299), .ZN(n7853) );
  INV_X1 U873 ( .A(n2380), .ZN(n7611) );
  INV_X1 U874 ( .A(n2300), .ZN(n7852) );
  INV_X1 U875 ( .A(n2376), .ZN(n7610) );
  INV_X1 U876 ( .A(n2301), .ZN(n7851) );
  INV_X1 U877 ( .A(n2372), .ZN(n7609) );
  INV_X1 U878 ( .A(n2302), .ZN(n7850) );
  INV_X1 U879 ( .A(n2368), .ZN(n7608) );
  INV_X1 U880 ( .A(n2303), .ZN(n7849) );
  INV_X1 U881 ( .A(n2364), .ZN(n7607) );
  INV_X1 U882 ( .A(n2304), .ZN(n7848) );
  INV_X1 U883 ( .A(n2360), .ZN(n7606) );
  INV_X1 U884 ( .A(n2305), .ZN(n7847) );
  INV_X1 U885 ( .A(n2356), .ZN(n7605) );
  INV_X1 U886 ( .A(n2306), .ZN(n7846) );
  INV_X1 U887 ( .A(n2352), .ZN(n7604) );
  INV_X1 U888 ( .A(n2307), .ZN(n7845) );
  INV_X1 U889 ( .A(n2348), .ZN(n7603) );
  INV_X1 U890 ( .A(n2308), .ZN(n7844) );
  INV_X1 U891 ( .A(n2344), .ZN(n7602) );
  INV_X1 U892 ( .A(n2309), .ZN(n7843) );
  INV_X1 U893 ( .A(n2340), .ZN(n7601) );
  INV_X1 U894 ( .A(n2310), .ZN(n7842) );
  INV_X1 U895 ( .A(n2336), .ZN(n7600) );
  INV_X1 U896 ( .A(n2311), .ZN(n7841) );
  INV_X1 U897 ( .A(n2332), .ZN(n7599) );
  INV_X1 U898 ( .A(n2312), .ZN(n7840) );
  INV_X1 U899 ( .A(n2328), .ZN(n7598) );
  INV_X1 U900 ( .A(n2313), .ZN(n7839) );
  INV_X1 U901 ( .A(n2324), .ZN(n7597) );
  INV_X1 U902 ( .A(n2314), .ZN(n7838) );
  INV_X1 U903 ( .A(n2320), .ZN(n7596) );
  INV_X1 U904 ( .A(n2029), .ZN(n7655) );
  INV_X1 U905 ( .A(n3743), .ZN(n7897) );
  INV_X1 U906 ( .A(n2030), .ZN(n7654) );
  INV_X1 U907 ( .A(n3744), .ZN(n7896) );
  INV_X1 U908 ( .A(n2031), .ZN(n7653) );
  INV_X1 U909 ( .A(n3745), .ZN(n7895) );
  INV_X1 U910 ( .A(n2032), .ZN(n7652) );
  INV_X1 U911 ( .A(n3746), .ZN(n7894) );
  INV_X1 U912 ( .A(n2033), .ZN(n7651) );
  INV_X1 U913 ( .A(n3747), .ZN(n7893) );
  INV_X1 U914 ( .A(n2034), .ZN(n7650) );
  INV_X1 U915 ( .A(n3748), .ZN(n7892) );
  INV_X1 U916 ( .A(n2035), .ZN(n7649) );
  INV_X1 U917 ( .A(n3749), .ZN(n7891) );
  INV_X1 U918 ( .A(n2036), .ZN(n7648) );
  INV_X1 U919 ( .A(n3750), .ZN(n7890) );
  INV_X1 U920 ( .A(n2037), .ZN(n7647) );
  INV_X1 U921 ( .A(n3751), .ZN(n7889) );
  INV_X1 U922 ( .A(n2038), .ZN(n7646) );
  INV_X1 U923 ( .A(n3752), .ZN(n7888) );
  INV_X1 U924 ( .A(n2039), .ZN(n7645) );
  INV_X1 U925 ( .A(n3753), .ZN(n7887) );
  INV_X1 U926 ( .A(n2040), .ZN(n7644) );
  INV_X1 U927 ( .A(n3754), .ZN(n7886) );
  INV_X1 U928 ( .A(n2041), .ZN(n7643) );
  INV_X1 U929 ( .A(n3755), .ZN(n7885) );
  INV_X1 U930 ( .A(n2042), .ZN(n7642) );
  INV_X1 U931 ( .A(n3756), .ZN(n7884) );
  INV_X1 U932 ( .A(n2043), .ZN(n7641) );
  INV_X1 U933 ( .A(n3757), .ZN(n7883) );
  INV_X1 U934 ( .A(n2044), .ZN(n7640) );
  INV_X1 U935 ( .A(n3758), .ZN(n7882) );
  INV_X1 U936 ( .A(n2045), .ZN(n7639) );
  INV_X1 U937 ( .A(n3759), .ZN(n7881) );
  INV_X1 U938 ( .A(n2046), .ZN(n7638) );
  INV_X1 U939 ( .A(n3760), .ZN(n7880) );
  INV_X1 U940 ( .A(n2047), .ZN(n7637) );
  INV_X1 U941 ( .A(n3761), .ZN(n7879) );
  INV_X1 U942 ( .A(n2048), .ZN(n7636) );
  INV_X1 U943 ( .A(n3762), .ZN(n7878) );
  INV_X1 U944 ( .A(n2049), .ZN(n7635) );
  INV_X1 U945 ( .A(n3763), .ZN(n7877) );
  INV_X1 U946 ( .A(n2050), .ZN(n7634) );
  INV_X1 U947 ( .A(n3764), .ZN(n7876) );
  INV_X1 U948 ( .A(n2051), .ZN(n7633) );
  INV_X1 U949 ( .A(n3765), .ZN(n7875) );
  INV_X1 U950 ( .A(n2052), .ZN(n7632) );
  INV_X1 U951 ( .A(n3766), .ZN(n7874) );
  INV_X1 U952 ( .A(n2053), .ZN(n7631) );
  INV_X1 U953 ( .A(n3767), .ZN(n7873) );
  INV_X1 U954 ( .A(n2054), .ZN(n7630) );
  INV_X1 U955 ( .A(n3768), .ZN(n7872) );
  INV_X1 U956 ( .A(n2055), .ZN(n7629) );
  INV_X1 U957 ( .A(n3769), .ZN(n7871) );
  INV_X1 U958 ( .A(n2056), .ZN(n7628) );
  INV_X1 U959 ( .A(n3770), .ZN(n7870) );
  INV_X1 U960 ( .A(n2057), .ZN(n7627) );
  INV_X1 U961 ( .A(n3771), .ZN(n7869) );
  INV_X1 U962 ( .A(n2058), .ZN(n7626) );
  INV_X1 U963 ( .A(n3772), .ZN(n7868) );
  AND2_X1 U964 ( .A1(WR), .A2(ENABLE), .ZN(n749) );
  INV_X1 U965 ( .A(n2220), .ZN(n4911) );
  INV_X1 U966 ( .A(n2060), .ZN(n4912) );
  INV_X1 U967 ( .A(n2282), .ZN(n4913) );
  INV_X1 U968 ( .A(n2281), .ZN(n4914) );
  INV_X1 U969 ( .A(n2280), .ZN(n4915) );
  INV_X1 U970 ( .A(n2279), .ZN(n4916) );
  INV_X1 U971 ( .A(n2278), .ZN(n4917) );
  INV_X1 U972 ( .A(n2277), .ZN(n4918) );
  INV_X1 U973 ( .A(n2276), .ZN(n4919) );
  INV_X1 U974 ( .A(n2275), .ZN(n4920) );
  INV_X1 U975 ( .A(n2274), .ZN(n4921) );
  INV_X1 U976 ( .A(n2273), .ZN(n4922) );
  INV_X1 U977 ( .A(n2272), .ZN(n4923) );
  INV_X1 U978 ( .A(n2271), .ZN(n4924) );
  INV_X1 U979 ( .A(n2270), .ZN(n4925) );
  INV_X1 U980 ( .A(n2269), .ZN(n4926) );
  INV_X1 U981 ( .A(n2268), .ZN(n4927) );
  INV_X1 U982 ( .A(n2267), .ZN(n4928) );
  INV_X1 U983 ( .A(n2266), .ZN(n4929) );
  INV_X1 U984 ( .A(n2265), .ZN(n4930) );
  INV_X1 U985 ( .A(n2264), .ZN(n4931) );
  INV_X1 U986 ( .A(n2263), .ZN(n4932) );
  INV_X1 U987 ( .A(n2262), .ZN(n4933) );
  INV_X1 U988 ( .A(n2261), .ZN(n4934) );
  INV_X1 U989 ( .A(n2260), .ZN(n4935) );
  INV_X1 U990 ( .A(n2259), .ZN(n4936) );
  INV_X1 U991 ( .A(n2258), .ZN(n4937) );
  INV_X1 U992 ( .A(n2257), .ZN(n4938) );
  INV_X1 U993 ( .A(n2256), .ZN(n4939) );
  INV_X1 U994 ( .A(n2255), .ZN(n4940) );
  INV_X1 U995 ( .A(n2254), .ZN(n4941) );
  INV_X1 U996 ( .A(n2253), .ZN(n4942) );
  INV_X1 U997 ( .A(n2717), .ZN(n4943) );
  INV_X1 U998 ( .A(n2716), .ZN(n4944) );
  INV_X1 U999 ( .A(n2715), .ZN(n4945) );
  INV_X1 U1000 ( .A(n2714), .ZN(n4946) );
  INV_X1 U1001 ( .A(n2713), .ZN(n4947) );
  INV_X1 U1002 ( .A(n2712), .ZN(n4948) );
  INV_X1 U1003 ( .A(n2711), .ZN(n4949) );
  INV_X1 U1004 ( .A(n2710), .ZN(n4950) );
  INV_X1 U1005 ( .A(n2709), .ZN(n4951) );
  INV_X1 U1006 ( .A(n2708), .ZN(n4952) );
  INV_X1 U1007 ( .A(n2707), .ZN(n4953) );
  INV_X1 U1008 ( .A(n2706), .ZN(n4954) );
  INV_X1 U1009 ( .A(n2705), .ZN(n4955) );
  INV_X1 U1010 ( .A(n2704), .ZN(n4956) );
  INV_X1 U1011 ( .A(n2703), .ZN(n4957) );
  INV_X1 U1012 ( .A(n2702), .ZN(n4958) );
  INV_X1 U1013 ( .A(n2701), .ZN(n4959) );
  INV_X1 U1014 ( .A(n2700), .ZN(n4960) );
  INV_X1 U1015 ( .A(n2699), .ZN(n4961) );
  INV_X1 U1016 ( .A(n2698), .ZN(n4962) );
  INV_X1 U1017 ( .A(n2697), .ZN(n4963) );
  INV_X1 U1018 ( .A(n2696), .ZN(n4964) );
  INV_X1 U1019 ( .A(n2695), .ZN(n4965) );
  INV_X1 U1020 ( .A(n2694), .ZN(n4966) );
  INV_X1 U1021 ( .A(n2693), .ZN(n4967) );
  INV_X1 U1022 ( .A(n2692), .ZN(n4968) );
  INV_X1 U1023 ( .A(n2691), .ZN(n4969) );
  INV_X1 U1024 ( .A(n2690), .ZN(n4970) );
  INV_X1 U1025 ( .A(n2942), .ZN(n4971) );
  INV_X1 U1026 ( .A(n2718), .ZN(n4972) );
  INV_X1 U1027 ( .A(n2250), .ZN(n4973) );
  INV_X1 U1028 ( .A(n2249), .ZN(n4974) );
  INV_X1 U1029 ( .A(n2248), .ZN(n4975) );
  INV_X1 U1030 ( .A(n2247), .ZN(n4976) );
  INV_X1 U1031 ( .A(n2246), .ZN(n4977) );
  INV_X1 U1032 ( .A(n2245), .ZN(n4978) );
  INV_X1 U1033 ( .A(n2244), .ZN(n4979) );
  INV_X1 U1034 ( .A(n2243), .ZN(n4980) );
  INV_X1 U1035 ( .A(n2242), .ZN(n4981) );
  INV_X1 U1036 ( .A(n2241), .ZN(n4982) );
  INV_X1 U1037 ( .A(n2240), .ZN(n4983) );
  INV_X1 U1038 ( .A(n2239), .ZN(n4984) );
  INV_X1 U1039 ( .A(n2238), .ZN(n4985) );
  INV_X1 U1040 ( .A(n2237), .ZN(n4986) );
  INV_X1 U1041 ( .A(n2236), .ZN(n4987) );
  INV_X1 U1042 ( .A(n2235), .ZN(n4988) );
  INV_X1 U1043 ( .A(n2234), .ZN(n4989) );
  INV_X1 U1044 ( .A(n2233), .ZN(n4990) );
  INV_X1 U1045 ( .A(n2232), .ZN(n4991) );
  INV_X1 U1046 ( .A(n2231), .ZN(n4992) );
  INV_X1 U1047 ( .A(n2230), .ZN(n4993) );
  INV_X1 U1048 ( .A(n2229), .ZN(n4994) );
  INV_X1 U1049 ( .A(n2228), .ZN(n4995) );
  INV_X1 U1050 ( .A(n2227), .ZN(n4996) );
  INV_X1 U1051 ( .A(n2226), .ZN(n4997) );
  INV_X1 U1052 ( .A(n2225), .ZN(n4998) );
  INV_X1 U1053 ( .A(n2224), .ZN(n4999) );
  INV_X1 U1054 ( .A(n2223), .ZN(n5000) );
  INV_X1 U1055 ( .A(n2222), .ZN(n5001) );
  INV_X1 U1056 ( .A(n2221), .ZN(n5002) );
  INV_X1 U1057 ( .A(n2219), .ZN(n5003) );
  INV_X1 U1058 ( .A(n2218), .ZN(n5004) );
  INV_X1 U1059 ( .A(n2217), .ZN(n5005) );
  INV_X1 U1060 ( .A(n2216), .ZN(n5006) );
  INV_X1 U1061 ( .A(n2215), .ZN(n5007) );
  INV_X1 U1062 ( .A(n2214), .ZN(n5008) );
  INV_X1 U1063 ( .A(n2213), .ZN(n5009) );
  INV_X1 U1064 ( .A(n2212), .ZN(n5010) );
  INV_X1 U1065 ( .A(n2211), .ZN(n5011) );
  INV_X1 U1066 ( .A(n2210), .ZN(n5012) );
  INV_X1 U1067 ( .A(n2209), .ZN(n5013) );
  INV_X1 U1068 ( .A(n2208), .ZN(n5014) );
  INV_X1 U1069 ( .A(n2207), .ZN(n5015) );
  INV_X1 U1070 ( .A(n2206), .ZN(n5016) );
  INV_X1 U1071 ( .A(n2205), .ZN(n5017) );
  INV_X1 U1072 ( .A(n2204), .ZN(n5018) );
  INV_X1 U1073 ( .A(n2203), .ZN(n5019) );
  INV_X1 U1074 ( .A(n2202), .ZN(n5020) );
  INV_X1 U1075 ( .A(n2201), .ZN(n5021) );
  INV_X1 U1076 ( .A(n2200), .ZN(n5022) );
  INV_X1 U1077 ( .A(n2199), .ZN(n5023) );
  INV_X1 U1078 ( .A(n2198), .ZN(n5024) );
  INV_X1 U1079 ( .A(n2197), .ZN(n5025) );
  INV_X1 U1080 ( .A(n2196), .ZN(n5026) );
  INV_X1 U1081 ( .A(n2195), .ZN(n5027) );
  INV_X1 U1082 ( .A(n2194), .ZN(n5028) );
  INV_X1 U1083 ( .A(n2193), .ZN(n5029) );
  INV_X1 U1084 ( .A(n2192), .ZN(n5030) );
  INV_X1 U1085 ( .A(n2191), .ZN(n5031) );
  INV_X1 U1086 ( .A(n2190), .ZN(n5032) );
  INV_X1 U1087 ( .A(n2189), .ZN(n5033) );
  INV_X1 U1088 ( .A(n987), .ZN(n5034) );
  INV_X1 U1089 ( .A(n971), .ZN(n5035) );
  INV_X1 U1090 ( .A(n955), .ZN(n5036) );
  INV_X1 U1091 ( .A(n2123), .ZN(n5037) );
  INV_X1 U1092 ( .A(n2122), .ZN(n5038) );
  INV_X1 U1093 ( .A(n2121), .ZN(n5039) );
  INV_X1 U1094 ( .A(n2120), .ZN(n5040) );
  INV_X1 U1095 ( .A(n2119), .ZN(n5041) );
  INV_X1 U1096 ( .A(n2118), .ZN(n5042) );
  INV_X1 U1097 ( .A(n2117), .ZN(n5043) );
  INV_X1 U1098 ( .A(n2116), .ZN(n5044) );
  INV_X1 U1099 ( .A(n2115), .ZN(n5045) );
  INV_X1 U1100 ( .A(n2114), .ZN(n5046) );
  INV_X1 U1101 ( .A(n2113), .ZN(n5047) );
  INV_X1 U1102 ( .A(n2112), .ZN(n5048) );
  INV_X1 U1103 ( .A(n2111), .ZN(n5049) );
  INV_X1 U1104 ( .A(n2110), .ZN(n5050) );
  INV_X1 U1105 ( .A(n2109), .ZN(n5051) );
  INV_X1 U1106 ( .A(n2108), .ZN(n5052) );
  INV_X1 U1107 ( .A(n2107), .ZN(n5053) );
  INV_X1 U1108 ( .A(n2106), .ZN(n5054) );
  INV_X1 U1109 ( .A(n2105), .ZN(n5055) );
  INV_X1 U1110 ( .A(n2104), .ZN(n5056) );
  INV_X1 U1111 ( .A(n2103), .ZN(n5057) );
  INV_X1 U1112 ( .A(n2102), .ZN(n5058) );
  INV_X1 U1113 ( .A(n2101), .ZN(n5059) );
  INV_X1 U1114 ( .A(n2100), .ZN(n5060) );
  INV_X1 U1115 ( .A(n2099), .ZN(n5061) );
  INV_X1 U1116 ( .A(n2098), .ZN(n5062) );
  INV_X1 U1117 ( .A(n2097), .ZN(n5063) );
  INV_X1 U1118 ( .A(n2096), .ZN(n5064) );
  INV_X1 U1119 ( .A(n2095), .ZN(n5065) );
  INV_X1 U1120 ( .A(n2094), .ZN(n5066) );
  INV_X1 U1121 ( .A(n2093), .ZN(n5067) );
  INV_X1 U1122 ( .A(n2092), .ZN(n5068) );
  INV_X1 U1123 ( .A(n3677), .ZN(n5069) );
  INV_X1 U1124 ( .A(n3676), .ZN(n5070) );
  INV_X1 U1125 ( .A(n3675), .ZN(n5071) );
  INV_X1 U1126 ( .A(n3674), .ZN(n5072) );
  INV_X1 U1127 ( .A(n3673), .ZN(n5073) );
  INV_X1 U1128 ( .A(n3672), .ZN(n5074) );
  INV_X1 U1129 ( .A(n3671), .ZN(n5075) );
  INV_X1 U1130 ( .A(n3670), .ZN(n5076) );
  INV_X1 U1131 ( .A(n3669), .ZN(n5077) );
  INV_X1 U1132 ( .A(n3668), .ZN(n5078) );
  INV_X1 U1133 ( .A(n3667), .ZN(n5079) );
  INV_X1 U1134 ( .A(n3666), .ZN(n5080) );
  INV_X1 U1135 ( .A(n3665), .ZN(n5081) );
  INV_X1 U1136 ( .A(n3664), .ZN(n5082) );
  INV_X1 U1137 ( .A(n3663), .ZN(n5083) );
  INV_X1 U1138 ( .A(n3662), .ZN(n5084) );
  INV_X1 U1139 ( .A(n3661), .ZN(n5085) );
  INV_X1 U1140 ( .A(n3660), .ZN(n5086) );
  INV_X1 U1141 ( .A(n3659), .ZN(n5087) );
  INV_X1 U1142 ( .A(n3658), .ZN(n5088) );
  INV_X1 U1143 ( .A(n3657), .ZN(n5089) );
  INV_X1 U1144 ( .A(n3656), .ZN(n5090) );
  INV_X1 U1145 ( .A(n3655), .ZN(n5091) );
  INV_X1 U1146 ( .A(n3654), .ZN(n5092) );
  INV_X1 U1147 ( .A(n3653), .ZN(n5093) );
  INV_X1 U1148 ( .A(n3652), .ZN(n5094) );
  INV_X1 U1149 ( .A(n3651), .ZN(n5095) );
  INV_X1 U1150 ( .A(n3650), .ZN(n5096) );
  INV_X1 U1151 ( .A(n3649), .ZN(n5097) );
  INV_X1 U1152 ( .A(n3648), .ZN(n5098) );
  INV_X1 U1153 ( .A(n3647), .ZN(n5099) );
  INV_X1 U1154 ( .A(n3646), .ZN(n5100) );
  INV_X1 U1155 ( .A(n3773), .ZN(n5101) );
  INV_X1 U1156 ( .A(n3742), .ZN(n5102) );
  INV_X1 U1157 ( .A(n2315), .ZN(n5103) );
  INV_X1 U1158 ( .A(n2284), .ZN(n5104) );
  OAI22_X1 U1159 ( .A1(n4029), .A2(n6305), .B1(n2317), .B2(n6302), .ZN(n1425)
         );
  OAI22_X1 U1160 ( .A1(n4029), .A2(n6270), .B1(n2317), .B2(n6267), .ZN(n1460)
         );
  OAI22_X1 U1161 ( .A1(n4028), .A2(n6305), .B1(n2321), .B2(n6302), .ZN(n1383)
         );
  OAI22_X1 U1162 ( .A1(n4028), .A2(n6270), .B1(n2321), .B2(n6267), .ZN(n1488)
         );
  OAI22_X1 U1163 ( .A1(n4027), .A2(n6305), .B1(n2325), .B2(n6302), .ZN(n1366)
         );
  OAI22_X1 U1164 ( .A1(n4027), .A2(n6270), .B1(n2325), .B2(n6267), .ZN(n1505)
         );
  OAI22_X1 U1165 ( .A1(n4026), .A2(n6305), .B1(n2329), .B2(n6302), .ZN(n1349)
         );
  OAI22_X1 U1166 ( .A1(n4026), .A2(n6270), .B1(n2329), .B2(n6267), .ZN(n1522)
         );
  OAI22_X1 U1167 ( .A1(n4025), .A2(n6305), .B1(n2333), .B2(n6302), .ZN(n1332)
         );
  OAI22_X1 U1168 ( .A1(n4025), .A2(n6270), .B1(n2333), .B2(n6267), .ZN(n1539)
         );
  OAI22_X1 U1169 ( .A1(n4024), .A2(n6305), .B1(n2337), .B2(n6302), .ZN(n1315)
         );
  OAI22_X1 U1170 ( .A1(n4024), .A2(n6270), .B1(n2337), .B2(n6267), .ZN(n1556)
         );
  OAI22_X1 U1171 ( .A1(n4023), .A2(n6305), .B1(n2341), .B2(n6302), .ZN(n1298)
         );
  OAI22_X1 U1172 ( .A1(n4023), .A2(n6270), .B1(n2341), .B2(n6267), .ZN(n1573)
         );
  OAI22_X1 U1173 ( .A1(n4022), .A2(n6305), .B1(n2345), .B2(n6302), .ZN(n1281)
         );
  OAI22_X1 U1174 ( .A1(n4022), .A2(n6270), .B1(n2345), .B2(n6267), .ZN(n1590)
         );
  OAI22_X1 U1175 ( .A1(n4021), .A2(n6305), .B1(n2349), .B2(n6302), .ZN(n1264)
         );
  OAI22_X1 U1176 ( .A1(n4021), .A2(n6269), .B1(n2349), .B2(n6266), .ZN(n1607)
         );
  OAI22_X1 U1177 ( .A1(n4020), .A2(n6305), .B1(n2353), .B2(n6302), .ZN(n1247)
         );
  OAI22_X1 U1178 ( .A1(n4020), .A2(n6269), .B1(n2353), .B2(n6266), .ZN(n1624)
         );
  OAI22_X1 U1179 ( .A1(n4019), .A2(n6305), .B1(n2357), .B2(n6302), .ZN(n1230)
         );
  OAI22_X1 U1180 ( .A1(n4019), .A2(n6269), .B1(n2357), .B2(n6266), .ZN(n1641)
         );
  OAI22_X1 U1181 ( .A1(n4018), .A2(n6305), .B1(n2361), .B2(n6302), .ZN(n1213)
         );
  OAI22_X1 U1182 ( .A1(n4018), .A2(n6269), .B1(n2361), .B2(n6266), .ZN(n1658)
         );
  OAI22_X1 U1183 ( .A1(n4017), .A2(n6306), .B1(n2365), .B2(n6303), .ZN(n1196)
         );
  OAI22_X1 U1184 ( .A1(n4017), .A2(n6269), .B1(n2365), .B2(n6266), .ZN(n1675)
         );
  OAI22_X1 U1185 ( .A1(n4016), .A2(n6306), .B1(n2369), .B2(n6303), .ZN(n1179)
         );
  OAI22_X1 U1186 ( .A1(n4016), .A2(n6269), .B1(n2369), .B2(n6266), .ZN(n1692)
         );
  OAI22_X1 U1187 ( .A1(n4015), .A2(n6306), .B1(n2373), .B2(n6303), .ZN(n1162)
         );
  OAI22_X1 U1188 ( .A1(n4015), .A2(n6269), .B1(n2373), .B2(n6266), .ZN(n1709)
         );
  OAI22_X1 U1189 ( .A1(n4014), .A2(n6306), .B1(n2377), .B2(n6303), .ZN(n1145)
         );
  OAI22_X1 U1190 ( .A1(n4014), .A2(n6269), .B1(n2377), .B2(n6266), .ZN(n1726)
         );
  OAI22_X1 U1191 ( .A1(n4013), .A2(n6306), .B1(n2381), .B2(n6303), .ZN(n1128)
         );
  OAI22_X1 U1192 ( .A1(n4013), .A2(n6269), .B1(n2381), .B2(n6266), .ZN(n1743)
         );
  OAI22_X1 U1193 ( .A1(n4012), .A2(n6306), .B1(n2385), .B2(n6303), .ZN(n1111)
         );
  OAI22_X1 U1194 ( .A1(n4012), .A2(n6269), .B1(n2385), .B2(n6266), .ZN(n1760)
         );
  OAI22_X1 U1195 ( .A1(n4011), .A2(n6306), .B1(n2389), .B2(n6303), .ZN(n1094)
         );
  OAI22_X1 U1196 ( .A1(n4011), .A2(n6269), .B1(n2389), .B2(n6266), .ZN(n1777)
         );
  OAI22_X1 U1197 ( .A1(n4010), .A2(n6306), .B1(n2393), .B2(n6303), .ZN(n1077)
         );
  OAI22_X1 U1198 ( .A1(n4010), .A2(n6269), .B1(n2393), .B2(n6266), .ZN(n1794)
         );
  OAI22_X1 U1199 ( .A1(n4009), .A2(n6306), .B1(n2397), .B2(n6303), .ZN(n1060)
         );
  OAI22_X1 U1200 ( .A1(n4009), .A2(n6268), .B1(n2397), .B2(n6265), .ZN(n1811)
         );
  OAI22_X1 U1201 ( .A1(n4008), .A2(n6306), .B1(n2401), .B2(n6303), .ZN(n1043)
         );
  OAI22_X1 U1202 ( .A1(n4008), .A2(n6268), .B1(n2401), .B2(n6265), .ZN(n1828)
         );
  OAI22_X1 U1203 ( .A1(n4007), .A2(n6306), .B1(n2405), .B2(n6303), .ZN(n1026)
         );
  OAI22_X1 U1204 ( .A1(n4007), .A2(n6268), .B1(n2405), .B2(n6265), .ZN(n1845)
         );
  OAI22_X1 U1205 ( .A1(n4006), .A2(n6306), .B1(n2409), .B2(n6303), .ZN(n1009)
         );
  OAI22_X1 U1206 ( .A1(n4006), .A2(n6268), .B1(n2409), .B2(n6265), .ZN(n1862)
         );
  OAI22_X1 U1207 ( .A1(n4005), .A2(n6307), .B1(n2413), .B2(n6304), .ZN(n991)
         );
  OAI22_X1 U1208 ( .A1(n4005), .A2(n6268), .B1(n2413), .B2(n6265), .ZN(n1879)
         );
  OAI22_X1 U1209 ( .A1(n4004), .A2(n6307), .B1(n2417), .B2(n6304), .ZN(n969)
         );
  OAI22_X1 U1210 ( .A1(n4004), .A2(n6268), .B1(n2417), .B2(n6265), .ZN(n1896)
         );
  OAI22_X1 U1211 ( .A1(n4003), .A2(n6307), .B1(n2421), .B2(n6304), .ZN(n948)
         );
  OAI22_X1 U1212 ( .A1(n4003), .A2(n6268), .B1(n2421), .B2(n6265), .ZN(n1913)
         );
  OAI22_X1 U1213 ( .A1(n4002), .A2(n6307), .B1(n2425), .B2(n6304), .ZN(n929)
         );
  OAI22_X1 U1214 ( .A1(n4002), .A2(n6268), .B1(n2425), .B2(n6265), .ZN(n1930)
         );
  OAI22_X1 U1215 ( .A1(n4001), .A2(n6307), .B1(n2429), .B2(n6304), .ZN(n912)
         );
  OAI22_X1 U1216 ( .A1(n4001), .A2(n6268), .B1(n2429), .B2(n6265), .ZN(n1947)
         );
  OAI22_X1 U1217 ( .A1(n4000), .A2(n6307), .B1(n2433), .B2(n6304), .ZN(n895)
         );
  OAI22_X1 U1218 ( .A1(n4000), .A2(n6268), .B1(n2433), .B2(n6265), .ZN(n1964)
         );
  OAI22_X1 U1219 ( .A1(n3999), .A2(n6307), .B1(n2437), .B2(n6304), .ZN(n878)
         );
  OAI22_X1 U1220 ( .A1(n3999), .A2(n6268), .B1(n2437), .B2(n6265), .ZN(n1981)
         );
  OAI22_X1 U1221 ( .A1(n3998), .A2(n6307), .B1(n2441), .B2(n6304), .ZN(n847)
         );
  OAI22_X1 U1222 ( .A1(n3998), .A2(n6268), .B1(n2441), .B2(n6265), .ZN(n2025)
         );
  OAI22_X1 U1223 ( .A1(n3901), .A2(n6330), .B1(n3933), .B2(n6327), .ZN(n1421)
         );
  OAI22_X1 U1224 ( .A1(n3901), .A2(n6295), .B1(n3933), .B2(n6292), .ZN(n1449)
         );
  OAI22_X1 U1225 ( .A1(n3900), .A2(n6330), .B1(n3932), .B2(n6327), .ZN(n1381)
         );
  OAI22_X1 U1226 ( .A1(n3900), .A2(n6295), .B1(n3932), .B2(n6292), .ZN(n1486)
         );
  OAI22_X1 U1227 ( .A1(n3899), .A2(n6330), .B1(n3931), .B2(n6327), .ZN(n1364)
         );
  OAI22_X1 U1228 ( .A1(n3899), .A2(n6295), .B1(n3931), .B2(n6292), .ZN(n1503)
         );
  OAI22_X1 U1229 ( .A1(n3898), .A2(n6330), .B1(n3930), .B2(n6327), .ZN(n1347)
         );
  OAI22_X1 U1230 ( .A1(n3898), .A2(n6295), .B1(n3930), .B2(n6292), .ZN(n1520)
         );
  OAI22_X1 U1231 ( .A1(n3897), .A2(n6330), .B1(n3929), .B2(n6327), .ZN(n1330)
         );
  OAI22_X1 U1232 ( .A1(n3897), .A2(n6295), .B1(n3929), .B2(n6292), .ZN(n1537)
         );
  OAI22_X1 U1233 ( .A1(n3896), .A2(n6330), .B1(n3928), .B2(n6327), .ZN(n1313)
         );
  OAI22_X1 U1234 ( .A1(n3896), .A2(n6295), .B1(n3928), .B2(n6292), .ZN(n1554)
         );
  OAI22_X1 U1235 ( .A1(n3895), .A2(n6330), .B1(n3927), .B2(n6327), .ZN(n1296)
         );
  OAI22_X1 U1236 ( .A1(n3895), .A2(n6295), .B1(n3927), .B2(n6292), .ZN(n1571)
         );
  OAI22_X1 U1237 ( .A1(n3894), .A2(n6330), .B1(n3926), .B2(n6327), .ZN(n1279)
         );
  OAI22_X1 U1238 ( .A1(n3894), .A2(n6295), .B1(n3926), .B2(n6292), .ZN(n1588)
         );
  OAI22_X1 U1239 ( .A1(n3893), .A2(n6330), .B1(n3925), .B2(n6327), .ZN(n1262)
         );
  OAI22_X1 U1240 ( .A1(n3893), .A2(n6294), .B1(n3925), .B2(n6291), .ZN(n1605)
         );
  OAI22_X1 U1241 ( .A1(n3892), .A2(n6330), .B1(n3924), .B2(n6327), .ZN(n1245)
         );
  OAI22_X1 U1242 ( .A1(n3892), .A2(n6294), .B1(n3924), .B2(n6291), .ZN(n1622)
         );
  OAI22_X1 U1243 ( .A1(n3891), .A2(n6330), .B1(n3923), .B2(n6327), .ZN(n1228)
         );
  OAI22_X1 U1244 ( .A1(n3891), .A2(n6294), .B1(n3923), .B2(n6291), .ZN(n1639)
         );
  OAI22_X1 U1245 ( .A1(n3890), .A2(n6330), .B1(n3922), .B2(n6327), .ZN(n1211)
         );
  OAI22_X1 U1246 ( .A1(n3890), .A2(n6294), .B1(n3922), .B2(n6291), .ZN(n1656)
         );
  OAI22_X1 U1247 ( .A1(n3889), .A2(n6331), .B1(n3921), .B2(n6328), .ZN(n1194)
         );
  OAI22_X1 U1248 ( .A1(n3889), .A2(n6294), .B1(n3921), .B2(n6291), .ZN(n1673)
         );
  OAI22_X1 U1249 ( .A1(n3888), .A2(n6331), .B1(n3920), .B2(n6328), .ZN(n1177)
         );
  OAI22_X1 U1250 ( .A1(n3888), .A2(n6294), .B1(n3920), .B2(n6291), .ZN(n1690)
         );
  OAI22_X1 U1251 ( .A1(n3887), .A2(n6331), .B1(n3919), .B2(n6328), .ZN(n1160)
         );
  OAI22_X1 U1252 ( .A1(n3887), .A2(n6294), .B1(n3919), .B2(n6291), .ZN(n1707)
         );
  OAI22_X1 U1253 ( .A1(n3886), .A2(n6331), .B1(n3918), .B2(n6328), .ZN(n1143)
         );
  OAI22_X1 U1254 ( .A1(n3886), .A2(n6294), .B1(n3918), .B2(n6291), .ZN(n1724)
         );
  OAI22_X1 U1255 ( .A1(n3885), .A2(n6331), .B1(n3917), .B2(n6328), .ZN(n1126)
         );
  OAI22_X1 U1256 ( .A1(n3885), .A2(n6294), .B1(n3917), .B2(n6291), .ZN(n1741)
         );
  OAI22_X1 U1257 ( .A1(n3884), .A2(n6331), .B1(n3916), .B2(n6328), .ZN(n1109)
         );
  OAI22_X1 U1258 ( .A1(n3884), .A2(n6294), .B1(n3916), .B2(n6291), .ZN(n1758)
         );
  OAI22_X1 U1259 ( .A1(n3883), .A2(n6331), .B1(n3915), .B2(n6328), .ZN(n1092)
         );
  OAI22_X1 U1260 ( .A1(n3883), .A2(n6294), .B1(n3915), .B2(n6291), .ZN(n1775)
         );
  OAI22_X1 U1261 ( .A1(n3882), .A2(n6331), .B1(n3914), .B2(n6328), .ZN(n1075)
         );
  OAI22_X1 U1262 ( .A1(n3882), .A2(n6294), .B1(n3914), .B2(n6291), .ZN(n1792)
         );
  OAI22_X1 U1263 ( .A1(n3881), .A2(n6331), .B1(n3913), .B2(n6328), .ZN(n1058)
         );
  OAI22_X1 U1264 ( .A1(n3881), .A2(n6293), .B1(n3913), .B2(n6290), .ZN(n1809)
         );
  OAI22_X1 U1265 ( .A1(n3880), .A2(n6331), .B1(n3912), .B2(n6328), .ZN(n1041)
         );
  OAI22_X1 U1266 ( .A1(n3880), .A2(n6293), .B1(n3912), .B2(n6290), .ZN(n1826)
         );
  OAI22_X1 U1267 ( .A1(n3879), .A2(n6331), .B1(n3911), .B2(n6328), .ZN(n1024)
         );
  OAI22_X1 U1268 ( .A1(n3879), .A2(n6293), .B1(n3911), .B2(n6290), .ZN(n1843)
         );
  OAI22_X1 U1269 ( .A1(n3878), .A2(n6331), .B1(n3910), .B2(n6328), .ZN(n1007)
         );
  OAI22_X1 U1270 ( .A1(n3878), .A2(n6293), .B1(n3910), .B2(n6290), .ZN(n1860)
         );
  OAI22_X1 U1271 ( .A1(n3877), .A2(n6332), .B1(n3909), .B2(n6329), .ZN(n989)
         );
  OAI22_X1 U1272 ( .A1(n3877), .A2(n6293), .B1(n3909), .B2(n6290), .ZN(n1877)
         );
  OAI22_X1 U1273 ( .A1(n3876), .A2(n6332), .B1(n3908), .B2(n6329), .ZN(n967)
         );
  OAI22_X1 U1274 ( .A1(n3876), .A2(n6293), .B1(n3908), .B2(n6290), .ZN(n1894)
         );
  OAI22_X1 U1275 ( .A1(n3875), .A2(n6332), .B1(n3907), .B2(n6329), .ZN(n946)
         );
  OAI22_X1 U1276 ( .A1(n3875), .A2(n6293), .B1(n3907), .B2(n6290), .ZN(n1911)
         );
  OAI22_X1 U1277 ( .A1(n3874), .A2(n6332), .B1(n3906), .B2(n6329), .ZN(n927)
         );
  OAI22_X1 U1278 ( .A1(n3874), .A2(n6293), .B1(n3906), .B2(n6290), .ZN(n1928)
         );
  OAI22_X1 U1279 ( .A1(n3873), .A2(n6332), .B1(n3905), .B2(n6329), .ZN(n910)
         );
  OAI22_X1 U1280 ( .A1(n3873), .A2(n6293), .B1(n3905), .B2(n6290), .ZN(n1945)
         );
  OAI22_X1 U1281 ( .A1(n3872), .A2(n6332), .B1(n3904), .B2(n6329), .ZN(n893)
         );
  OAI22_X1 U1282 ( .A1(n3872), .A2(n6293), .B1(n3904), .B2(n6290), .ZN(n1962)
         );
  OAI22_X1 U1283 ( .A1(n3871), .A2(n6332), .B1(n3903), .B2(n6329), .ZN(n876)
         );
  OAI22_X1 U1284 ( .A1(n3871), .A2(n6293), .B1(n3903), .B2(n6290), .ZN(n1979)
         );
  OAI22_X1 U1285 ( .A1(n3870), .A2(n6332), .B1(n3902), .B2(n6329), .ZN(n836)
         );
  OAI22_X1 U1286 ( .A1(n3870), .A2(n6293), .B1(n3902), .B2(n6290), .ZN(n2021)
         );
  OAI222_X1 U1287 ( .A1(n2319), .A2(n6319), .B1(n2318), .B2(n6316), .C1(n3805), 
        .C2(n6313), .ZN(n1424) );
  OAI222_X1 U1288 ( .A1(n2319), .A2(n6284), .B1(n2318), .B2(n6281), .C1(n3805), 
        .C2(n6278), .ZN(n1454) );
  OAI222_X1 U1289 ( .A1(n2323), .A2(n6319), .B1(n2322), .B2(n6316), .C1(n3804), 
        .C2(n6313), .ZN(n1382) );
  OAI222_X1 U1290 ( .A1(n2323), .A2(n6284), .B1(n2322), .B2(n6281), .C1(n3804), 
        .C2(n6278), .ZN(n1487) );
  OAI222_X1 U1291 ( .A1(n2327), .A2(n6319), .B1(n2326), .B2(n6316), .C1(n3803), 
        .C2(n6313), .ZN(n1365) );
  OAI222_X1 U1292 ( .A1(n2327), .A2(n6284), .B1(n2326), .B2(n6281), .C1(n3803), 
        .C2(n6278), .ZN(n1504) );
  OAI222_X1 U1293 ( .A1(n2331), .A2(n6319), .B1(n2330), .B2(n6316), .C1(n3802), 
        .C2(n6313), .ZN(n1348) );
  OAI222_X1 U1294 ( .A1(n2331), .A2(n6284), .B1(n2330), .B2(n6281), .C1(n3802), 
        .C2(n6278), .ZN(n1521) );
  OAI222_X1 U1295 ( .A1(n2335), .A2(n6319), .B1(n2334), .B2(n6316), .C1(n3801), 
        .C2(n6313), .ZN(n1331) );
  OAI222_X1 U1296 ( .A1(n2335), .A2(n6284), .B1(n2334), .B2(n6281), .C1(n3801), 
        .C2(n6278), .ZN(n1538) );
  OAI222_X1 U1297 ( .A1(n2339), .A2(n6319), .B1(n2338), .B2(n6316), .C1(n3800), 
        .C2(n6313), .ZN(n1314) );
  OAI222_X1 U1298 ( .A1(n2339), .A2(n6284), .B1(n2338), .B2(n6281), .C1(n3800), 
        .C2(n6278), .ZN(n1555) );
  OAI222_X1 U1299 ( .A1(n2343), .A2(n6319), .B1(n2342), .B2(n6316), .C1(n3799), 
        .C2(n6313), .ZN(n1297) );
  OAI222_X1 U1300 ( .A1(n2343), .A2(n6284), .B1(n2342), .B2(n6281), .C1(n3799), 
        .C2(n6278), .ZN(n1572) );
  OAI222_X1 U1301 ( .A1(n2347), .A2(n6319), .B1(n2346), .B2(n6316), .C1(n3798), 
        .C2(n6313), .ZN(n1280) );
  OAI222_X1 U1302 ( .A1(n2347), .A2(n6284), .B1(n2346), .B2(n6281), .C1(n3798), 
        .C2(n6278), .ZN(n1589) );
  OAI222_X1 U1303 ( .A1(n2351), .A2(n6319), .B1(n2350), .B2(n6316), .C1(n3797), 
        .C2(n6313), .ZN(n1263) );
  OAI222_X1 U1304 ( .A1(n2351), .A2(n6283), .B1(n2350), .B2(n6280), .C1(n3797), 
        .C2(n6277), .ZN(n1606) );
  OAI222_X1 U1305 ( .A1(n2355), .A2(n6319), .B1(n2354), .B2(n6316), .C1(n3796), 
        .C2(n6313), .ZN(n1246) );
  OAI222_X1 U1306 ( .A1(n2355), .A2(n6283), .B1(n2354), .B2(n6280), .C1(n3796), 
        .C2(n6277), .ZN(n1623) );
  OAI222_X1 U1307 ( .A1(n2359), .A2(n6319), .B1(n2358), .B2(n6316), .C1(n3795), 
        .C2(n6313), .ZN(n1229) );
  OAI222_X1 U1308 ( .A1(n2359), .A2(n6283), .B1(n2358), .B2(n6280), .C1(n3795), 
        .C2(n6277), .ZN(n1640) );
  OAI222_X1 U1309 ( .A1(n2363), .A2(n6319), .B1(n2362), .B2(n6316), .C1(n3794), 
        .C2(n6313), .ZN(n1212) );
  OAI222_X1 U1310 ( .A1(n2363), .A2(n6283), .B1(n2362), .B2(n6280), .C1(n3794), 
        .C2(n6277), .ZN(n1657) );
  OAI222_X1 U1311 ( .A1(n2367), .A2(n6320), .B1(n2366), .B2(n6317), .C1(n3793), 
        .C2(n6314), .ZN(n1195) );
  OAI222_X1 U1312 ( .A1(n2367), .A2(n6283), .B1(n2366), .B2(n6280), .C1(n3793), 
        .C2(n6277), .ZN(n1674) );
  OAI222_X1 U1313 ( .A1(n2371), .A2(n6320), .B1(n2370), .B2(n6317), .C1(n3792), 
        .C2(n6314), .ZN(n1178) );
  OAI222_X1 U1314 ( .A1(n2371), .A2(n6283), .B1(n2370), .B2(n6280), .C1(n3792), 
        .C2(n6277), .ZN(n1691) );
  OAI222_X1 U1315 ( .A1(n2375), .A2(n6320), .B1(n2374), .B2(n6317), .C1(n3791), 
        .C2(n6314), .ZN(n1161) );
  OAI222_X1 U1316 ( .A1(n2375), .A2(n6283), .B1(n2374), .B2(n6280), .C1(n3791), 
        .C2(n6277), .ZN(n1708) );
  OAI222_X1 U1317 ( .A1(n2379), .A2(n6320), .B1(n2378), .B2(n6317), .C1(n3790), 
        .C2(n6314), .ZN(n1144) );
  OAI222_X1 U1318 ( .A1(n2379), .A2(n6283), .B1(n2378), .B2(n6280), .C1(n3790), 
        .C2(n6277), .ZN(n1725) );
  OAI222_X1 U1319 ( .A1(n2383), .A2(n6320), .B1(n2382), .B2(n6317), .C1(n3789), 
        .C2(n6314), .ZN(n1127) );
  OAI222_X1 U1320 ( .A1(n2383), .A2(n6283), .B1(n2382), .B2(n6280), .C1(n3789), 
        .C2(n6277), .ZN(n1742) );
  OAI222_X1 U1321 ( .A1(n2387), .A2(n6320), .B1(n2386), .B2(n6317), .C1(n3788), 
        .C2(n6314), .ZN(n1110) );
  OAI222_X1 U1322 ( .A1(n2387), .A2(n6283), .B1(n2386), .B2(n6280), .C1(n3788), 
        .C2(n6277), .ZN(n1759) );
  OAI222_X1 U1323 ( .A1(n2391), .A2(n6320), .B1(n2390), .B2(n6317), .C1(n3787), 
        .C2(n6314), .ZN(n1093) );
  OAI222_X1 U1324 ( .A1(n2391), .A2(n6283), .B1(n2390), .B2(n6280), .C1(n3787), 
        .C2(n6277), .ZN(n1776) );
  OAI222_X1 U1325 ( .A1(n2395), .A2(n6320), .B1(n2394), .B2(n6317), .C1(n3786), 
        .C2(n6314), .ZN(n1076) );
  OAI222_X1 U1326 ( .A1(n2395), .A2(n6283), .B1(n2394), .B2(n6280), .C1(n3786), 
        .C2(n6277), .ZN(n1793) );
  OAI222_X1 U1327 ( .A1(n2399), .A2(n6320), .B1(n2398), .B2(n6317), .C1(n3785), 
        .C2(n6314), .ZN(n1059) );
  OAI222_X1 U1328 ( .A1(n2399), .A2(n6282), .B1(n2398), .B2(n6279), .C1(n3785), 
        .C2(n6276), .ZN(n1810) );
  OAI222_X1 U1329 ( .A1(n2403), .A2(n6320), .B1(n2402), .B2(n6317), .C1(n3784), 
        .C2(n6314), .ZN(n1042) );
  OAI222_X1 U1330 ( .A1(n2403), .A2(n6282), .B1(n2402), .B2(n6279), .C1(n3784), 
        .C2(n6276), .ZN(n1827) );
  OAI222_X1 U1331 ( .A1(n2407), .A2(n6320), .B1(n2406), .B2(n6317), .C1(n3783), 
        .C2(n6314), .ZN(n1025) );
  OAI222_X1 U1332 ( .A1(n2407), .A2(n6282), .B1(n2406), .B2(n6279), .C1(n3783), 
        .C2(n6276), .ZN(n1844) );
  OAI222_X1 U1333 ( .A1(n2411), .A2(n6320), .B1(n2410), .B2(n6317), .C1(n3782), 
        .C2(n6314), .ZN(n1008) );
  OAI222_X1 U1334 ( .A1(n2411), .A2(n6282), .B1(n2410), .B2(n6279), .C1(n3782), 
        .C2(n6276), .ZN(n1861) );
  OAI222_X1 U1335 ( .A1(n2415), .A2(n6321), .B1(n2414), .B2(n6318), .C1(n3781), 
        .C2(n6315), .ZN(n990) );
  OAI222_X1 U1336 ( .A1(n2415), .A2(n6282), .B1(n2414), .B2(n6279), .C1(n3781), 
        .C2(n6276), .ZN(n1878) );
  OAI222_X1 U1337 ( .A1(n2419), .A2(n6321), .B1(n2418), .B2(n6318), .C1(n3780), 
        .C2(n6315), .ZN(n968) );
  OAI222_X1 U1338 ( .A1(n2419), .A2(n6282), .B1(n2418), .B2(n6279), .C1(n3780), 
        .C2(n6276), .ZN(n1895) );
  OAI222_X1 U1339 ( .A1(n2423), .A2(n6321), .B1(n2422), .B2(n6318), .C1(n3779), 
        .C2(n6315), .ZN(n947) );
  OAI222_X1 U1340 ( .A1(n2423), .A2(n6282), .B1(n2422), .B2(n6279), .C1(n3779), 
        .C2(n6276), .ZN(n1912) );
  OAI222_X1 U1341 ( .A1(n2427), .A2(n6321), .B1(n2426), .B2(n6318), .C1(n3778), 
        .C2(n6315), .ZN(n928) );
  OAI222_X1 U1342 ( .A1(n2427), .A2(n6282), .B1(n2426), .B2(n6279), .C1(n3778), 
        .C2(n6276), .ZN(n1929) );
  OAI222_X1 U1343 ( .A1(n2431), .A2(n6321), .B1(n2430), .B2(n6318), .C1(n3777), 
        .C2(n6315), .ZN(n911) );
  OAI222_X1 U1344 ( .A1(n2431), .A2(n6282), .B1(n2430), .B2(n6279), .C1(n3777), 
        .C2(n6276), .ZN(n1946) );
  OAI222_X1 U1345 ( .A1(n2435), .A2(n6321), .B1(n2434), .B2(n6318), .C1(n3776), 
        .C2(n6315), .ZN(n894) );
  OAI222_X1 U1346 ( .A1(n2435), .A2(n6282), .B1(n2434), .B2(n6279), .C1(n3776), 
        .C2(n6276), .ZN(n1963) );
  OAI222_X1 U1347 ( .A1(n2439), .A2(n6321), .B1(n2438), .B2(n6318), .C1(n3775), 
        .C2(n6315), .ZN(n877) );
  OAI222_X1 U1348 ( .A1(n2439), .A2(n6282), .B1(n2438), .B2(n6279), .C1(n3775), 
        .C2(n6276), .ZN(n1980) );
  OAI222_X1 U1349 ( .A1(n2443), .A2(n6321), .B1(n2442), .B2(n6318), .C1(n3774), 
        .C2(n6315), .ZN(n841) );
  OAI222_X1 U1350 ( .A1(n2443), .A2(n6282), .B1(n2442), .B2(n6279), .C1(n3774), 
        .C2(n6276), .ZN(n2024) );
  AOI221_X1 U1351 ( .B1(n6338), .B2(n4060), .C1(n6335), .C2(n4092), .A(n1381), 
        .ZN(n1378) );
  AOI221_X1 U1352 ( .B1(n6299), .B2(n4060), .C1(n6296), .C2(n4092), .A(n1486), 
        .ZN(n1483) );
  AOI221_X1 U1353 ( .B1(n6338), .B2(n4059), .C1(n6335), .C2(n4091), .A(n1364), 
        .ZN(n1361) );
  AOI221_X1 U1354 ( .B1(n6299), .B2(n4059), .C1(n6296), .C2(n4091), .A(n1503), 
        .ZN(n1500) );
  AOI221_X1 U1355 ( .B1(n6338), .B2(n4058), .C1(n6335), .C2(n4090), .A(n1347), 
        .ZN(n1344) );
  AOI221_X1 U1356 ( .B1(n6299), .B2(n4058), .C1(n6296), .C2(n4090), .A(n1520), 
        .ZN(n1517) );
  AOI221_X1 U1357 ( .B1(n6338), .B2(n4057), .C1(n6335), .C2(n4089), .A(n1330), 
        .ZN(n1327) );
  AOI221_X1 U1358 ( .B1(n6299), .B2(n4057), .C1(n6296), .C2(n4089), .A(n1537), 
        .ZN(n1534) );
  AOI221_X1 U1359 ( .B1(n6338), .B2(n4056), .C1(n6335), .C2(n4088), .A(n1313), 
        .ZN(n1310) );
  AOI221_X1 U1360 ( .B1(n6299), .B2(n4056), .C1(n6296), .C2(n4088), .A(n1554), 
        .ZN(n1551) );
  AOI221_X1 U1361 ( .B1(n6338), .B2(n4055), .C1(n6335), .C2(n4087), .A(n1296), 
        .ZN(n1293) );
  AOI221_X1 U1362 ( .B1(n6299), .B2(n4055), .C1(n6296), .C2(n4087), .A(n1571), 
        .ZN(n1568) );
  AOI221_X1 U1363 ( .B1(n6338), .B2(n4054), .C1(n6335), .C2(n4086), .A(n1279), 
        .ZN(n1276) );
  AOI221_X1 U1364 ( .B1(n6299), .B2(n4054), .C1(n6296), .C2(n4086), .A(n1588), 
        .ZN(n1585) );
  AOI221_X1 U1365 ( .B1(n6337), .B2(n4053), .C1(n6334), .C2(n4085), .A(n1262), 
        .ZN(n1259) );
  AOI221_X1 U1366 ( .B1(n6299), .B2(n4053), .C1(n6296), .C2(n4085), .A(n1605), 
        .ZN(n1602) );
  AOI221_X1 U1367 ( .B1(n6337), .B2(n4052), .C1(n6334), .C2(n4084), .A(n1245), 
        .ZN(n1242) );
  AOI221_X1 U1368 ( .B1(n6299), .B2(n4052), .C1(n6296), .C2(n4084), .A(n1622), 
        .ZN(n1619) );
  AOI221_X1 U1369 ( .B1(n6337), .B2(n4051), .C1(n6334), .C2(n4083), .A(n1228), 
        .ZN(n1225) );
  AOI221_X1 U1370 ( .B1(n6299), .B2(n4051), .C1(n6296), .C2(n4083), .A(n1639), 
        .ZN(n1636) );
  AOI221_X1 U1371 ( .B1(n6337), .B2(n4050), .C1(n6334), .C2(n4082), .A(n1211), 
        .ZN(n1208) );
  AOI221_X1 U1372 ( .B1(n6299), .B2(n4050), .C1(n6296), .C2(n4082), .A(n1656), 
        .ZN(n1653) );
  AOI221_X1 U1373 ( .B1(n6337), .B2(n4049), .C1(n6334), .C2(n4081), .A(n1194), 
        .ZN(n1191) );
  AOI221_X1 U1374 ( .B1(n6300), .B2(n4049), .C1(n6297), .C2(n4081), .A(n1673), 
        .ZN(n1670) );
  AOI221_X1 U1375 ( .B1(n6337), .B2(n4048), .C1(n6334), .C2(n4080), .A(n1177), 
        .ZN(n1174) );
  AOI221_X1 U1376 ( .B1(n6300), .B2(n4048), .C1(n6297), .C2(n4080), .A(n1690), 
        .ZN(n1687) );
  AOI221_X1 U1377 ( .B1(n6337), .B2(n4047), .C1(n6334), .C2(n4079), .A(n1160), 
        .ZN(n1157) );
  AOI221_X1 U1378 ( .B1(n6300), .B2(n4047), .C1(n6297), .C2(n4079), .A(n1707), 
        .ZN(n1704) );
  AOI221_X1 U1379 ( .B1(n6337), .B2(n4046), .C1(n6334), .C2(n4078), .A(n1143), 
        .ZN(n1140) );
  AOI221_X1 U1380 ( .B1(n6300), .B2(n4046), .C1(n6297), .C2(n4078), .A(n1724), 
        .ZN(n1721) );
  AOI221_X1 U1381 ( .B1(n6337), .B2(n4045), .C1(n6334), .C2(n4077), .A(n1126), 
        .ZN(n1123) );
  AOI221_X1 U1382 ( .B1(n6300), .B2(n4045), .C1(n6297), .C2(n4077), .A(n1741), 
        .ZN(n1738) );
  AOI221_X1 U1383 ( .B1(n6337), .B2(n4044), .C1(n6334), .C2(n4076), .A(n1109), 
        .ZN(n1106) );
  AOI221_X1 U1384 ( .B1(n6300), .B2(n4044), .C1(n6297), .C2(n4076), .A(n1758), 
        .ZN(n1755) );
  AOI221_X1 U1385 ( .B1(n6337), .B2(n4043), .C1(n6334), .C2(n4075), .A(n1092), 
        .ZN(n1089) );
  AOI221_X1 U1386 ( .B1(n6300), .B2(n4043), .C1(n6297), .C2(n4075), .A(n1775), 
        .ZN(n1772) );
  AOI221_X1 U1387 ( .B1(n6337), .B2(n4042), .C1(n6334), .C2(n4074), .A(n1075), 
        .ZN(n1072) );
  AOI221_X1 U1388 ( .B1(n6300), .B2(n4042), .C1(n6297), .C2(n4074), .A(n1792), 
        .ZN(n1789) );
  AOI221_X1 U1389 ( .B1(n6336), .B2(n4041), .C1(n6333), .C2(n4073), .A(n1058), 
        .ZN(n1055) );
  AOI221_X1 U1390 ( .B1(n6300), .B2(n4041), .C1(n6297), .C2(n4073), .A(n1809), 
        .ZN(n1806) );
  AOI221_X1 U1391 ( .B1(n6336), .B2(n4040), .C1(n6333), .C2(n4072), .A(n1041), 
        .ZN(n1038) );
  AOI221_X1 U1392 ( .B1(n6300), .B2(n4040), .C1(n6297), .C2(n4072), .A(n1826), 
        .ZN(n1823) );
  AOI221_X1 U1393 ( .B1(n6336), .B2(n4039), .C1(n6333), .C2(n4071), .A(n1024), 
        .ZN(n1021) );
  AOI221_X1 U1394 ( .B1(n6300), .B2(n4039), .C1(n6297), .C2(n4071), .A(n1843), 
        .ZN(n1840) );
  AOI221_X1 U1395 ( .B1(n6336), .B2(n4038), .C1(n6333), .C2(n4070), .A(n1007), 
        .ZN(n1004) );
  AOI221_X1 U1396 ( .B1(n6300), .B2(n4038), .C1(n6297), .C2(n4070), .A(n1860), 
        .ZN(n1857) );
  AOI221_X1 U1397 ( .B1(n6336), .B2(n4037), .C1(n6333), .C2(n4069), .A(n989), 
        .ZN(n984) );
  AOI221_X1 U1398 ( .B1(n6301), .B2(n4037), .C1(n6298), .C2(n4069), .A(n1877), 
        .ZN(n1874) );
  AOI221_X1 U1399 ( .B1(n6336), .B2(n4036), .C1(n6333), .C2(n4068), .A(n967), 
        .ZN(n963) );
  AOI221_X1 U1400 ( .B1(n6301), .B2(n4036), .C1(n6298), .C2(n4068), .A(n1894), 
        .ZN(n1891) );
  AOI221_X1 U1401 ( .B1(n6336), .B2(n4035), .C1(n6333), .C2(n4067), .A(n946), 
        .ZN(n943) );
  AOI221_X1 U1402 ( .B1(n6301), .B2(n4035), .C1(n6298), .C2(n4067), .A(n1911), 
        .ZN(n1908) );
  AOI221_X1 U1403 ( .B1(n6336), .B2(n4034), .C1(n6333), .C2(n4066), .A(n927), 
        .ZN(n924) );
  AOI221_X1 U1404 ( .B1(n6301), .B2(n4034), .C1(n6298), .C2(n4066), .A(n1928), 
        .ZN(n1925) );
  AOI221_X1 U1405 ( .B1(n6336), .B2(n4033), .C1(n6333), .C2(n4065), .A(n910), 
        .ZN(n907) );
  AOI221_X1 U1406 ( .B1(n6301), .B2(n4033), .C1(n6298), .C2(n4065), .A(n1945), 
        .ZN(n1942) );
  AOI221_X1 U1407 ( .B1(n6336), .B2(n4032), .C1(n6333), .C2(n4064), .A(n893), 
        .ZN(n890) );
  AOI221_X1 U1408 ( .B1(n6301), .B2(n4032), .C1(n6298), .C2(n4064), .A(n1962), 
        .ZN(n1959) );
  AOI221_X1 U1409 ( .B1(n6336), .B2(n4031), .C1(n6333), .C2(n4063), .A(n876), 
        .ZN(n873) );
  AOI221_X1 U1410 ( .B1(n6301), .B2(n4031), .C1(n6298), .C2(n4063), .A(n1979), 
        .ZN(n1976) );
  INV_X1 U1411 ( .A(n6084), .ZN(n6083) );
  INV_X1 U1412 ( .A(n6093), .ZN(n6092) );
  INV_X1 U1413 ( .A(DATAIN[0]), .ZN(n6339) );
  INV_X1 U1414 ( .A(DATAIN[0]), .ZN(n6340) );
  INV_X1 U1415 ( .A(DATAIN[1]), .ZN(n6341) );
  INV_X1 U1416 ( .A(DATAIN[1]), .ZN(n6342) );
  INV_X1 U1417 ( .A(DATAIN[2]), .ZN(n6343) );
  INV_X1 U1418 ( .A(DATAIN[2]), .ZN(n6344) );
  INV_X1 U1419 ( .A(DATAIN[3]), .ZN(n6345) );
  INV_X1 U1420 ( .A(DATAIN[3]), .ZN(n6346) );
  CLKBUF_X1 U1421 ( .A(n6478), .Z(n6382) );
  CLKBUF_X1 U1422 ( .A(n6478), .Z(n6383) );
  CLKBUF_X1 U1423 ( .A(n6478), .Z(n6384) );
  CLKBUF_X1 U1424 ( .A(n6478), .Z(n6385) );
  CLKBUF_X1 U1425 ( .A(n6478), .Z(n6386) );
  CLKBUF_X1 U1426 ( .A(n6477), .Z(n6387) );
  CLKBUF_X1 U1427 ( .A(n6477), .Z(n6388) );
  CLKBUF_X1 U1428 ( .A(n6477), .Z(n6389) );
  CLKBUF_X1 U1429 ( .A(n6477), .Z(n6390) );
  CLKBUF_X1 U1430 ( .A(n6477), .Z(n6391) );
  CLKBUF_X1 U1431 ( .A(n6477), .Z(n6392) );
  CLKBUF_X1 U1432 ( .A(n6476), .Z(n6393) );
  CLKBUF_X1 U1433 ( .A(n6476), .Z(n6394) );
  CLKBUF_X1 U1434 ( .A(n6476), .Z(n6395) );
  CLKBUF_X1 U1435 ( .A(n6476), .Z(n6396) );
  CLKBUF_X1 U1436 ( .A(n6476), .Z(n6397) );
  CLKBUF_X1 U1437 ( .A(n6476), .Z(n6398) );
  CLKBUF_X1 U1438 ( .A(n6475), .Z(n6399) );
  CLKBUF_X1 U1439 ( .A(n6475), .Z(n6400) );
  CLKBUF_X1 U1440 ( .A(n6475), .Z(n6401) );
  CLKBUF_X1 U1441 ( .A(n6475), .Z(n6402) );
  CLKBUF_X1 U1442 ( .A(n6475), .Z(n6403) );
  CLKBUF_X1 U1443 ( .A(n6475), .Z(n6404) );
  CLKBUF_X1 U1444 ( .A(n6474), .Z(n6405) );
  CLKBUF_X1 U1445 ( .A(n6474), .Z(n6406) );
  CLKBUF_X1 U1446 ( .A(n6474), .Z(n6407) );
  CLKBUF_X1 U1447 ( .A(n6474), .Z(n6408) );
  CLKBUF_X1 U1448 ( .A(n6474), .Z(n6409) );
  CLKBUF_X1 U1449 ( .A(n6474), .Z(n6410) );
  CLKBUF_X1 U1450 ( .A(n6473), .Z(n6411) );
  CLKBUF_X1 U1451 ( .A(n6473), .Z(n6412) );
  CLKBUF_X1 U1452 ( .A(n6473), .Z(n6413) );
  CLKBUF_X1 U1453 ( .A(n6473), .Z(n6414) );
  CLKBUF_X1 U1454 ( .A(n6473), .Z(n6415) );
  CLKBUF_X1 U1455 ( .A(n6473), .Z(n6416) );
  CLKBUF_X1 U1456 ( .A(n6472), .Z(n6417) );
  CLKBUF_X1 U1457 ( .A(n6472), .Z(n6418) );
  CLKBUF_X1 U1458 ( .A(n6472), .Z(n6419) );
  CLKBUF_X1 U1459 ( .A(n6472), .Z(n6420) );
  CLKBUF_X1 U1460 ( .A(n6472), .Z(n6421) );
  CLKBUF_X1 U1461 ( .A(n6472), .Z(n6422) );
  CLKBUF_X1 U1462 ( .A(n6471), .Z(n6423) );
  CLKBUF_X1 U1463 ( .A(n6471), .Z(n6424) );
  CLKBUF_X1 U1464 ( .A(n6471), .Z(n6425) );
  CLKBUF_X1 U1465 ( .A(n6471), .Z(n6426) );
  CLKBUF_X1 U1466 ( .A(n6471), .Z(n6427) );
  CLKBUF_X1 U1467 ( .A(n6471), .Z(n6428) );
  CLKBUF_X1 U1468 ( .A(n6470), .Z(n6429) );
  CLKBUF_X1 U1469 ( .A(n6470), .Z(n6430) );
  CLKBUF_X1 U1470 ( .A(n6470), .Z(n6431) );
  CLKBUF_X1 U1471 ( .A(n6470), .Z(n6432) );
  CLKBUF_X1 U1472 ( .A(n6470), .Z(n6433) );
  CLKBUF_X1 U1473 ( .A(n6470), .Z(n6434) );
  CLKBUF_X1 U1474 ( .A(n6469), .Z(n6435) );
  CLKBUF_X1 U1475 ( .A(n6469), .Z(n6436) );
  CLKBUF_X1 U1476 ( .A(n6469), .Z(n6437) );
  CLKBUF_X1 U1477 ( .A(n6469), .Z(n6438) );
  CLKBUF_X1 U1478 ( .A(n6469), .Z(n6439) );
  CLKBUF_X1 U1479 ( .A(n6469), .Z(n6440) );
  CLKBUF_X1 U1480 ( .A(n6468), .Z(n6441) );
  CLKBUF_X1 U1481 ( .A(n6468), .Z(n6442) );
  CLKBUF_X1 U1482 ( .A(n6468), .Z(n6443) );
  CLKBUF_X1 U1483 ( .A(n6468), .Z(n6444) );
  CLKBUF_X1 U1484 ( .A(n6468), .Z(n6445) );
  CLKBUF_X1 U1485 ( .A(n6468), .Z(n6446) );
  CLKBUF_X1 U1486 ( .A(n6467), .Z(n6447) );
  CLKBUF_X1 U1487 ( .A(n6467), .Z(n6448) );
  CLKBUF_X1 U1488 ( .A(n6467), .Z(n6449) );
  CLKBUF_X1 U1489 ( .A(n6467), .Z(n6450) );
  CLKBUF_X1 U1490 ( .A(n6467), .Z(n6451) );
  CLKBUF_X1 U1491 ( .A(n6467), .Z(n6452) );
  CLKBUF_X1 U1492 ( .A(n6466), .Z(n6453) );
  CLKBUF_X1 U1493 ( .A(n6466), .Z(n6454) );
  CLKBUF_X1 U1494 ( .A(n6466), .Z(n6455) );
  CLKBUF_X1 U1495 ( .A(n6466), .Z(n6456) );
  CLKBUF_X1 U1496 ( .A(n6466), .Z(n6457) );
  CLKBUF_X1 U1497 ( .A(n6466), .Z(n6458) );
  CLKBUF_X1 U1498 ( .A(n6465), .Z(n6459) );
  CLKBUF_X1 U1499 ( .A(n6465), .Z(n6460) );
  CLKBUF_X1 U1500 ( .A(n6465), .Z(n6461) );
  CLKBUF_X1 U1501 ( .A(n6465), .Z(n6462) );
  CLKBUF_X1 U1502 ( .A(n6465), .Z(n6463) );
  INV_X1 U1503 ( .A(ADD_WR[2]), .ZN(n7591) );
  INV_X1 U1504 ( .A(ADD_WR[3]), .ZN(n7590) );
  INV_X1 U1505 ( .A(ADD_WR[4]), .ZN(n7589) );
  INV_X1 U1506 ( .A(ADD_RS1[3]), .ZN(n7592) );
  INV_X1 U1507 ( .A(ADD_RS1[0]), .ZN(n7593) );
  INV_X1 U1508 ( .A(ADD_RS1[4]), .ZN(n7901) );
  INV_X1 U1509 ( .A(ADD_RS1[1]), .ZN(n6479) );
  INV_X1 U1510 ( .A(n2059), .ZN(n7587) );
  INV_X1 U1511 ( .A(n2316), .ZN(n7585) );
  INV_X1 U1512 ( .A(ADD_RS2[3]), .ZN(n7594) );
  INV_X1 U1513 ( .A(ADD_RS2[0]), .ZN(n7595) );
  INV_X1 U1514 ( .A(ADD_RS2[4]), .ZN(n7899) );
  INV_X1 U1515 ( .A(ADD_RS2[1]), .ZN(n6480) );
  INV_X1 U1516 ( .A(n2028), .ZN(n7588) );
  INV_X1 U1517 ( .A(n2440), .ZN(n7586) );
  INV_X1 U1518 ( .A(n4125), .ZN(n6938) );
  NAND3_X1 U1519 ( .A1(n749), .A2(n7589), .A3(n7590), .ZN(n6481) );
  INV_X1 U1520 ( .A(n6481), .ZN(n6489) );
  INV_X1 U1521 ( .A(ADD_WR[1]), .ZN(n6482) );
  INV_X1 U1522 ( .A(n4124), .ZN(n6957) );
  INV_X1 U1523 ( .A(n4123), .ZN(n6975) );
  INV_X1 U1524 ( .A(n4122), .ZN(n6993) );
  INV_X1 U1525 ( .A(n4121), .ZN(n7012) );
  INV_X1 U1526 ( .A(n4120), .ZN(n7031) );
  INV_X1 U1527 ( .A(n4119), .ZN(n7050) );
  INV_X1 U1528 ( .A(n4118), .ZN(n7069) );
  INV_X1 U1529 ( .A(n4117), .ZN(n7088) );
  INV_X1 U1530 ( .A(n4116), .ZN(n7107) );
  INV_X1 U1531 ( .A(n4115), .ZN(n7126) );
  INV_X1 U1532 ( .A(n4114), .ZN(n7145) );
  INV_X1 U1533 ( .A(n4113), .ZN(n7164) );
  INV_X1 U1534 ( .A(n4112), .ZN(n7183) );
  INV_X1 U1535 ( .A(n4111), .ZN(n7202) );
  INV_X1 U1536 ( .A(n4110), .ZN(n7221) );
  INV_X1 U1537 ( .A(n4109), .ZN(n7240) );
  INV_X1 U1538 ( .A(n4108), .ZN(n7259) );
  INV_X1 U1539 ( .A(n4107), .ZN(n7278) );
  INV_X1 U1540 ( .A(n4106), .ZN(n7297) );
  INV_X1 U1541 ( .A(n4105), .ZN(n7316) );
  INV_X1 U1542 ( .A(n4104), .ZN(n7335) );
  INV_X1 U1543 ( .A(n4103), .ZN(n7354) );
  INV_X1 U1544 ( .A(n4102), .ZN(n7373) );
  MUX2_X1 U1545 ( .A(n5210), .B(DATAIN[23]), .S(n6006), .Z(n4277) );
  INV_X1 U1546 ( .A(n4101), .ZN(n7392) );
  INV_X1 U1547 ( .A(n4100), .ZN(n7411) );
  INV_X1 U1548 ( .A(n4099), .ZN(n7430) );
  INV_X1 U1549 ( .A(n4098), .ZN(n7449) );
  INV_X1 U1550 ( .A(n4097), .ZN(n7468) );
  INV_X1 U1551 ( .A(n4096), .ZN(n7487) );
  MUX2_X1 U1552 ( .A(n5204), .B(DATAIN[29]), .S(n6007), .Z(n4283) );
  INV_X1 U1553 ( .A(n4095), .ZN(n7506) );
  MUX2_X1 U1554 ( .A(n5203), .B(DATAIN[30]), .S(n6007), .Z(n4284) );
  INV_X1 U1555 ( .A(n4094), .ZN(n7531) );
  MUX2_X1 U1556 ( .A(n5169), .B(DATAIN[31]), .S(n6007), .Z(n4285) );
  MUX2_X1 U1557 ( .A(n5872), .B(DATAIN[0]), .S(n6008), .Z(n4158) );
  MUX2_X1 U1558 ( .A(n5871), .B(DATAIN[1]), .S(n6008), .Z(n4159) );
  MUX2_X1 U1559 ( .A(n5870), .B(DATAIN[2]), .S(n6008), .Z(n4160) );
  MUX2_X1 U1560 ( .A(n5869), .B(DATAIN[3]), .S(n6008), .Z(n4161) );
  MUX2_X1 U1561 ( .A(n5868), .B(DATAIN[4]), .S(n6008), .Z(n4162) );
  MUX2_X1 U1562 ( .A(n5867), .B(DATAIN[5]), .S(n6008), .Z(n4163) );
  MUX2_X1 U1563 ( .A(n5866), .B(DATAIN[6]), .S(n6008), .Z(n4164) );
  MUX2_X1 U1564 ( .A(n5865), .B(DATAIN[7]), .S(n6008), .Z(n4165) );
  MUX2_X1 U1565 ( .A(n5864), .B(DATAIN[8]), .S(n6008), .Z(n4166) );
  MUX2_X1 U1566 ( .A(n5863), .B(DATAIN[9]), .S(n6008), .Z(n4167) );
  MUX2_X1 U1567 ( .A(n5862), .B(DATAIN[10]), .S(n6008), .Z(n4168) );
  MUX2_X1 U1568 ( .A(n5861), .B(DATAIN[11]), .S(n6008), .Z(n4169) );
  MUX2_X1 U1569 ( .A(n5860), .B(DATAIN[12]), .S(n6009), .Z(n4170) );
  MUX2_X1 U1570 ( .A(n5859), .B(DATAIN[13]), .S(n6009), .Z(n4171) );
  MUX2_X1 U1571 ( .A(n5858), .B(DATAIN[14]), .S(n6009), .Z(n4172) );
  MUX2_X1 U1572 ( .A(n5857), .B(DATAIN[15]), .S(n6009), .Z(n4173) );
  MUX2_X1 U1573 ( .A(n5856), .B(DATAIN[16]), .S(n6009), .Z(n4174) );
  MUX2_X1 U1574 ( .A(n5855), .B(DATAIN[17]), .S(n6009), .Z(n4175) );
  MUX2_X1 U1575 ( .A(n5854), .B(DATAIN[18]), .S(n6009), .Z(n4176) );
  MUX2_X1 U1576 ( .A(n5853), .B(DATAIN[19]), .S(n6009), .Z(n4177) );
  MUX2_X1 U1577 ( .A(n5852), .B(DATAIN[20]), .S(n6009), .Z(n4178) );
  MUX2_X1 U1578 ( .A(n5851), .B(DATAIN[21]), .S(n6009), .Z(n4179) );
  MUX2_X1 U1579 ( .A(n5850), .B(DATAIN[22]), .S(n6009), .Z(n4180) );
  MUX2_X1 U1580 ( .A(n5849), .B(DATAIN[23]), .S(n6009), .Z(n4181) );
  MUX2_X1 U1581 ( .A(n5848), .B(DATAIN[24]), .S(n6010), .Z(n4182) );
  MUX2_X1 U1582 ( .A(n5847), .B(DATAIN[25]), .S(n6010), .Z(n4183) );
  MUX2_X1 U1583 ( .A(n5846), .B(DATAIN[26]), .S(n6010), .Z(n4184) );
  MUX2_X1 U1584 ( .A(n5845), .B(DATAIN[27]), .S(n6010), .Z(n4185) );
  MUX2_X1 U1585 ( .A(n5844), .B(DATAIN[28]), .S(n6010), .Z(n4186) );
  MUX2_X1 U1586 ( .A(n5843), .B(DATAIN[29]), .S(n6010), .Z(n4187) );
  MUX2_X1 U1587 ( .A(n5842), .B(DATAIN[30]), .S(n6010), .Z(n4188) );
  MUX2_X1 U1588 ( .A(n5841), .B(DATAIN[31]), .S(n6010), .Z(n4189) );
  MUX2_X1 U1589 ( .A(n5874), .B(DATAIN[0]), .S(n6011), .Z(n4222) );
  MUX2_X1 U1590 ( .A(n5357), .B(DATAIN[1]), .S(n6011), .Z(n4223) );
  MUX2_X1 U1591 ( .A(n5356), .B(DATAIN[2]), .S(n6011), .Z(n4224) );
  MUX2_X1 U1592 ( .A(n5355), .B(DATAIN[3]), .S(n6011), .Z(n4225) );
  MUX2_X1 U1593 ( .A(n5354), .B(DATAIN[4]), .S(n6011), .Z(n4226) );
  MUX2_X1 U1594 ( .A(n5353), .B(DATAIN[5]), .S(n6011), .Z(n4227) );
  MUX2_X1 U1595 ( .A(n5352), .B(DATAIN[6]), .S(n6011), .Z(n4228) );
  MUX2_X1 U1596 ( .A(n5351), .B(DATAIN[7]), .S(n6011), .Z(n4229) );
  MUX2_X1 U1597 ( .A(n5350), .B(DATAIN[8]), .S(n6011), .Z(n4230) );
  MUX2_X1 U1598 ( .A(n5349), .B(DATAIN[9]), .S(n6011), .Z(n4231) );
  MUX2_X1 U1599 ( .A(n5348), .B(DATAIN[10]), .S(n6011), .Z(n4232) );
  MUX2_X1 U1600 ( .A(n5347), .B(DATAIN[11]), .S(n6011), .Z(n4233) );
  MUX2_X1 U1601 ( .A(n5346), .B(DATAIN[12]), .S(n6012), .Z(n4234) );
  MUX2_X1 U1602 ( .A(n5345), .B(DATAIN[13]), .S(n6012), .Z(n4235) );
  MUX2_X1 U1603 ( .A(n5344), .B(DATAIN[14]), .S(n6012), .Z(n4236) );
  MUX2_X1 U1604 ( .A(n5343), .B(DATAIN[15]), .S(n6012), .Z(n4237) );
  MUX2_X1 U1605 ( .A(n5342), .B(DATAIN[16]), .S(n6012), .Z(n4238) );
  MUX2_X1 U1606 ( .A(n5341), .B(DATAIN[17]), .S(n6012), .Z(n4239) );
  MUX2_X1 U1607 ( .A(n5340), .B(DATAIN[18]), .S(n6012), .Z(n4240) );
  MUX2_X1 U1608 ( .A(n5339), .B(DATAIN[19]), .S(n6012), .Z(n4241) );
  MUX2_X1 U1609 ( .A(n5338), .B(DATAIN[20]), .S(n6012), .Z(n4242) );
  MUX2_X1 U1610 ( .A(n5337), .B(DATAIN[21]), .S(n6012), .Z(n4243) );
  MUX2_X1 U1611 ( .A(n5336), .B(DATAIN[22]), .S(n6012), .Z(n4244) );
  MUX2_X1 U1612 ( .A(n5335), .B(DATAIN[23]), .S(n6012), .Z(n4245) );
  MUX2_X1 U1613 ( .A(n5334), .B(DATAIN[24]), .S(n6013), .Z(n4246) );
  MUX2_X1 U1614 ( .A(n5333), .B(DATAIN[25]), .S(n6013), .Z(n4247) );
  MUX2_X1 U1615 ( .A(n5332), .B(DATAIN[26]), .S(n6013), .Z(n4248) );
  MUX2_X1 U1616 ( .A(n5331), .B(DATAIN[27]), .S(n6013), .Z(n4249) );
  MUX2_X1 U1617 ( .A(n5330), .B(DATAIN[28]), .S(n6013), .Z(n4250) );
  MUX2_X1 U1618 ( .A(n5329), .B(DATAIN[29]), .S(n6013), .Z(n4251) );
  MUX2_X1 U1619 ( .A(n5328), .B(DATAIN[30]), .S(n6013), .Z(n4252) );
  MUX2_X1 U1620 ( .A(n5873), .B(DATAIN[31]), .S(n6013), .Z(n4253) );
  INV_X1 U1621 ( .A(ADD_WR[0]), .ZN(n6485) );
  MUX2_X1 U1622 ( .A(n5547), .B(DATAIN[0]), .S(n6014), .Z(n4350) );
  MUX2_X1 U1623 ( .A(n5452), .B(DATAIN[1]), .S(n6014), .Z(n4351) );
  MUX2_X1 U1624 ( .A(n5451), .B(DATAIN[2]), .S(n6014), .Z(n4352) );
  MUX2_X1 U1625 ( .A(n5450), .B(DATAIN[3]), .S(n6014), .Z(n4353) );
  MUX2_X1 U1626 ( .A(n5449), .B(DATAIN[4]), .S(n6014), .Z(n4354) );
  MUX2_X1 U1627 ( .A(n5448), .B(DATAIN[5]), .S(n6014), .Z(n4355) );
  MUX2_X1 U1628 ( .A(n5447), .B(DATAIN[6]), .S(n6014), .Z(n4356) );
  MUX2_X1 U1629 ( .A(n5446), .B(DATAIN[7]), .S(n6014), .Z(n4357) );
  MUX2_X1 U1630 ( .A(n5445), .B(DATAIN[8]), .S(n6014), .Z(n4358) );
  MUX2_X1 U1631 ( .A(n5444), .B(DATAIN[9]), .S(n6014), .Z(n4359) );
  MUX2_X1 U1632 ( .A(n5443), .B(DATAIN[10]), .S(n6014), .Z(n4360) );
  MUX2_X1 U1633 ( .A(n5442), .B(DATAIN[11]), .S(n6014), .Z(n4361) );
  MUX2_X1 U1634 ( .A(n5441), .B(DATAIN[12]), .S(n6015), .Z(n4362) );
  MUX2_X1 U1635 ( .A(n5440), .B(DATAIN[13]), .S(n6015), .Z(n4363) );
  MUX2_X1 U1636 ( .A(n5439), .B(DATAIN[14]), .S(n6015), .Z(n4364) );
  MUX2_X1 U1637 ( .A(n5438), .B(DATAIN[15]), .S(n6015), .Z(n4365) );
  MUX2_X1 U1638 ( .A(n5437), .B(DATAIN[16]), .S(n6015), .Z(n4366) );
  MUX2_X1 U1639 ( .A(n5436), .B(DATAIN[17]), .S(n6015), .Z(n4367) );
  MUX2_X1 U1640 ( .A(n5435), .B(DATAIN[18]), .S(n6015), .Z(n4368) );
  MUX2_X1 U1641 ( .A(n5434), .B(DATAIN[19]), .S(n6015), .Z(n4369) );
  MUX2_X1 U1642 ( .A(n5433), .B(DATAIN[20]), .S(n6015), .Z(n4370) );
  MUX2_X1 U1643 ( .A(n5432), .B(DATAIN[21]), .S(n6015), .Z(n4371) );
  MUX2_X1 U1644 ( .A(n5431), .B(DATAIN[22]), .S(n6015), .Z(n4372) );
  MUX2_X1 U1645 ( .A(n5430), .B(DATAIN[23]), .S(n6015), .Z(n4373) );
  MUX2_X1 U1646 ( .A(n5429), .B(DATAIN[24]), .S(n6016), .Z(n4374) );
  MUX2_X1 U1647 ( .A(n5428), .B(DATAIN[25]), .S(n6016), .Z(n4375) );
  MUX2_X1 U1648 ( .A(n5427), .B(DATAIN[26]), .S(n6016), .Z(n4376) );
  MUX2_X1 U1649 ( .A(n5426), .B(DATAIN[27]), .S(n6016), .Z(n4377) );
  MUX2_X1 U1650 ( .A(n5425), .B(DATAIN[28]), .S(n6016), .Z(n4378) );
  MUX2_X1 U1651 ( .A(n5424), .B(DATAIN[29]), .S(n6016), .Z(n4379) );
  MUX2_X1 U1652 ( .A(n5423), .B(DATAIN[30]), .S(n6016), .Z(n4380) );
  MUX2_X1 U1653 ( .A(n5422), .B(DATAIN[31]), .S(n6016), .Z(n4381) );
  INV_X1 U1654 ( .A(n2974), .ZN(n6934) );
  MUX2_X1 U1655 ( .A(n5136), .B(DATAIN[0]), .S(n6017), .Z(n4414) );
  INV_X1 U1656 ( .A(n2975), .ZN(n6953) );
  MUX2_X1 U1657 ( .A(n5135), .B(DATAIN[1]), .S(n6017), .Z(n4415) );
  INV_X1 U1658 ( .A(n2976), .ZN(n6971) );
  MUX2_X1 U1659 ( .A(n5134), .B(DATAIN[2]), .S(n6017), .Z(n4416) );
  INV_X1 U1660 ( .A(n2977), .ZN(n6989) );
  MUX2_X1 U1661 ( .A(n5133), .B(DATAIN[3]), .S(n6017), .Z(n4417) );
  INV_X1 U1662 ( .A(n2978), .ZN(n7008) );
  MUX2_X1 U1663 ( .A(n5132), .B(DATAIN[4]), .S(n6017), .Z(n4418) );
  INV_X1 U1664 ( .A(n2979), .ZN(n7027) );
  MUX2_X1 U1665 ( .A(n5131), .B(DATAIN[5]), .S(n6017), .Z(n4419) );
  INV_X1 U1666 ( .A(n2980), .ZN(n7046) );
  MUX2_X1 U1667 ( .A(n5130), .B(DATAIN[6]), .S(n6017), .Z(n4420) );
  INV_X1 U1668 ( .A(n2981), .ZN(n7065) );
  MUX2_X1 U1669 ( .A(n5129), .B(DATAIN[7]), .S(n6017), .Z(n4421) );
  INV_X1 U1670 ( .A(n2982), .ZN(n7084) );
  MUX2_X1 U1671 ( .A(n5128), .B(DATAIN[8]), .S(n6017), .Z(n4422) );
  INV_X1 U1672 ( .A(n3559), .ZN(n7103) );
  MUX2_X1 U1673 ( .A(n5127), .B(DATAIN[9]), .S(n6017), .Z(n4423) );
  INV_X1 U1674 ( .A(n3560), .ZN(n7122) );
  MUX2_X1 U1675 ( .A(n5126), .B(DATAIN[10]), .S(n6017), .Z(n4424) );
  INV_X1 U1676 ( .A(n3561), .ZN(n7141) );
  MUX2_X1 U1677 ( .A(n5125), .B(DATAIN[11]), .S(n6017), .Z(n4425) );
  INV_X1 U1678 ( .A(n3562), .ZN(n7160) );
  MUX2_X1 U1679 ( .A(n5124), .B(DATAIN[12]), .S(n6018), .Z(n4426) );
  INV_X1 U1680 ( .A(n3563), .ZN(n7179) );
  MUX2_X1 U1681 ( .A(n5123), .B(DATAIN[13]), .S(n6018), .Z(n4427) );
  INV_X1 U1682 ( .A(n3564), .ZN(n7198) );
  MUX2_X1 U1683 ( .A(n5122), .B(DATAIN[14]), .S(n6018), .Z(n4428) );
  INV_X1 U1684 ( .A(n3565), .ZN(n7217) );
  MUX2_X1 U1685 ( .A(n5121), .B(DATAIN[15]), .S(n6018), .Z(n4429) );
  INV_X1 U1686 ( .A(n3566), .ZN(n7236) );
  MUX2_X1 U1687 ( .A(n5120), .B(DATAIN[16]), .S(n6018), .Z(n4430) );
  INV_X1 U1688 ( .A(n3567), .ZN(n7255) );
  MUX2_X1 U1689 ( .A(n5119), .B(DATAIN[17]), .S(n6018), .Z(n4431) );
  INV_X1 U1690 ( .A(n3568), .ZN(n7274) );
  MUX2_X1 U1691 ( .A(n5118), .B(DATAIN[18]), .S(n6018), .Z(n4432) );
  INV_X1 U1692 ( .A(n3569), .ZN(n7293) );
  MUX2_X1 U1693 ( .A(n5117), .B(DATAIN[19]), .S(n6018), .Z(n4433) );
  INV_X1 U1694 ( .A(n3570), .ZN(n7312) );
  MUX2_X1 U1695 ( .A(n5116), .B(DATAIN[20]), .S(n6018), .Z(n4434) );
  INV_X1 U1696 ( .A(n3571), .ZN(n7331) );
  MUX2_X1 U1697 ( .A(n5115), .B(DATAIN[21]), .S(n6018), .Z(n4435) );
  INV_X1 U1698 ( .A(n3572), .ZN(n7350) );
  MUX2_X1 U1699 ( .A(n5114), .B(DATAIN[22]), .S(n6018), .Z(n4436) );
  INV_X1 U1700 ( .A(n3573), .ZN(n7369) );
  MUX2_X1 U1701 ( .A(n5113), .B(DATAIN[23]), .S(n6018), .Z(n4437) );
  INV_X1 U1702 ( .A(n3574), .ZN(n7388) );
  MUX2_X1 U1703 ( .A(n5112), .B(DATAIN[24]), .S(n6019), .Z(n4438) );
  INV_X1 U1704 ( .A(n3575), .ZN(n7407) );
  MUX2_X1 U1705 ( .A(n5111), .B(DATAIN[25]), .S(n6019), .Z(n4439) );
  INV_X1 U1706 ( .A(n3576), .ZN(n7426) );
  MUX2_X1 U1707 ( .A(n5110), .B(DATAIN[26]), .S(n6019), .Z(n4440) );
  INV_X1 U1708 ( .A(n3577), .ZN(n7445) );
  MUX2_X1 U1709 ( .A(n5109), .B(DATAIN[27]), .S(n6019), .Z(n4441) );
  INV_X1 U1710 ( .A(n3578), .ZN(n7464) );
  MUX2_X1 U1711 ( .A(n5108), .B(DATAIN[28]), .S(n6019), .Z(n4442) );
  INV_X1 U1712 ( .A(n3579), .ZN(n7483) );
  MUX2_X1 U1713 ( .A(n5107), .B(DATAIN[29]), .S(n6019), .Z(n4443) );
  INV_X1 U1714 ( .A(n3580), .ZN(n7502) );
  MUX2_X1 U1715 ( .A(n5106), .B(DATAIN[30]), .S(n6019), .Z(n4444) );
  INV_X1 U1716 ( .A(n3581), .ZN(n7532) );
  MUX2_X1 U1717 ( .A(n5105), .B(DATAIN[31]), .S(n6019), .Z(n4445) );
  MUX2_X1 U1718 ( .A(n5360), .B(DATAIN[0]), .S(n6020), .Z(n4542) );
  MUX2_X1 U1719 ( .A(n5614), .B(DATAIN[1]), .S(n6020), .Z(n4543) );
  MUX2_X1 U1720 ( .A(n5613), .B(DATAIN[2]), .S(n6020), .Z(n4544) );
  MUX2_X1 U1721 ( .A(n5612), .B(DATAIN[3]), .S(n6020), .Z(n4545) );
  MUX2_X1 U1722 ( .A(n5611), .B(DATAIN[4]), .S(n6020), .Z(n4546) );
  MUX2_X1 U1723 ( .A(n5610), .B(DATAIN[5]), .S(n6020), .Z(n4547) );
  MUX2_X1 U1724 ( .A(n5609), .B(DATAIN[6]), .S(n6020), .Z(n4548) );
  MUX2_X1 U1725 ( .A(n5608), .B(DATAIN[7]), .S(n6020), .Z(n4549) );
  MUX2_X1 U1726 ( .A(n5607), .B(DATAIN[8]), .S(n6020), .Z(n4550) );
  MUX2_X1 U1727 ( .A(n5606), .B(DATAIN[9]), .S(n6020), .Z(n4551) );
  MUX2_X1 U1728 ( .A(n5605), .B(DATAIN[10]), .S(n6020), .Z(n4552) );
  MUX2_X1 U1729 ( .A(n5604), .B(DATAIN[11]), .S(n6020), .Z(n4553) );
  MUX2_X1 U1730 ( .A(n5603), .B(DATAIN[12]), .S(n6021), .Z(n4554) );
  MUX2_X1 U1731 ( .A(n5602), .B(DATAIN[13]), .S(n6021), .Z(n4555) );
  MUX2_X1 U1732 ( .A(n5601), .B(DATAIN[14]), .S(n6021), .Z(n4556) );
  MUX2_X1 U1733 ( .A(n5600), .B(DATAIN[15]), .S(n6021), .Z(n4557) );
  MUX2_X1 U1734 ( .A(n5599), .B(DATAIN[16]), .S(n6021), .Z(n4558) );
  MUX2_X1 U1735 ( .A(n5598), .B(DATAIN[17]), .S(n6021), .Z(n4559) );
  MUX2_X1 U1736 ( .A(n5597), .B(DATAIN[18]), .S(n6021), .Z(n4560) );
  MUX2_X1 U1737 ( .A(n5596), .B(DATAIN[19]), .S(n6021), .Z(n4561) );
  MUX2_X1 U1738 ( .A(n5595), .B(DATAIN[20]), .S(n6021), .Z(n4562) );
  MUX2_X1 U1739 ( .A(n5594), .B(DATAIN[21]), .S(n6021), .Z(n4563) );
  MUX2_X1 U1740 ( .A(n5593), .B(DATAIN[22]), .S(n6021), .Z(n4564) );
  MUX2_X1 U1741 ( .A(n5592), .B(DATAIN[23]), .S(n6021), .Z(n4565) );
  MUX2_X1 U1742 ( .A(n5591), .B(DATAIN[24]), .S(n6022), .Z(n4566) );
  MUX2_X1 U1743 ( .A(n5590), .B(DATAIN[25]), .S(n6022), .Z(n4567) );
  MUX2_X1 U1744 ( .A(n5589), .B(DATAIN[26]), .S(n6022), .Z(n4568) );
  MUX2_X1 U1745 ( .A(n5588), .B(DATAIN[27]), .S(n6022), .Z(n4569) );
  MUX2_X1 U1746 ( .A(n5587), .B(DATAIN[28]), .S(n6022), .Z(n4570) );
  MUX2_X1 U1747 ( .A(n5586), .B(DATAIN[29]), .S(n6022), .Z(n4571) );
  MUX2_X1 U1748 ( .A(n5585), .B(DATAIN[30]), .S(n6022), .Z(n4572) );
  MUX2_X1 U1749 ( .A(n5584), .B(DATAIN[31]), .S(n6022), .Z(n4573) );
  MUX2_X1 U1750 ( .A(n5808), .B(DATAIN[0]), .S(n6023), .Z(n4126) );
  MUX2_X1 U1751 ( .A(n5807), .B(DATAIN[1]), .S(n6023), .Z(n4127) );
  MUX2_X1 U1752 ( .A(n5806), .B(DATAIN[2]), .S(n6023), .Z(n4128) );
  MUX2_X1 U1753 ( .A(n5805), .B(DATAIN[3]), .S(n6023), .Z(n4129) );
  MUX2_X1 U1754 ( .A(n5804), .B(DATAIN[4]), .S(n6023), .Z(n4130) );
  MUX2_X1 U1755 ( .A(n5803), .B(DATAIN[5]), .S(n6023), .Z(n4131) );
  MUX2_X1 U1756 ( .A(n5802), .B(DATAIN[6]), .S(n6023), .Z(n4132) );
  MUX2_X1 U1757 ( .A(n5801), .B(DATAIN[7]), .S(n6023), .Z(n4133) );
  MUX2_X1 U1758 ( .A(n5800), .B(DATAIN[8]), .S(n6023), .Z(n4134) );
  MUX2_X1 U1759 ( .A(n5799), .B(DATAIN[9]), .S(n6023), .Z(n4135) );
  MUX2_X1 U1760 ( .A(n5798), .B(DATAIN[10]), .S(n6023), .Z(n4136) );
  MUX2_X1 U1761 ( .A(n5797), .B(DATAIN[11]), .S(n6023), .Z(n4137) );
  MUX2_X1 U1762 ( .A(n5796), .B(DATAIN[12]), .S(n6024), .Z(n4138) );
  MUX2_X1 U1763 ( .A(n5795), .B(DATAIN[13]), .S(n6024), .Z(n4139) );
  MUX2_X1 U1764 ( .A(n5794), .B(DATAIN[14]), .S(n6024), .Z(n4140) );
  MUX2_X1 U1765 ( .A(n5793), .B(DATAIN[15]), .S(n6024), .Z(n4141) );
  MUX2_X1 U1766 ( .A(n5792), .B(DATAIN[16]), .S(n6024), .Z(n4142) );
  MUX2_X1 U1767 ( .A(n5791), .B(DATAIN[17]), .S(n6024), .Z(n4143) );
  MUX2_X1 U1768 ( .A(n5790), .B(DATAIN[18]), .S(n6024), .Z(n4144) );
  MUX2_X1 U1769 ( .A(n5789), .B(DATAIN[19]), .S(n6024), .Z(n4145) );
  MUX2_X1 U1770 ( .A(n5788), .B(DATAIN[20]), .S(n6024), .Z(n4146) );
  MUX2_X1 U1771 ( .A(n5787), .B(DATAIN[21]), .S(n6024), .Z(n4147) );
  MUX2_X1 U1772 ( .A(n5786), .B(DATAIN[22]), .S(n6024), .Z(n4148) );
  MUX2_X1 U1773 ( .A(n5785), .B(DATAIN[23]), .S(n6024), .Z(n4149) );
  MUX2_X1 U1774 ( .A(n5784), .B(DATAIN[24]), .S(n6025), .Z(n4150) );
  MUX2_X1 U1775 ( .A(n5783), .B(DATAIN[25]), .S(n6025), .Z(n4151) );
  MUX2_X1 U1776 ( .A(n5782), .B(DATAIN[26]), .S(n6025), .Z(n4152) );
  MUX2_X1 U1777 ( .A(n5781), .B(DATAIN[27]), .S(n6025), .Z(n4153) );
  MUX2_X1 U1778 ( .A(n5780), .B(DATAIN[28]), .S(n6025), .Z(n4154) );
  MUX2_X1 U1779 ( .A(n5779), .B(DATAIN[29]), .S(n6025), .Z(n4155) );
  MUX2_X1 U1780 ( .A(n5778), .B(DATAIN[30]), .S(n6025), .Z(n4156) );
  MUX2_X1 U1781 ( .A(n5777), .B(DATAIN[31]), .S(n6025), .Z(n4157) );
  MUX2_X1 U1782 ( .A(n5646), .B(DATAIN[0]), .S(n6026), .Z(n4190) );
  MUX2_X1 U1783 ( .A(n5645), .B(DATAIN[1]), .S(n6026), .Z(n4191) );
  MUX2_X1 U1784 ( .A(n5644), .B(DATAIN[2]), .S(n6026), .Z(n4192) );
  MUX2_X1 U1785 ( .A(n5643), .B(DATAIN[3]), .S(n6026), .Z(n4193) );
  MUX2_X1 U1786 ( .A(n5642), .B(DATAIN[4]), .S(n6026), .Z(n4194) );
  MUX2_X1 U1787 ( .A(n5641), .B(DATAIN[5]), .S(n6026), .Z(n4195) );
  MUX2_X1 U1788 ( .A(n5640), .B(DATAIN[6]), .S(n6026), .Z(n4196) );
  MUX2_X1 U1789 ( .A(n5639), .B(DATAIN[7]), .S(n6026), .Z(n4197) );
  MUX2_X1 U1790 ( .A(n5638), .B(DATAIN[8]), .S(n6026), .Z(n4198) );
  MUX2_X1 U1791 ( .A(n5637), .B(DATAIN[9]), .S(n6026), .Z(n4199) );
  MUX2_X1 U1792 ( .A(n5636), .B(DATAIN[10]), .S(n6026), .Z(n4200) );
  MUX2_X1 U1793 ( .A(n5635), .B(DATAIN[11]), .S(n6026), .Z(n4201) );
  MUX2_X1 U1794 ( .A(n5634), .B(DATAIN[12]), .S(n6027), .Z(n4202) );
  MUX2_X1 U1795 ( .A(n5633), .B(DATAIN[13]), .S(n6027), .Z(n4203) );
  MUX2_X1 U1796 ( .A(n5632), .B(DATAIN[14]), .S(n6027), .Z(n4204) );
  MUX2_X1 U1797 ( .A(n5631), .B(DATAIN[15]), .S(n6027), .Z(n4205) );
  MUX2_X1 U1798 ( .A(n5630), .B(DATAIN[16]), .S(n6027), .Z(n4206) );
  MUX2_X1 U1799 ( .A(n5629), .B(DATAIN[17]), .S(n6027), .Z(n4207) );
  MUX2_X1 U1800 ( .A(n5628), .B(DATAIN[18]), .S(n6027), .Z(n4208) );
  MUX2_X1 U1801 ( .A(n5627), .B(DATAIN[19]), .S(n6027), .Z(n4209) );
  MUX2_X1 U1802 ( .A(n5626), .B(DATAIN[20]), .S(n6027), .Z(n4210) );
  MUX2_X1 U1803 ( .A(n5625), .B(DATAIN[21]), .S(n6027), .Z(n4211) );
  MUX2_X1 U1804 ( .A(n5624), .B(DATAIN[22]), .S(n6027), .Z(n4212) );
  MUX2_X1 U1805 ( .A(n5623), .B(DATAIN[23]), .S(n6027), .Z(n4213) );
  MUX2_X1 U1806 ( .A(n5622), .B(DATAIN[24]), .S(n6028), .Z(n4214) );
  MUX2_X1 U1807 ( .A(n5621), .B(DATAIN[25]), .S(n6028), .Z(n4215) );
  MUX2_X1 U1808 ( .A(n5620), .B(DATAIN[26]), .S(n6028), .Z(n4216) );
  MUX2_X1 U1809 ( .A(n5619), .B(DATAIN[27]), .S(n6028), .Z(n4217) );
  MUX2_X1 U1810 ( .A(n5618), .B(DATAIN[28]), .S(n6028), .Z(n4218) );
  MUX2_X1 U1811 ( .A(n5617), .B(DATAIN[29]), .S(n6028), .Z(n4219) );
  MUX2_X1 U1812 ( .A(n5616), .B(DATAIN[30]), .S(n6028), .Z(n4220) );
  MUX2_X1 U1813 ( .A(n5615), .B(DATAIN[31]), .S(n6028), .Z(n4221) );
  MUX2_X1 U1814 ( .A(n5359), .B(DATAIN[0]), .S(n6029), .Z(n4446) );
  INV_X1 U1815 ( .A(n2943), .ZN(n6951) );
  MUX2_X1 U1816 ( .A(n5202), .B(DATAIN[1]), .S(n6029), .Z(n4447) );
  INV_X1 U1817 ( .A(n2944), .ZN(n6969) );
  MUX2_X1 U1818 ( .A(n5201), .B(DATAIN[2]), .S(n6029), .Z(n4448) );
  INV_X1 U1819 ( .A(n2945), .ZN(n6987) );
  MUX2_X1 U1820 ( .A(n5200), .B(DATAIN[3]), .S(n6029), .Z(n4449) );
  INV_X1 U1821 ( .A(n2946), .ZN(n7006) );
  MUX2_X1 U1822 ( .A(n5199), .B(DATAIN[4]), .S(n6029), .Z(n4450) );
  INV_X1 U1823 ( .A(n2947), .ZN(n7025) );
  MUX2_X1 U1824 ( .A(n5198), .B(DATAIN[5]), .S(n6029), .Z(n4451) );
  INV_X1 U1825 ( .A(n2948), .ZN(n7044) );
  MUX2_X1 U1826 ( .A(n5197), .B(DATAIN[6]), .S(n6029), .Z(n4452) );
  INV_X1 U1827 ( .A(n2949), .ZN(n7063) );
  MUX2_X1 U1828 ( .A(n5196), .B(DATAIN[7]), .S(n6029), .Z(n4453) );
  INV_X1 U1829 ( .A(n2950), .ZN(n7082) );
  MUX2_X1 U1830 ( .A(n5195), .B(DATAIN[8]), .S(n6029), .Z(n4454) );
  INV_X1 U1831 ( .A(n2951), .ZN(n7101) );
  MUX2_X1 U1832 ( .A(n5194), .B(DATAIN[9]), .S(n6029), .Z(n4455) );
  INV_X1 U1833 ( .A(n2952), .ZN(n7120) );
  MUX2_X1 U1834 ( .A(n5193), .B(DATAIN[10]), .S(n6029), .Z(n4456) );
  INV_X1 U1835 ( .A(n2953), .ZN(n7139) );
  MUX2_X1 U1836 ( .A(n5192), .B(DATAIN[11]), .S(n6029), .Z(n4457) );
  INV_X1 U1837 ( .A(n2954), .ZN(n7158) );
  MUX2_X1 U1838 ( .A(n5191), .B(DATAIN[12]), .S(n6030), .Z(n4458) );
  INV_X1 U1839 ( .A(n2955), .ZN(n7177) );
  MUX2_X1 U1840 ( .A(n5190), .B(DATAIN[13]), .S(n6030), .Z(n4459) );
  INV_X1 U1841 ( .A(n2956), .ZN(n7196) );
  MUX2_X1 U1842 ( .A(n5189), .B(DATAIN[14]), .S(n6030), .Z(n4460) );
  INV_X1 U1843 ( .A(n2957), .ZN(n7215) );
  MUX2_X1 U1844 ( .A(n5188), .B(DATAIN[15]), .S(n6030), .Z(n4461) );
  INV_X1 U1845 ( .A(n2958), .ZN(n7234) );
  MUX2_X1 U1846 ( .A(n5187), .B(DATAIN[16]), .S(n6030), .Z(n4462) );
  INV_X1 U1847 ( .A(n2959), .ZN(n7253) );
  MUX2_X1 U1848 ( .A(n5186), .B(DATAIN[17]), .S(n6030), .Z(n4463) );
  INV_X1 U1849 ( .A(n2960), .ZN(n7272) );
  MUX2_X1 U1850 ( .A(n5185), .B(DATAIN[18]), .S(n6030), .Z(n4464) );
  INV_X1 U1851 ( .A(n2961), .ZN(n7291) );
  MUX2_X1 U1852 ( .A(n5184), .B(DATAIN[19]), .S(n6030), .Z(n4465) );
  INV_X1 U1853 ( .A(n2962), .ZN(n7310) );
  MUX2_X1 U1854 ( .A(n5183), .B(DATAIN[20]), .S(n6030), .Z(n4466) );
  INV_X1 U1855 ( .A(n2963), .ZN(n7329) );
  MUX2_X1 U1856 ( .A(n5182), .B(DATAIN[21]), .S(n6030), .Z(n4467) );
  INV_X1 U1857 ( .A(n2964), .ZN(n7348) );
  MUX2_X1 U1858 ( .A(n5181), .B(DATAIN[22]), .S(n6030), .Z(n4468) );
  INV_X1 U1859 ( .A(n2965), .ZN(n7367) );
  MUX2_X1 U1860 ( .A(n5180), .B(DATAIN[23]), .S(n6030), .Z(n4469) );
  INV_X1 U1861 ( .A(n2966), .ZN(n7386) );
  MUX2_X1 U1862 ( .A(n5179), .B(DATAIN[24]), .S(n6031), .Z(n4470) );
  INV_X1 U1863 ( .A(n2967), .ZN(n7405) );
  MUX2_X1 U1864 ( .A(n5178), .B(DATAIN[25]), .S(n6031), .Z(n4471) );
  INV_X1 U1865 ( .A(n2968), .ZN(n7424) );
  MUX2_X1 U1866 ( .A(n5177), .B(DATAIN[26]), .S(n6031), .Z(n4472) );
  INV_X1 U1867 ( .A(n2969), .ZN(n7443) );
  MUX2_X1 U1868 ( .A(n5176), .B(DATAIN[27]), .S(n6031), .Z(n4473) );
  INV_X1 U1869 ( .A(n2970), .ZN(n7462) );
  MUX2_X1 U1870 ( .A(n5175), .B(DATAIN[28]), .S(n6031), .Z(n4474) );
  INV_X1 U1871 ( .A(n2971), .ZN(n7481) );
  MUX2_X1 U1872 ( .A(n5174), .B(DATAIN[29]), .S(n6031), .Z(n4475) );
  INV_X1 U1873 ( .A(n2972), .ZN(n7500) );
  MUX2_X1 U1874 ( .A(n5173), .B(DATAIN[30]), .S(n6031), .Z(n4476) );
  INV_X1 U1875 ( .A(n2973), .ZN(n7526) );
  MUX2_X1 U1876 ( .A(n5172), .B(DATAIN[31]), .S(n6031), .Z(n4477) );
  NAND2_X1 U1877 ( .A1(n4606), .A2(n4611), .ZN(n6483) );
  INV_X1 U1878 ( .A(n6483), .ZN(n6484) );
  OAI22_X1 U1879 ( .A1(n6034), .A2(n5908), .B1(n6339), .B2(n6483), .ZN(n4574)
         );
  OAI22_X1 U1880 ( .A1(n6034), .A2(n5879), .B1(n6341), .B2(n6483), .ZN(n4575)
         );
  OAI22_X1 U1881 ( .A1(n6034), .A2(n5878), .B1(n6343), .B2(n6483), .ZN(n4576)
         );
  OAI22_X1 U1882 ( .A1(n6034), .A2(n5877), .B1(n6345), .B2(n6483), .ZN(n4577)
         );
  MUX2_X1 U1883 ( .A(n5514), .B(DATAIN[4]), .S(n6034), .Z(n4578) );
  MUX2_X1 U1884 ( .A(n5513), .B(DATAIN[5]), .S(n6034), .Z(n4579) );
  MUX2_X1 U1885 ( .A(n5512), .B(DATAIN[6]), .S(n6034), .Z(n4580) );
  MUX2_X1 U1886 ( .A(n5511), .B(DATAIN[7]), .S(n6034), .Z(n4581) );
  MUX2_X1 U1887 ( .A(n5510), .B(DATAIN[8]), .S(n6033), .Z(n4582) );
  MUX2_X1 U1888 ( .A(n5509), .B(DATAIN[9]), .S(n6033), .Z(n4583) );
  MUX2_X1 U1889 ( .A(n5508), .B(DATAIN[10]), .S(n6033), .Z(n4584) );
  MUX2_X1 U1890 ( .A(n5507), .B(DATAIN[11]), .S(n6033), .Z(n4585) );
  MUX2_X1 U1891 ( .A(n5506), .B(DATAIN[12]), .S(n6033), .Z(n4586) );
  MUX2_X1 U1892 ( .A(n5505), .B(DATAIN[13]), .S(n6033), .Z(n4587) );
  MUX2_X1 U1893 ( .A(n5504), .B(DATAIN[14]), .S(n6033), .Z(n4588) );
  MUX2_X1 U1894 ( .A(n5503), .B(DATAIN[15]), .S(n6033), .Z(n4589) );
  MUX2_X1 U1895 ( .A(n5502), .B(DATAIN[16]), .S(n6033), .Z(n4590) );
  MUX2_X1 U1896 ( .A(n5501), .B(DATAIN[17]), .S(n6033), .Z(n4591) );
  MUX2_X1 U1897 ( .A(n5500), .B(DATAIN[18]), .S(n6033), .Z(n4592) );
  MUX2_X1 U1898 ( .A(n5499), .B(DATAIN[19]), .S(n6033), .Z(n4593) );
  MUX2_X1 U1899 ( .A(n5498), .B(DATAIN[20]), .S(n6032), .Z(n4594) );
  MUX2_X1 U1900 ( .A(n5497), .B(DATAIN[21]), .S(n6032), .Z(n4595) );
  MUX2_X1 U1901 ( .A(n5496), .B(DATAIN[22]), .S(n6032), .Z(n4596) );
  MUX2_X1 U1902 ( .A(n5495), .B(DATAIN[23]), .S(n6032), .Z(n4597) );
  MUX2_X1 U1903 ( .A(n5494), .B(DATAIN[24]), .S(n6032), .Z(n4598) );
  MUX2_X1 U1904 ( .A(n5493), .B(DATAIN[25]), .S(n6032), .Z(n4599) );
  MUX2_X1 U1905 ( .A(n5492), .B(DATAIN[26]), .S(n6032), .Z(n4600) );
  MUX2_X1 U1906 ( .A(n5491), .B(DATAIN[27]), .S(n6032), .Z(n4601) );
  MUX2_X1 U1907 ( .A(n5490), .B(DATAIN[28]), .S(n6032), .Z(n4602) );
  MUX2_X1 U1908 ( .A(n5489), .B(DATAIN[29]), .S(n6032), .Z(n4603) );
  MUX2_X1 U1909 ( .A(n5488), .B(DATAIN[30]), .S(n6032), .Z(n4604) );
  MUX2_X1 U1910 ( .A(n5487), .B(DATAIN[31]), .S(n6032), .Z(n4605) );
  MUX2_X1 U1911 ( .A(n5840), .B(DATAIN[0]), .S(n6035), .Z(n4318) );
  MUX2_X1 U1912 ( .A(n5839), .B(DATAIN[1]), .S(n6035), .Z(n4319) );
  MUX2_X1 U1913 ( .A(n5838), .B(DATAIN[2]), .S(n6035), .Z(n4320) );
  MUX2_X1 U1914 ( .A(n5837), .B(DATAIN[3]), .S(n6035), .Z(n4321) );
  MUX2_X1 U1915 ( .A(n5836), .B(DATAIN[4]), .S(n6035), .Z(n4322) );
  MUX2_X1 U1916 ( .A(n5835), .B(DATAIN[5]), .S(n6035), .Z(n4323) );
  MUX2_X1 U1917 ( .A(n5834), .B(DATAIN[6]), .S(n6035), .Z(n4324) );
  MUX2_X1 U1918 ( .A(n5833), .B(DATAIN[7]), .S(n6035), .Z(n4325) );
  MUX2_X1 U1919 ( .A(n5832), .B(DATAIN[8]), .S(n6035), .Z(n4326) );
  MUX2_X1 U1920 ( .A(n5831), .B(DATAIN[9]), .S(n6035), .Z(n4327) );
  MUX2_X1 U1921 ( .A(n5830), .B(DATAIN[10]), .S(n6035), .Z(n4328) );
  MUX2_X1 U1922 ( .A(n5829), .B(DATAIN[11]), .S(n6035), .Z(n4329) );
  MUX2_X1 U1923 ( .A(n5828), .B(DATAIN[12]), .S(n6036), .Z(n4330) );
  MUX2_X1 U1924 ( .A(n5827), .B(DATAIN[13]), .S(n6036), .Z(n4331) );
  MUX2_X1 U1925 ( .A(n5826), .B(DATAIN[14]), .S(n6036), .Z(n4332) );
  MUX2_X1 U1926 ( .A(n5825), .B(DATAIN[15]), .S(n6036), .Z(n4333) );
  MUX2_X1 U1927 ( .A(n5824), .B(DATAIN[16]), .S(n6036), .Z(n4334) );
  MUX2_X1 U1928 ( .A(n5823), .B(DATAIN[17]), .S(n6036), .Z(n4335) );
  MUX2_X1 U1929 ( .A(n5822), .B(DATAIN[18]), .S(n6036), .Z(n4336) );
  MUX2_X1 U1930 ( .A(n5821), .B(DATAIN[19]), .S(n6036), .Z(n4337) );
  MUX2_X1 U1931 ( .A(n5820), .B(DATAIN[20]), .S(n6036), .Z(n4338) );
  MUX2_X1 U1932 ( .A(n5819), .B(DATAIN[21]), .S(n6036), .Z(n4339) );
  MUX2_X1 U1933 ( .A(n5818), .B(DATAIN[22]), .S(n6036), .Z(n4340) );
  MUX2_X1 U1934 ( .A(n5817), .B(DATAIN[23]), .S(n6036), .Z(n4341) );
  MUX2_X1 U1935 ( .A(n5816), .B(DATAIN[24]), .S(n6037), .Z(n4342) );
  MUX2_X1 U1936 ( .A(n5815), .B(DATAIN[25]), .S(n6037), .Z(n4343) );
  MUX2_X1 U1937 ( .A(n5814), .B(DATAIN[26]), .S(n6037), .Z(n4344) );
  MUX2_X1 U1938 ( .A(n5813), .B(DATAIN[27]), .S(n6037), .Z(n4345) );
  MUX2_X1 U1939 ( .A(n5812), .B(DATAIN[28]), .S(n6037), .Z(n4346) );
  MUX2_X1 U1940 ( .A(n5811), .B(DATAIN[29]), .S(n6037), .Z(n4347) );
  MUX2_X1 U1941 ( .A(n5810), .B(DATAIN[30]), .S(n6037), .Z(n4348) );
  MUX2_X1 U1942 ( .A(n5809), .B(DATAIN[31]), .S(n6037), .Z(n4349) );
  INV_X1 U1943 ( .A(n2252), .ZN(n6942) );
  MUX2_X1 U1944 ( .A(n5233), .B(DATAIN[0]), .S(n6038), .Z(n4382) );
  MUX2_X1 U1945 ( .A(n5390), .B(DATAIN[1]), .S(n6038), .Z(n4383) );
  MUX2_X1 U1946 ( .A(n5389), .B(DATAIN[2]), .S(n6038), .Z(n4384) );
  MUX2_X1 U1947 ( .A(n5388), .B(DATAIN[3]), .S(n6038), .Z(n4385) );
  MUX2_X1 U1948 ( .A(n5387), .B(DATAIN[4]), .S(n6038), .Z(n4386) );
  MUX2_X1 U1949 ( .A(n5386), .B(DATAIN[5]), .S(n6038), .Z(n4387) );
  MUX2_X1 U1950 ( .A(n5385), .B(DATAIN[6]), .S(n6038), .Z(n4388) );
  MUX2_X1 U1951 ( .A(n5384), .B(DATAIN[7]), .S(n6038), .Z(n4389) );
  MUX2_X1 U1952 ( .A(n5383), .B(DATAIN[8]), .S(n6038), .Z(n4390) );
  MUX2_X1 U1953 ( .A(n5382), .B(DATAIN[9]), .S(n6038), .Z(n4391) );
  MUX2_X1 U1954 ( .A(n5381), .B(DATAIN[10]), .S(n6038), .Z(n4392) );
  MUX2_X1 U1955 ( .A(n5380), .B(DATAIN[11]), .S(n6038), .Z(n4393) );
  MUX2_X1 U1956 ( .A(n5379), .B(DATAIN[12]), .S(n6039), .Z(n4394) );
  MUX2_X1 U1957 ( .A(n5378), .B(DATAIN[13]), .S(n6039), .Z(n4395) );
  MUX2_X1 U1958 ( .A(n5377), .B(DATAIN[14]), .S(n6039), .Z(n4396) );
  MUX2_X1 U1959 ( .A(n5376), .B(DATAIN[15]), .S(n6039), .Z(n4397) );
  MUX2_X1 U1960 ( .A(n5375), .B(DATAIN[16]), .S(n6039), .Z(n4398) );
  MUX2_X1 U1961 ( .A(n5374), .B(DATAIN[17]), .S(n6039), .Z(n4399) );
  MUX2_X1 U1962 ( .A(n5373), .B(DATAIN[18]), .S(n6039), .Z(n4400) );
  MUX2_X1 U1963 ( .A(n5372), .B(DATAIN[19]), .S(n6039), .Z(n4401) );
  MUX2_X1 U1964 ( .A(n5371), .B(DATAIN[20]), .S(n6039), .Z(n4402) );
  MUX2_X1 U1965 ( .A(n5370), .B(DATAIN[21]), .S(n6039), .Z(n4403) );
  MUX2_X1 U1966 ( .A(n5369), .B(DATAIN[22]), .S(n6039), .Z(n4404) );
  MUX2_X1 U1967 ( .A(n5368), .B(DATAIN[23]), .S(n6039), .Z(n4405) );
  MUX2_X1 U1968 ( .A(n5367), .B(DATAIN[24]), .S(n6040), .Z(n4406) );
  MUX2_X1 U1969 ( .A(n5366), .B(DATAIN[25]), .S(n6040), .Z(n4407) );
  MUX2_X1 U1970 ( .A(n5365), .B(DATAIN[26]), .S(n6040), .Z(n4408) );
  MUX2_X1 U1971 ( .A(n5364), .B(DATAIN[27]), .S(n6040), .Z(n4409) );
  MUX2_X1 U1972 ( .A(n5363), .B(DATAIN[28]), .S(n6040), .Z(n4410) );
  MUX2_X1 U1973 ( .A(n5362), .B(DATAIN[29]), .S(n6040), .Z(n4411) );
  MUX2_X1 U1974 ( .A(n5361), .B(DATAIN[30]), .S(n6040), .Z(n4412) );
  INV_X1 U1975 ( .A(n2283), .ZN(n7540) );
  MUX2_X1 U1976 ( .A(n5168), .B(DATAIN[31]), .S(n6040), .Z(n4413) );
  MUX2_X1 U1977 ( .A(n5648), .B(DATAIN[0]), .S(n6041), .Z(n4478) );
  MUX2_X1 U1978 ( .A(n5679), .B(DATAIN[1]), .S(n6041), .Z(n4479) );
  MUX2_X1 U1979 ( .A(n5678), .B(DATAIN[2]), .S(n6041), .Z(n4480) );
  MUX2_X1 U1980 ( .A(n5677), .B(DATAIN[3]), .S(n6041), .Z(n4481) );
  MUX2_X1 U1981 ( .A(n5676), .B(DATAIN[4]), .S(n6041), .Z(n4482) );
  MUX2_X1 U1982 ( .A(n5675), .B(DATAIN[5]), .S(n6041), .Z(n4483) );
  MUX2_X1 U1983 ( .A(n5674), .B(DATAIN[6]), .S(n6041), .Z(n4484) );
  MUX2_X1 U1984 ( .A(n5673), .B(DATAIN[7]), .S(n6041), .Z(n4485) );
  MUX2_X1 U1985 ( .A(n5672), .B(DATAIN[8]), .S(n6041), .Z(n4486) );
  MUX2_X1 U1986 ( .A(n5671), .B(DATAIN[9]), .S(n6041), .Z(n4487) );
  MUX2_X1 U1987 ( .A(n5670), .B(DATAIN[10]), .S(n6041), .Z(n4488) );
  MUX2_X1 U1988 ( .A(n5669), .B(DATAIN[11]), .S(n6041), .Z(n4489) );
  MUX2_X1 U1989 ( .A(n5668), .B(DATAIN[12]), .S(n6042), .Z(n4490) );
  MUX2_X1 U1990 ( .A(n5667), .B(DATAIN[13]), .S(n6042), .Z(n4491) );
  MUX2_X1 U1991 ( .A(n5666), .B(DATAIN[14]), .S(n6042), .Z(n4492) );
  MUX2_X1 U1992 ( .A(n5665), .B(DATAIN[15]), .S(n6042), .Z(n4493) );
  MUX2_X1 U1993 ( .A(n5664), .B(DATAIN[16]), .S(n6042), .Z(n4494) );
  MUX2_X1 U1994 ( .A(n5663), .B(DATAIN[17]), .S(n6042), .Z(n4495) );
  MUX2_X1 U1995 ( .A(n5662), .B(DATAIN[18]), .S(n6042), .Z(n4496) );
  MUX2_X1 U1996 ( .A(n5661), .B(DATAIN[19]), .S(n6042), .Z(n4497) );
  MUX2_X1 U1997 ( .A(n5660), .B(DATAIN[20]), .S(n6042), .Z(n4498) );
  MUX2_X1 U1998 ( .A(n5659), .B(DATAIN[21]), .S(n6042), .Z(n4499) );
  MUX2_X1 U1999 ( .A(n5658), .B(DATAIN[22]), .S(n6042), .Z(n4500) );
  MUX2_X1 U2000 ( .A(n5657), .B(DATAIN[23]), .S(n6042), .Z(n4501) );
  MUX2_X1 U2001 ( .A(n5656), .B(DATAIN[24]), .S(n6043), .Z(n4502) );
  MUX2_X1 U2002 ( .A(n5655), .B(DATAIN[25]), .S(n6043), .Z(n4503) );
  MUX2_X1 U2003 ( .A(n5654), .B(DATAIN[26]), .S(n6043), .Z(n4504) );
  MUX2_X1 U2004 ( .A(n5653), .B(DATAIN[27]), .S(n6043), .Z(n4505) );
  MUX2_X1 U2005 ( .A(n5652), .B(DATAIN[28]), .S(n6043), .Z(n4506) );
  MUX2_X1 U2006 ( .A(n5651), .B(DATAIN[29]), .S(n6043), .Z(n4507) );
  MUX2_X1 U2007 ( .A(n5650), .B(DATAIN[30]), .S(n6043), .Z(n4508) );
  MUX2_X1 U2008 ( .A(n5649), .B(DATAIN[31]), .S(n6043), .Z(n4509) );
  MUX2_X1 U2009 ( .A(n5876), .B(DATAIN[0]), .S(n6044), .Z(n4286) );
  MUX2_X1 U2010 ( .A(n5327), .B(DATAIN[1]), .S(n6044), .Z(n4287) );
  MUX2_X1 U2011 ( .A(n5326), .B(DATAIN[2]), .S(n6044), .Z(n4288) );
  MUX2_X1 U2012 ( .A(n5325), .B(DATAIN[3]), .S(n6044), .Z(n4289) );
  MUX2_X1 U2013 ( .A(n5324), .B(DATAIN[4]), .S(n6044), .Z(n4290) );
  MUX2_X1 U2014 ( .A(n5323), .B(DATAIN[5]), .S(n6044), .Z(n4291) );
  MUX2_X1 U2015 ( .A(n5322), .B(DATAIN[6]), .S(n6044), .Z(n4292) );
  MUX2_X1 U2016 ( .A(n5321), .B(DATAIN[7]), .S(n6044), .Z(n4293) );
  MUX2_X1 U2017 ( .A(n5320), .B(DATAIN[8]), .S(n6044), .Z(n4294) );
  MUX2_X1 U2018 ( .A(n5319), .B(DATAIN[9]), .S(n6044), .Z(n4295) );
  MUX2_X1 U2019 ( .A(n5318), .B(DATAIN[10]), .S(n6044), .Z(n4296) );
  MUX2_X1 U2020 ( .A(n5317), .B(DATAIN[11]), .S(n6044), .Z(n4297) );
  MUX2_X1 U2021 ( .A(n5316), .B(DATAIN[12]), .S(n6045), .Z(n4298) );
  MUX2_X1 U2022 ( .A(n5315), .B(DATAIN[13]), .S(n6045), .Z(n4299) );
  MUX2_X1 U2023 ( .A(n5314), .B(DATAIN[14]), .S(n6045), .Z(n4300) );
  MUX2_X1 U2024 ( .A(n5313), .B(DATAIN[15]), .S(n6045), .Z(n4301) );
  MUX2_X1 U2025 ( .A(n5312), .B(DATAIN[16]), .S(n6045), .Z(n4302) );
  MUX2_X1 U2026 ( .A(n5311), .B(DATAIN[17]), .S(n6045), .Z(n4303) );
  MUX2_X1 U2027 ( .A(n5310), .B(DATAIN[18]), .S(n6045), .Z(n4304) );
  MUX2_X1 U2028 ( .A(n5309), .B(DATAIN[19]), .S(n6045), .Z(n4305) );
  MUX2_X1 U2029 ( .A(n5308), .B(DATAIN[20]), .S(n6045), .Z(n4306) );
  MUX2_X1 U2030 ( .A(n5307), .B(DATAIN[21]), .S(n6045), .Z(n4307) );
  MUX2_X1 U2031 ( .A(n5306), .B(DATAIN[22]), .S(n6045), .Z(n4308) );
  MUX2_X1 U2032 ( .A(n5305), .B(DATAIN[23]), .S(n6045), .Z(n4309) );
  MUX2_X1 U2033 ( .A(n5304), .B(DATAIN[24]), .S(n6046), .Z(n4310) );
  MUX2_X1 U2034 ( .A(n5303), .B(DATAIN[25]), .S(n6046), .Z(n4311) );
  MUX2_X1 U2035 ( .A(n5302), .B(DATAIN[26]), .S(n6046), .Z(n4312) );
  MUX2_X1 U2036 ( .A(n5301), .B(DATAIN[27]), .S(n6046), .Z(n4313) );
  MUX2_X1 U2037 ( .A(n5300), .B(DATAIN[28]), .S(n6046), .Z(n4314) );
  MUX2_X1 U2038 ( .A(n5299), .B(DATAIN[29]), .S(n6046), .Z(n4315) );
  MUX2_X1 U2039 ( .A(n5298), .B(DATAIN[30]), .S(n6046), .Z(n4316) );
  MUX2_X1 U2040 ( .A(n5875), .B(DATAIN[31]), .S(n6046), .Z(n4317) );
  MUX2_X1 U2041 ( .A(n5546), .B(DATAIN[0]), .S(n6047), .Z(n4510) );
  MUX2_X1 U2042 ( .A(n5421), .B(DATAIN[1]), .S(n6047), .Z(n4511) );
  MUX2_X1 U2043 ( .A(n5420), .B(DATAIN[2]), .S(n6047), .Z(n4512) );
  MUX2_X1 U2044 ( .A(n5419), .B(DATAIN[3]), .S(n6047), .Z(n4513) );
  MUX2_X1 U2045 ( .A(n5418), .B(DATAIN[4]), .S(n6047), .Z(n4514) );
  MUX2_X1 U2046 ( .A(n5417), .B(DATAIN[5]), .S(n6047), .Z(n4515) );
  MUX2_X1 U2047 ( .A(n5416), .B(DATAIN[6]), .S(n6047), .Z(n4516) );
  MUX2_X1 U2048 ( .A(n5415), .B(DATAIN[7]), .S(n6047), .Z(n4517) );
  MUX2_X1 U2049 ( .A(n5414), .B(DATAIN[8]), .S(n6047), .Z(n4518) );
  MUX2_X1 U2050 ( .A(n5413), .B(DATAIN[9]), .S(n6047), .Z(n4519) );
  MUX2_X1 U2051 ( .A(n5412), .B(DATAIN[10]), .S(n6047), .Z(n4520) );
  MUX2_X1 U2052 ( .A(n5411), .B(DATAIN[11]), .S(n6047), .Z(n4521) );
  MUX2_X1 U2053 ( .A(n5410), .B(DATAIN[12]), .S(n6048), .Z(n4522) );
  MUX2_X1 U2054 ( .A(n5409), .B(DATAIN[13]), .S(n6048), .Z(n4523) );
  MUX2_X1 U2055 ( .A(n5408), .B(DATAIN[14]), .S(n6048), .Z(n4524) );
  MUX2_X1 U2056 ( .A(n5407), .B(DATAIN[15]), .S(n6048), .Z(n4525) );
  MUX2_X1 U2057 ( .A(n5406), .B(DATAIN[16]), .S(n6048), .Z(n4526) );
  MUX2_X1 U2058 ( .A(n5405), .B(DATAIN[17]), .S(n6048), .Z(n4527) );
  MUX2_X1 U2059 ( .A(n5404), .B(DATAIN[18]), .S(n6048), .Z(n4528) );
  MUX2_X1 U2060 ( .A(n5403), .B(DATAIN[19]), .S(n6048), .Z(n4529) );
  MUX2_X1 U2061 ( .A(n5402), .B(DATAIN[20]), .S(n6048), .Z(n4530) );
  MUX2_X1 U2062 ( .A(n5401), .B(DATAIN[21]), .S(n6048), .Z(n4531) );
  MUX2_X1 U2063 ( .A(n5400), .B(DATAIN[22]), .S(n6048), .Z(n4532) );
  MUX2_X1 U2064 ( .A(n5399), .B(DATAIN[23]), .S(n6048), .Z(n4533) );
  MUX2_X1 U2065 ( .A(n5398), .B(DATAIN[24]), .S(n6049), .Z(n4534) );
  MUX2_X1 U2066 ( .A(n5397), .B(DATAIN[25]), .S(n6049), .Z(n4535) );
  MUX2_X1 U2067 ( .A(n5396), .B(DATAIN[26]), .S(n6049), .Z(n4536) );
  MUX2_X1 U2068 ( .A(n5395), .B(DATAIN[27]), .S(n6049), .Z(n4537) );
  MUX2_X1 U2069 ( .A(n5394), .B(DATAIN[28]), .S(n6049), .Z(n4538) );
  MUX2_X1 U2070 ( .A(n5393), .B(DATAIN[29]), .S(n6049), .Z(n4539) );
  MUX2_X1 U2071 ( .A(n5392), .B(DATAIN[30]), .S(n6049), .Z(n4540) );
  MUX2_X1 U2072 ( .A(n5391), .B(DATAIN[31]), .S(n6049), .Z(n4541) );
  MUX2_X1 U2073 ( .A(n5744), .B(DATAIN[31]), .S(n6250), .Z(n3302) );
  MUX2_X1 U2074 ( .A(n5358), .B(DATAIN[0]), .S(n6050), .Z(n3079) );
  MUX2_X1 U2075 ( .A(n5711), .B(DATAIN[1]), .S(n6050), .Z(n3080) );
  MUX2_X1 U2076 ( .A(n5710), .B(DATAIN[2]), .S(n6050), .Z(n3081) );
  MUX2_X1 U2077 ( .A(n5709), .B(DATAIN[3]), .S(n6050), .Z(n3082) );
  MUX2_X1 U2078 ( .A(n5708), .B(DATAIN[4]), .S(n6050), .Z(n3083) );
  MUX2_X1 U2079 ( .A(n5707), .B(DATAIN[5]), .S(n6050), .Z(n3084) );
  MUX2_X1 U2080 ( .A(n5706), .B(DATAIN[6]), .S(n6050), .Z(n3085) );
  MUX2_X1 U2081 ( .A(n5705), .B(DATAIN[7]), .S(n6050), .Z(n3086) );
  MUX2_X1 U2082 ( .A(n5704), .B(DATAIN[8]), .S(n6050), .Z(n3087) );
  MUX2_X1 U2083 ( .A(n5703), .B(DATAIN[9]), .S(n6050), .Z(n3088) );
  MUX2_X1 U2084 ( .A(n5702), .B(DATAIN[10]), .S(n6050), .Z(n3089) );
  MUX2_X1 U2085 ( .A(n5701), .B(DATAIN[11]), .S(n6050), .Z(n3090) );
  MUX2_X1 U2086 ( .A(n5700), .B(DATAIN[12]), .S(n6051), .Z(n3091) );
  MUX2_X1 U2087 ( .A(n5699), .B(DATAIN[13]), .S(n6051), .Z(n3092) );
  MUX2_X1 U2088 ( .A(n5698), .B(DATAIN[14]), .S(n6051), .Z(n3093) );
  MUX2_X1 U2089 ( .A(n5697), .B(DATAIN[15]), .S(n6051), .Z(n3094) );
  MUX2_X1 U2090 ( .A(n5696), .B(DATAIN[16]), .S(n6051), .Z(n3095) );
  MUX2_X1 U2091 ( .A(n5695), .B(DATAIN[17]), .S(n6051), .Z(n3096) );
  MUX2_X1 U2092 ( .A(n5694), .B(DATAIN[18]), .S(n6051), .Z(n3097) );
  MUX2_X1 U2093 ( .A(n5693), .B(DATAIN[19]), .S(n6051), .Z(n3098) );
  MUX2_X1 U2094 ( .A(n5692), .B(DATAIN[20]), .S(n6051), .Z(n3099) );
  MUX2_X1 U2095 ( .A(n5691), .B(DATAIN[21]), .S(n6051), .Z(n3100) );
  MUX2_X1 U2096 ( .A(n5690), .B(DATAIN[22]), .S(n6051), .Z(n3101) );
  MUX2_X1 U2097 ( .A(n5689), .B(DATAIN[23]), .S(n6051), .Z(n3102) );
  MUX2_X1 U2098 ( .A(n5688), .B(DATAIN[24]), .S(n6052), .Z(n3103) );
  MUX2_X1 U2099 ( .A(n5687), .B(DATAIN[25]), .S(n6052), .Z(n3104) );
  MUX2_X1 U2100 ( .A(n5686), .B(DATAIN[26]), .S(n6052), .Z(n3105) );
  MUX2_X1 U2101 ( .A(n5685), .B(DATAIN[27]), .S(n6052), .Z(n3106) );
  MUX2_X1 U2102 ( .A(n5684), .B(DATAIN[28]), .S(n6052), .Z(n3107) );
  MUX2_X1 U2103 ( .A(n5683), .B(DATAIN[29]), .S(n6052), .Z(n3108) );
  MUX2_X1 U2104 ( .A(n5682), .B(DATAIN[30]), .S(n6052), .Z(n3109) );
  MUX2_X1 U2105 ( .A(n5681), .B(DATAIN[31]), .S(n6052), .Z(n3110) );
  NAND2_X1 U2106 ( .A1(n6489), .A2(n4619), .ZN(n6486) );
  OAI22_X1 U2107 ( .A1(n6056), .A2(n5974), .B1(n6340), .B2(n6057), .ZN(n7837)
         );
  OAI22_X1 U2108 ( .A1(n6055), .A2(n6004), .B1(n6342), .B2(n6057), .ZN(n7836)
         );
  OAI22_X1 U2109 ( .A1(n6056), .A2(n6003), .B1(n6344), .B2(n6057), .ZN(n7835)
         );
  OAI22_X1 U2110 ( .A1(n6055), .A2(n6002), .B1(n6346), .B2(n6057), .ZN(n7834)
         );
  OAI22_X1 U2111 ( .A1(n6056), .A2(n6001), .B1(n6347), .B2(n6058), .ZN(n7833)
         );
  OAI22_X1 U2112 ( .A1(n6055), .A2(n6000), .B1(n6348), .B2(n6058), .ZN(n7832)
         );
  OAI22_X1 U2113 ( .A1(n6056), .A2(n5999), .B1(n6349), .B2(n6058), .ZN(n7831)
         );
  OAI22_X1 U2114 ( .A1(n6055), .A2(n5998), .B1(n6350), .B2(n6058), .ZN(n7830)
         );
  OAI22_X1 U2115 ( .A1(n6056), .A2(n5997), .B1(n6351), .B2(n6058), .ZN(n7829)
         );
  OAI22_X1 U2116 ( .A1(n6056), .A2(n5996), .B1(n6352), .B2(n6058), .ZN(n7828)
         );
  OAI22_X1 U2117 ( .A1(n6056), .A2(n5995), .B1(n6353), .B2(n6058), .ZN(n7827)
         );
  OAI22_X1 U2118 ( .A1(n6056), .A2(n5994), .B1(n6354), .B2(n6059), .ZN(n7826)
         );
  OAI22_X1 U2119 ( .A1(n6056), .A2(n5993), .B1(n6355), .B2(n6059), .ZN(n7825)
         );
  OAI22_X1 U2120 ( .A1(n6056), .A2(n5992), .B1(n6356), .B2(n6059), .ZN(n7824)
         );
  OAI22_X1 U2121 ( .A1(n6056), .A2(n5991), .B1(n6357), .B2(n6059), .ZN(n7823)
         );
  OAI22_X1 U2122 ( .A1(n6056), .A2(n5990), .B1(n6358), .B2(n6059), .ZN(n7822)
         );
  OAI22_X1 U2123 ( .A1(n6056), .A2(n5989), .B1(n6359), .B2(n6059), .ZN(n7821)
         );
  OAI22_X1 U2124 ( .A1(n6056), .A2(n5988), .B1(n6360), .B2(n6059), .ZN(n7820)
         );
  OAI22_X1 U2125 ( .A1(n6056), .A2(n5987), .B1(n6361), .B2(n6060), .ZN(n7819)
         );
  OAI22_X1 U2126 ( .A1(n6056), .A2(n5986), .B1(n6362), .B2(n6060), .ZN(n7818)
         );
  OAI22_X1 U2127 ( .A1(n6055), .A2(n5985), .B1(n6363), .B2(n6060), .ZN(n7817)
         );
  OAI22_X1 U2128 ( .A1(n6055), .A2(n5984), .B1(n6364), .B2(n6060), .ZN(n7816)
         );
  OAI22_X1 U2129 ( .A1(n6055), .A2(n5983), .B1(n6365), .B2(n6060), .ZN(n7815)
         );
  OAI22_X1 U2130 ( .A1(n6055), .A2(n5982), .B1(n6366), .B2(n6060), .ZN(n7814)
         );
  OAI22_X1 U2131 ( .A1(n6055), .A2(n5981), .B1(n6367), .B2(n6060), .ZN(n7813)
         );
  OAI22_X1 U2132 ( .A1(n6055), .A2(n5980), .B1(n6368), .B2(n6061), .ZN(n7812)
         );
  OAI22_X1 U2133 ( .A1(n6055), .A2(n5979), .B1(n6369), .B2(n6061), .ZN(n7811)
         );
  OAI22_X1 U2134 ( .A1(n6055), .A2(n5978), .B1(n6370), .B2(n6061), .ZN(n7810)
         );
  OAI22_X1 U2135 ( .A1(n6055), .A2(n5977), .B1(n6371), .B2(n6061), .ZN(n7809)
         );
  OAI22_X1 U2136 ( .A1(n6055), .A2(n5976), .B1(n6372), .B2(n6061), .ZN(n7808)
         );
  OAI22_X1 U2137 ( .A1(n6055), .A2(n5975), .B1(n6373), .B2(n6061), .ZN(n7807)
         );
  OAI22_X1 U2138 ( .A1(n6055), .A2(n5973), .B1(n6374), .B2(n6061), .ZN(n7806)
         );
  NAND2_X1 U2139 ( .A1(n6489), .A2(n4620), .ZN(n6487) );
  OAI22_X1 U2140 ( .A1(n6065), .A2(n5910), .B1(n6340), .B2(n6066), .ZN(n7805)
         );
  OAI22_X1 U2141 ( .A1(n6064), .A2(n5940), .B1(n6342), .B2(n6066), .ZN(n7804)
         );
  OAI22_X1 U2142 ( .A1(n6065), .A2(n5939), .B1(n6344), .B2(n6066), .ZN(n7803)
         );
  OAI22_X1 U2143 ( .A1(n6064), .A2(n5938), .B1(n6346), .B2(n6066), .ZN(n7802)
         );
  OAI22_X1 U2144 ( .A1(n6065), .A2(n5937), .B1(n6347), .B2(n6067), .ZN(n7801)
         );
  OAI22_X1 U2145 ( .A1(n6064), .A2(n5936), .B1(n6348), .B2(n6067), .ZN(n7800)
         );
  OAI22_X1 U2146 ( .A1(n6065), .A2(n5935), .B1(n6349), .B2(n6067), .ZN(n7799)
         );
  OAI22_X1 U2147 ( .A1(n6064), .A2(n5934), .B1(n6350), .B2(n6067), .ZN(n7798)
         );
  OAI22_X1 U2148 ( .A1(n6065), .A2(n5933), .B1(n6351), .B2(n6067), .ZN(n7797)
         );
  OAI22_X1 U2149 ( .A1(n6065), .A2(n5932), .B1(n6352), .B2(n6067), .ZN(n7796)
         );
  OAI22_X1 U2150 ( .A1(n6065), .A2(n5931), .B1(n6353), .B2(n6067), .ZN(n7795)
         );
  OAI22_X1 U2151 ( .A1(n6065), .A2(n5930), .B1(n6354), .B2(n6068), .ZN(n7794)
         );
  OAI22_X1 U2152 ( .A1(n6065), .A2(n5929), .B1(n6355), .B2(n6068), .ZN(n7793)
         );
  OAI22_X1 U2153 ( .A1(n6065), .A2(n5928), .B1(n6356), .B2(n6068), .ZN(n7792)
         );
  OAI22_X1 U2154 ( .A1(n6065), .A2(n5927), .B1(n6357), .B2(n6068), .ZN(n7791)
         );
  OAI22_X1 U2155 ( .A1(n6065), .A2(n5926), .B1(n6358), .B2(n6068), .ZN(n7790)
         );
  OAI22_X1 U2156 ( .A1(n6065), .A2(n5925), .B1(n6359), .B2(n6068), .ZN(n7789)
         );
  OAI22_X1 U2157 ( .A1(n6065), .A2(n5924), .B1(n6360), .B2(n6068), .ZN(n7788)
         );
  OAI22_X1 U2158 ( .A1(n6065), .A2(n5923), .B1(n6361), .B2(n6069), .ZN(n7787)
         );
  OAI22_X1 U2159 ( .A1(n6065), .A2(n5922), .B1(n6362), .B2(n6069), .ZN(n7786)
         );
  OAI22_X1 U2160 ( .A1(n6064), .A2(n5921), .B1(n6363), .B2(n6069), .ZN(n7785)
         );
  OAI22_X1 U2161 ( .A1(n6064), .A2(n5920), .B1(n6364), .B2(n6069), .ZN(n7784)
         );
  OAI22_X1 U2162 ( .A1(n6064), .A2(n5919), .B1(n6365), .B2(n6069), .ZN(n7783)
         );
  OAI22_X1 U2163 ( .A1(n6064), .A2(n5918), .B1(n6366), .B2(n6069), .ZN(n7782)
         );
  OAI22_X1 U2164 ( .A1(n6064), .A2(n5917), .B1(n6367), .B2(n6069), .ZN(n7781)
         );
  OAI22_X1 U2165 ( .A1(n6064), .A2(n5916), .B1(n6368), .B2(n6070), .ZN(n7780)
         );
  OAI22_X1 U2166 ( .A1(n6064), .A2(n5915), .B1(n6369), .B2(n6070), .ZN(n7779)
         );
  OAI22_X1 U2167 ( .A1(n6064), .A2(n5914), .B1(n6370), .B2(n6070), .ZN(n7778)
         );
  OAI22_X1 U2168 ( .A1(n6064), .A2(n5913), .B1(n6371), .B2(n6070), .ZN(n7777)
         );
  OAI22_X1 U2169 ( .A1(n6064), .A2(n5912), .B1(n6372), .B2(n6070), .ZN(n7776)
         );
  OAI22_X1 U2170 ( .A1(n6064), .A2(n5911), .B1(n6373), .B2(n6070), .ZN(n7775)
         );
  OAI22_X1 U2171 ( .A1(n6064), .A2(n5909), .B1(n6374), .B2(n6070), .ZN(n7774)
         );
  NAND2_X1 U2172 ( .A1(n6489), .A2(n4614), .ZN(n6488) );
  OAI22_X1 U2173 ( .A1(n6074), .A2(n6936), .B1(n6340), .B2(n6075), .ZN(n7773)
         );
  OAI22_X1 U2174 ( .A1(n6073), .A2(n6955), .B1(n6342), .B2(n6075), .ZN(n7772)
         );
  OAI22_X1 U2175 ( .A1(n6074), .A2(n6973), .B1(n6344), .B2(n6075), .ZN(n7771)
         );
  OAI22_X1 U2176 ( .A1(n6073), .A2(n6991), .B1(n6346), .B2(n6075), .ZN(n7770)
         );
  OAI22_X1 U2177 ( .A1(n6074), .A2(n7010), .B1(n6347), .B2(n6076), .ZN(n7769)
         );
  OAI22_X1 U2178 ( .A1(n6073), .A2(n7029), .B1(n6348), .B2(n6076), .ZN(n7768)
         );
  OAI22_X1 U2179 ( .A1(n6074), .A2(n7048), .B1(n6349), .B2(n6076), .ZN(n7767)
         );
  OAI22_X1 U2180 ( .A1(n6073), .A2(n7067), .B1(n6350), .B2(n6076), .ZN(n7766)
         );
  OAI22_X1 U2181 ( .A1(n6074), .A2(n7086), .B1(n6351), .B2(n6076), .ZN(n7765)
         );
  OAI22_X1 U2182 ( .A1(n6074), .A2(n7105), .B1(n6352), .B2(n6076), .ZN(n7764)
         );
  OAI22_X1 U2183 ( .A1(n6074), .A2(n7124), .B1(n6353), .B2(n6076), .ZN(n7763)
         );
  OAI22_X1 U2184 ( .A1(n6074), .A2(n7143), .B1(n6354), .B2(n6077), .ZN(n7762)
         );
  OAI22_X1 U2185 ( .A1(n6074), .A2(n7162), .B1(n6355), .B2(n6077), .ZN(n7761)
         );
  OAI22_X1 U2186 ( .A1(n6074), .A2(n7181), .B1(n6356), .B2(n6077), .ZN(n7760)
         );
  OAI22_X1 U2187 ( .A1(n6074), .A2(n7200), .B1(n6357), .B2(n6077), .ZN(n7759)
         );
  OAI22_X1 U2188 ( .A1(n6074), .A2(n7219), .B1(n6358), .B2(n6077), .ZN(n7758)
         );
  OAI22_X1 U2189 ( .A1(n6074), .A2(n7238), .B1(n6359), .B2(n6077), .ZN(n7757)
         );
  OAI22_X1 U2190 ( .A1(n6074), .A2(n7257), .B1(n6360), .B2(n6077), .ZN(n7756)
         );
  OAI22_X1 U2191 ( .A1(n6074), .A2(n7276), .B1(n6361), .B2(n6078), .ZN(n7755)
         );
  OAI22_X1 U2192 ( .A1(n6074), .A2(n7295), .B1(n6362), .B2(n6078), .ZN(n7754)
         );
  OAI22_X1 U2193 ( .A1(n6073), .A2(n7314), .B1(n6363), .B2(n6078), .ZN(n7753)
         );
  OAI22_X1 U2194 ( .A1(n6073), .A2(n7333), .B1(n6364), .B2(n6078), .ZN(n7752)
         );
  OAI22_X1 U2195 ( .A1(n6073), .A2(n7352), .B1(n6365), .B2(n6078), .ZN(n7751)
         );
  OAI22_X1 U2196 ( .A1(n6073), .A2(n7371), .B1(n6366), .B2(n6078), .ZN(n7750)
         );
  OAI22_X1 U2197 ( .A1(n6073), .A2(n7390), .B1(n6367), .B2(n6078), .ZN(n7749)
         );
  OAI22_X1 U2198 ( .A1(n6073), .A2(n7409), .B1(n6368), .B2(n6079), .ZN(n7748)
         );
  OAI22_X1 U2199 ( .A1(n6073), .A2(n7428), .B1(n6369), .B2(n6079), .ZN(n7747)
         );
  OAI22_X1 U2200 ( .A1(n6073), .A2(n7447), .B1(n6370), .B2(n6079), .ZN(n7746)
         );
  OAI22_X1 U2201 ( .A1(n6073), .A2(n7466), .B1(n6371), .B2(n6079), .ZN(n7745)
         );
  OAI22_X1 U2202 ( .A1(n6073), .A2(n7485), .B1(n6372), .B2(n6079), .ZN(n7744)
         );
  OAI22_X1 U2203 ( .A1(n6073), .A2(n7504), .B1(n6373), .B2(n6079), .ZN(n7743)
         );
  OAI22_X1 U2204 ( .A1(n6073), .A2(n7534), .B1(n6374), .B2(n6079), .ZN(n7742)
         );
  NAND2_X1 U2205 ( .A1(n6489), .A2(n4611), .ZN(n6490) );
  OAI22_X1 U2206 ( .A1(n6083), .A2(n6937), .B1(n6339), .B2(n6084), .ZN(n7741)
         );
  OAI22_X1 U2207 ( .A1(n6083), .A2(n6956), .B1(n6341), .B2(n6084), .ZN(n7740)
         );
  OAI22_X1 U2208 ( .A1(n6083), .A2(n6974), .B1(n6343), .B2(n6084), .ZN(n7739)
         );
  OAI22_X1 U2209 ( .A1(n6083), .A2(n6992), .B1(n6345), .B2(n6084), .ZN(n7738)
         );
  OAI22_X1 U2210 ( .A1(n6083), .A2(n7011), .B1(n6347), .B2(n6085), .ZN(n7737)
         );
  OAI22_X1 U2211 ( .A1(n6083), .A2(n7030), .B1(n6348), .B2(n6085), .ZN(n7736)
         );
  OAI22_X1 U2212 ( .A1(n6083), .A2(n7049), .B1(n6349), .B2(n6085), .ZN(n7735)
         );
  OAI22_X1 U2213 ( .A1(n6083), .A2(n7068), .B1(n6350), .B2(n6085), .ZN(n7734)
         );
  OAI22_X1 U2214 ( .A1(n6082), .A2(n7087), .B1(n6351), .B2(n6085), .ZN(n7733)
         );
  OAI22_X1 U2215 ( .A1(n6082), .A2(n7106), .B1(n6352), .B2(n6085), .ZN(n7732)
         );
  OAI22_X1 U2216 ( .A1(n6082), .A2(n7125), .B1(n6353), .B2(n6085), .ZN(n7731)
         );
  OAI22_X1 U2217 ( .A1(n6082), .A2(n7144), .B1(n6354), .B2(n6086), .ZN(n7730)
         );
  OAI22_X1 U2218 ( .A1(n6082), .A2(n7163), .B1(n6355), .B2(n6086), .ZN(n7729)
         );
  OAI22_X1 U2219 ( .A1(n6082), .A2(n7182), .B1(n6356), .B2(n6086), .ZN(n7728)
         );
  OAI22_X1 U2220 ( .A1(n6082), .A2(n7201), .B1(n6357), .B2(n6086), .ZN(n7727)
         );
  OAI22_X1 U2221 ( .A1(n6082), .A2(n7220), .B1(n6358), .B2(n6086), .ZN(n7726)
         );
  OAI22_X1 U2222 ( .A1(n6082), .A2(n7239), .B1(n6359), .B2(n6086), .ZN(n7725)
         );
  OAI22_X1 U2223 ( .A1(n6082), .A2(n7258), .B1(n6360), .B2(n6086), .ZN(n7724)
         );
  OAI22_X1 U2224 ( .A1(n6082), .A2(n7277), .B1(n6361), .B2(n6087), .ZN(n7723)
         );
  OAI22_X1 U2225 ( .A1(n6082), .A2(n7296), .B1(n6362), .B2(n6087), .ZN(n7722)
         );
  OAI22_X1 U2226 ( .A1(n6083), .A2(n7315), .B1(n6363), .B2(n6087), .ZN(n7721)
         );
  OAI22_X1 U2227 ( .A1(n6083), .A2(n7334), .B1(n6364), .B2(n6087), .ZN(n7720)
         );
  OAI22_X1 U2228 ( .A1(n6083), .A2(n7353), .B1(n6365), .B2(n6087), .ZN(n7719)
         );
  OAI22_X1 U2229 ( .A1(n6083), .A2(n7372), .B1(n6366), .B2(n6087), .ZN(n7718)
         );
  OAI22_X1 U2230 ( .A1(n6082), .A2(n7391), .B1(n6367), .B2(n6087), .ZN(n7717)
         );
  OAI22_X1 U2231 ( .A1(n6083), .A2(n7410), .B1(n6368), .B2(n6088), .ZN(n7716)
         );
  OAI22_X1 U2232 ( .A1(n6082), .A2(n7429), .B1(n6369), .B2(n6088), .ZN(n7715)
         );
  OAI22_X1 U2233 ( .A1(n6083), .A2(n7448), .B1(n6370), .B2(n6088), .ZN(n7714)
         );
  OAI22_X1 U2234 ( .A1(n6082), .A2(n7467), .B1(n6371), .B2(n6088), .ZN(n7713)
         );
  OAI22_X1 U2235 ( .A1(n6083), .A2(n7486), .B1(n6372), .B2(n6088), .ZN(n7712)
         );
  OAI22_X1 U2236 ( .A1(n6082), .A2(n7505), .B1(n6373), .B2(n6088), .ZN(n7711)
         );
  OAI22_X1 U2237 ( .A1(n6083), .A2(n7535), .B1(n6374), .B2(n6088), .ZN(n7710)
         );
  NAND2_X1 U2238 ( .A1(n4607), .A2(n4614), .ZN(n6491) );
  OAI22_X1 U2239 ( .A1(n6092), .A2(n5972), .B1(n6340), .B2(n6093), .ZN(n3207)
         );
  OAI22_X1 U2240 ( .A1(n6092), .A2(n5971), .B1(n6342), .B2(n6093), .ZN(n3208)
         );
  OAI22_X1 U2241 ( .A1(n6092), .A2(n5970), .B1(n6344), .B2(n6093), .ZN(n3209)
         );
  OAI22_X1 U2242 ( .A1(n6092), .A2(n5969), .B1(n6346), .B2(n6093), .ZN(n3210)
         );
  OAI22_X1 U2243 ( .A1(n6092), .A2(n5968), .B1(n6347), .B2(n6094), .ZN(n3211)
         );
  OAI22_X1 U2244 ( .A1(n6092), .A2(n5967), .B1(n6348), .B2(n6094), .ZN(n3212)
         );
  OAI22_X1 U2245 ( .A1(n6092), .A2(n5966), .B1(n6349), .B2(n6094), .ZN(n3213)
         );
  OAI22_X1 U2246 ( .A1(n6092), .A2(n5965), .B1(n6350), .B2(n6094), .ZN(n3214)
         );
  OAI22_X1 U2247 ( .A1(n6091), .A2(n5964), .B1(n6351), .B2(n6094), .ZN(n3215)
         );
  OAI22_X1 U2248 ( .A1(n6091), .A2(n5963), .B1(n6352), .B2(n6094), .ZN(n3216)
         );
  OAI22_X1 U2249 ( .A1(n6091), .A2(n5962), .B1(n6353), .B2(n6094), .ZN(n3217)
         );
  OAI22_X1 U2250 ( .A1(n6091), .A2(n5961), .B1(n6354), .B2(n6095), .ZN(n3218)
         );
  OAI22_X1 U2251 ( .A1(n6091), .A2(n5960), .B1(n6355), .B2(n6095), .ZN(n3219)
         );
  OAI22_X1 U2252 ( .A1(n6091), .A2(n5959), .B1(n6356), .B2(n6095), .ZN(n3220)
         );
  OAI22_X1 U2253 ( .A1(n6091), .A2(n5958), .B1(n6357), .B2(n6095), .ZN(n3221)
         );
  OAI22_X1 U2254 ( .A1(n6091), .A2(n5957), .B1(n6358), .B2(n6095), .ZN(n3222)
         );
  OAI22_X1 U2255 ( .A1(n6091), .A2(n5956), .B1(n6359), .B2(n6095), .ZN(n3223)
         );
  OAI22_X1 U2256 ( .A1(n6091), .A2(n5955), .B1(n6360), .B2(n6095), .ZN(n3224)
         );
  OAI22_X1 U2257 ( .A1(n6091), .A2(n5954), .B1(n6361), .B2(n6096), .ZN(n3225)
         );
  OAI22_X1 U2258 ( .A1(n6091), .A2(n5953), .B1(n6362), .B2(n6096), .ZN(n3226)
         );
  OAI22_X1 U2259 ( .A1(n6092), .A2(n5952), .B1(n6363), .B2(n6096), .ZN(n3227)
         );
  OAI22_X1 U2260 ( .A1(n6092), .A2(n5951), .B1(n6364), .B2(n6096), .ZN(n3228)
         );
  OAI22_X1 U2261 ( .A1(n6092), .A2(n5950), .B1(n6365), .B2(n6096), .ZN(n3229)
         );
  OAI22_X1 U2262 ( .A1(n6092), .A2(n5949), .B1(n6366), .B2(n6096), .ZN(n3230)
         );
  OAI22_X1 U2263 ( .A1(n6091), .A2(n5948), .B1(n6367), .B2(n6096), .ZN(n3231)
         );
  OAI22_X1 U2264 ( .A1(n6092), .A2(n5947), .B1(n6368), .B2(n6097), .ZN(n3232)
         );
  OAI22_X1 U2265 ( .A1(n6091), .A2(n5946), .B1(n6369), .B2(n6097), .ZN(n3233)
         );
  OAI22_X1 U2266 ( .A1(n6092), .A2(n5945), .B1(n6370), .B2(n6097), .ZN(n3234)
         );
  OAI22_X1 U2267 ( .A1(n6091), .A2(n5944), .B1(n6371), .B2(n6097), .ZN(n3235)
         );
  OAI22_X1 U2268 ( .A1(n6092), .A2(n5943), .B1(n6372), .B2(n6097), .ZN(n3236)
         );
  OAI22_X1 U2269 ( .A1(n6091), .A2(n5942), .B1(n6373), .B2(n6097), .ZN(n3237)
         );
  OAI22_X1 U2270 ( .A1(n6092), .A2(n5941), .B1(n6374), .B2(n6097), .ZN(n3238)
         );
  NAND2_X1 U2271 ( .A1(n4607), .A2(n4611), .ZN(n6492) );
  MUX2_X1 U2272 ( .A(n5647), .B(DATAIN[0]), .S(n6100), .Z(n3175) );
  MUX2_X1 U2273 ( .A(n5582), .B(DATAIN[1]), .S(n6100), .Z(n3176) );
  MUX2_X1 U2274 ( .A(n5581), .B(DATAIN[2]), .S(n6100), .Z(n3177) );
  MUX2_X1 U2275 ( .A(n5580), .B(DATAIN[3]), .S(n6100), .Z(n3178) );
  OAI22_X1 U2276 ( .A1(n6100), .A2(n7004), .B1(n6347), .B2(n6102), .ZN(n7709)
         );
  OAI22_X1 U2277 ( .A1(n6100), .A2(n7023), .B1(n6348), .B2(n6102), .ZN(n7708)
         );
  OAI22_X1 U2278 ( .A1(n6100), .A2(n7042), .B1(n6349), .B2(n6102), .ZN(n7707)
         );
  OAI22_X1 U2279 ( .A1(n6100), .A2(n7061), .B1(n6350), .B2(n6102), .ZN(n7706)
         );
  OAI22_X1 U2280 ( .A1(n6100), .A2(n7080), .B1(n6351), .B2(n6103), .ZN(n7705)
         );
  OAI22_X1 U2281 ( .A1(n6100), .A2(n7099), .B1(n6352), .B2(n6103), .ZN(n7704)
         );
  OAI22_X1 U2282 ( .A1(n6100), .A2(n7118), .B1(n6353), .B2(n6103), .ZN(n7703)
         );
  OAI22_X1 U2283 ( .A1(n6100), .A2(n7137), .B1(n6354), .B2(n6103), .ZN(n7702)
         );
  OAI22_X1 U2284 ( .A1(n6100), .A2(n7156), .B1(n6355), .B2(n6103), .ZN(n7701)
         );
  OAI22_X1 U2285 ( .A1(n6101), .A2(n7175), .B1(n6356), .B2(n6103), .ZN(n7700)
         );
  OAI22_X1 U2286 ( .A1(n6101), .A2(n7194), .B1(n6357), .B2(n6103), .ZN(n7699)
         );
  OAI22_X1 U2287 ( .A1(n6101), .A2(n7213), .B1(n6358), .B2(n6104), .ZN(n7698)
         );
  OAI22_X1 U2288 ( .A1(n6101), .A2(n7232), .B1(n6359), .B2(n6104), .ZN(n7697)
         );
  OAI22_X1 U2289 ( .A1(n6101), .A2(n7251), .B1(n6360), .B2(n6104), .ZN(n7696)
         );
  OAI22_X1 U2290 ( .A1(n6101), .A2(n7270), .B1(n6361), .B2(n6104), .ZN(n7695)
         );
  OAI22_X1 U2291 ( .A1(n6101), .A2(n7289), .B1(n6362), .B2(n6104), .ZN(n7694)
         );
  OAI22_X1 U2292 ( .A1(n6101), .A2(n7308), .B1(n6363), .B2(n6104), .ZN(n7693)
         );
  OAI22_X1 U2293 ( .A1(n6101), .A2(n7327), .B1(n6364), .B2(n6104), .ZN(n7692)
         );
  OAI22_X1 U2294 ( .A1(n6101), .A2(n7346), .B1(n6365), .B2(n6105), .ZN(n7691)
         );
  OAI22_X1 U2295 ( .A1(n6101), .A2(n7365), .B1(n6366), .B2(n6105), .ZN(n7690)
         );
  OAI22_X1 U2296 ( .A1(n6101), .A2(n7384), .B1(n6367), .B2(n6105), .ZN(n7689)
         );
  OAI22_X1 U2297 ( .A1(n6101), .A2(n7403), .B1(n6368), .B2(n6105), .ZN(n7688)
         );
  OAI22_X1 U2298 ( .A1(n6100), .A2(n7422), .B1(n6369), .B2(n6105), .ZN(n7687)
         );
  OAI22_X1 U2299 ( .A1(n6101), .A2(n7441), .B1(n6370), .B2(n6105), .ZN(n7686)
         );
  OAI22_X1 U2300 ( .A1(n6100), .A2(n7460), .B1(n6371), .B2(n6105), .ZN(n7685)
         );
  OAI22_X1 U2301 ( .A1(n6101), .A2(n7479), .B1(n6372), .B2(n6106), .ZN(n7684)
         );
  OAI22_X1 U2302 ( .A1(n6100), .A2(n7498), .B1(n6373), .B2(n6106), .ZN(n7683)
         );
  OAI22_X1 U2303 ( .A1(n6101), .A2(n7521), .B1(n6374), .B2(n6106), .ZN(n3206)
         );
  NAND2_X1 U2304 ( .A1(n4625), .A2(n4606), .ZN(n6493) );
  MUX2_X1 U2305 ( .A(n5583), .B(DATAIN[0]), .S(n6109), .Z(n3143) );
  MUX2_X1 U2306 ( .A(n5485), .B(DATAIN[1]), .S(n6109), .Z(n3144) );
  MUX2_X1 U2307 ( .A(n5484), .B(DATAIN[2]), .S(n6109), .Z(n3145) );
  MUX2_X1 U2308 ( .A(n5483), .B(DATAIN[3]), .S(n6109), .Z(n3146) );
  OAI22_X1 U2309 ( .A1(n6109), .A2(n5907), .B1(n6347), .B2(n6111), .ZN(n7682)
         );
  OAI22_X1 U2310 ( .A1(n6109), .A2(n5906), .B1(n6348), .B2(n6111), .ZN(n7681)
         );
  OAI22_X1 U2311 ( .A1(n6109), .A2(n5905), .B1(n6349), .B2(n6111), .ZN(n7680)
         );
  OAI22_X1 U2312 ( .A1(n6109), .A2(n5904), .B1(n6350), .B2(n6111), .ZN(n7679)
         );
  OAI22_X1 U2313 ( .A1(n6109), .A2(n5903), .B1(n6351), .B2(n6112), .ZN(n7678)
         );
  OAI22_X1 U2314 ( .A1(n6109), .A2(n5902), .B1(n6352), .B2(n6112), .ZN(n7677)
         );
  OAI22_X1 U2315 ( .A1(n6109), .A2(n5901), .B1(n6353), .B2(n6112), .ZN(n7676)
         );
  OAI22_X1 U2316 ( .A1(n6109), .A2(n5900), .B1(n6354), .B2(n6112), .ZN(n7675)
         );
  OAI22_X1 U2317 ( .A1(n6109), .A2(n5899), .B1(n6355), .B2(n6112), .ZN(n7674)
         );
  OAI22_X1 U2318 ( .A1(n6110), .A2(n5898), .B1(n6356), .B2(n6112), .ZN(n7673)
         );
  OAI22_X1 U2319 ( .A1(n6110), .A2(n5897), .B1(n6357), .B2(n6112), .ZN(n7672)
         );
  OAI22_X1 U2320 ( .A1(n6110), .A2(n5896), .B1(n6358), .B2(n6113), .ZN(n7671)
         );
  OAI22_X1 U2321 ( .A1(n6110), .A2(n5895), .B1(n6359), .B2(n6113), .ZN(n7670)
         );
  OAI22_X1 U2322 ( .A1(n6110), .A2(n5894), .B1(n6360), .B2(n6113), .ZN(n7669)
         );
  OAI22_X1 U2323 ( .A1(n6110), .A2(n5893), .B1(n6361), .B2(n6113), .ZN(n7668)
         );
  OAI22_X1 U2324 ( .A1(n6110), .A2(n5892), .B1(n6362), .B2(n6113), .ZN(n7667)
         );
  OAI22_X1 U2325 ( .A1(n6110), .A2(n5891), .B1(n6363), .B2(n6113), .ZN(n7666)
         );
  OAI22_X1 U2326 ( .A1(n6110), .A2(n5890), .B1(n6364), .B2(n6113), .ZN(n7665)
         );
  OAI22_X1 U2327 ( .A1(n6110), .A2(n5889), .B1(n6365), .B2(n6114), .ZN(n7664)
         );
  OAI22_X1 U2328 ( .A1(n6110), .A2(n5888), .B1(n6366), .B2(n6114), .ZN(n7663)
         );
  OAI22_X1 U2329 ( .A1(n6110), .A2(n5887), .B1(n6367), .B2(n6114), .ZN(n7662)
         );
  OAI22_X1 U2330 ( .A1(n6110), .A2(n5886), .B1(n6368), .B2(n6114), .ZN(n7661)
         );
  OAI22_X1 U2331 ( .A1(n6109), .A2(n5885), .B1(n6369), .B2(n6114), .ZN(n7660)
         );
  OAI22_X1 U2332 ( .A1(n6110), .A2(n5884), .B1(n6370), .B2(n6114), .ZN(n7659)
         );
  OAI22_X1 U2333 ( .A1(n6109), .A2(n5883), .B1(n6371), .B2(n6114), .ZN(n7658)
         );
  OAI22_X1 U2334 ( .A1(n6110), .A2(n5882), .B1(n6372), .B2(n6115), .ZN(n7657)
         );
  OAI22_X1 U2335 ( .A1(n6109), .A2(n5881), .B1(n6373), .B2(n6115), .ZN(n7656)
         );
  OAI22_X1 U2336 ( .A1(n6110), .A2(n5880), .B1(n6374), .B2(n6115), .ZN(n3174)
         );
  INV_X1 U2337 ( .A(n2002), .ZN(n6494) );
  NAND4_X1 U2338 ( .A1(n1997), .A2(n2027), .A3(n1998), .A4(n6494), .ZN(n6495)
         );
  NAND2_X1 U2339 ( .A1(n6173), .A2(n6495), .ZN(n6502) );
  INV_X1 U2340 ( .A(n6502), .ZN(n6916) );
  NAND2_X1 U2341 ( .A1(n4612), .A2(n4618), .ZN(n6906) );
  NAND2_X1 U2342 ( .A1(n4626), .A2(n4610), .ZN(n6907) );
  OAI22_X1 U2343 ( .A1(n3742), .A2(n4902), .B1(n2284), .B2(n4900), .ZN(n6496)
         );
  AOI221_X1 U2344 ( .B1(n6160), .B2(n6938), .C1(n6275), .C2(n7588), .A(n6496), 
        .ZN(n6501) );
  AOI222_X1 U2345 ( .A1(n6298), .A2(n4062), .B1(n6287), .B2(n7586), .C1(n6301), 
        .C2(n4030), .ZN(n6500) );
  AOI22_X1 U2346 ( .A1(n2910), .A2(n6149), .B1(n6934), .B2(n6146), .ZN(n6497)
         );
  OAI221_X1 U2347 ( .B1(n4813), .B2(n6155), .C1(n6936), .C2(n6152), .A(n6497), 
        .ZN(n6498) );
  NOR4_X1 U2348 ( .A1(n6498), .A2(n2025), .A3(n2024), .A4(n2021), .ZN(n6499)
         );
  AND3_X1 U2349 ( .A1(n6501), .A2(n6500), .A3(n6499), .ZN(n6503) );
  OAI222_X1 U2350 ( .A1(n2124), .A2(n6116), .B1(n939), .B2(n6121), .C1(n6503), 
        .C2(n6502), .ZN(n6510) );
  NAND2_X1 U2351 ( .A1(n2006), .A2(n4618), .ZN(n6910) );
  NAND2_X1 U2352 ( .A1(n4612), .A2(n4621), .ZN(n6513) );
  INV_X1 U2353 ( .A(n2156), .ZN(n7553) );
  AOI22_X1 U2354 ( .A1(n6124), .A2(n7553), .B1(n4897), .B2(n4972), .ZN(n6504)
         );
  OAI221_X1 U2355 ( .B1(n2092), .B2(n6130), .C1(n938), .C2(n6513), .A(n6504), 
        .ZN(n6509) );
  NAND2_X1 U2356 ( .A1(n4621), .A2(n1993), .ZN(n6913) );
  NAND2_X1 U2357 ( .A1(n4610), .A2(n4618), .ZN(n6515) );
  AOI22_X1 U2358 ( .A1(n6135), .A2(n950), .B1(n4898), .B2(n4912), .ZN(n6505)
         );
  OAI221_X1 U2359 ( .B1(n3646), .B2(n6141), .C1(n2188), .C2(n6515), .A(n6505), 
        .ZN(n6508) );
  NAND2_X1 U2360 ( .A1(n1993), .A2(n4618), .ZN(n6922) );
  NAND2_X1 U2361 ( .A1(n4661), .A2(n4610), .ZN(n6521) );
  AOI22_X1 U2362 ( .A1(n6164), .A2(n6942), .B1(n4616), .B2(DATAIN[0]), .ZN(
        n6506) );
  OAI221_X1 U2363 ( .B1(n2220), .B2(n6170), .C1(n2942), .C2(n6521), .A(n6506), 
        .ZN(n6507) );
  NOR4_X1 U2364 ( .A1(n6510), .A2(n6509), .A3(n6508), .A4(n6507), .ZN(n6511)
         );
  OAI21_X1 U2365 ( .B1(n6173), .B2(n6512), .A(n6511), .ZN(n2983) );
  OAI222_X1 U2366 ( .A1(n956), .A2(n6121), .B1(n2719), .B2(n6119), .C1(n2125), 
        .C2(n6116), .ZN(n6527) );
  INV_X1 U2367 ( .A(n6513), .ZN(n6908) );
  INV_X1 U2368 ( .A(n2157), .ZN(n7554) );
  AOI22_X1 U2369 ( .A1(n6127), .A2(n5036), .B1(n6124), .B2(n7554), .ZN(n6514)
         );
  OAI221_X1 U2370 ( .B1(n2061), .B2(n6133), .C1(n2093), .C2(n6130), .A(n6514), 
        .ZN(n6526) );
  INV_X1 U2371 ( .A(n6515), .ZN(n6911) );
  AOI22_X1 U2372 ( .A1(n6138), .A2(n5033), .B1(n6135), .B2(n966), .ZN(n6516)
         );
  OAI221_X1 U2373 ( .B1(n6342), .B2(n6144), .C1(n3647), .C2(n6141), .A(n6516), 
        .ZN(n6525) );
  AOI22_X1 U2374 ( .A1(n2911), .A2(n6149), .B1(n6953), .B2(n6146), .ZN(n6517)
         );
  OAI221_X1 U2375 ( .B1(n4811), .B2(n6155), .C1(n6955), .C2(n6152), .A(n6517), 
        .ZN(n6520) );
  NAND2_X1 U2376 ( .A1(n6160), .A2(n6957), .ZN(n6518) );
  NAND4_X1 U2377 ( .A1(n1975), .A2(n1976), .A3(n1974), .A4(n6518), .ZN(n6519)
         );
  OAI21_X1 U2378 ( .B1(n6520), .B2(n6519), .A(n6163), .ZN(n6523) );
  INV_X1 U2379 ( .A(n6521), .ZN(n6919) );
  AOI22_X1 U2380 ( .A1(n6167), .A2(n6951), .B1(n6164), .B2(n4942), .ZN(n6522)
         );
  OAI211_X1 U2381 ( .C1(n2221), .C2(n6170), .A(n6523), .B(n6522), .ZN(n6524)
         );
  NOR4_X1 U2382 ( .A1(n6527), .A2(n6526), .A3(n6525), .A4(n6524), .ZN(n6528)
         );
  OAI21_X1 U2383 ( .B1(n2623), .B2(n6173), .A(n6528), .ZN(n2984) );
  OAI222_X1 U2384 ( .A1(n972), .A2(n6121), .B1(n2720), .B2(n6119), .C1(n2126), 
        .C2(n6116), .ZN(n6540) );
  INV_X1 U2385 ( .A(n2158), .ZN(n7555) );
  AOI22_X1 U2386 ( .A1(n6127), .A2(n5035), .B1(n6124), .B2(n7555), .ZN(n6529)
         );
  OAI221_X1 U2387 ( .B1(n2062), .B2(n6133), .C1(n2094), .C2(n6130), .A(n6529), 
        .ZN(n6539) );
  AOI22_X1 U2388 ( .A1(n6138), .A2(n5032), .B1(n6135), .B2(n982), .ZN(n6530)
         );
  OAI221_X1 U2389 ( .B1(n6344), .B2(n6144), .C1(n3648), .C2(n6141), .A(n6530), 
        .ZN(n6538) );
  AOI22_X1 U2390 ( .A1(n2912), .A2(n6149), .B1(n6971), .B2(n6146), .ZN(n6531)
         );
  OAI221_X1 U2391 ( .B1(n4809), .B2(n6155), .C1(n6973), .C2(n6152), .A(n6531), 
        .ZN(n6534) );
  NAND2_X1 U2392 ( .A1(n6160), .A2(n6975), .ZN(n6532) );
  NAND4_X1 U2393 ( .A1(n1958), .A2(n1959), .A3(n1957), .A4(n6532), .ZN(n6533)
         );
  OAI21_X1 U2394 ( .B1(n6534), .B2(n6533), .A(n6163), .ZN(n6536) );
  AOI22_X1 U2395 ( .A1(n6167), .A2(n6969), .B1(n6164), .B2(n4941), .ZN(n6535)
         );
  OAI211_X1 U2396 ( .C1(n2222), .C2(n6170), .A(n6536), .B(n6535), .ZN(n6537)
         );
  NOR4_X1 U2397 ( .A1(n6540), .A2(n6539), .A3(n6538), .A4(n6537), .ZN(n6541)
         );
  OAI21_X1 U2398 ( .B1(n2624), .B2(n6175), .A(n6541), .ZN(n2985) );
  OAI222_X1 U2399 ( .A1(n988), .A2(n6121), .B1(n2721), .B2(n6119), .C1(n2127), 
        .C2(n6116), .ZN(n6553) );
  INV_X1 U2400 ( .A(n2159), .ZN(n7556) );
  AOI22_X1 U2401 ( .A1(n6127), .A2(n5034), .B1(n6124), .B2(n7556), .ZN(n6542)
         );
  OAI221_X1 U2402 ( .B1(n2063), .B2(n6133), .C1(n2095), .C2(n6130), .A(n6542), 
        .ZN(n6552) );
  AOI22_X1 U2403 ( .A1(n6138), .A2(n5031), .B1(n6135), .B2(n998), .ZN(n6543)
         );
  OAI221_X1 U2404 ( .B1(n6346), .B2(n6144), .C1(n3649), .C2(n6141), .A(n6543), 
        .ZN(n6551) );
  AOI22_X1 U2405 ( .A1(n2913), .A2(n6149), .B1(n6989), .B2(n6146), .ZN(n6544)
         );
  OAI221_X1 U2406 ( .B1(n4807), .B2(n6155), .C1(n6991), .C2(n6152), .A(n6544), 
        .ZN(n6547) );
  NAND2_X1 U2407 ( .A1(n6160), .A2(n6993), .ZN(n6545) );
  NAND4_X1 U2408 ( .A1(n1941), .A2(n1942), .A3(n1940), .A4(n6545), .ZN(n6546)
         );
  OAI21_X1 U2409 ( .B1(n6547), .B2(n6546), .A(n6163), .ZN(n6549) );
  AOI22_X1 U2410 ( .A1(n6167), .A2(n6987), .B1(n6164), .B2(n4940), .ZN(n6548)
         );
  OAI211_X1 U2411 ( .C1(n2223), .C2(n6170), .A(n6549), .B(n6548), .ZN(n6550)
         );
  NOR4_X1 U2412 ( .A1(n6553), .A2(n6552), .A3(n6551), .A4(n6550), .ZN(n6554)
         );
  OAI21_X1 U2413 ( .B1(n2625), .B2(n6175), .A(n6554), .ZN(n2986) );
  OAI222_X1 U2414 ( .A1(n4699), .A2(n6121), .B1(n2722), .B2(n6119), .C1(n2128), 
        .C2(n6116), .ZN(n6566) );
  INV_X1 U2415 ( .A(n2160), .ZN(n7557) );
  AOI22_X1 U2416 ( .A1(n6127), .A2(n2850), .B1(n6124), .B2(n7557), .ZN(n6555)
         );
  OAI221_X1 U2417 ( .B1(n2064), .B2(n6133), .C1(n2096), .C2(n6130), .A(n6555), 
        .ZN(n6565) );
  AOI22_X1 U2418 ( .A1(n6138), .A2(n5030), .B1(n6135), .B2(n4970), .ZN(n6556)
         );
  OAI221_X1 U2419 ( .B1(n6347), .B2(n6144), .C1(n3650), .C2(n6141), .A(n6556), 
        .ZN(n6564) );
  AOI22_X1 U2420 ( .A1(n2914), .A2(n6149), .B1(n7008), .B2(n6146), .ZN(n6557)
         );
  OAI221_X1 U2421 ( .B1(n4805), .B2(n6155), .C1(n7010), .C2(n6152), .A(n6557), 
        .ZN(n6560) );
  NAND2_X1 U2422 ( .A1(n6160), .A2(n7012), .ZN(n6558) );
  NAND4_X1 U2423 ( .A1(n1924), .A2(n1925), .A3(n1923), .A4(n6558), .ZN(n6559)
         );
  OAI21_X1 U2424 ( .B1(n6560), .B2(n6559), .A(n6163), .ZN(n6562) );
  AOI22_X1 U2425 ( .A1(n6167), .A2(n7006), .B1(n6164), .B2(n4939), .ZN(n6561)
         );
  OAI211_X1 U2426 ( .C1(n2224), .C2(n6170), .A(n6562), .B(n6561), .ZN(n6563)
         );
  NOR4_X1 U2427 ( .A1(n6566), .A2(n6565), .A3(n6564), .A4(n6563), .ZN(n6567)
         );
  OAI21_X1 U2428 ( .B1(n2626), .B2(n6175), .A(n6567), .ZN(n2987) );
  OAI222_X1 U2429 ( .A1(n4697), .A2(n6121), .B1(n2723), .B2(n6119), .C1(n2129), 
        .C2(n6116), .ZN(n6579) );
  INV_X1 U2430 ( .A(n2161), .ZN(n7558) );
  AOI22_X1 U2431 ( .A1(n6127), .A2(n2851), .B1(n6124), .B2(n7558), .ZN(n6568)
         );
  OAI221_X1 U2432 ( .B1(n2065), .B2(n6133), .C1(n2097), .C2(n6130), .A(n6568), 
        .ZN(n6578) );
  AOI22_X1 U2433 ( .A1(n6138), .A2(n5029), .B1(n6135), .B2(n4969), .ZN(n6569)
         );
  OAI221_X1 U2434 ( .B1(n6348), .B2(n6144), .C1(n3651), .C2(n6141), .A(n6569), 
        .ZN(n6577) );
  AOI22_X1 U2435 ( .A1(n2915), .A2(n6149), .B1(n7027), .B2(n6146), .ZN(n6570)
         );
  OAI221_X1 U2436 ( .B1(n4803), .B2(n6155), .C1(n7029), .C2(n6152), .A(n6570), 
        .ZN(n6573) );
  NAND2_X1 U2437 ( .A1(n6160), .A2(n7031), .ZN(n6571) );
  NAND4_X1 U2438 ( .A1(n1907), .A2(n1908), .A3(n1906), .A4(n6571), .ZN(n6572)
         );
  OAI21_X1 U2439 ( .B1(n6573), .B2(n6572), .A(n6163), .ZN(n6575) );
  AOI22_X1 U2440 ( .A1(n6167), .A2(n7025), .B1(n6164), .B2(n4938), .ZN(n6574)
         );
  OAI211_X1 U2441 ( .C1(n2225), .C2(n6170), .A(n6575), .B(n6574), .ZN(n6576)
         );
  NOR4_X1 U2442 ( .A1(n6579), .A2(n6578), .A3(n6577), .A4(n6576), .ZN(n6580)
         );
  OAI21_X1 U2443 ( .B1(n2627), .B2(n6175), .A(n6580), .ZN(n2988) );
  OAI222_X1 U2444 ( .A1(n4705), .A2(n6121), .B1(n2724), .B2(n6119), .C1(n2130), 
        .C2(n6116), .ZN(n6592) );
  INV_X1 U2445 ( .A(n2162), .ZN(n7559) );
  AOI22_X1 U2446 ( .A1(n6127), .A2(n2852), .B1(n6124), .B2(n7559), .ZN(n6581)
         );
  OAI221_X1 U2447 ( .B1(n2066), .B2(n6133), .C1(n2098), .C2(n6130), .A(n6581), 
        .ZN(n6591) );
  AOI22_X1 U2448 ( .A1(n6138), .A2(n5028), .B1(n6135), .B2(n4968), .ZN(n6582)
         );
  OAI221_X1 U2449 ( .B1(n6349), .B2(n6144), .C1(n3652), .C2(n6141), .A(n6582), 
        .ZN(n6590) );
  AOI22_X1 U2450 ( .A1(n2916), .A2(n6149), .B1(n7046), .B2(n6146), .ZN(n6583)
         );
  OAI221_X1 U2451 ( .B1(n4801), .B2(n6155), .C1(n7048), .C2(n6152), .A(n6583), 
        .ZN(n6586) );
  NAND2_X1 U2452 ( .A1(n6160), .A2(n7050), .ZN(n6584) );
  NAND4_X1 U2453 ( .A1(n1890), .A2(n1891), .A3(n1889), .A4(n6584), .ZN(n6585)
         );
  OAI21_X1 U2454 ( .B1(n6586), .B2(n6585), .A(n6163), .ZN(n6588) );
  AOI22_X1 U2455 ( .A1(n6167), .A2(n7044), .B1(n6164), .B2(n4937), .ZN(n6587)
         );
  OAI211_X1 U2456 ( .C1(n2226), .C2(n6170), .A(n6588), .B(n6587), .ZN(n6589)
         );
  NOR4_X1 U2457 ( .A1(n6592), .A2(n6591), .A3(n6590), .A4(n6589), .ZN(n6593)
         );
  OAI21_X1 U2458 ( .B1(n2628), .B2(n6175), .A(n6593), .ZN(n2989) );
  OAI222_X1 U2459 ( .A1(n4703), .A2(n6121), .B1(n2725), .B2(n6119), .C1(n2131), 
        .C2(n6116), .ZN(n6605) );
  INV_X1 U2460 ( .A(n2163), .ZN(n7560) );
  AOI22_X1 U2461 ( .A1(n6127), .A2(n2853), .B1(n6124), .B2(n7560), .ZN(n6594)
         );
  OAI221_X1 U2462 ( .B1(n2067), .B2(n6133), .C1(n2099), .C2(n6130), .A(n6594), 
        .ZN(n6604) );
  AOI22_X1 U2463 ( .A1(n6138), .A2(n5027), .B1(n6135), .B2(n4967), .ZN(n6595)
         );
  OAI221_X1 U2464 ( .B1(n6350), .B2(n6144), .C1(n3653), .C2(n6141), .A(n6595), 
        .ZN(n6603) );
  AOI22_X1 U2465 ( .A1(n2917), .A2(n6149), .B1(n7065), .B2(n6146), .ZN(n6596)
         );
  OAI221_X1 U2466 ( .B1(n4799), .B2(n6155), .C1(n7067), .C2(n6152), .A(n6596), 
        .ZN(n6599) );
  NAND2_X1 U2467 ( .A1(n6160), .A2(n7069), .ZN(n6597) );
  NAND4_X1 U2468 ( .A1(n1873), .A2(n1874), .A3(n1872), .A4(n6597), .ZN(n6598)
         );
  OAI21_X1 U2469 ( .B1(n6599), .B2(n6598), .A(n6163), .ZN(n6601) );
  AOI22_X1 U2470 ( .A1(n6167), .A2(n7063), .B1(n6164), .B2(n4936), .ZN(n6600)
         );
  OAI211_X1 U2471 ( .C1(n2227), .C2(n6170), .A(n6601), .B(n6600), .ZN(n6602)
         );
  NOR4_X1 U2472 ( .A1(n6605), .A2(n6604), .A3(n6603), .A4(n6602), .ZN(n6606)
         );
  OAI21_X1 U2473 ( .B1(n2629), .B2(n6175), .A(n6606), .ZN(n2990) );
  OAI222_X1 U2474 ( .A1(n4701), .A2(n6121), .B1(n2726), .B2(n6119), .C1(n2132), 
        .C2(n6116), .ZN(n6618) );
  INV_X1 U2475 ( .A(n2164), .ZN(n7561) );
  AOI22_X1 U2476 ( .A1(n6127), .A2(n2854), .B1(n6124), .B2(n7561), .ZN(n6607)
         );
  OAI221_X1 U2477 ( .B1(n2068), .B2(n6133), .C1(n2100), .C2(n6130), .A(n6607), 
        .ZN(n6617) );
  AOI22_X1 U2478 ( .A1(n6138), .A2(n5026), .B1(n6135), .B2(n4966), .ZN(n6608)
         );
  OAI221_X1 U2479 ( .B1(n6351), .B2(n6144), .C1(n3654), .C2(n6141), .A(n6608), 
        .ZN(n6616) );
  AOI22_X1 U2480 ( .A1(n2918), .A2(n6149), .B1(n7084), .B2(n6146), .ZN(n6609)
         );
  OAI221_X1 U2481 ( .B1(n4797), .B2(n6155), .C1(n7086), .C2(n6152), .A(n6609), 
        .ZN(n6612) );
  NAND2_X1 U2482 ( .A1(n6159), .A2(n7088), .ZN(n6610) );
  NAND4_X1 U2483 ( .A1(n1856), .A2(n1857), .A3(n1855), .A4(n6610), .ZN(n6611)
         );
  OAI21_X1 U2484 ( .B1(n6612), .B2(n6611), .A(n6162), .ZN(n6614) );
  AOI22_X1 U2485 ( .A1(n6167), .A2(n7082), .B1(n6164), .B2(n4935), .ZN(n6613)
         );
  OAI211_X1 U2486 ( .C1(n2228), .C2(n6170), .A(n6614), .B(n6613), .ZN(n6615)
         );
  NOR4_X1 U2487 ( .A1(n6618), .A2(n6617), .A3(n6616), .A4(n6615), .ZN(n6619)
         );
  OAI21_X1 U2488 ( .B1(n2630), .B2(n6175), .A(n6619), .ZN(n2991) );
  OAI222_X1 U2489 ( .A1(n4711), .A2(n6121), .B1(n2727), .B2(n6119), .C1(n2133), 
        .C2(n6116), .ZN(n6631) );
  INV_X1 U2490 ( .A(n2165), .ZN(n7562) );
  AOI22_X1 U2491 ( .A1(n6127), .A2(n2855), .B1(n6124), .B2(n7562), .ZN(n6620)
         );
  OAI221_X1 U2492 ( .B1(n2069), .B2(n6133), .C1(n2101), .C2(n6130), .A(n6620), 
        .ZN(n6630) );
  AOI22_X1 U2493 ( .A1(n6138), .A2(n5025), .B1(n6135), .B2(n4965), .ZN(n6621)
         );
  OAI221_X1 U2494 ( .B1(n6352), .B2(n6144), .C1(n3655), .C2(n6141), .A(n6621), 
        .ZN(n6629) );
  AOI22_X1 U2495 ( .A1(n2919), .A2(n6149), .B1(n7103), .B2(n6146), .ZN(n6622)
         );
  OAI221_X1 U2496 ( .B1(n4795), .B2(n6155), .C1(n7105), .C2(n6152), .A(n6622), 
        .ZN(n6625) );
  NAND2_X1 U2497 ( .A1(n6159), .A2(n7107), .ZN(n6623) );
  NAND4_X1 U2498 ( .A1(n1839), .A2(n1840), .A3(n1838), .A4(n6623), .ZN(n6624)
         );
  OAI21_X1 U2499 ( .B1(n6625), .B2(n6624), .A(n6162), .ZN(n6627) );
  AOI22_X1 U2500 ( .A1(n6167), .A2(n7101), .B1(n6164), .B2(n4934), .ZN(n6626)
         );
  OAI211_X1 U2501 ( .C1(n2229), .C2(n6170), .A(n6627), .B(n6626), .ZN(n6628)
         );
  NOR4_X1 U2502 ( .A1(n6631), .A2(n6630), .A3(n6629), .A4(n6628), .ZN(n6632)
         );
  OAI21_X1 U2503 ( .B1(n2631), .B2(n6175), .A(n6632), .ZN(n2992) );
  OAI222_X1 U2504 ( .A1(n4709), .A2(n6121), .B1(n2728), .B2(n6119), .C1(n2134), 
        .C2(n6116), .ZN(n6644) );
  INV_X1 U2505 ( .A(n2166), .ZN(n7563) );
  AOI22_X1 U2506 ( .A1(n6127), .A2(n2856), .B1(n6124), .B2(n7563), .ZN(n6633)
         );
  OAI221_X1 U2507 ( .B1(n2070), .B2(n6133), .C1(n2102), .C2(n6130), .A(n6633), 
        .ZN(n6643) );
  AOI22_X1 U2508 ( .A1(n6138), .A2(n5024), .B1(n6135), .B2(n4964), .ZN(n6634)
         );
  OAI221_X1 U2509 ( .B1(n6353), .B2(n6144), .C1(n3656), .C2(n6141), .A(n6634), 
        .ZN(n6642) );
  AOI22_X1 U2510 ( .A1(n2920), .A2(n6149), .B1(n7122), .B2(n6146), .ZN(n6635)
         );
  OAI221_X1 U2511 ( .B1(n4793), .B2(n6155), .C1(n7124), .C2(n6152), .A(n6635), 
        .ZN(n6638) );
  NAND2_X1 U2512 ( .A1(n6159), .A2(n7126), .ZN(n6636) );
  NAND4_X1 U2513 ( .A1(n1822), .A2(n1823), .A3(n1821), .A4(n6636), .ZN(n6637)
         );
  OAI21_X1 U2514 ( .B1(n6638), .B2(n6637), .A(n6162), .ZN(n6640) );
  AOI22_X1 U2515 ( .A1(n6167), .A2(n7120), .B1(n6164), .B2(n4933), .ZN(n6639)
         );
  OAI211_X1 U2516 ( .C1(n2230), .C2(n6170), .A(n6640), .B(n6639), .ZN(n6641)
         );
  NOR4_X1 U2517 ( .A1(n6644), .A2(n6643), .A3(n6642), .A4(n6641), .ZN(n6645)
         );
  OAI21_X1 U2518 ( .B1(n2632), .B2(n6175), .A(n6645), .ZN(n2993) );
  OAI222_X1 U2519 ( .A1(n4707), .A2(n6121), .B1(n2729), .B2(n6119), .C1(n2135), 
        .C2(n6116), .ZN(n6657) );
  INV_X1 U2520 ( .A(n2167), .ZN(n7564) );
  AOI22_X1 U2521 ( .A1(n6127), .A2(n2857), .B1(n6124), .B2(n7564), .ZN(n6646)
         );
  OAI221_X1 U2522 ( .B1(n2071), .B2(n6133), .C1(n2103), .C2(n6130), .A(n6646), 
        .ZN(n6656) );
  AOI22_X1 U2523 ( .A1(n6138), .A2(n5023), .B1(n6135), .B2(n4963), .ZN(n6647)
         );
  OAI221_X1 U2524 ( .B1(n6354), .B2(n6144), .C1(n3657), .C2(n6141), .A(n6647), 
        .ZN(n6655) );
  AOI22_X1 U2525 ( .A1(n2921), .A2(n6149), .B1(n7141), .B2(n6146), .ZN(n6648)
         );
  OAI221_X1 U2526 ( .B1(n4791), .B2(n6155), .C1(n7143), .C2(n6152), .A(n6648), 
        .ZN(n6651) );
  NAND2_X1 U2527 ( .A1(n6159), .A2(n7145), .ZN(n6649) );
  NAND4_X1 U2528 ( .A1(n1805), .A2(n1806), .A3(n1804), .A4(n6649), .ZN(n6650)
         );
  OAI21_X1 U2529 ( .B1(n6651), .B2(n6650), .A(n6162), .ZN(n6653) );
  AOI22_X1 U2530 ( .A1(n6167), .A2(n7139), .B1(n6164), .B2(n4932), .ZN(n6652)
         );
  OAI211_X1 U2531 ( .C1(n2231), .C2(n6170), .A(n6653), .B(n6652), .ZN(n6654)
         );
  NOR4_X1 U2532 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(n6658)
         );
  OAI21_X1 U2533 ( .B1(n2633), .B2(n6175), .A(n6658), .ZN(n2994) );
  OAI222_X1 U2534 ( .A1(n4717), .A2(n6122), .B1(n2730), .B2(n6119), .C1(n2136), 
        .C2(n6117), .ZN(n6670) );
  INV_X1 U2535 ( .A(n2168), .ZN(n7565) );
  AOI22_X1 U2536 ( .A1(n6127), .A2(n2858), .B1(n6125), .B2(n7565), .ZN(n6659)
         );
  OAI221_X1 U2537 ( .B1(n2072), .B2(n6133), .C1(n2104), .C2(n6131), .A(n6659), 
        .ZN(n6669) );
  AOI22_X1 U2538 ( .A1(n6138), .A2(n5022), .B1(n6136), .B2(n4962), .ZN(n6660)
         );
  OAI221_X1 U2539 ( .B1(n6355), .B2(n6144), .C1(n3658), .C2(n6142), .A(n6660), 
        .ZN(n6668) );
  AOI22_X1 U2540 ( .A1(n2922), .A2(n6150), .B1(n7160), .B2(n6147), .ZN(n6661)
         );
  OAI221_X1 U2541 ( .B1(n4789), .B2(n6156), .C1(n7162), .C2(n6153), .A(n6661), 
        .ZN(n6664) );
  NAND2_X1 U2542 ( .A1(n6159), .A2(n7164), .ZN(n6662) );
  NAND4_X1 U2543 ( .A1(n1788), .A2(n1789), .A3(n1787), .A4(n6662), .ZN(n6663)
         );
  OAI21_X1 U2544 ( .B1(n6664), .B2(n6663), .A(n6162), .ZN(n6666) );
  AOI22_X1 U2545 ( .A1(n6167), .A2(n7158), .B1(n6165), .B2(n4931), .ZN(n6665)
         );
  OAI211_X1 U2546 ( .C1(n2232), .C2(n6171), .A(n6666), .B(n6665), .ZN(n6667)
         );
  NOR4_X1 U2547 ( .A1(n6670), .A2(n6669), .A3(n6668), .A4(n6667), .ZN(n6671)
         );
  OAI21_X1 U2548 ( .B1(n2634), .B2(n6174), .A(n6671), .ZN(n2995) );
  OAI222_X1 U2549 ( .A1(n4715), .A2(n6122), .B1(n2731), .B2(n6120), .C1(n2137), 
        .C2(n6117), .ZN(n6683) );
  INV_X1 U2550 ( .A(n2169), .ZN(n7566) );
  AOI22_X1 U2551 ( .A1(n6128), .A2(n2859), .B1(n6125), .B2(n7566), .ZN(n6672)
         );
  OAI221_X1 U2552 ( .B1(n2073), .B2(n6134), .C1(n2105), .C2(n6131), .A(n6672), 
        .ZN(n6682) );
  AOI22_X1 U2553 ( .A1(n6139), .A2(n5021), .B1(n6136), .B2(n4961), .ZN(n6673)
         );
  OAI221_X1 U2554 ( .B1(n6356), .B2(n6145), .C1(n3659), .C2(n6142), .A(n6673), 
        .ZN(n6681) );
  AOI22_X1 U2555 ( .A1(n2923), .A2(n6150), .B1(n7179), .B2(n6147), .ZN(n6674)
         );
  OAI221_X1 U2556 ( .B1(n4787), .B2(n6156), .C1(n7181), .C2(n6153), .A(n6674), 
        .ZN(n6677) );
  NAND2_X1 U2557 ( .A1(n6159), .A2(n7183), .ZN(n6675) );
  NAND4_X1 U2558 ( .A1(n1771), .A2(n1772), .A3(n1770), .A4(n6675), .ZN(n6676)
         );
  OAI21_X1 U2559 ( .B1(n6677), .B2(n6676), .A(n6162), .ZN(n6679) );
  AOI22_X1 U2560 ( .A1(n6168), .A2(n7177), .B1(n6165), .B2(n4930), .ZN(n6678)
         );
  OAI211_X1 U2561 ( .C1(n2233), .C2(n6171), .A(n6679), .B(n6678), .ZN(n6680)
         );
  NOR4_X1 U2562 ( .A1(n6683), .A2(n6682), .A3(n6681), .A4(n6680), .ZN(n6684)
         );
  OAI21_X1 U2563 ( .B1(n2635), .B2(n6174), .A(n6684), .ZN(n2996) );
  OAI222_X1 U2564 ( .A1(n4713), .A2(n6122), .B1(n2732), .B2(n6120), .C1(n2138), 
        .C2(n6117), .ZN(n6696) );
  INV_X1 U2565 ( .A(n2170), .ZN(n7567) );
  AOI22_X1 U2566 ( .A1(n6128), .A2(n2860), .B1(n6125), .B2(n7567), .ZN(n6685)
         );
  OAI221_X1 U2567 ( .B1(n2074), .B2(n6134), .C1(n2106), .C2(n6131), .A(n6685), 
        .ZN(n6695) );
  AOI22_X1 U2568 ( .A1(n6139), .A2(n5020), .B1(n6136), .B2(n4960), .ZN(n6686)
         );
  OAI221_X1 U2569 ( .B1(n6357), .B2(n6145), .C1(n3660), .C2(n6142), .A(n6686), 
        .ZN(n6694) );
  AOI22_X1 U2570 ( .A1(n2924), .A2(n6150), .B1(n7198), .B2(n6147), .ZN(n6687)
         );
  OAI221_X1 U2571 ( .B1(n4785), .B2(n6156), .C1(n7200), .C2(n6153), .A(n6687), 
        .ZN(n6690) );
  NAND2_X1 U2572 ( .A1(n6159), .A2(n7202), .ZN(n6688) );
  NAND4_X1 U2573 ( .A1(n1754), .A2(n1755), .A3(n1753), .A4(n6688), .ZN(n6689)
         );
  OAI21_X1 U2574 ( .B1(n6690), .B2(n6689), .A(n6162), .ZN(n6692) );
  AOI22_X1 U2575 ( .A1(n6168), .A2(n7196), .B1(n6165), .B2(n4929), .ZN(n6691)
         );
  OAI211_X1 U2576 ( .C1(n2234), .C2(n6171), .A(n6692), .B(n6691), .ZN(n6693)
         );
  NOR4_X1 U2577 ( .A1(n6696), .A2(n6695), .A3(n6694), .A4(n6693), .ZN(n6697)
         );
  OAI21_X1 U2578 ( .B1(n2636), .B2(n6174), .A(n6697), .ZN(n2997) );
  OAI222_X1 U2579 ( .A1(n4723), .A2(n6122), .B1(n2733), .B2(n6120), .C1(n2139), 
        .C2(n6117), .ZN(n6709) );
  INV_X1 U2580 ( .A(n2171), .ZN(n7568) );
  AOI22_X1 U2581 ( .A1(n6128), .A2(n2861), .B1(n6125), .B2(n7568), .ZN(n6698)
         );
  OAI221_X1 U2582 ( .B1(n2075), .B2(n6134), .C1(n2107), .C2(n6131), .A(n6698), 
        .ZN(n6708) );
  AOI22_X1 U2583 ( .A1(n6139), .A2(n5019), .B1(n6136), .B2(n4959), .ZN(n6699)
         );
  OAI221_X1 U2584 ( .B1(n6358), .B2(n6145), .C1(n3661), .C2(n6142), .A(n6699), 
        .ZN(n6707) );
  AOI22_X1 U2585 ( .A1(n2925), .A2(n6150), .B1(n7217), .B2(n6147), .ZN(n6700)
         );
  OAI221_X1 U2586 ( .B1(n4783), .B2(n6156), .C1(n7219), .C2(n6153), .A(n6700), 
        .ZN(n6703) );
  NAND2_X1 U2587 ( .A1(n6159), .A2(n7221), .ZN(n6701) );
  NAND4_X1 U2588 ( .A1(n1737), .A2(n1738), .A3(n1736), .A4(n6701), .ZN(n6702)
         );
  OAI21_X1 U2589 ( .B1(n6703), .B2(n6702), .A(n6162), .ZN(n6705) );
  AOI22_X1 U2590 ( .A1(n6168), .A2(n7215), .B1(n6165), .B2(n4928), .ZN(n6704)
         );
  OAI211_X1 U2591 ( .C1(n2235), .C2(n6171), .A(n6705), .B(n6704), .ZN(n6706)
         );
  NOR4_X1 U2592 ( .A1(n6709), .A2(n6708), .A3(n6707), .A4(n6706), .ZN(n6710)
         );
  OAI21_X1 U2593 ( .B1(n2637), .B2(n6174), .A(n6710), .ZN(n2998) );
  OAI222_X1 U2594 ( .A1(n4721), .A2(n6122), .B1(n2734), .B2(n6120), .C1(n2140), 
        .C2(n6117), .ZN(n6722) );
  INV_X1 U2595 ( .A(n2172), .ZN(n7569) );
  AOI22_X1 U2596 ( .A1(n6128), .A2(n2862), .B1(n6125), .B2(n7569), .ZN(n6711)
         );
  OAI221_X1 U2597 ( .B1(n2076), .B2(n6134), .C1(n2108), .C2(n6131), .A(n6711), 
        .ZN(n6721) );
  AOI22_X1 U2598 ( .A1(n6139), .A2(n5018), .B1(n6136), .B2(n4958), .ZN(n6712)
         );
  OAI221_X1 U2599 ( .B1(n6359), .B2(n6145), .C1(n3662), .C2(n6142), .A(n6712), 
        .ZN(n6720) );
  AOI22_X1 U2600 ( .A1(n2926), .A2(n6150), .B1(n7236), .B2(n6147), .ZN(n6713)
         );
  OAI221_X1 U2601 ( .B1(n4753), .B2(n6156), .C1(n7238), .C2(n6153), .A(n6713), 
        .ZN(n6716) );
  NAND2_X1 U2602 ( .A1(n6159), .A2(n7240), .ZN(n6714) );
  NAND4_X1 U2603 ( .A1(n1720), .A2(n1721), .A3(n1719), .A4(n6714), .ZN(n6715)
         );
  OAI21_X1 U2604 ( .B1(n6716), .B2(n6715), .A(n6162), .ZN(n6718) );
  AOI22_X1 U2605 ( .A1(n6168), .A2(n7234), .B1(n6165), .B2(n4927), .ZN(n6717)
         );
  OAI211_X1 U2606 ( .C1(n2236), .C2(n6171), .A(n6718), .B(n6717), .ZN(n6719)
         );
  NOR4_X1 U2607 ( .A1(n6722), .A2(n6721), .A3(n6720), .A4(n6719), .ZN(n6723)
         );
  OAI21_X1 U2608 ( .B1(n2638), .B2(n6174), .A(n6723), .ZN(n2999) );
  OAI222_X1 U2609 ( .A1(n4719), .A2(n6122), .B1(n2735), .B2(n6120), .C1(n2141), 
        .C2(n6117), .ZN(n6735) );
  INV_X1 U2610 ( .A(n2173), .ZN(n7570) );
  AOI22_X1 U2611 ( .A1(n6128), .A2(n2863), .B1(n6125), .B2(n7570), .ZN(n6724)
         );
  OAI221_X1 U2612 ( .B1(n2077), .B2(n6134), .C1(n2109), .C2(n6131), .A(n6724), 
        .ZN(n6734) );
  AOI22_X1 U2613 ( .A1(n6139), .A2(n5017), .B1(n6136), .B2(n4957), .ZN(n6725)
         );
  OAI221_X1 U2614 ( .B1(n6360), .B2(n6145), .C1(n3663), .C2(n6142), .A(n6725), 
        .ZN(n6733) );
  AOI22_X1 U2615 ( .A1(n2927), .A2(n6150), .B1(n7255), .B2(n6147), .ZN(n6726)
         );
  OAI221_X1 U2616 ( .B1(n4763), .B2(n6156), .C1(n7257), .C2(n6153), .A(n6726), 
        .ZN(n6729) );
  NAND2_X1 U2617 ( .A1(n6159), .A2(n7259), .ZN(n6727) );
  NAND4_X1 U2618 ( .A1(n1703), .A2(n1704), .A3(n1702), .A4(n6727), .ZN(n6728)
         );
  OAI21_X1 U2619 ( .B1(n6729), .B2(n6728), .A(n6162), .ZN(n6731) );
  AOI22_X1 U2620 ( .A1(n6168), .A2(n7253), .B1(n6165), .B2(n4926), .ZN(n6730)
         );
  OAI211_X1 U2621 ( .C1(n2237), .C2(n6171), .A(n6731), .B(n6730), .ZN(n6732)
         );
  NOR4_X1 U2622 ( .A1(n6735), .A2(n6734), .A3(n6733), .A4(n6732), .ZN(n6736)
         );
  OAI21_X1 U2623 ( .B1(n2639), .B2(n6174), .A(n6736), .ZN(n3000) );
  OAI222_X1 U2624 ( .A1(n4729), .A2(n6122), .B1(n2736), .B2(n6120), .C1(n2142), 
        .C2(n6117), .ZN(n6748) );
  INV_X1 U2625 ( .A(n2174), .ZN(n7571) );
  AOI22_X1 U2626 ( .A1(n6128), .A2(n2864), .B1(n6125), .B2(n7571), .ZN(n6737)
         );
  OAI221_X1 U2627 ( .B1(n2078), .B2(n6134), .C1(n2110), .C2(n6131), .A(n6737), 
        .ZN(n6747) );
  AOI22_X1 U2628 ( .A1(n6139), .A2(n5016), .B1(n6136), .B2(n4956), .ZN(n6738)
         );
  OAI221_X1 U2629 ( .B1(n6361), .B2(n6145), .C1(n3664), .C2(n6142), .A(n6738), 
        .ZN(n6746) );
  AOI22_X1 U2630 ( .A1(n2928), .A2(n6150), .B1(n7274), .B2(n6147), .ZN(n6739)
         );
  OAI221_X1 U2631 ( .B1(n4757), .B2(n6156), .C1(n7276), .C2(n6153), .A(n6739), 
        .ZN(n6742) );
  NAND2_X1 U2632 ( .A1(n6159), .A2(n7278), .ZN(n6740) );
  NAND4_X1 U2633 ( .A1(n1686), .A2(n1687), .A3(n1685), .A4(n6740), .ZN(n6741)
         );
  OAI21_X1 U2634 ( .B1(n6742), .B2(n6741), .A(n6162), .ZN(n6744) );
  AOI22_X1 U2635 ( .A1(n6168), .A2(n7272), .B1(n6165), .B2(n4925), .ZN(n6743)
         );
  OAI211_X1 U2636 ( .C1(n2238), .C2(n6171), .A(n6744), .B(n6743), .ZN(n6745)
         );
  NOR4_X1 U2637 ( .A1(n6748), .A2(n6747), .A3(n6746), .A4(n6745), .ZN(n6749)
         );
  OAI21_X1 U2638 ( .B1(n2640), .B2(n6174), .A(n6749), .ZN(n3001) );
  OAI222_X1 U2639 ( .A1(n4727), .A2(n6122), .B1(n2737), .B2(n6120), .C1(n2143), 
        .C2(n6117), .ZN(n6761) );
  INV_X1 U2640 ( .A(n2175), .ZN(n7572) );
  AOI22_X1 U2641 ( .A1(n6128), .A2(n2865), .B1(n6125), .B2(n7572), .ZN(n6750)
         );
  OAI221_X1 U2642 ( .B1(n2079), .B2(n6134), .C1(n2111), .C2(n6131), .A(n6750), 
        .ZN(n6760) );
  AOI22_X1 U2643 ( .A1(n6139), .A2(n5015), .B1(n6136), .B2(n4955), .ZN(n6751)
         );
  OAI221_X1 U2644 ( .B1(n6362), .B2(n6145), .C1(n3665), .C2(n6142), .A(n6751), 
        .ZN(n6759) );
  AOI22_X1 U2645 ( .A1(n2929), .A2(n6150), .B1(n7293), .B2(n6147), .ZN(n6752)
         );
  OAI221_X1 U2646 ( .B1(n4759), .B2(n6156), .C1(n7295), .C2(n6153), .A(n6752), 
        .ZN(n6755) );
  NAND2_X1 U2647 ( .A1(n6159), .A2(n7297), .ZN(n6753) );
  NAND4_X1 U2648 ( .A1(n1669), .A2(n1670), .A3(n1668), .A4(n6753), .ZN(n6754)
         );
  OAI21_X1 U2649 ( .B1(n6755), .B2(n6754), .A(n6161), .ZN(n6757) );
  AOI22_X1 U2650 ( .A1(n6168), .A2(n7291), .B1(n6165), .B2(n4924), .ZN(n6756)
         );
  OAI211_X1 U2651 ( .C1(n2239), .C2(n6171), .A(n6757), .B(n6756), .ZN(n6758)
         );
  NOR4_X1 U2652 ( .A1(n6761), .A2(n6760), .A3(n6759), .A4(n6758), .ZN(n6762)
         );
  OAI21_X1 U2653 ( .B1(n2641), .B2(n6174), .A(n6762), .ZN(n3002) );
  OAI222_X1 U2654 ( .A1(n4725), .A2(n6122), .B1(n2738), .B2(n6120), .C1(n2144), 
        .C2(n6117), .ZN(n6774) );
  INV_X1 U2655 ( .A(n2176), .ZN(n7573) );
  AOI22_X1 U2656 ( .A1(n6128), .A2(n2866), .B1(n6125), .B2(n7573), .ZN(n6763)
         );
  OAI221_X1 U2657 ( .B1(n2080), .B2(n6134), .C1(n2112), .C2(n6131), .A(n6763), 
        .ZN(n6773) );
  AOI22_X1 U2658 ( .A1(n6139), .A2(n5014), .B1(n6136), .B2(n4954), .ZN(n6764)
         );
  OAI221_X1 U2659 ( .B1(n6363), .B2(n6145), .C1(n3666), .C2(n6142), .A(n6764), 
        .ZN(n6772) );
  AOI22_X1 U2660 ( .A1(n2930), .A2(n6150), .B1(n7312), .B2(n6147), .ZN(n6765)
         );
  OAI221_X1 U2661 ( .B1(n4769), .B2(n6156), .C1(n7314), .C2(n6153), .A(n6765), 
        .ZN(n6768) );
  NAND2_X1 U2662 ( .A1(n6158), .A2(n7316), .ZN(n6766) );
  NAND4_X1 U2663 ( .A1(n1652), .A2(n1653), .A3(n1651), .A4(n6766), .ZN(n6767)
         );
  OAI21_X1 U2664 ( .B1(n6768), .B2(n6767), .A(n6161), .ZN(n6770) );
  AOI22_X1 U2665 ( .A1(n6168), .A2(n7310), .B1(n6165), .B2(n4923), .ZN(n6769)
         );
  OAI211_X1 U2666 ( .C1(n2240), .C2(n6171), .A(n6770), .B(n6769), .ZN(n6771)
         );
  NOR4_X1 U2667 ( .A1(n6774), .A2(n6773), .A3(n6772), .A4(n6771), .ZN(n6775)
         );
  OAI21_X1 U2668 ( .B1(n2642), .B2(n6174), .A(n6775), .ZN(n3003) );
  OAI222_X1 U2669 ( .A1(n4735), .A2(n6122), .B1(n2739), .B2(n6120), .C1(n2145), 
        .C2(n6117), .ZN(n6787) );
  INV_X1 U2670 ( .A(n2177), .ZN(n7574) );
  AOI22_X1 U2671 ( .A1(n6128), .A2(n2867), .B1(n6125), .B2(n7574), .ZN(n6776)
         );
  OAI221_X1 U2672 ( .B1(n2081), .B2(n6134), .C1(n2113), .C2(n6131), .A(n6776), 
        .ZN(n6786) );
  AOI22_X1 U2673 ( .A1(n6139), .A2(n5013), .B1(n6136), .B2(n4953), .ZN(n6777)
         );
  OAI221_X1 U2674 ( .B1(n6364), .B2(n6145), .C1(n3667), .C2(n6142), .A(n6777), 
        .ZN(n6785) );
  AOI22_X1 U2675 ( .A1(n2931), .A2(n6150), .B1(n7331), .B2(n6147), .ZN(n6778)
         );
  OAI221_X1 U2676 ( .B1(n4761), .B2(n6156), .C1(n7333), .C2(n6153), .A(n6778), 
        .ZN(n6781) );
  NAND2_X1 U2677 ( .A1(n6158), .A2(n7335), .ZN(n6779) );
  NAND4_X1 U2678 ( .A1(n1635), .A2(n1636), .A3(n1634), .A4(n6779), .ZN(n6780)
         );
  OAI21_X1 U2679 ( .B1(n6781), .B2(n6780), .A(n6161), .ZN(n6783) );
  AOI22_X1 U2680 ( .A1(n6168), .A2(n7329), .B1(n6165), .B2(n4922), .ZN(n6782)
         );
  OAI211_X1 U2681 ( .C1(n2241), .C2(n6171), .A(n6783), .B(n6782), .ZN(n6784)
         );
  NOR4_X1 U2682 ( .A1(n6787), .A2(n6786), .A3(n6785), .A4(n6784), .ZN(n6788)
         );
  OAI21_X1 U2683 ( .B1(n2643), .B2(n6174), .A(n6788), .ZN(n3004) );
  OAI222_X1 U2684 ( .A1(n4733), .A2(n6122), .B1(n2740), .B2(n6120), .C1(n2146), 
        .C2(n6117), .ZN(n6800) );
  INV_X1 U2685 ( .A(n2178), .ZN(n7575) );
  AOI22_X1 U2686 ( .A1(n6128), .A2(n2868), .B1(n6125), .B2(n7575), .ZN(n6789)
         );
  OAI221_X1 U2687 ( .B1(n2082), .B2(n6134), .C1(n2114), .C2(n6131), .A(n6789), 
        .ZN(n6799) );
  AOI22_X1 U2688 ( .A1(n6139), .A2(n5012), .B1(n6136), .B2(n4952), .ZN(n6790)
         );
  OAI221_X1 U2689 ( .B1(n6365), .B2(n6145), .C1(n3668), .C2(n6142), .A(n6790), 
        .ZN(n6798) );
  AOI22_X1 U2690 ( .A1(n2932), .A2(n6150), .B1(n7350), .B2(n6147), .ZN(n6791)
         );
  OAI221_X1 U2691 ( .B1(n4765), .B2(n6156), .C1(n7352), .C2(n6153), .A(n6791), 
        .ZN(n6794) );
  NAND2_X1 U2692 ( .A1(n6158), .A2(n7354), .ZN(n6792) );
  NAND4_X1 U2693 ( .A1(n1618), .A2(n1619), .A3(n1617), .A4(n6792), .ZN(n6793)
         );
  OAI21_X1 U2694 ( .B1(n6794), .B2(n6793), .A(n6161), .ZN(n6796) );
  AOI22_X1 U2695 ( .A1(n6168), .A2(n7348), .B1(n6165), .B2(n4921), .ZN(n6795)
         );
  OAI211_X1 U2696 ( .C1(n2242), .C2(n6171), .A(n6796), .B(n6795), .ZN(n6797)
         );
  NOR4_X1 U2697 ( .A1(n6800), .A2(n6799), .A3(n6798), .A4(n6797), .ZN(n6801)
         );
  OAI21_X1 U2698 ( .B1(n2644), .B2(n6174), .A(n6801), .ZN(n3005) );
  OAI222_X1 U2699 ( .A1(n4731), .A2(n6122), .B1(n2741), .B2(n6120), .C1(n2147), 
        .C2(n6117), .ZN(n6813) );
  INV_X1 U2700 ( .A(n2179), .ZN(n7576) );
  AOI22_X1 U2701 ( .A1(n6128), .A2(n2869), .B1(n6125), .B2(n7576), .ZN(n6802)
         );
  OAI221_X1 U2702 ( .B1(n2083), .B2(n6134), .C1(n2115), .C2(n6131), .A(n6802), 
        .ZN(n6812) );
  AOI22_X1 U2703 ( .A1(n6139), .A2(n5011), .B1(n6136), .B2(n4951), .ZN(n6803)
         );
  OAI221_X1 U2704 ( .B1(n6366), .B2(n6145), .C1(n3669), .C2(n6142), .A(n6803), 
        .ZN(n6811) );
  AOI22_X1 U2705 ( .A1(n2933), .A2(n6150), .B1(n7369), .B2(n6147), .ZN(n6804)
         );
  OAI221_X1 U2706 ( .B1(n4771), .B2(n6156), .C1(n7371), .C2(n6153), .A(n6804), 
        .ZN(n6807) );
  NAND2_X1 U2707 ( .A1(n6158), .A2(n7373), .ZN(n6805) );
  NAND4_X1 U2708 ( .A1(n1601), .A2(n1602), .A3(n1600), .A4(n6805), .ZN(n6806)
         );
  OAI21_X1 U2709 ( .B1(n6807), .B2(n6806), .A(n6161), .ZN(n6809) );
  AOI22_X1 U2710 ( .A1(n6168), .A2(n7367), .B1(n6165), .B2(n4920), .ZN(n6808)
         );
  OAI211_X1 U2711 ( .C1(n2243), .C2(n6171), .A(n6809), .B(n6808), .ZN(n6810)
         );
  NOR4_X1 U2712 ( .A1(n6813), .A2(n6812), .A3(n6811), .A4(n6810), .ZN(n6814)
         );
  OAI21_X1 U2713 ( .B1(n2645), .B2(n6173), .A(n6814), .ZN(n3006) );
  OAI222_X1 U2714 ( .A1(n4741), .A2(n6123), .B1(n2742), .B2(n6120), .C1(n2148), 
        .C2(n6118), .ZN(n6826) );
  INV_X1 U2715 ( .A(n2180), .ZN(n7577) );
  AOI22_X1 U2716 ( .A1(n6128), .A2(n2870), .B1(n6126), .B2(n7577), .ZN(n6815)
         );
  OAI221_X1 U2717 ( .B1(n2084), .B2(n6134), .C1(n2116), .C2(n6132), .A(n6815), 
        .ZN(n6825) );
  AOI22_X1 U2718 ( .A1(n6139), .A2(n5010), .B1(n6137), .B2(n4950), .ZN(n6816)
         );
  OAI221_X1 U2719 ( .B1(n6367), .B2(n6145), .C1(n3670), .C2(n6143), .A(n6816), 
        .ZN(n6824) );
  AOI22_X1 U2720 ( .A1(n2934), .A2(n6151), .B1(n7388), .B2(n6148), .ZN(n6817)
         );
  OAI221_X1 U2721 ( .B1(n4767), .B2(n6157), .C1(n7390), .C2(n6154), .A(n6817), 
        .ZN(n6820) );
  NAND2_X1 U2722 ( .A1(n6158), .A2(n7392), .ZN(n6818) );
  NAND4_X1 U2723 ( .A1(n1584), .A2(n1585), .A3(n1583), .A4(n6818), .ZN(n6819)
         );
  OAI21_X1 U2724 ( .B1(n6820), .B2(n6819), .A(n6161), .ZN(n6822) );
  AOI22_X1 U2725 ( .A1(n6168), .A2(n7386), .B1(n6166), .B2(n4919), .ZN(n6821)
         );
  OAI211_X1 U2726 ( .C1(n2244), .C2(n6172), .A(n6822), .B(n6821), .ZN(n6823)
         );
  NOR4_X1 U2727 ( .A1(n6826), .A2(n6825), .A3(n6824), .A4(n6823), .ZN(n6827)
         );
  OAI21_X1 U2728 ( .B1(n2646), .B2(n6173), .A(n6827), .ZN(n3007) );
  OAI222_X1 U2729 ( .A1(n4739), .A2(n6123), .B1(n2743), .B2(n6119), .C1(n2149), 
        .C2(n6118), .ZN(n6839) );
  INV_X1 U2730 ( .A(n2181), .ZN(n7578) );
  AOI22_X1 U2731 ( .A1(n6129), .A2(n2871), .B1(n6126), .B2(n7578), .ZN(n6828)
         );
  OAI221_X1 U2732 ( .B1(n2085), .B2(n6133), .C1(n2117), .C2(n6132), .A(n6828), 
        .ZN(n6838) );
  AOI22_X1 U2733 ( .A1(n6140), .A2(n5009), .B1(n6137), .B2(n4949), .ZN(n6829)
         );
  OAI221_X1 U2734 ( .B1(n6368), .B2(n6144), .C1(n3671), .C2(n6143), .A(n6829), 
        .ZN(n6837) );
  AOI22_X1 U2735 ( .A1(n2935), .A2(n6151), .B1(n7407), .B2(n6148), .ZN(n6830)
         );
  OAI221_X1 U2736 ( .B1(n4775), .B2(n6157), .C1(n7409), .C2(n6154), .A(n6830), 
        .ZN(n6833) );
  NAND2_X1 U2737 ( .A1(n6158), .A2(n7411), .ZN(n6831) );
  NAND4_X1 U2738 ( .A1(n1567), .A2(n1568), .A3(n1566), .A4(n6831), .ZN(n6832)
         );
  OAI21_X1 U2739 ( .B1(n6833), .B2(n6832), .A(n6161), .ZN(n6835) );
  AOI22_X1 U2740 ( .A1(n6169), .A2(n7405), .B1(n6166), .B2(n4918), .ZN(n6834)
         );
  OAI211_X1 U2741 ( .C1(n2245), .C2(n6172), .A(n6835), .B(n6834), .ZN(n6836)
         );
  NOR4_X1 U2742 ( .A1(n6839), .A2(n6838), .A3(n6837), .A4(n6836), .ZN(n6840)
         );
  OAI21_X1 U2743 ( .B1(n2647), .B2(n6173), .A(n6840), .ZN(n3008) );
  OAI222_X1 U2744 ( .A1(n4737), .A2(n6123), .B1(n2744), .B2(n6120), .C1(n2150), 
        .C2(n6118), .ZN(n6852) );
  INV_X1 U2745 ( .A(n2182), .ZN(n7579) );
  AOI22_X1 U2746 ( .A1(n6129), .A2(n2872), .B1(n6126), .B2(n7579), .ZN(n6841)
         );
  OAI221_X1 U2747 ( .B1(n2086), .B2(n6134), .C1(n2118), .C2(n6132), .A(n6841), 
        .ZN(n6851) );
  AOI22_X1 U2748 ( .A1(n6140), .A2(n5008), .B1(n6137), .B2(n4948), .ZN(n6842)
         );
  OAI221_X1 U2749 ( .B1(n6369), .B2(n6145), .C1(n3672), .C2(n6143), .A(n6842), 
        .ZN(n6850) );
  AOI22_X1 U2750 ( .A1(n2936), .A2(n6151), .B1(n7426), .B2(n6148), .ZN(n6843)
         );
  OAI221_X1 U2751 ( .B1(n4773), .B2(n6157), .C1(n7428), .C2(n6154), .A(n6843), 
        .ZN(n6846) );
  NAND2_X1 U2752 ( .A1(n6158), .A2(n7430), .ZN(n6844) );
  NAND4_X1 U2753 ( .A1(n1550), .A2(n1551), .A3(n1549), .A4(n6844), .ZN(n6845)
         );
  OAI21_X1 U2754 ( .B1(n6846), .B2(n6845), .A(n6161), .ZN(n6848) );
  AOI22_X1 U2755 ( .A1(n6169), .A2(n7424), .B1(n6166), .B2(n4917), .ZN(n6847)
         );
  OAI211_X1 U2756 ( .C1(n2246), .C2(n6172), .A(n6848), .B(n6847), .ZN(n6849)
         );
  NOR4_X1 U2757 ( .A1(n6852), .A2(n6851), .A3(n6850), .A4(n6849), .ZN(n6853)
         );
  OAI21_X1 U2758 ( .B1(n2648), .B2(n6173), .A(n6853), .ZN(n3009) );
  OAI222_X1 U2759 ( .A1(n4747), .A2(n6123), .B1(n2745), .B2(n6119), .C1(n2151), 
        .C2(n6118), .ZN(n6865) );
  INV_X1 U2760 ( .A(n2183), .ZN(n7580) );
  AOI22_X1 U2761 ( .A1(n6129), .A2(n2873), .B1(n6126), .B2(n7580), .ZN(n6854)
         );
  OAI221_X1 U2762 ( .B1(n2087), .B2(n6133), .C1(n2119), .C2(n6132), .A(n6854), 
        .ZN(n6864) );
  AOI22_X1 U2763 ( .A1(n6140), .A2(n5007), .B1(n6137), .B2(n4947), .ZN(n6855)
         );
  OAI221_X1 U2764 ( .B1(n6370), .B2(n6144), .C1(n3673), .C2(n6143), .A(n6855), 
        .ZN(n6863) );
  AOI22_X1 U2765 ( .A1(n2937), .A2(n6151), .B1(n7445), .B2(n6148), .ZN(n6856)
         );
  OAI221_X1 U2766 ( .B1(n4755), .B2(n6157), .C1(n7447), .C2(n6154), .A(n6856), 
        .ZN(n6859) );
  NAND2_X1 U2767 ( .A1(n6158), .A2(n7449), .ZN(n6857) );
  NAND4_X1 U2768 ( .A1(n1533), .A2(n1534), .A3(n1532), .A4(n6857), .ZN(n6858)
         );
  OAI21_X1 U2769 ( .B1(n6859), .B2(n6858), .A(n6161), .ZN(n6861) );
  AOI22_X1 U2770 ( .A1(n6169), .A2(n7443), .B1(n6166), .B2(n4916), .ZN(n6860)
         );
  OAI211_X1 U2771 ( .C1(n2247), .C2(n6172), .A(n6861), .B(n6860), .ZN(n6862)
         );
  NOR4_X1 U2772 ( .A1(n6865), .A2(n6864), .A3(n6863), .A4(n6862), .ZN(n6866)
         );
  OAI21_X1 U2773 ( .B1(n2649), .B2(n6173), .A(n6866), .ZN(n3010) );
  OAI222_X1 U2774 ( .A1(n4745), .A2(n6123), .B1(n2746), .B2(n6120), .C1(n2152), 
        .C2(n6118), .ZN(n6878) );
  INV_X1 U2775 ( .A(n2184), .ZN(n7581) );
  AOI22_X1 U2776 ( .A1(n6129), .A2(n2874), .B1(n6126), .B2(n7581), .ZN(n6867)
         );
  OAI221_X1 U2777 ( .B1(n2088), .B2(n6134), .C1(n2120), .C2(n6132), .A(n6867), 
        .ZN(n6877) );
  AOI22_X1 U2778 ( .A1(n6140), .A2(n5006), .B1(n6137), .B2(n4946), .ZN(n6868)
         );
  OAI221_X1 U2779 ( .B1(n6371), .B2(n6145), .C1(n3674), .C2(n6143), .A(n6868), 
        .ZN(n6876) );
  AOI22_X1 U2780 ( .A1(n2938), .A2(n6151), .B1(n7464), .B2(n6148), .ZN(n6869)
         );
  OAI221_X1 U2781 ( .B1(n4779), .B2(n6157), .C1(n7466), .C2(n6154), .A(n6869), 
        .ZN(n6872) );
  NAND2_X1 U2782 ( .A1(n6158), .A2(n7468), .ZN(n6870) );
  NAND4_X1 U2783 ( .A1(n1516), .A2(n1517), .A3(n1515), .A4(n6870), .ZN(n6871)
         );
  OAI21_X1 U2784 ( .B1(n6872), .B2(n6871), .A(n6161), .ZN(n6874) );
  AOI22_X1 U2785 ( .A1(n6169), .A2(n7462), .B1(n6166), .B2(n4915), .ZN(n6873)
         );
  OAI211_X1 U2786 ( .C1(n2248), .C2(n6172), .A(n6874), .B(n6873), .ZN(n6875)
         );
  NOR4_X1 U2787 ( .A1(n6878), .A2(n6877), .A3(n6876), .A4(n6875), .ZN(n6879)
         );
  OAI21_X1 U2788 ( .B1(n2650), .B2(n6173), .A(n6879), .ZN(n3011) );
  OAI222_X1 U2789 ( .A1(n4743), .A2(n6123), .B1(n2747), .B2(n6119), .C1(n2153), 
        .C2(n6118), .ZN(n6891) );
  INV_X1 U2790 ( .A(n2185), .ZN(n7582) );
  AOI22_X1 U2791 ( .A1(n6129), .A2(n2875), .B1(n6126), .B2(n7582), .ZN(n6880)
         );
  OAI221_X1 U2792 ( .B1(n2089), .B2(n6133), .C1(n2121), .C2(n6132), .A(n6880), 
        .ZN(n6890) );
  AOI22_X1 U2793 ( .A1(n6140), .A2(n5005), .B1(n6137), .B2(n4945), .ZN(n6881)
         );
  OAI221_X1 U2794 ( .B1(n6372), .B2(n6144), .C1(n3675), .C2(n6143), .A(n6881), 
        .ZN(n6889) );
  AOI22_X1 U2795 ( .A1(n2939), .A2(n6151), .B1(n7483), .B2(n6148), .ZN(n6882)
         );
  OAI221_X1 U2796 ( .B1(n4777), .B2(n6157), .C1(n7485), .C2(n6154), .A(n6882), 
        .ZN(n6885) );
  NAND2_X1 U2797 ( .A1(n6158), .A2(n7487), .ZN(n6883) );
  NAND4_X1 U2798 ( .A1(n1499), .A2(n1500), .A3(n1498), .A4(n6883), .ZN(n6884)
         );
  OAI21_X1 U2799 ( .B1(n6885), .B2(n6884), .A(n6161), .ZN(n6887) );
  AOI22_X1 U2800 ( .A1(n6169), .A2(n7481), .B1(n6166), .B2(n4914), .ZN(n6886)
         );
  OAI211_X1 U2801 ( .C1(n2249), .C2(n6172), .A(n6887), .B(n6886), .ZN(n6888)
         );
  NOR4_X1 U2802 ( .A1(n6891), .A2(n6890), .A3(n6889), .A4(n6888), .ZN(n6892)
         );
  OAI21_X1 U2803 ( .B1(n2651), .B2(n6173), .A(n6892), .ZN(n3012) );
  OAI222_X1 U2804 ( .A1(n4749), .A2(n6123), .B1(n2748), .B2(n6120), .C1(n2154), 
        .C2(n6118), .ZN(n6904) );
  INV_X1 U2805 ( .A(n2186), .ZN(n7583) );
  AOI22_X1 U2806 ( .A1(n6129), .A2(n2876), .B1(n6126), .B2(n7583), .ZN(n6893)
         );
  OAI221_X1 U2807 ( .B1(n2090), .B2(n6134), .C1(n2122), .C2(n6132), .A(n6893), 
        .ZN(n6903) );
  AOI22_X1 U2808 ( .A1(n6140), .A2(n5004), .B1(n6137), .B2(n4944), .ZN(n6894)
         );
  OAI221_X1 U2809 ( .B1(n6373), .B2(n6145), .C1(n3676), .C2(n6143), .A(n6894), 
        .ZN(n6902) );
  AOI22_X1 U2810 ( .A1(n2940), .A2(n6151), .B1(n7502), .B2(n6148), .ZN(n6895)
         );
  OAI221_X1 U2811 ( .B1(n4781), .B2(n6157), .C1(n7504), .C2(n6154), .A(n6895), 
        .ZN(n6898) );
  NAND2_X1 U2812 ( .A1(n6158), .A2(n7506), .ZN(n6896) );
  NAND4_X1 U2813 ( .A1(n1482), .A2(n1483), .A3(n1481), .A4(n6896), .ZN(n6897)
         );
  OAI21_X1 U2814 ( .B1(n6898), .B2(n6897), .A(n6161), .ZN(n6900) );
  AOI22_X1 U2815 ( .A1(n6169), .A2(n7500), .B1(n6166), .B2(n4913), .ZN(n6899)
         );
  OAI211_X1 U2816 ( .C1(n2250), .C2(n6172), .A(n6900), .B(n6899), .ZN(n6901)
         );
  NOR4_X1 U2817 ( .A1(n6904), .A2(n6903), .A3(n6902), .A4(n6901), .ZN(n6905)
         );
  OAI21_X1 U2818 ( .B1(n2652), .B2(n6173), .A(n6905), .ZN(n3013) );
  OAI222_X1 U2819 ( .A1(n4751), .A2(n6123), .B1(n2749), .B2(n6119), .C1(n2155), 
        .C2(n6118), .ZN(n6926) );
  INV_X1 U2820 ( .A(n2187), .ZN(n7584) );
  AOI22_X1 U2821 ( .A1(n6129), .A2(n2877), .B1(n6126), .B2(n7584), .ZN(n6909)
         );
  OAI221_X1 U2822 ( .B1(n2091), .B2(n6133), .C1(n2123), .C2(n6132), .A(n6909), 
        .ZN(n6925) );
  AOI22_X1 U2823 ( .A1(n6140), .A2(n5003), .B1(n6137), .B2(n4943), .ZN(n6912)
         );
  OAI221_X1 U2824 ( .B1(n6374), .B2(n6144), .C1(n3677), .C2(n6143), .A(n6912), 
        .ZN(n6924) );
  AOI22_X1 U2825 ( .A1(n2941), .A2(n6151), .B1(n7532), .B2(n6148), .ZN(n6914)
         );
  OAI221_X1 U2826 ( .B1(n4815), .B2(n6157), .C1(n7534), .C2(n6154), .A(n6914), 
        .ZN(n6918) );
  NAND2_X1 U2827 ( .A1(n6158), .A2(n7531), .ZN(n6915) );
  NAND4_X1 U2828 ( .A1(n1438), .A2(n1439), .A3(n1437), .A4(n6915), .ZN(n6917)
         );
  OAI21_X1 U2829 ( .B1(n6918), .B2(n6917), .A(n6162), .ZN(n6921) );
  AOI22_X1 U2830 ( .A1(n6169), .A2(n7526), .B1(n6166), .B2(n7540), .ZN(n6920)
         );
  OAI211_X1 U2831 ( .C1(n2251), .C2(n6172), .A(n6921), .B(n6920), .ZN(n6923)
         );
  NOR4_X1 U2832 ( .A1(n6926), .A2(n6925), .A3(n6924), .A4(n6923), .ZN(n6927)
         );
  OAI21_X1 U2833 ( .B1(n2653), .B2(n6174), .A(n6927), .ZN(n3014) );
  NAND2_X1 U2834 ( .A1(RD2), .A2(n4657), .ZN(n6929) );
  INV_X1 U2835 ( .A(n6929), .ZN(n7552) );
  NAND2_X1 U2836 ( .A1(n1412), .A2(n4617), .ZN(n7522) );
  NAND2_X1 U2837 ( .A1(n4615), .A2(n1413), .ZN(n7520) );
  NAND2_X1 U2838 ( .A1(n4615), .A2(n4608), .ZN(n7519) );
  OAI222_X1 U2839 ( .A1(n939), .A2(n6190), .B1(n2124), .B2(n6187), .C1(n938), 
        .C2(n6186), .ZN(n6948) );
  NAND3_X1 U2840 ( .A1(n1406), .A2(n1412), .A3(n6237), .ZN(n7525) );
  NAND2_X1 U2841 ( .A1(n1412), .A2(n4615), .ZN(n7524) );
  AOI22_X1 U2842 ( .A1(n6196), .A2(n5068), .B1(n6193), .B2(n7553), .ZN(n6932)
         );
  OAI221_X1 U2843 ( .B1(n6202), .B2(n4695), .C1(n2718), .C2(n6199), .A(n6932), 
        .ZN(n6947) );
  NAND2_X1 U2844 ( .A1(n1413), .A2(n4617), .ZN(n7529) );
  NAND2_X1 U2845 ( .A1(n1394), .A2(n4615), .ZN(n7528) );
  AOI22_X1 U2846 ( .A1(n6208), .A2(n5100), .B1(n6205), .B2(n4971), .ZN(n6933)
         );
  OAI221_X1 U2847 ( .B1(n2188), .B2(n6214), .C1(n2060), .C2(n6211), .A(n6933), 
        .ZN(n6946) );
  NAND4_X1 U2848 ( .A1(n1399), .A2(n1397), .A3(n6238), .A4(n1398), .ZN(n7544)
         );
  AOI22_X1 U2849 ( .A1(n2910), .A2(n6223), .B1(n6934), .B2(n6220), .ZN(n6935)
         );
  OAI221_X1 U2850 ( .B1(n6229), .B2(n4813), .C1(n6228), .C2(n6936), .A(n6935), 
        .ZN(n6941) );
  NAND2_X1 U2851 ( .A1(n6217), .A2(n6938), .ZN(n6939) );
  NAND4_X1 U2852 ( .A1(n825), .A2(n826), .A3(n824), .A4(n6939), .ZN(n6940) );
  OAI21_X1 U2853 ( .B1(n6941), .B2(n6940), .A(n6236), .ZN(n6944) );
  NAND3_X1 U2854 ( .A1(n1413), .A2(n1393), .A3(n6236), .ZN(n7545) );
  INV_X1 U2855 ( .A(n7545), .ZN(n7511) );
  AOI22_X1 U2856 ( .A1(n4896), .A2(n6942), .B1(n6181), .B2(n4911), .ZN(n6943)
         );
  OAI211_X1 U2857 ( .C1(n7544), .C2(n6340), .A(n6944), .B(n6943), .ZN(n6945)
         );
  NOR4_X1 U2858 ( .A1(n6948), .A2(n6947), .A3(n6946), .A4(n6945), .ZN(n6949)
         );
  OAI21_X1 U2859 ( .B1(n2685), .B2(n6238), .A(n6949), .ZN(n3046) );
  OAI222_X1 U2860 ( .A1(n956), .A2(n6190), .B1(n2125), .B2(n6187), .C1(n955), 
        .C2(n6186), .ZN(n6966) );
  AOI22_X1 U2861 ( .A1(n6196), .A2(n5067), .B1(n6193), .B2(n7554), .ZN(n6950)
         );
  OAI221_X1 U2862 ( .B1(n6202), .B2(n4694), .C1(n2719), .C2(n6199), .A(n6950), 
        .ZN(n6965) );
  AOI22_X1 U2863 ( .A1(n6208), .A2(n5099), .B1(n6205), .B2(n6951), .ZN(n6952)
         );
  OAI221_X1 U2864 ( .B1(n2189), .B2(n6214), .C1(n2061), .C2(n6211), .A(n6952), 
        .ZN(n6964) );
  AOI22_X1 U2865 ( .A1(n2911), .A2(n6223), .B1(n6953), .B2(n6220), .ZN(n6954)
         );
  OAI221_X1 U2866 ( .B1(n6229), .B2(n4811), .C1(n6228), .C2(n6955), .A(n6954), 
        .ZN(n6960) );
  NAND2_X1 U2867 ( .A1(n6217), .A2(n6957), .ZN(n6958) );
  NAND4_X1 U2868 ( .A1(n872), .A2(n873), .A3(n871), .A4(n6958), .ZN(n6959) );
  OAI21_X1 U2869 ( .B1(n6960), .B2(n6959), .A(n6236), .ZN(n6962) );
  INV_X1 U2870 ( .A(n7544), .ZN(n7510) );
  AOI22_X1 U2871 ( .A1(n6181), .A2(n5002), .B1(DATAIN[1]), .B2(n6176), .ZN(
        n6961) );
  OAI211_X1 U2872 ( .C1(n2253), .C2(n6182), .A(n6962), .B(n6961), .ZN(n6963)
         );
  NOR4_X1 U2873 ( .A1(n6966), .A2(n6965), .A3(n6964), .A4(n6963), .ZN(n6967)
         );
  OAI21_X1 U2874 ( .B1(n2684), .B2(n6240), .A(n6967), .ZN(n3045) );
  OAI222_X1 U2875 ( .A1(n972), .A2(n6190), .B1(n2126), .B2(n6187), .C1(n971), 
        .C2(n6186), .ZN(n6984) );
  AOI22_X1 U2876 ( .A1(n6196), .A2(n5066), .B1(n6193), .B2(n7555), .ZN(n6968)
         );
  OAI221_X1 U2877 ( .B1(n6202), .B2(n4693), .C1(n2720), .C2(n6199), .A(n6968), 
        .ZN(n6983) );
  AOI22_X1 U2878 ( .A1(n6208), .A2(n5098), .B1(n6205), .B2(n6969), .ZN(n6970)
         );
  OAI221_X1 U2879 ( .B1(n2190), .B2(n6214), .C1(n2062), .C2(n6211), .A(n6970), 
        .ZN(n6982) );
  AOI22_X1 U2880 ( .A1(n2912), .A2(n6223), .B1(n6971), .B2(n6220), .ZN(n6972)
         );
  OAI221_X1 U2881 ( .B1(n6229), .B2(n4809), .C1(n6228), .C2(n6973), .A(n6972), 
        .ZN(n6978) );
  NAND2_X1 U2882 ( .A1(n6217), .A2(n6975), .ZN(n6976) );
  NAND4_X1 U2883 ( .A1(n889), .A2(n890), .A3(n888), .A4(n6976), .ZN(n6977) );
  OAI21_X1 U2884 ( .B1(n6978), .B2(n6977), .A(n6236), .ZN(n6980) );
  AOI22_X1 U2885 ( .A1(n6181), .A2(n5001), .B1(DATAIN[2]), .B2(n6176), .ZN(
        n6979) );
  OAI211_X1 U2886 ( .C1(n2254), .C2(n6182), .A(n6980), .B(n6979), .ZN(n6981)
         );
  NOR4_X1 U2887 ( .A1(n6984), .A2(n6983), .A3(n6982), .A4(n6981), .ZN(n6985)
         );
  OAI21_X1 U2888 ( .B1(n2683), .B2(n6240), .A(n6985), .ZN(n3044) );
  OAI222_X1 U2889 ( .A1(n988), .A2(n6190), .B1(n2127), .B2(n6187), .C1(n987), 
        .C2(n6186), .ZN(n7002) );
  AOI22_X1 U2890 ( .A1(n6196), .A2(n5065), .B1(n6193), .B2(n7556), .ZN(n6986)
         );
  OAI221_X1 U2891 ( .B1(n6202), .B2(n4692), .C1(n2721), .C2(n6199), .A(n6986), 
        .ZN(n7001) );
  AOI22_X1 U2892 ( .A1(n6208), .A2(n5097), .B1(n6205), .B2(n6987), .ZN(n6988)
         );
  OAI221_X1 U2893 ( .B1(n2191), .B2(n6214), .C1(n2063), .C2(n6211), .A(n6988), 
        .ZN(n7000) );
  AOI22_X1 U2894 ( .A1(n2913), .A2(n6223), .B1(n6989), .B2(n6220), .ZN(n6990)
         );
  OAI221_X1 U2895 ( .B1(n6229), .B2(n4807), .C1(n6228), .C2(n6991), .A(n6990), 
        .ZN(n6996) );
  NAND2_X1 U2896 ( .A1(n6217), .A2(n6993), .ZN(n6994) );
  NAND4_X1 U2897 ( .A1(n906), .A2(n907), .A3(n905), .A4(n6994), .ZN(n6995) );
  OAI21_X1 U2898 ( .B1(n6996), .B2(n6995), .A(n6236), .ZN(n6998) );
  AOI22_X1 U2899 ( .A1(n6181), .A2(n5000), .B1(DATAIN[3]), .B2(n6176), .ZN(
        n6997) );
  OAI211_X1 U2900 ( .C1(n2255), .C2(n6182), .A(n6998), .B(n6997), .ZN(n6999)
         );
  NOR4_X1 U2901 ( .A1(n7002), .A2(n7001), .A3(n7000), .A4(n6999), .ZN(n7003)
         );
  OAI21_X1 U2902 ( .B1(n2682), .B2(n6240), .A(n7003), .ZN(n3043) );
  OAI222_X1 U2903 ( .A1(n6190), .A2(n4699), .B1(n2128), .B2(n6187), .C1(n6186), 
        .C2(n4691), .ZN(n7021) );
  AOI22_X1 U2904 ( .A1(n6196), .A2(n5064), .B1(n6193), .B2(n7557), .ZN(n7005)
         );
  OAI221_X1 U2905 ( .B1(n2690), .B2(n6202), .C1(n2722), .C2(n6199), .A(n7005), 
        .ZN(n7020) );
  AOI22_X1 U2906 ( .A1(n6208), .A2(n5096), .B1(n6205), .B2(n7006), .ZN(n7007)
         );
  OAI221_X1 U2907 ( .B1(n2192), .B2(n6214), .C1(n2064), .C2(n6211), .A(n7007), 
        .ZN(n7019) );
  AOI22_X1 U2908 ( .A1(n2914), .A2(n6223), .B1(n7008), .B2(n6220), .ZN(n7009)
         );
  OAI221_X1 U2909 ( .B1(n6229), .B2(n4805), .C1(n6228), .C2(n7010), .A(n7009), 
        .ZN(n7015) );
  NAND2_X1 U2910 ( .A1(n6217), .A2(n7012), .ZN(n7013) );
  NAND4_X1 U2911 ( .A1(n923), .A2(n924), .A3(n922), .A4(n7013), .ZN(n7014) );
  OAI21_X1 U2912 ( .B1(n7015), .B2(n7014), .A(n6236), .ZN(n7017) );
  AOI22_X1 U2913 ( .A1(n6181), .A2(n4999), .B1(DATAIN[4]), .B2(n6176), .ZN(
        n7016) );
  OAI211_X1 U2914 ( .C1(n2256), .C2(n6182), .A(n7017), .B(n7016), .ZN(n7018)
         );
  NOR4_X1 U2915 ( .A1(n7021), .A2(n7020), .A3(n7019), .A4(n7018), .ZN(n7022)
         );
  OAI21_X1 U2916 ( .B1(n2681), .B2(n6240), .A(n7022), .ZN(n3042) );
  OAI222_X1 U2917 ( .A1(n6190), .A2(n4697), .B1(n2129), .B2(n6187), .C1(n6186), 
        .C2(n4690), .ZN(n7040) );
  AOI22_X1 U2918 ( .A1(n6196), .A2(n5063), .B1(n6193), .B2(n7558), .ZN(n7024)
         );
  OAI221_X1 U2919 ( .B1(n2691), .B2(n6202), .C1(n2723), .C2(n6199), .A(n7024), 
        .ZN(n7039) );
  AOI22_X1 U2920 ( .A1(n6208), .A2(n5095), .B1(n6205), .B2(n7025), .ZN(n7026)
         );
  OAI221_X1 U2921 ( .B1(n2193), .B2(n6214), .C1(n2065), .C2(n6211), .A(n7026), 
        .ZN(n7038) );
  AOI22_X1 U2922 ( .A1(n2915), .A2(n6223), .B1(n7027), .B2(n6220), .ZN(n7028)
         );
  OAI221_X1 U2923 ( .B1(n6229), .B2(n4803), .C1(n6228), .C2(n7029), .A(n7028), 
        .ZN(n7034) );
  NAND2_X1 U2924 ( .A1(n6217), .A2(n7031), .ZN(n7032) );
  NAND4_X1 U2925 ( .A1(n942), .A2(n943), .A3(n941), .A4(n7032), .ZN(n7033) );
  OAI21_X1 U2926 ( .B1(n7034), .B2(n7033), .A(n6236), .ZN(n7036) );
  AOI22_X1 U2927 ( .A1(n6181), .A2(n4998), .B1(DATAIN[5]), .B2(n6176), .ZN(
        n7035) );
  OAI211_X1 U2928 ( .C1(n2257), .C2(n6182), .A(n7036), .B(n7035), .ZN(n7037)
         );
  NOR4_X1 U2929 ( .A1(n7040), .A2(n7039), .A3(n7038), .A4(n7037), .ZN(n7041)
         );
  OAI21_X1 U2930 ( .B1(n2680), .B2(n6240), .A(n7041), .ZN(n3041) );
  OAI222_X1 U2931 ( .A1(n6190), .A2(n4705), .B1(n2130), .B2(n6187), .C1(n6186), 
        .C2(n4689), .ZN(n7059) );
  AOI22_X1 U2932 ( .A1(n6196), .A2(n5062), .B1(n6193), .B2(n7559), .ZN(n7043)
         );
  OAI221_X1 U2933 ( .B1(n2692), .B2(n6202), .C1(n2724), .C2(n6199), .A(n7043), 
        .ZN(n7058) );
  AOI22_X1 U2934 ( .A1(n6208), .A2(n5094), .B1(n6205), .B2(n7044), .ZN(n7045)
         );
  OAI221_X1 U2935 ( .B1(n2194), .B2(n6214), .C1(n2066), .C2(n6211), .A(n7045), 
        .ZN(n7057) );
  AOI22_X1 U2936 ( .A1(n2916), .A2(n6223), .B1(n7046), .B2(n6220), .ZN(n7047)
         );
  OAI221_X1 U2937 ( .B1(n6229), .B2(n4801), .C1(n6228), .C2(n7048), .A(n7047), 
        .ZN(n7053) );
  NAND2_X1 U2938 ( .A1(n6217), .A2(n7050), .ZN(n7051) );
  NAND4_X1 U2939 ( .A1(n962), .A2(n963), .A3(n961), .A4(n7051), .ZN(n7052) );
  OAI21_X1 U2940 ( .B1(n7053), .B2(n7052), .A(n6236), .ZN(n7055) );
  AOI22_X1 U2941 ( .A1(n6181), .A2(n4997), .B1(DATAIN[6]), .B2(n6176), .ZN(
        n7054) );
  OAI211_X1 U2942 ( .C1(n2258), .C2(n6182), .A(n7055), .B(n7054), .ZN(n7056)
         );
  NOR4_X1 U2943 ( .A1(n7059), .A2(n7058), .A3(n7057), .A4(n7056), .ZN(n7060)
         );
  OAI21_X1 U2944 ( .B1(n2679), .B2(n6240), .A(n7060), .ZN(n3040) );
  OAI222_X1 U2945 ( .A1(n6190), .A2(n4703), .B1(n2131), .B2(n6187), .C1(n6186), 
        .C2(n4688), .ZN(n7078) );
  AOI22_X1 U2946 ( .A1(n6196), .A2(n5061), .B1(n6193), .B2(n7560), .ZN(n7062)
         );
  OAI221_X1 U2947 ( .B1(n2693), .B2(n6202), .C1(n2725), .C2(n6199), .A(n7062), 
        .ZN(n7077) );
  AOI22_X1 U2948 ( .A1(n6208), .A2(n5093), .B1(n6205), .B2(n7063), .ZN(n7064)
         );
  OAI221_X1 U2949 ( .B1(n2195), .B2(n6214), .C1(n2067), .C2(n6211), .A(n7064), 
        .ZN(n7076) );
  AOI22_X1 U2950 ( .A1(n2917), .A2(n6223), .B1(n7065), .B2(n6220), .ZN(n7066)
         );
  OAI221_X1 U2951 ( .B1(n6229), .B2(n4799), .C1(n6228), .C2(n7067), .A(n7066), 
        .ZN(n7072) );
  NAND2_X1 U2952 ( .A1(n6217), .A2(n7069), .ZN(n7070) );
  NAND4_X1 U2953 ( .A1(n983), .A2(n984), .A3(n981), .A4(n7070), .ZN(n7071) );
  OAI21_X1 U2954 ( .B1(n7072), .B2(n7071), .A(n6236), .ZN(n7074) );
  AOI22_X1 U2955 ( .A1(n6180), .A2(n4996), .B1(DATAIN[7]), .B2(n6176), .ZN(
        n7073) );
  OAI211_X1 U2956 ( .C1(n2259), .C2(n6182), .A(n7074), .B(n7073), .ZN(n7075)
         );
  NOR4_X1 U2957 ( .A1(n7078), .A2(n7077), .A3(n7076), .A4(n7075), .ZN(n7079)
         );
  OAI21_X1 U2958 ( .B1(n2678), .B2(n6240), .A(n7079), .ZN(n3039) );
  OAI222_X1 U2959 ( .A1(n6190), .A2(n4701), .B1(n2132), .B2(n6187), .C1(n6185), 
        .C2(n4687), .ZN(n7097) );
  AOI22_X1 U2960 ( .A1(n6196), .A2(n5060), .B1(n6193), .B2(n7561), .ZN(n7081)
         );
  OAI221_X1 U2961 ( .B1(n2694), .B2(n6202), .C1(n2726), .C2(n6199), .A(n7081), 
        .ZN(n7096) );
  AOI22_X1 U2962 ( .A1(n6208), .A2(n5092), .B1(n6205), .B2(n7082), .ZN(n7083)
         );
  OAI221_X1 U2963 ( .B1(n2196), .B2(n6214), .C1(n2068), .C2(n6211), .A(n7083), 
        .ZN(n7095) );
  AOI22_X1 U2964 ( .A1(n2918), .A2(n6223), .B1(n7084), .B2(n6220), .ZN(n7085)
         );
  OAI221_X1 U2965 ( .B1(n6229), .B2(n4797), .C1(n6227), .C2(n7086), .A(n7085), 
        .ZN(n7091) );
  NAND2_X1 U2966 ( .A1(n6217), .A2(n7088), .ZN(n7089) );
  NAND4_X1 U2967 ( .A1(n1003), .A2(n1004), .A3(n1002), .A4(n7089), .ZN(n7090)
         );
  OAI21_X1 U2968 ( .B1(n7091), .B2(n7090), .A(n6235), .ZN(n7093) );
  AOI22_X1 U2969 ( .A1(n6180), .A2(n4995), .B1(DATAIN[8]), .B2(n6176), .ZN(
        n7092) );
  OAI211_X1 U2970 ( .C1(n2260), .C2(n6182), .A(n7093), .B(n7092), .ZN(n7094)
         );
  NOR4_X1 U2971 ( .A1(n7097), .A2(n7096), .A3(n7095), .A4(n7094), .ZN(n7098)
         );
  OAI21_X1 U2972 ( .B1(n2677), .B2(n6240), .A(n7098), .ZN(n3038) );
  OAI222_X1 U2973 ( .A1(n6190), .A2(n4711), .B1(n2133), .B2(n6187), .C1(n6185), 
        .C2(n4686), .ZN(n7116) );
  AOI22_X1 U2974 ( .A1(n6196), .A2(n5059), .B1(n6193), .B2(n7562), .ZN(n7100)
         );
  OAI221_X1 U2975 ( .B1(n2695), .B2(n6202), .C1(n2727), .C2(n6199), .A(n7100), 
        .ZN(n7115) );
  AOI22_X1 U2976 ( .A1(n6208), .A2(n5091), .B1(n6205), .B2(n7101), .ZN(n7102)
         );
  OAI221_X1 U2977 ( .B1(n2197), .B2(n6214), .C1(n2069), .C2(n6211), .A(n7102), 
        .ZN(n7114) );
  AOI22_X1 U2978 ( .A1(n2919), .A2(n6223), .B1(n7103), .B2(n6220), .ZN(n7104)
         );
  OAI221_X1 U2979 ( .B1(n6229), .B2(n4795), .C1(n6227), .C2(n7105), .A(n7104), 
        .ZN(n7110) );
  NAND2_X1 U2980 ( .A1(n6217), .A2(n7107), .ZN(n7108) );
  NAND4_X1 U2981 ( .A1(n1020), .A2(n1021), .A3(n1019), .A4(n7108), .ZN(n7109)
         );
  OAI21_X1 U2982 ( .B1(n7110), .B2(n7109), .A(n6235), .ZN(n7112) );
  AOI22_X1 U2983 ( .A1(n6180), .A2(n4994), .B1(DATAIN[9]), .B2(n6176), .ZN(
        n7111) );
  OAI211_X1 U2984 ( .C1(n2261), .C2(n6182), .A(n7112), .B(n7111), .ZN(n7113)
         );
  NOR4_X1 U2985 ( .A1(n7116), .A2(n7115), .A3(n7114), .A4(n7113), .ZN(n7117)
         );
  OAI21_X1 U2986 ( .B1(n2676), .B2(n6240), .A(n7117), .ZN(n3037) );
  OAI222_X1 U2987 ( .A1(n6190), .A2(n4709), .B1(n2134), .B2(n6187), .C1(n6185), 
        .C2(n4685), .ZN(n7135) );
  AOI22_X1 U2988 ( .A1(n6196), .A2(n5058), .B1(n6193), .B2(n7563), .ZN(n7119)
         );
  OAI221_X1 U2989 ( .B1(n2696), .B2(n6202), .C1(n2728), .C2(n6199), .A(n7119), 
        .ZN(n7134) );
  AOI22_X1 U2990 ( .A1(n6208), .A2(n5090), .B1(n6205), .B2(n7120), .ZN(n7121)
         );
  OAI221_X1 U2991 ( .B1(n2198), .B2(n6214), .C1(n2070), .C2(n6211), .A(n7121), 
        .ZN(n7133) );
  AOI22_X1 U2992 ( .A1(n2920), .A2(n6223), .B1(n7122), .B2(n6220), .ZN(n7123)
         );
  OAI221_X1 U2993 ( .B1(n6229), .B2(n4793), .C1(n6227), .C2(n7124), .A(n7123), 
        .ZN(n7129) );
  NAND2_X1 U2994 ( .A1(n6217), .A2(n7126), .ZN(n7127) );
  NAND4_X1 U2995 ( .A1(n1037), .A2(n1038), .A3(n1036), .A4(n7127), .ZN(n7128)
         );
  OAI21_X1 U2996 ( .B1(n7129), .B2(n7128), .A(n6235), .ZN(n7131) );
  AOI22_X1 U2997 ( .A1(n6180), .A2(n4993), .B1(DATAIN[10]), .B2(n6176), .ZN(
        n7130) );
  OAI211_X1 U2998 ( .C1(n2262), .C2(n6182), .A(n7131), .B(n7130), .ZN(n7132)
         );
  NOR4_X1 U2999 ( .A1(n7135), .A2(n7134), .A3(n7133), .A4(n7132), .ZN(n7136)
         );
  OAI21_X1 U3000 ( .B1(n2675), .B2(n6239), .A(n7136), .ZN(n3036) );
  OAI222_X1 U3001 ( .A1(n6190), .A2(n4707), .B1(n2135), .B2(n6187), .C1(n6185), 
        .C2(n4684), .ZN(n7154) );
  AOI22_X1 U3002 ( .A1(n6196), .A2(n5057), .B1(n6193), .B2(n7564), .ZN(n7138)
         );
  OAI221_X1 U3003 ( .B1(n2697), .B2(n6202), .C1(n2729), .C2(n6199), .A(n7138), 
        .ZN(n7153) );
  AOI22_X1 U3004 ( .A1(n6208), .A2(n5089), .B1(n6205), .B2(n7139), .ZN(n7140)
         );
  OAI221_X1 U3005 ( .B1(n2199), .B2(n6214), .C1(n2071), .C2(n6211), .A(n7140), 
        .ZN(n7152) );
  AOI22_X1 U3006 ( .A1(n2921), .A2(n6223), .B1(n7141), .B2(n6220), .ZN(n7142)
         );
  OAI221_X1 U3007 ( .B1(n6229), .B2(n4791), .C1(n6227), .C2(n7143), .A(n7142), 
        .ZN(n7148) );
  NAND2_X1 U3008 ( .A1(n6217), .A2(n7145), .ZN(n7146) );
  NAND4_X1 U3009 ( .A1(n1054), .A2(n1055), .A3(n1053), .A4(n7146), .ZN(n7147)
         );
  OAI21_X1 U3010 ( .B1(n7148), .B2(n7147), .A(n6235), .ZN(n7150) );
  AOI22_X1 U3011 ( .A1(n6180), .A2(n4992), .B1(DATAIN[11]), .B2(n6176), .ZN(
        n7149) );
  OAI211_X1 U3012 ( .C1(n2263), .C2(n6182), .A(n7150), .B(n7149), .ZN(n7151)
         );
  NOR4_X1 U3013 ( .A1(n7154), .A2(n7153), .A3(n7152), .A4(n7151), .ZN(n7155)
         );
  OAI21_X1 U3014 ( .B1(n2674), .B2(n6239), .A(n7155), .ZN(n3035) );
  OAI222_X1 U3015 ( .A1(n6191), .A2(n4717), .B1(n2136), .B2(n6188), .C1(n6185), 
        .C2(n4683), .ZN(n7173) );
  AOI22_X1 U3016 ( .A1(n6197), .A2(n5056), .B1(n6194), .B2(n7565), .ZN(n7157)
         );
  OAI221_X1 U3017 ( .B1(n2698), .B2(n6203), .C1(n2730), .C2(n6200), .A(n7157), 
        .ZN(n7172) );
  AOI22_X1 U3018 ( .A1(n6209), .A2(n5088), .B1(n6206), .B2(n7158), .ZN(n7159)
         );
  OAI221_X1 U3019 ( .B1(n2200), .B2(n6215), .C1(n2072), .C2(n6212), .A(n7159), 
        .ZN(n7171) );
  AOI22_X1 U3020 ( .A1(n2922), .A2(n6224), .B1(n7160), .B2(n6221), .ZN(n7161)
         );
  OAI221_X1 U3021 ( .B1(n6230), .B2(n4789), .C1(n6227), .C2(n7162), .A(n7161), 
        .ZN(n7167) );
  NAND2_X1 U3022 ( .A1(n6218), .A2(n7164), .ZN(n7165) );
  NAND4_X1 U3023 ( .A1(n1071), .A2(n1072), .A3(n1070), .A4(n7165), .ZN(n7166)
         );
  OAI21_X1 U3024 ( .B1(n7167), .B2(n7166), .A(n6235), .ZN(n7169) );
  AOI22_X1 U3025 ( .A1(n6180), .A2(n4991), .B1(DATAIN[12]), .B2(n6176), .ZN(
        n7168) );
  OAI211_X1 U3026 ( .C1(n2264), .C2(n6182), .A(n7169), .B(n7168), .ZN(n7170)
         );
  NOR4_X1 U3027 ( .A1(n7173), .A2(n7172), .A3(n7171), .A4(n7170), .ZN(n7174)
         );
  OAI21_X1 U3028 ( .B1(n2673), .B2(n6239), .A(n7174), .ZN(n3034) );
  OAI222_X1 U3029 ( .A1(n6191), .A2(n4715), .B1(n2137), .B2(n6188), .C1(n6185), 
        .C2(n4682), .ZN(n7192) );
  AOI22_X1 U3030 ( .A1(n6197), .A2(n5055), .B1(n6194), .B2(n7566), .ZN(n7176)
         );
  OAI221_X1 U3031 ( .B1(n2699), .B2(n6203), .C1(n2731), .C2(n6200), .A(n7176), 
        .ZN(n7191) );
  AOI22_X1 U3032 ( .A1(n6209), .A2(n5087), .B1(n6206), .B2(n7177), .ZN(n7178)
         );
  OAI221_X1 U3033 ( .B1(n2201), .B2(n6215), .C1(n2073), .C2(n6212), .A(n7178), 
        .ZN(n7190) );
  AOI22_X1 U3034 ( .A1(n2923), .A2(n6224), .B1(n7179), .B2(n6221), .ZN(n7180)
         );
  OAI221_X1 U3035 ( .B1(n6230), .B2(n4787), .C1(n6227), .C2(n7181), .A(n7180), 
        .ZN(n7186) );
  NAND2_X1 U3036 ( .A1(n6218), .A2(n7183), .ZN(n7184) );
  NAND4_X1 U3037 ( .A1(n1088), .A2(n1089), .A3(n1087), .A4(n7184), .ZN(n7185)
         );
  OAI21_X1 U3038 ( .B1(n7186), .B2(n7185), .A(n6235), .ZN(n7188) );
  AOI22_X1 U3039 ( .A1(n6180), .A2(n4990), .B1(DATAIN[13]), .B2(n6177), .ZN(
        n7187) );
  OAI211_X1 U3040 ( .C1(n2265), .C2(n6183), .A(n7188), .B(n7187), .ZN(n7189)
         );
  NOR4_X1 U3041 ( .A1(n7192), .A2(n7191), .A3(n7190), .A4(n7189), .ZN(n7193)
         );
  OAI21_X1 U3042 ( .B1(n2672), .B2(n6239), .A(n7193), .ZN(n3033) );
  OAI222_X1 U3043 ( .A1(n6191), .A2(n4713), .B1(n2138), .B2(n6188), .C1(n6185), 
        .C2(n4681), .ZN(n7211) );
  AOI22_X1 U3044 ( .A1(n6197), .A2(n5054), .B1(n6194), .B2(n7567), .ZN(n7195)
         );
  OAI221_X1 U3045 ( .B1(n2700), .B2(n6203), .C1(n2732), .C2(n6200), .A(n7195), 
        .ZN(n7210) );
  AOI22_X1 U3046 ( .A1(n6209), .A2(n5086), .B1(n6206), .B2(n7196), .ZN(n7197)
         );
  OAI221_X1 U3047 ( .B1(n2202), .B2(n6215), .C1(n2074), .C2(n6212), .A(n7197), 
        .ZN(n7209) );
  AOI22_X1 U3048 ( .A1(n2924), .A2(n6224), .B1(n7198), .B2(n6221), .ZN(n7199)
         );
  OAI221_X1 U3049 ( .B1(n6230), .B2(n4785), .C1(n6227), .C2(n7200), .A(n7199), 
        .ZN(n7205) );
  NAND2_X1 U3050 ( .A1(n6218), .A2(n7202), .ZN(n7203) );
  NAND4_X1 U3051 ( .A1(n1105), .A2(n1106), .A3(n1104), .A4(n7203), .ZN(n7204)
         );
  OAI21_X1 U3052 ( .B1(n7205), .B2(n7204), .A(n6235), .ZN(n7207) );
  AOI22_X1 U3053 ( .A1(n6180), .A2(n4989), .B1(DATAIN[14]), .B2(n6177), .ZN(
        n7206) );
  OAI211_X1 U3054 ( .C1(n2266), .C2(n6183), .A(n7207), .B(n7206), .ZN(n7208)
         );
  NOR4_X1 U3055 ( .A1(n7211), .A2(n7210), .A3(n7209), .A4(n7208), .ZN(n7212)
         );
  OAI21_X1 U3056 ( .B1(n2671), .B2(n6239), .A(n7212), .ZN(n3032) );
  OAI222_X1 U3057 ( .A1(n6191), .A2(n4723), .B1(n2139), .B2(n6188), .C1(n6185), 
        .C2(n4680), .ZN(n7230) );
  AOI22_X1 U3058 ( .A1(n6197), .A2(n5053), .B1(n6194), .B2(n7568), .ZN(n7214)
         );
  OAI221_X1 U3059 ( .B1(n2701), .B2(n6203), .C1(n2733), .C2(n6200), .A(n7214), 
        .ZN(n7229) );
  AOI22_X1 U3060 ( .A1(n6209), .A2(n5085), .B1(n6206), .B2(n7215), .ZN(n7216)
         );
  OAI221_X1 U3061 ( .B1(n2203), .B2(n6215), .C1(n2075), .C2(n6212), .A(n7216), 
        .ZN(n7228) );
  AOI22_X1 U3062 ( .A1(n2925), .A2(n6224), .B1(n7217), .B2(n6221), .ZN(n7218)
         );
  OAI221_X1 U3063 ( .B1(n6230), .B2(n4783), .C1(n6227), .C2(n7219), .A(n7218), 
        .ZN(n7224) );
  NAND2_X1 U3064 ( .A1(n6218), .A2(n7221), .ZN(n7222) );
  NAND4_X1 U3065 ( .A1(n1122), .A2(n1123), .A3(n1121), .A4(n7222), .ZN(n7223)
         );
  OAI21_X1 U3066 ( .B1(n7224), .B2(n7223), .A(n6235), .ZN(n7226) );
  AOI22_X1 U3067 ( .A1(n6180), .A2(n4988), .B1(DATAIN[15]), .B2(n6177), .ZN(
        n7225) );
  OAI211_X1 U3068 ( .C1(n2267), .C2(n6183), .A(n7226), .B(n7225), .ZN(n7227)
         );
  NOR4_X1 U3069 ( .A1(n7230), .A2(n7229), .A3(n7228), .A4(n7227), .ZN(n7231)
         );
  OAI21_X1 U3070 ( .B1(n2670), .B2(n6239), .A(n7231), .ZN(n3031) );
  OAI222_X1 U3071 ( .A1(n6191), .A2(n4721), .B1(n2140), .B2(n6188), .C1(n6185), 
        .C2(n4679), .ZN(n7249) );
  AOI22_X1 U3072 ( .A1(n6197), .A2(n5052), .B1(n6194), .B2(n7569), .ZN(n7233)
         );
  OAI221_X1 U3073 ( .B1(n2702), .B2(n6203), .C1(n2734), .C2(n6200), .A(n7233), 
        .ZN(n7248) );
  AOI22_X1 U3074 ( .A1(n6209), .A2(n5084), .B1(n6206), .B2(n7234), .ZN(n7235)
         );
  OAI221_X1 U3075 ( .B1(n2204), .B2(n6215), .C1(n2076), .C2(n6212), .A(n7235), 
        .ZN(n7247) );
  AOI22_X1 U3076 ( .A1(n2926), .A2(n6224), .B1(n7236), .B2(n6221), .ZN(n7237)
         );
  OAI221_X1 U3077 ( .B1(n6230), .B2(n4753), .C1(n6227), .C2(n7238), .A(n7237), 
        .ZN(n7243) );
  NAND2_X1 U3078 ( .A1(n6218), .A2(n7240), .ZN(n7241) );
  NAND4_X1 U3079 ( .A1(n1139), .A2(n1140), .A3(n1138), .A4(n7241), .ZN(n7242)
         );
  OAI21_X1 U3080 ( .B1(n7243), .B2(n7242), .A(n6235), .ZN(n7245) );
  AOI22_X1 U3081 ( .A1(n6180), .A2(n4987), .B1(DATAIN[16]), .B2(n6177), .ZN(
        n7244) );
  OAI211_X1 U3082 ( .C1(n2268), .C2(n6183), .A(n7245), .B(n7244), .ZN(n7246)
         );
  NOR4_X1 U3083 ( .A1(n7249), .A2(n7248), .A3(n7247), .A4(n7246), .ZN(n7250)
         );
  OAI21_X1 U3084 ( .B1(n2669), .B2(n6239), .A(n7250), .ZN(n3030) );
  OAI222_X1 U3085 ( .A1(n6191), .A2(n4719), .B1(n2141), .B2(n6188), .C1(n6185), 
        .C2(n4678), .ZN(n7268) );
  AOI22_X1 U3086 ( .A1(n6197), .A2(n5051), .B1(n6194), .B2(n7570), .ZN(n7252)
         );
  OAI221_X1 U3087 ( .B1(n2703), .B2(n6203), .C1(n2735), .C2(n6200), .A(n7252), 
        .ZN(n7267) );
  AOI22_X1 U3088 ( .A1(n6209), .A2(n5083), .B1(n6206), .B2(n7253), .ZN(n7254)
         );
  OAI221_X1 U3089 ( .B1(n2205), .B2(n6215), .C1(n2077), .C2(n6212), .A(n7254), 
        .ZN(n7266) );
  AOI22_X1 U3090 ( .A1(n2927), .A2(n6224), .B1(n7255), .B2(n6221), .ZN(n7256)
         );
  OAI221_X1 U3091 ( .B1(n6230), .B2(n4763), .C1(n6227), .C2(n7257), .A(n7256), 
        .ZN(n7262) );
  NAND2_X1 U3092 ( .A1(n6218), .A2(n7259), .ZN(n7260) );
  NAND4_X1 U3093 ( .A1(n1156), .A2(n1157), .A3(n1155), .A4(n7260), .ZN(n7261)
         );
  OAI21_X1 U3094 ( .B1(n7262), .B2(n7261), .A(n6235), .ZN(n7264) );
  AOI22_X1 U3095 ( .A1(n6180), .A2(n4986), .B1(DATAIN[17]), .B2(n6177), .ZN(
        n7263) );
  OAI211_X1 U3096 ( .C1(n2269), .C2(n6183), .A(n7264), .B(n7263), .ZN(n7265)
         );
  NOR4_X1 U3097 ( .A1(n7268), .A2(n7267), .A3(n7266), .A4(n7265), .ZN(n7269)
         );
  OAI21_X1 U3098 ( .B1(n2668), .B2(n6239), .A(n7269), .ZN(n3029) );
  OAI222_X1 U3099 ( .A1(n6191), .A2(n4729), .B1(n2142), .B2(n6188), .C1(n6185), 
        .C2(n4677), .ZN(n7287) );
  AOI22_X1 U3100 ( .A1(n6197), .A2(n5050), .B1(n6194), .B2(n7571), .ZN(n7271)
         );
  OAI221_X1 U3101 ( .B1(n2704), .B2(n6203), .C1(n2736), .C2(n6200), .A(n7271), 
        .ZN(n7286) );
  AOI22_X1 U3102 ( .A1(n6209), .A2(n5082), .B1(n6206), .B2(n7272), .ZN(n7273)
         );
  OAI221_X1 U3103 ( .B1(n2206), .B2(n6215), .C1(n2078), .C2(n6212), .A(n7273), 
        .ZN(n7285) );
  AOI22_X1 U3104 ( .A1(n2928), .A2(n6224), .B1(n7274), .B2(n6221), .ZN(n7275)
         );
  OAI221_X1 U3105 ( .B1(n6230), .B2(n4757), .C1(n6227), .C2(n7276), .A(n7275), 
        .ZN(n7281) );
  NAND2_X1 U3106 ( .A1(n6218), .A2(n7278), .ZN(n7279) );
  NAND4_X1 U3107 ( .A1(n1173), .A2(n1174), .A3(n1172), .A4(n7279), .ZN(n7280)
         );
  OAI21_X1 U3108 ( .B1(n7281), .B2(n7280), .A(n6235), .ZN(n7283) );
  AOI22_X1 U3109 ( .A1(n6180), .A2(n4985), .B1(DATAIN[18]), .B2(n6177), .ZN(
        n7282) );
  OAI211_X1 U3110 ( .C1(n2270), .C2(n6183), .A(n7283), .B(n7282), .ZN(n7284)
         );
  NOR4_X1 U3111 ( .A1(n7287), .A2(n7286), .A3(n7285), .A4(n7284), .ZN(n7288)
         );
  OAI21_X1 U3112 ( .B1(n2667), .B2(n6239), .A(n7288), .ZN(n3028) );
  OAI222_X1 U3113 ( .A1(n6191), .A2(n4727), .B1(n2143), .B2(n6188), .C1(n6185), 
        .C2(n4676), .ZN(n7306) );
  AOI22_X1 U3114 ( .A1(n6197), .A2(n5049), .B1(n6194), .B2(n7572), .ZN(n7290)
         );
  OAI221_X1 U3115 ( .B1(n2705), .B2(n6203), .C1(n2737), .C2(n6200), .A(n7290), 
        .ZN(n7305) );
  AOI22_X1 U3116 ( .A1(n6209), .A2(n5081), .B1(n6206), .B2(n7291), .ZN(n7292)
         );
  OAI221_X1 U3117 ( .B1(n2207), .B2(n6215), .C1(n2079), .C2(n6212), .A(n7292), 
        .ZN(n7304) );
  AOI22_X1 U3118 ( .A1(n2929), .A2(n6224), .B1(n7293), .B2(n6221), .ZN(n7294)
         );
  OAI221_X1 U3119 ( .B1(n6230), .B2(n4759), .C1(n6227), .C2(n7295), .A(n7294), 
        .ZN(n7300) );
  NAND2_X1 U3120 ( .A1(n6218), .A2(n7297), .ZN(n7298) );
  NAND4_X1 U3121 ( .A1(n1190), .A2(n1191), .A3(n1189), .A4(n7298), .ZN(n7299)
         );
  OAI21_X1 U3122 ( .B1(n7300), .B2(n7299), .A(n6234), .ZN(n7302) );
  AOI22_X1 U3123 ( .A1(n6179), .A2(n4984), .B1(DATAIN[19]), .B2(n6177), .ZN(
        n7301) );
  OAI211_X1 U3124 ( .C1(n2271), .C2(n6183), .A(n7302), .B(n7301), .ZN(n7303)
         );
  NOR4_X1 U3125 ( .A1(n7306), .A2(n7305), .A3(n7304), .A4(n7303), .ZN(n7307)
         );
  OAI21_X1 U3126 ( .B1(n2666), .B2(n6239), .A(n7307), .ZN(n3027) );
  OAI222_X1 U3127 ( .A1(n6191), .A2(n4725), .B1(n2144), .B2(n6188), .C1(n6184), 
        .C2(n4675), .ZN(n7325) );
  AOI22_X1 U3128 ( .A1(n6197), .A2(n5048), .B1(n6194), .B2(n7573), .ZN(n7309)
         );
  OAI221_X1 U3129 ( .B1(n2706), .B2(n6203), .C1(n2738), .C2(n6200), .A(n7309), 
        .ZN(n7324) );
  AOI22_X1 U3130 ( .A1(n6209), .A2(n5080), .B1(n6206), .B2(n7310), .ZN(n7311)
         );
  OAI221_X1 U3131 ( .B1(n2208), .B2(n6215), .C1(n2080), .C2(n6212), .A(n7311), 
        .ZN(n7323) );
  AOI22_X1 U3132 ( .A1(n2930), .A2(n6224), .B1(n7312), .B2(n6221), .ZN(n7313)
         );
  OAI221_X1 U3133 ( .B1(n6230), .B2(n4769), .C1(n6226), .C2(n7314), .A(n7313), 
        .ZN(n7319) );
  NAND2_X1 U3134 ( .A1(n6218), .A2(n7316), .ZN(n7317) );
  NAND4_X1 U3135 ( .A1(n1207), .A2(n1208), .A3(n1206), .A4(n7317), .ZN(n7318)
         );
  OAI21_X1 U3136 ( .B1(n7319), .B2(n7318), .A(n6235), .ZN(n7321) );
  AOI22_X1 U3137 ( .A1(n6179), .A2(n4983), .B1(DATAIN[20]), .B2(n6177), .ZN(
        n7320) );
  OAI211_X1 U3138 ( .C1(n2272), .C2(n6183), .A(n7321), .B(n7320), .ZN(n7322)
         );
  NOR4_X1 U3139 ( .A1(n7325), .A2(n7324), .A3(n7323), .A4(n7322), .ZN(n7326)
         );
  OAI21_X1 U3140 ( .B1(n2665), .B2(n6239), .A(n7326), .ZN(n3026) );
  OAI222_X1 U3141 ( .A1(n6191), .A2(n4735), .B1(n2145), .B2(n6188), .C1(n6184), 
        .C2(n4674), .ZN(n7344) );
  AOI22_X1 U3142 ( .A1(n6197), .A2(n5047), .B1(n6194), .B2(n7574), .ZN(n7328)
         );
  OAI221_X1 U3143 ( .B1(n2707), .B2(n6203), .C1(n2739), .C2(n6200), .A(n7328), 
        .ZN(n7343) );
  AOI22_X1 U3144 ( .A1(n6209), .A2(n5079), .B1(n6206), .B2(n7329), .ZN(n7330)
         );
  OAI221_X1 U3145 ( .B1(n2209), .B2(n6215), .C1(n2081), .C2(n6212), .A(n7330), 
        .ZN(n7342) );
  AOI22_X1 U3146 ( .A1(n2931), .A2(n6224), .B1(n7331), .B2(n6221), .ZN(n7332)
         );
  OAI221_X1 U3147 ( .B1(n6230), .B2(n4761), .C1(n6226), .C2(n7333), .A(n7332), 
        .ZN(n7338) );
  NAND2_X1 U3148 ( .A1(n6218), .A2(n7335), .ZN(n7336) );
  NAND4_X1 U3149 ( .A1(n1224), .A2(n1225), .A3(n1223), .A4(n7336), .ZN(n7337)
         );
  OAI21_X1 U3150 ( .B1(n7338), .B2(n7337), .A(n6234), .ZN(n7340) );
  AOI22_X1 U3151 ( .A1(n6179), .A2(n4982), .B1(DATAIN[21]), .B2(n6177), .ZN(
        n7339) );
  OAI211_X1 U3152 ( .C1(n2273), .C2(n6183), .A(n7340), .B(n7339), .ZN(n7341)
         );
  NOR4_X1 U3153 ( .A1(n7344), .A2(n7343), .A3(n7342), .A4(n7341), .ZN(n7345)
         );
  OAI21_X1 U3154 ( .B1(n2664), .B2(n6238), .A(n7345), .ZN(n3025) );
  OAI222_X1 U3155 ( .A1(n6191), .A2(n4733), .B1(n2146), .B2(n6188), .C1(n6184), 
        .C2(n4673), .ZN(n7363) );
  AOI22_X1 U3156 ( .A1(n6197), .A2(n5046), .B1(n6194), .B2(n7575), .ZN(n7347)
         );
  OAI221_X1 U3157 ( .B1(n2708), .B2(n6203), .C1(n2740), .C2(n6200), .A(n7347), 
        .ZN(n7362) );
  AOI22_X1 U3158 ( .A1(n6209), .A2(n5078), .B1(n6206), .B2(n7348), .ZN(n7349)
         );
  OAI221_X1 U3159 ( .B1(n2210), .B2(n6215), .C1(n2082), .C2(n6212), .A(n7349), 
        .ZN(n7361) );
  AOI22_X1 U3160 ( .A1(n2932), .A2(n6224), .B1(n7350), .B2(n6221), .ZN(n7351)
         );
  OAI221_X1 U3161 ( .B1(n6230), .B2(n4765), .C1(n6226), .C2(n7352), .A(n7351), 
        .ZN(n7357) );
  NAND2_X1 U3162 ( .A1(n6218), .A2(n7354), .ZN(n7355) );
  NAND4_X1 U3163 ( .A1(n1241), .A2(n1242), .A3(n1240), .A4(n7355), .ZN(n7356)
         );
  OAI21_X1 U3164 ( .B1(n7357), .B2(n7356), .A(n6234), .ZN(n7359) );
  AOI22_X1 U3165 ( .A1(n6179), .A2(n4981), .B1(DATAIN[22]), .B2(n6177), .ZN(
        n7358) );
  OAI211_X1 U3166 ( .C1(n2274), .C2(n6183), .A(n7359), .B(n7358), .ZN(n7360)
         );
  NOR4_X1 U3167 ( .A1(n7363), .A2(n7362), .A3(n7361), .A4(n7360), .ZN(n7364)
         );
  OAI21_X1 U3168 ( .B1(n2663), .B2(n6238), .A(n7364), .ZN(n3024) );
  OAI222_X1 U3169 ( .A1(n6191), .A2(n4731), .B1(n2147), .B2(n6188), .C1(n6184), 
        .C2(n4672), .ZN(n7382) );
  AOI22_X1 U3170 ( .A1(n6197), .A2(n5045), .B1(n6194), .B2(n7576), .ZN(n7366)
         );
  OAI221_X1 U3171 ( .B1(n2709), .B2(n6203), .C1(n2741), .C2(n6200), .A(n7366), 
        .ZN(n7381) );
  AOI22_X1 U3172 ( .A1(n6209), .A2(n5077), .B1(n6206), .B2(n7367), .ZN(n7368)
         );
  OAI221_X1 U3173 ( .B1(n2211), .B2(n6215), .C1(n2083), .C2(n6212), .A(n7368), 
        .ZN(n7380) );
  AOI22_X1 U3174 ( .A1(n2933), .A2(n6224), .B1(n7369), .B2(n6221), .ZN(n7370)
         );
  OAI221_X1 U3175 ( .B1(n6230), .B2(n4771), .C1(n6226), .C2(n7371), .A(n7370), 
        .ZN(n7376) );
  NAND2_X1 U3176 ( .A1(n6218), .A2(n7373), .ZN(n7374) );
  NAND4_X1 U3177 ( .A1(n1258), .A2(n1259), .A3(n1257), .A4(n7374), .ZN(n7375)
         );
  OAI21_X1 U3178 ( .B1(n7376), .B2(n7375), .A(n6234), .ZN(n7378) );
  AOI22_X1 U3179 ( .A1(n6179), .A2(n4980), .B1(DATAIN[23]), .B2(n6177), .ZN(
        n7377) );
  OAI211_X1 U3180 ( .C1(n2275), .C2(n6183), .A(n7378), .B(n7377), .ZN(n7379)
         );
  NOR4_X1 U3181 ( .A1(n7382), .A2(n7381), .A3(n7380), .A4(n7379), .ZN(n7383)
         );
  OAI21_X1 U3182 ( .B1(n2662), .B2(n6239), .A(n7383), .ZN(n3023) );
  OAI222_X1 U3183 ( .A1(n6192), .A2(n4741), .B1(n2148), .B2(n6189), .C1(n6184), 
        .C2(n4671), .ZN(n7401) );
  AOI22_X1 U3184 ( .A1(n6198), .A2(n5044), .B1(n6195), .B2(n7577), .ZN(n7385)
         );
  OAI221_X1 U3185 ( .B1(n2710), .B2(n6204), .C1(n2742), .C2(n6201), .A(n7385), 
        .ZN(n7400) );
  AOI22_X1 U3186 ( .A1(n6210), .A2(n5076), .B1(n6207), .B2(n7386), .ZN(n7387)
         );
  OAI221_X1 U3187 ( .B1(n2212), .B2(n6216), .C1(n2084), .C2(n6213), .A(n7387), 
        .ZN(n7399) );
  AOI22_X1 U3188 ( .A1(n2934), .A2(n6225), .B1(n7388), .B2(n6222), .ZN(n7389)
         );
  OAI221_X1 U3189 ( .B1(n6231), .B2(n4767), .C1(n6226), .C2(n7390), .A(n7389), 
        .ZN(n7395) );
  NAND2_X1 U3190 ( .A1(n6219), .A2(n7392), .ZN(n7393) );
  NAND4_X1 U3191 ( .A1(n1275), .A2(n1276), .A3(n1274), .A4(n7393), .ZN(n7394)
         );
  OAI21_X1 U3192 ( .B1(n7395), .B2(n7394), .A(n6234), .ZN(n7397) );
  AOI22_X1 U3193 ( .A1(n6179), .A2(n4979), .B1(DATAIN[24]), .B2(n6177), .ZN(
        n7396) );
  OAI211_X1 U3194 ( .C1(n2276), .C2(n6183), .A(n7397), .B(n7396), .ZN(n7398)
         );
  NOR4_X1 U3195 ( .A1(n7401), .A2(n7400), .A3(n7399), .A4(n7398), .ZN(n7402)
         );
  OAI21_X1 U3196 ( .B1(n2661), .B2(n6238), .A(n7402), .ZN(n3022) );
  OAI222_X1 U3197 ( .A1(n6192), .A2(n4739), .B1(n2149), .B2(n6189), .C1(n6184), 
        .C2(n4670), .ZN(n7420) );
  AOI22_X1 U3198 ( .A1(n6198), .A2(n5043), .B1(n6195), .B2(n7578), .ZN(n7404)
         );
  OAI221_X1 U3199 ( .B1(n2711), .B2(n6204), .C1(n2743), .C2(n6201), .A(n7404), 
        .ZN(n7419) );
  AOI22_X1 U3200 ( .A1(n6210), .A2(n5075), .B1(n6207), .B2(n7405), .ZN(n7406)
         );
  OAI221_X1 U3201 ( .B1(n2213), .B2(n6216), .C1(n2085), .C2(n6213), .A(n7406), 
        .ZN(n7418) );
  AOI22_X1 U3202 ( .A1(n2935), .A2(n6225), .B1(n7407), .B2(n6222), .ZN(n7408)
         );
  OAI221_X1 U3203 ( .B1(n6231), .B2(n4775), .C1(n6226), .C2(n7409), .A(n7408), 
        .ZN(n7414) );
  NAND2_X1 U3204 ( .A1(n6219), .A2(n7411), .ZN(n7412) );
  NAND4_X1 U3205 ( .A1(n1292), .A2(n1293), .A3(n1291), .A4(n7412), .ZN(n7413)
         );
  OAI21_X1 U3206 ( .B1(n7414), .B2(n7413), .A(n6234), .ZN(n7416) );
  AOI22_X1 U3207 ( .A1(n6179), .A2(n4978), .B1(DATAIN[25]), .B2(n6178), .ZN(
        n7415) );
  OAI211_X1 U3208 ( .C1(n2277), .C2(n6183), .A(n7416), .B(n7415), .ZN(n7417)
         );
  NOR4_X1 U3209 ( .A1(n7420), .A2(n7419), .A3(n7418), .A4(n7417), .ZN(n7421)
         );
  OAI21_X1 U3210 ( .B1(n2660), .B2(n6238), .A(n7421), .ZN(n3021) );
  OAI222_X1 U3211 ( .A1(n6192), .A2(n4737), .B1(n2150), .B2(n6189), .C1(n6184), 
        .C2(n4669), .ZN(n7439) );
  AOI22_X1 U3212 ( .A1(n6198), .A2(n5042), .B1(n6195), .B2(n7579), .ZN(n7423)
         );
  OAI221_X1 U3213 ( .B1(n2712), .B2(n6204), .C1(n2744), .C2(n6201), .A(n7423), 
        .ZN(n7438) );
  AOI22_X1 U3214 ( .A1(n6210), .A2(n5074), .B1(n6207), .B2(n7424), .ZN(n7425)
         );
  OAI221_X1 U3215 ( .B1(n2214), .B2(n6216), .C1(n2086), .C2(n6213), .A(n7425), 
        .ZN(n7437) );
  AOI22_X1 U3216 ( .A1(n2936), .A2(n6225), .B1(n7426), .B2(n6222), .ZN(n7427)
         );
  OAI221_X1 U3217 ( .B1(n6231), .B2(n4773), .C1(n6226), .C2(n7428), .A(n7427), 
        .ZN(n7433) );
  NAND2_X1 U3218 ( .A1(n6219), .A2(n7430), .ZN(n7431) );
  NAND4_X1 U3219 ( .A1(n1309), .A2(n1310), .A3(n1308), .A4(n7431), .ZN(n7432)
         );
  OAI21_X1 U3220 ( .B1(n7433), .B2(n7432), .A(n6234), .ZN(n7435) );
  AOI22_X1 U3221 ( .A1(n6179), .A2(n4977), .B1(DATAIN[26]), .B2(n6178), .ZN(
        n7434) );
  OAI211_X1 U3222 ( .C1(n2278), .C2(n6182), .A(n7435), .B(n7434), .ZN(n7436)
         );
  NOR4_X1 U3223 ( .A1(n7439), .A2(n7438), .A3(n7437), .A4(n7436), .ZN(n7440)
         );
  OAI21_X1 U3224 ( .B1(n2659), .B2(n6238), .A(n7440), .ZN(n3020) );
  OAI222_X1 U3225 ( .A1(n6192), .A2(n4747), .B1(n2151), .B2(n6189), .C1(n6184), 
        .C2(n4668), .ZN(n7458) );
  AOI22_X1 U3226 ( .A1(n6198), .A2(n5041), .B1(n6195), .B2(n7580), .ZN(n7442)
         );
  OAI221_X1 U3227 ( .B1(n2713), .B2(n6204), .C1(n2745), .C2(n6201), .A(n7442), 
        .ZN(n7457) );
  AOI22_X1 U3228 ( .A1(n6210), .A2(n5073), .B1(n6207), .B2(n7443), .ZN(n7444)
         );
  OAI221_X1 U3229 ( .B1(n2215), .B2(n6216), .C1(n2087), .C2(n6213), .A(n7444), 
        .ZN(n7456) );
  AOI22_X1 U3230 ( .A1(n2937), .A2(n6225), .B1(n7445), .B2(n6222), .ZN(n7446)
         );
  OAI221_X1 U3231 ( .B1(n6231), .B2(n4755), .C1(n6226), .C2(n7447), .A(n7446), 
        .ZN(n7452) );
  NAND2_X1 U3232 ( .A1(n6219), .A2(n7449), .ZN(n7450) );
  NAND4_X1 U3233 ( .A1(n1326), .A2(n1327), .A3(n1325), .A4(n7450), .ZN(n7451)
         );
  OAI21_X1 U3234 ( .B1(n7452), .B2(n7451), .A(n6234), .ZN(n7454) );
  AOI22_X1 U3235 ( .A1(n6179), .A2(n4976), .B1(DATAIN[27]), .B2(n6178), .ZN(
        n7453) );
  OAI211_X1 U3236 ( .C1(n2279), .C2(n6183), .A(n7454), .B(n7453), .ZN(n7455)
         );
  NOR4_X1 U3237 ( .A1(n7458), .A2(n7457), .A3(n7456), .A4(n7455), .ZN(n7459)
         );
  OAI21_X1 U3238 ( .B1(n2658), .B2(n6238), .A(n7459), .ZN(n3019) );
  OAI222_X1 U3239 ( .A1(n6192), .A2(n4745), .B1(n2152), .B2(n6189), .C1(n6184), 
        .C2(n4667), .ZN(n7477) );
  AOI22_X1 U3240 ( .A1(n6198), .A2(n5040), .B1(n6195), .B2(n7581), .ZN(n7461)
         );
  OAI221_X1 U3241 ( .B1(n2714), .B2(n6204), .C1(n2746), .C2(n6201), .A(n7461), 
        .ZN(n7476) );
  AOI22_X1 U3242 ( .A1(n6210), .A2(n5072), .B1(n6207), .B2(n7462), .ZN(n7463)
         );
  OAI221_X1 U3243 ( .B1(n2216), .B2(n6216), .C1(n2088), .C2(n6213), .A(n7463), 
        .ZN(n7475) );
  AOI22_X1 U3244 ( .A1(n2938), .A2(n6225), .B1(n7464), .B2(n6222), .ZN(n7465)
         );
  OAI221_X1 U3245 ( .B1(n6231), .B2(n4779), .C1(n6226), .C2(n7466), .A(n7465), 
        .ZN(n7471) );
  NAND2_X1 U3246 ( .A1(n6219), .A2(n7468), .ZN(n7469) );
  NAND4_X1 U3247 ( .A1(n1343), .A2(n1344), .A3(n1342), .A4(n7469), .ZN(n7470)
         );
  OAI21_X1 U3248 ( .B1(n7471), .B2(n7470), .A(n6234), .ZN(n7473) );
  AOI22_X1 U3249 ( .A1(n6179), .A2(n4975), .B1(DATAIN[28]), .B2(n6178), .ZN(
        n7472) );
  OAI211_X1 U3250 ( .C1(n2280), .C2(n6182), .A(n7473), .B(n7472), .ZN(n7474)
         );
  NOR4_X1 U3251 ( .A1(n7477), .A2(n7476), .A3(n7475), .A4(n7474), .ZN(n7478)
         );
  OAI21_X1 U3252 ( .B1(n2657), .B2(n6238), .A(n7478), .ZN(n3018) );
  OAI222_X1 U3253 ( .A1(n6192), .A2(n4743), .B1(n2153), .B2(n6189), .C1(n6184), 
        .C2(n4666), .ZN(n7496) );
  AOI22_X1 U3254 ( .A1(n6198), .A2(n5039), .B1(n6195), .B2(n7582), .ZN(n7480)
         );
  OAI221_X1 U3255 ( .B1(n2715), .B2(n6204), .C1(n2747), .C2(n6201), .A(n7480), 
        .ZN(n7495) );
  AOI22_X1 U3256 ( .A1(n6210), .A2(n5071), .B1(n6207), .B2(n7481), .ZN(n7482)
         );
  OAI221_X1 U3257 ( .B1(n2217), .B2(n6216), .C1(n2089), .C2(n6213), .A(n7482), 
        .ZN(n7494) );
  AOI22_X1 U3258 ( .A1(n2939), .A2(n6225), .B1(n7483), .B2(n6222), .ZN(n7484)
         );
  OAI221_X1 U3259 ( .B1(n6231), .B2(n4777), .C1(n6226), .C2(n7485), .A(n7484), 
        .ZN(n7490) );
  NAND2_X1 U3260 ( .A1(n6219), .A2(n7487), .ZN(n7488) );
  NAND4_X1 U3261 ( .A1(n1360), .A2(n1361), .A3(n1359), .A4(n7488), .ZN(n7489)
         );
  OAI21_X1 U3262 ( .B1(n7490), .B2(n7489), .A(n6234), .ZN(n7492) );
  AOI22_X1 U3263 ( .A1(n6179), .A2(n4974), .B1(DATAIN[29]), .B2(n6178), .ZN(
        n7491) );
  OAI211_X1 U3264 ( .C1(n2281), .C2(n6183), .A(n7492), .B(n7491), .ZN(n7493)
         );
  NOR4_X1 U3265 ( .A1(n7496), .A2(n7495), .A3(n7494), .A4(n7493), .ZN(n7497)
         );
  OAI21_X1 U3266 ( .B1(n2656), .B2(n6238), .A(n7497), .ZN(n3017) );
  OAI222_X1 U3267 ( .A1(n6192), .A2(n4749), .B1(n2154), .B2(n6189), .C1(n6184), 
        .C2(n4665), .ZN(n7517) );
  AOI22_X1 U3268 ( .A1(n6198), .A2(n5038), .B1(n6195), .B2(n7583), .ZN(n7499)
         );
  OAI221_X1 U3269 ( .B1(n2716), .B2(n6204), .C1(n2748), .C2(n6201), .A(n7499), 
        .ZN(n7516) );
  AOI22_X1 U3270 ( .A1(n6210), .A2(n5070), .B1(n6207), .B2(n7500), .ZN(n7501)
         );
  OAI221_X1 U3271 ( .B1(n2218), .B2(n6216), .C1(n2090), .C2(n6213), .A(n7501), 
        .ZN(n7515) );
  AOI22_X1 U3272 ( .A1(n2940), .A2(n6225), .B1(n7502), .B2(n6222), .ZN(n7503)
         );
  OAI221_X1 U3273 ( .B1(n6231), .B2(n4781), .C1(n6226), .C2(n7504), .A(n7503), 
        .ZN(n7509) );
  NAND2_X1 U3274 ( .A1(n6219), .A2(n7506), .ZN(n7507) );
  NAND4_X1 U3275 ( .A1(n1377), .A2(n1378), .A3(n1376), .A4(n7507), .ZN(n7508)
         );
  OAI21_X1 U3276 ( .B1(n7509), .B2(n7508), .A(n6234), .ZN(n7513) );
  AOI22_X1 U3277 ( .A1(n6179), .A2(n4973), .B1(DATAIN[30]), .B2(n6178), .ZN(
        n7512) );
  OAI211_X1 U3278 ( .C1(n2282), .C2(n6182), .A(n7513), .B(n7512), .ZN(n7514)
         );
  NOR4_X1 U3279 ( .A1(n7517), .A2(n7516), .A3(n7515), .A4(n7514), .ZN(n7518)
         );
  OAI21_X1 U3280 ( .B1(n2655), .B2(n6238), .A(n7518), .ZN(n3016) );
  OAI222_X1 U3281 ( .A1(n6192), .A2(n4751), .B1(n2155), .B2(n6189), .C1(n6184), 
        .C2(n4664), .ZN(n7549) );
  AOI22_X1 U3282 ( .A1(n6198), .A2(n5037), .B1(n6195), .B2(n7584), .ZN(n7523)
         );
  OAI221_X1 U3283 ( .B1(n2717), .B2(n6204), .C1(n2749), .C2(n6201), .A(n7523), 
        .ZN(n7548) );
  AOI22_X1 U3284 ( .A1(n6210), .A2(n5069), .B1(n6207), .B2(n7526), .ZN(n7527)
         );
  OAI221_X1 U3285 ( .B1(n2219), .B2(n6216), .C1(n2091), .C2(n6213), .A(n7527), 
        .ZN(n7547) );
  OAI22_X1 U3286 ( .A1(n3773), .A2(n4901), .B1(n2315), .B2(n4899), .ZN(n7530)
         );
  AOI221_X1 U3287 ( .B1(n6219), .B2(n7531), .C1(n6312), .C2(n7587), .A(n7530), 
        .ZN(n7539) );
  AOI222_X1 U3288 ( .A1(n6335), .A2(n4093), .B1(n6324), .B2(n7585), .C1(n6338), 
        .C2(n4061), .ZN(n7538) );
  AOI22_X1 U3289 ( .A1(n2941), .A2(n6225), .B1(n7532), .B2(n6222), .ZN(n7533)
         );
  OAI221_X1 U3290 ( .B1(n4815), .B2(n6231), .C1(n7534), .C2(n6226), .A(n7533), 
        .ZN(n7536) );
  NOR4_X1 U3291 ( .A1(n7536), .A2(n1425), .A3(n1424), .A4(n1421), .ZN(n7537)
         );
  NAND3_X1 U3292 ( .A1(n7539), .A2(n7538), .A3(n7537), .ZN(n7541) );
  AOI22_X1 U3293 ( .A1(n6234), .A2(n7541), .B1(n4896), .B2(n7540), .ZN(n7543)
         );
  OAI221_X1 U3294 ( .B1(n2251), .B2(n7545), .C1(n7544), .C2(n6374), .A(n7543), 
        .ZN(n7546) );
  NOR4_X1 U3295 ( .A1(n7549), .A2(n7548), .A3(n7547), .A4(n7546), .ZN(n7550)
         );
  OAI21_X1 U3296 ( .B1(n6238), .B2(n7551), .A(n7550), .ZN(n3015) );
  MUX2_X1 U3297 ( .A(n5235), .B(DATAIN[0]), .S(n6241), .Z(n3047) );
  MUX2_X1 U3298 ( .A(n5297), .B(DATAIN[1]), .S(n6241), .Z(n3048) );
  MUX2_X1 U3299 ( .A(n5296), .B(DATAIN[2]), .S(n6241), .Z(n3049) );
  MUX2_X1 U3300 ( .A(n5295), .B(DATAIN[3]), .S(n6241), .Z(n3050) );
  MUX2_X1 U3301 ( .A(n5294), .B(DATAIN[4]), .S(n6241), .Z(n3051) );
  MUX2_X1 U3302 ( .A(n5293), .B(DATAIN[5]), .S(n6241), .Z(n3052) );
  MUX2_X1 U3303 ( .A(n5292), .B(DATAIN[6]), .S(n6241), .Z(n3053) );
  MUX2_X1 U3304 ( .A(n5291), .B(DATAIN[7]), .S(n6241), .Z(n3054) );
  MUX2_X1 U3305 ( .A(n5290), .B(DATAIN[8]), .S(n6241), .Z(n3055) );
  MUX2_X1 U3306 ( .A(n5289), .B(DATAIN[9]), .S(n6241), .Z(n3056) );
  MUX2_X1 U3307 ( .A(n5288), .B(DATAIN[10]), .S(n6241), .Z(n3057) );
  MUX2_X1 U3308 ( .A(n5287), .B(DATAIN[11]), .S(n6241), .Z(n3058) );
  MUX2_X1 U3309 ( .A(n5286), .B(DATAIN[12]), .S(n6242), .Z(n3059) );
  MUX2_X1 U3310 ( .A(n5285), .B(DATAIN[13]), .S(n6242), .Z(n3060) );
  MUX2_X1 U3311 ( .A(n5284), .B(DATAIN[14]), .S(n6242), .Z(n3061) );
  MUX2_X1 U3312 ( .A(n5283), .B(DATAIN[15]), .S(n6242), .Z(n3062) );
  MUX2_X1 U3313 ( .A(n5282), .B(DATAIN[16]), .S(n6242), .Z(n3063) );
  MUX2_X1 U3314 ( .A(n5281), .B(DATAIN[17]), .S(n6242), .Z(n3064) );
  MUX2_X1 U3315 ( .A(n5280), .B(DATAIN[18]), .S(n6242), .Z(n3065) );
  MUX2_X1 U3316 ( .A(n5279), .B(DATAIN[19]), .S(n6242), .Z(n3066) );
  MUX2_X1 U3317 ( .A(n5278), .B(DATAIN[20]), .S(n6242), .Z(n3067) );
  MUX2_X1 U3318 ( .A(n5277), .B(DATAIN[21]), .S(n6242), .Z(n3068) );
  MUX2_X1 U3319 ( .A(n5276), .B(DATAIN[22]), .S(n6242), .Z(n3069) );
  MUX2_X1 U3320 ( .A(n5275), .B(DATAIN[23]), .S(n6242), .Z(n3070) );
  MUX2_X1 U3321 ( .A(n5274), .B(DATAIN[24]), .S(n6243), .Z(n3071) );
  MUX2_X1 U3322 ( .A(n5273), .B(DATAIN[25]), .S(n6243), .Z(n3072) );
  MUX2_X1 U3323 ( .A(n5272), .B(DATAIN[26]), .S(n6243), .Z(n3073) );
  MUX2_X1 U3324 ( .A(n5271), .B(DATAIN[27]), .S(n6243), .Z(n3074) );
  MUX2_X1 U3325 ( .A(n5270), .B(DATAIN[28]), .S(n6243), .Z(n3075) );
  MUX2_X1 U3326 ( .A(n5269), .B(DATAIN[29]), .S(n6243), .Z(n3076) );
  MUX2_X1 U3327 ( .A(n5268), .B(DATAIN[30]), .S(n6243), .Z(n3077) );
  MUX2_X1 U3328 ( .A(n5234), .B(DATAIN[31]), .S(n6243), .Z(n3078) );
  MUX2_X1 U3329 ( .A(n5171), .B(DATAIN[0]), .S(n6244), .Z(n3111) );
  MUX2_X1 U3330 ( .A(n5167), .B(DATAIN[1]), .S(n6244), .Z(n3112) );
  MUX2_X1 U3331 ( .A(n5166), .B(DATAIN[2]), .S(n6244), .Z(n3113) );
  MUX2_X1 U3332 ( .A(n5165), .B(DATAIN[3]), .S(n6244), .Z(n3114) );
  MUX2_X1 U3333 ( .A(n5164), .B(DATAIN[4]), .S(n6244), .Z(n3115) );
  MUX2_X1 U3334 ( .A(n5163), .B(DATAIN[5]), .S(n6244), .Z(n3116) );
  MUX2_X1 U3335 ( .A(n5162), .B(DATAIN[6]), .S(n6244), .Z(n3117) );
  MUX2_X1 U3336 ( .A(n5161), .B(DATAIN[7]), .S(n6244), .Z(n3118) );
  MUX2_X1 U3337 ( .A(n5160), .B(DATAIN[8]), .S(n6244), .Z(n3119) );
  MUX2_X1 U3338 ( .A(n5159), .B(DATAIN[9]), .S(n6244), .Z(n3120) );
  MUX2_X1 U3339 ( .A(n5158), .B(DATAIN[10]), .S(n6244), .Z(n3121) );
  MUX2_X1 U3340 ( .A(n5157), .B(DATAIN[11]), .S(n6244), .Z(n3122) );
  MUX2_X1 U3341 ( .A(n5156), .B(DATAIN[12]), .S(n6245), .Z(n3123) );
  MUX2_X1 U3342 ( .A(n5155), .B(DATAIN[13]), .S(n6245), .Z(n3124) );
  MUX2_X1 U3343 ( .A(n5154), .B(DATAIN[14]), .S(n6245), .Z(n3125) );
  MUX2_X1 U3344 ( .A(n5153), .B(DATAIN[15]), .S(n6245), .Z(n3126) );
  MUX2_X1 U3345 ( .A(n5152), .B(DATAIN[16]), .S(n6245), .Z(n3127) );
  MUX2_X1 U3346 ( .A(n5151), .B(DATAIN[17]), .S(n6245), .Z(n3128) );
  MUX2_X1 U3347 ( .A(n5150), .B(DATAIN[18]), .S(n6245), .Z(n3129) );
  MUX2_X1 U3348 ( .A(n5149), .B(DATAIN[19]), .S(n6245), .Z(n3130) );
  MUX2_X1 U3349 ( .A(n5148), .B(DATAIN[20]), .S(n6245), .Z(n3131) );
  MUX2_X1 U3350 ( .A(n5147), .B(DATAIN[21]), .S(n6245), .Z(n3132) );
  MUX2_X1 U3351 ( .A(n5146), .B(DATAIN[22]), .S(n6245), .Z(n3133) );
  MUX2_X1 U3352 ( .A(n5145), .B(DATAIN[23]), .S(n6245), .Z(n3134) );
  MUX2_X1 U3353 ( .A(n5144), .B(DATAIN[24]), .S(n6246), .Z(n3135) );
  MUX2_X1 U3354 ( .A(n5143), .B(DATAIN[25]), .S(n6246), .Z(n3136) );
  MUX2_X1 U3355 ( .A(n5142), .B(DATAIN[26]), .S(n6246), .Z(n3137) );
  MUX2_X1 U3356 ( .A(n5141), .B(DATAIN[27]), .S(n6246), .Z(n3138) );
  MUX2_X1 U3357 ( .A(n5140), .B(DATAIN[28]), .S(n6246), .Z(n3139) );
  MUX2_X1 U3358 ( .A(n5139), .B(DATAIN[29]), .S(n6246), .Z(n3140) );
  MUX2_X1 U3359 ( .A(n5138), .B(DATAIN[30]), .S(n6246), .Z(n3141) );
  MUX2_X1 U3360 ( .A(n5137), .B(DATAIN[31]), .S(n6246), .Z(n3142) );
  MUX2_X1 U3361 ( .A(n5680), .B(DATAIN[0]), .S(n6247), .Z(n3239) );
  MUX2_X1 U3362 ( .A(n5545), .B(DATAIN[1]), .S(n6247), .Z(n3240) );
  MUX2_X1 U3363 ( .A(n5544), .B(DATAIN[2]), .S(n6247), .Z(n3241) );
  MUX2_X1 U3364 ( .A(n5543), .B(DATAIN[3]), .S(n6247), .Z(n3242) );
  MUX2_X1 U3365 ( .A(n5542), .B(DATAIN[4]), .S(n6247), .Z(n3243) );
  MUX2_X1 U3366 ( .A(n5541), .B(DATAIN[5]), .S(n6247), .Z(n3244) );
  MUX2_X1 U3367 ( .A(n5540), .B(DATAIN[6]), .S(n6247), .Z(n3245) );
  MUX2_X1 U3368 ( .A(n5539), .B(DATAIN[7]), .S(n6247), .Z(n3246) );
  MUX2_X1 U3369 ( .A(n5538), .B(DATAIN[8]), .S(n6247), .Z(n3247) );
  MUX2_X1 U3370 ( .A(n5537), .B(DATAIN[9]), .S(n6247), .Z(n3248) );
  MUX2_X1 U3371 ( .A(n5536), .B(DATAIN[10]), .S(n6247), .Z(n3249) );
  MUX2_X1 U3372 ( .A(n5535), .B(DATAIN[11]), .S(n6247), .Z(n3250) );
  MUX2_X1 U3373 ( .A(n5534), .B(DATAIN[12]), .S(n6248), .Z(n3251) );
  MUX2_X1 U3374 ( .A(n5533), .B(DATAIN[13]), .S(n6248), .Z(n3252) );
  MUX2_X1 U3375 ( .A(n5532), .B(DATAIN[14]), .S(n6248), .Z(n3253) );
  MUX2_X1 U3376 ( .A(n5531), .B(DATAIN[15]), .S(n6248), .Z(n3254) );
  MUX2_X1 U3377 ( .A(n5530), .B(DATAIN[16]), .S(n6248), .Z(n3255) );
  MUX2_X1 U3378 ( .A(n5529), .B(DATAIN[17]), .S(n6248), .Z(n3256) );
  MUX2_X1 U3379 ( .A(n5528), .B(DATAIN[18]), .S(n6248), .Z(n3257) );
  MUX2_X1 U3380 ( .A(n5527), .B(DATAIN[19]), .S(n6248), .Z(n3258) );
  MUX2_X1 U3381 ( .A(n5526), .B(DATAIN[20]), .S(n6248), .Z(n3259) );
  MUX2_X1 U3382 ( .A(n5525), .B(DATAIN[21]), .S(n6248), .Z(n3260) );
  MUX2_X1 U3383 ( .A(n5524), .B(DATAIN[22]), .S(n6248), .Z(n3261) );
  MUX2_X1 U3384 ( .A(n5523), .B(DATAIN[23]), .S(n6248), .Z(n3262) );
  MUX2_X1 U3385 ( .A(n5522), .B(DATAIN[24]), .S(n6249), .Z(n3263) );
  MUX2_X1 U3386 ( .A(n5521), .B(DATAIN[25]), .S(n6249), .Z(n3264) );
  MUX2_X1 U3387 ( .A(n5520), .B(DATAIN[26]), .S(n6249), .Z(n3265) );
  MUX2_X1 U3388 ( .A(n5519), .B(DATAIN[27]), .S(n6249), .Z(n3266) );
  MUX2_X1 U3389 ( .A(n5518), .B(DATAIN[28]), .S(n6249), .Z(n3267) );
  MUX2_X1 U3390 ( .A(n5517), .B(DATAIN[29]), .S(n6249), .Z(n3268) );
  MUX2_X1 U3391 ( .A(n5516), .B(DATAIN[30]), .S(n6249), .Z(n3269) );
  MUX2_X1 U3392 ( .A(n5515), .B(DATAIN[31]), .S(n6249), .Z(n3270) );
  MUX2_X1 U3393 ( .A(n5486), .B(DATAIN[0]), .S(n6250), .Z(n3271) );
  MUX2_X1 U3394 ( .A(n5482), .B(DATAIN[1]), .S(n6250), .Z(n3272) );
  MUX2_X1 U3395 ( .A(n5481), .B(DATAIN[2]), .S(n6250), .Z(n3273) );
  MUX2_X1 U3396 ( .A(n5480), .B(DATAIN[3]), .S(n6250), .Z(n3274) );
  MUX2_X1 U3397 ( .A(n5479), .B(DATAIN[4]), .S(n6250), .Z(n3275) );
  MUX2_X1 U3398 ( .A(n5478), .B(DATAIN[5]), .S(n6250), .Z(n3276) );
  MUX2_X1 U3399 ( .A(n5477), .B(DATAIN[6]), .S(n6250), .Z(n3277) );
  MUX2_X1 U3400 ( .A(n5476), .B(DATAIN[7]), .S(n6250), .Z(n3278) );
  MUX2_X1 U3401 ( .A(n5475), .B(DATAIN[8]), .S(n6250), .Z(n3279) );
  MUX2_X1 U3402 ( .A(n5474), .B(DATAIN[9]), .S(n6250), .Z(n3280) );
  MUX2_X1 U3403 ( .A(n5473), .B(DATAIN[10]), .S(n6250), .Z(n3281) );
  MUX2_X1 U3404 ( .A(n5472), .B(DATAIN[11]), .S(n6251), .Z(n3282) );
  MUX2_X1 U3405 ( .A(n5471), .B(DATAIN[12]), .S(n6251), .Z(n3283) );
  MUX2_X1 U3406 ( .A(n5470), .B(DATAIN[13]), .S(n6251), .Z(n3284) );
  MUX2_X1 U3407 ( .A(n5469), .B(DATAIN[14]), .S(n6251), .Z(n3285) );
  MUX2_X1 U3408 ( .A(n5468), .B(DATAIN[15]), .S(n6251), .Z(n3286) );
  MUX2_X1 U3409 ( .A(n5467), .B(DATAIN[16]), .S(n6251), .Z(n3287) );
  MUX2_X1 U3410 ( .A(n5466), .B(DATAIN[17]), .S(n6251), .Z(n3288) );
  MUX2_X1 U3411 ( .A(n5465), .B(DATAIN[18]), .S(n6251), .Z(n3289) );
  MUX2_X1 U3412 ( .A(n5464), .B(DATAIN[19]), .S(n6251), .Z(n3290) );
  MUX2_X1 U3413 ( .A(n5463), .B(DATAIN[20]), .S(n6251), .Z(n3291) );
  MUX2_X1 U3414 ( .A(n5462), .B(DATAIN[21]), .S(n6251), .Z(n3292) );
  MUX2_X1 U3415 ( .A(n5461), .B(DATAIN[22]), .S(n6251), .Z(n3293) );
  MUX2_X1 U3416 ( .A(n5460), .B(DATAIN[23]), .S(n6252), .Z(n3294) );
  MUX2_X1 U3417 ( .A(n5459), .B(DATAIN[24]), .S(n6252), .Z(n3295) );
  MUX2_X1 U3418 ( .A(n5458), .B(DATAIN[25]), .S(n6252), .Z(n3296) );
  MUX2_X1 U3419 ( .A(n5457), .B(DATAIN[26]), .S(n6252), .Z(n3297) );
  MUX2_X1 U3420 ( .A(n5456), .B(DATAIN[27]), .S(n6252), .Z(n3298) );
  MUX2_X1 U3421 ( .A(n5455), .B(DATAIN[28]), .S(n6252), .Z(n3299) );
  MUX2_X1 U3422 ( .A(n5454), .B(DATAIN[29]), .S(n6252), .Z(n3300) );
  MUX2_X1 U3423 ( .A(n5453), .B(DATAIN[30]), .S(n6252), .Z(n3301) );
  MUX2_X1 U3424 ( .A(n5776), .B(DATAIN[0]), .S(n6253), .Z(n3303) );
  MUX2_X1 U3425 ( .A(n5775), .B(DATAIN[1]), .S(n6253), .Z(n3304) );
  MUX2_X1 U3426 ( .A(n5774), .B(DATAIN[2]), .S(n6253), .Z(n3305) );
  MUX2_X1 U3427 ( .A(n5773), .B(DATAIN[3]), .S(n6253), .Z(n3306) );
  MUX2_X1 U3428 ( .A(n5772), .B(DATAIN[4]), .S(n6253), .Z(n3307) );
  MUX2_X1 U3429 ( .A(n5771), .B(DATAIN[5]), .S(n6253), .Z(n3308) );
  MUX2_X1 U3430 ( .A(n5770), .B(DATAIN[6]), .S(n6253), .Z(n3309) );
  MUX2_X1 U3431 ( .A(n5769), .B(DATAIN[7]), .S(n6253), .Z(n3310) );
  MUX2_X1 U3432 ( .A(n5768), .B(DATAIN[8]), .S(n6253), .Z(n3311) );
  MUX2_X1 U3433 ( .A(n5767), .B(DATAIN[9]), .S(n6253), .Z(n3312) );
  MUX2_X1 U3434 ( .A(n5766), .B(DATAIN[10]), .S(n6253), .Z(n3313) );
  MUX2_X1 U3435 ( .A(n5765), .B(DATAIN[11]), .S(n6253), .Z(n3314) );
  MUX2_X1 U3436 ( .A(n5764), .B(DATAIN[12]), .S(n6254), .Z(n3315) );
  MUX2_X1 U3437 ( .A(n5763), .B(DATAIN[13]), .S(n6254), .Z(n3316) );
  MUX2_X1 U3438 ( .A(n5762), .B(DATAIN[14]), .S(n6254), .Z(n3317) );
  MUX2_X1 U3439 ( .A(n5761), .B(DATAIN[15]), .S(n6254), .Z(n3318) );
  MUX2_X1 U3440 ( .A(n5760), .B(DATAIN[16]), .S(n6254), .Z(n3319) );
  MUX2_X1 U3441 ( .A(n5759), .B(DATAIN[17]), .S(n6254), .Z(n3320) );
  MUX2_X1 U3442 ( .A(n5758), .B(DATAIN[18]), .S(n6254), .Z(n3321) );
  MUX2_X1 U3443 ( .A(n5757), .B(DATAIN[19]), .S(n6254), .Z(n3322) );
  MUX2_X1 U3444 ( .A(n5756), .B(DATAIN[20]), .S(n6254), .Z(n3323) );
  MUX2_X1 U3445 ( .A(n5755), .B(DATAIN[21]), .S(n6254), .Z(n3324) );
  MUX2_X1 U3446 ( .A(n5754), .B(DATAIN[22]), .S(n6254), .Z(n3325) );
  MUX2_X1 U3447 ( .A(n5753), .B(DATAIN[23]), .S(n6254), .Z(n3326) );
  MUX2_X1 U3448 ( .A(n5752), .B(DATAIN[24]), .S(n6255), .Z(n3327) );
  MUX2_X1 U3449 ( .A(n5751), .B(DATAIN[25]), .S(n6255), .Z(n3328) );
  MUX2_X1 U3450 ( .A(n5750), .B(DATAIN[26]), .S(n6255), .Z(n3329) );
  MUX2_X1 U3451 ( .A(n5749), .B(DATAIN[27]), .S(n6255), .Z(n3330) );
  MUX2_X1 U3452 ( .A(n5748), .B(DATAIN[28]), .S(n6255), .Z(n3331) );
  MUX2_X1 U3453 ( .A(n5747), .B(DATAIN[29]), .S(n6255), .Z(n3332) );
  MUX2_X1 U3454 ( .A(n5746), .B(DATAIN[30]), .S(n6255), .Z(n3333) );
  MUX2_X1 U3455 ( .A(n5745), .B(DATAIN[31]), .S(n6255), .Z(n3334) );
  MUX2_X1 U3456 ( .A(n5237), .B(DATAIN[0]), .S(n6256), .Z(n3335) );
  MUX2_X1 U3457 ( .A(n5267), .B(DATAIN[1]), .S(n6256), .Z(n3336) );
  MUX2_X1 U3458 ( .A(n5266), .B(DATAIN[2]), .S(n6256), .Z(n3337) );
  MUX2_X1 U3459 ( .A(n5265), .B(DATAIN[3]), .S(n6256), .Z(n3338) );
  MUX2_X1 U3460 ( .A(n5264), .B(DATAIN[4]), .S(n6256), .Z(n3339) );
  MUX2_X1 U3461 ( .A(n5263), .B(DATAIN[5]), .S(n6256), .Z(n3340) );
  MUX2_X1 U3462 ( .A(n5262), .B(DATAIN[6]), .S(n6256), .Z(n3341) );
  MUX2_X1 U3463 ( .A(n5261), .B(DATAIN[7]), .S(n6256), .Z(n3342) );
  MUX2_X1 U3464 ( .A(n5260), .B(DATAIN[8]), .S(n6256), .Z(n3343) );
  MUX2_X1 U3465 ( .A(n5259), .B(DATAIN[9]), .S(n6256), .Z(n3344) );
  MUX2_X1 U3466 ( .A(n5258), .B(DATAIN[10]), .S(n6256), .Z(n3345) );
  MUX2_X1 U3467 ( .A(n5257), .B(DATAIN[11]), .S(n6256), .Z(n3346) );
  MUX2_X1 U3468 ( .A(n5256), .B(DATAIN[12]), .S(n6257), .Z(n3347) );
  MUX2_X1 U3469 ( .A(n5255), .B(DATAIN[13]), .S(n6257), .Z(n3348) );
  MUX2_X1 U3470 ( .A(n5254), .B(DATAIN[14]), .S(n6257), .Z(n3349) );
  MUX2_X1 U3471 ( .A(n5253), .B(DATAIN[15]), .S(n6257), .Z(n3350) );
  MUX2_X1 U3472 ( .A(n5252), .B(DATAIN[16]), .S(n6257), .Z(n3351) );
  MUX2_X1 U3473 ( .A(n5251), .B(DATAIN[17]), .S(n6257), .Z(n3352) );
  MUX2_X1 U3474 ( .A(n5250), .B(DATAIN[18]), .S(n6257), .Z(n3353) );
  MUX2_X1 U3475 ( .A(n5249), .B(DATAIN[19]), .S(n6257), .Z(n3354) );
  MUX2_X1 U3476 ( .A(n5248), .B(DATAIN[20]), .S(n6257), .Z(n3355) );
  MUX2_X1 U3477 ( .A(n5247), .B(DATAIN[21]), .S(n6257), .Z(n3356) );
  MUX2_X1 U3478 ( .A(n5246), .B(DATAIN[22]), .S(n6257), .Z(n3357) );
  MUX2_X1 U3479 ( .A(n5245), .B(DATAIN[23]), .S(n6257), .Z(n3358) );
  MUX2_X1 U3480 ( .A(n5244), .B(DATAIN[24]), .S(n6258), .Z(n3359) );
  MUX2_X1 U3481 ( .A(n5243), .B(DATAIN[25]), .S(n6258), .Z(n3360) );
  MUX2_X1 U3482 ( .A(n5242), .B(DATAIN[26]), .S(n6258), .Z(n3361) );
  MUX2_X1 U3483 ( .A(n5241), .B(DATAIN[27]), .S(n6258), .Z(n3362) );
  MUX2_X1 U3484 ( .A(n5240), .B(DATAIN[28]), .S(n6258), .Z(n3363) );
  MUX2_X1 U3485 ( .A(n5239), .B(DATAIN[29]), .S(n6258), .Z(n3364) );
  MUX2_X1 U3486 ( .A(n5238), .B(DATAIN[30]), .S(n6258), .Z(n3365) );
  MUX2_X1 U3487 ( .A(n5236), .B(DATAIN[31]), .S(n6258), .Z(n3366) );
  MUX2_X1 U3488 ( .A(n5579), .B(DATAIN[0]), .S(n6259), .Z(n3367) );
  MUX2_X1 U3489 ( .A(n5578), .B(DATAIN[1]), .S(n6259), .Z(n3368) );
  MUX2_X1 U3490 ( .A(n5577), .B(DATAIN[2]), .S(n6259), .Z(n3369) );
  MUX2_X1 U3491 ( .A(n5576), .B(DATAIN[3]), .S(n6259), .Z(n3370) );
  MUX2_X1 U3492 ( .A(n5575), .B(DATAIN[4]), .S(n6259), .Z(n3371) );
  MUX2_X1 U3493 ( .A(n5574), .B(DATAIN[5]), .S(n6259), .Z(n3372) );
  MUX2_X1 U3494 ( .A(n5573), .B(DATAIN[6]), .S(n6259), .Z(n3373) );
  MUX2_X1 U3495 ( .A(n5572), .B(DATAIN[7]), .S(n6259), .Z(n3374) );
  MUX2_X1 U3496 ( .A(n5571), .B(DATAIN[8]), .S(n6259), .Z(n3375) );
  MUX2_X1 U3497 ( .A(n5570), .B(DATAIN[9]), .S(n6259), .Z(n3376) );
  MUX2_X1 U3498 ( .A(n5569), .B(DATAIN[10]), .S(n6259), .Z(n3377) );
  MUX2_X1 U3499 ( .A(n5568), .B(DATAIN[11]), .S(n6259), .Z(n3378) );
  MUX2_X1 U3500 ( .A(n5567), .B(DATAIN[12]), .S(n6260), .Z(n3379) );
  MUX2_X1 U3501 ( .A(n5566), .B(DATAIN[13]), .S(n6260), .Z(n3380) );
  MUX2_X1 U3502 ( .A(n5565), .B(DATAIN[14]), .S(n6260), .Z(n3381) );
  MUX2_X1 U3503 ( .A(n5564), .B(DATAIN[15]), .S(n6260), .Z(n3382) );
  MUX2_X1 U3504 ( .A(n5563), .B(DATAIN[16]), .S(n6260), .Z(n3383) );
  MUX2_X1 U3505 ( .A(n5562), .B(DATAIN[17]), .S(n6260), .Z(n3384) );
  MUX2_X1 U3506 ( .A(n5561), .B(DATAIN[18]), .S(n6260), .Z(n3385) );
  MUX2_X1 U3507 ( .A(n5560), .B(DATAIN[19]), .S(n6260), .Z(n3386) );
  MUX2_X1 U3508 ( .A(n5559), .B(DATAIN[20]), .S(n6260), .Z(n3387) );
  MUX2_X1 U3509 ( .A(n5558), .B(DATAIN[21]), .S(n6260), .Z(n3388) );
  MUX2_X1 U3510 ( .A(n5557), .B(DATAIN[22]), .S(n6260), .Z(n3389) );
  MUX2_X1 U3511 ( .A(n5556), .B(DATAIN[23]), .S(n6260), .Z(n3390) );
  MUX2_X1 U3512 ( .A(n5555), .B(DATAIN[24]), .S(n6261), .Z(n3391) );
  MUX2_X1 U3513 ( .A(n5554), .B(DATAIN[25]), .S(n6261), .Z(n3392) );
  MUX2_X1 U3514 ( .A(n5553), .B(DATAIN[26]), .S(n6261), .Z(n3393) );
  MUX2_X1 U3515 ( .A(n5552), .B(DATAIN[27]), .S(n6261), .Z(n3394) );
  MUX2_X1 U3516 ( .A(n5551), .B(DATAIN[28]), .S(n6261), .Z(n3395) );
  MUX2_X1 U3517 ( .A(n5550), .B(DATAIN[29]), .S(n6261), .Z(n3396) );
  MUX2_X1 U3518 ( .A(n5549), .B(DATAIN[30]), .S(n6261), .Z(n3397) );
  MUX2_X1 U3519 ( .A(n5548), .B(DATAIN[31]), .S(n6261), .Z(n3398) );
  MUX2_X1 U3520 ( .A(n5743), .B(DATAIN[0]), .S(n6262), .Z(n3399) );
  MUX2_X1 U3521 ( .A(n5742), .B(DATAIN[1]), .S(n6262), .Z(n3400) );
  MUX2_X1 U3522 ( .A(n5741), .B(DATAIN[2]), .S(n6262), .Z(n3401) );
  MUX2_X1 U3523 ( .A(n5740), .B(DATAIN[3]), .S(n6262), .Z(n3402) );
  MUX2_X1 U3524 ( .A(n5739), .B(DATAIN[4]), .S(n6262), .Z(n3403) );
  MUX2_X1 U3525 ( .A(n5738), .B(DATAIN[5]), .S(n6262), .Z(n3404) );
  MUX2_X1 U3526 ( .A(n5737), .B(DATAIN[6]), .S(n6262), .Z(n3405) );
  MUX2_X1 U3527 ( .A(n5736), .B(DATAIN[7]), .S(n6262), .Z(n3406) );
  MUX2_X1 U3528 ( .A(n5735), .B(DATAIN[8]), .S(n6262), .Z(n3407) );
  MUX2_X1 U3529 ( .A(n5734), .B(DATAIN[9]), .S(n6262), .Z(n3408) );
  MUX2_X1 U3530 ( .A(n5733), .B(DATAIN[10]), .S(n6262), .Z(n3409) );
  MUX2_X1 U3531 ( .A(n5732), .B(DATAIN[11]), .S(n6262), .Z(n3410) );
  MUX2_X1 U3532 ( .A(n5731), .B(DATAIN[12]), .S(n6263), .Z(n3411) );
  MUX2_X1 U3533 ( .A(n5730), .B(DATAIN[13]), .S(n6263), .Z(n3412) );
  MUX2_X1 U3534 ( .A(n5729), .B(DATAIN[14]), .S(n6263), .Z(n3413) );
  MUX2_X1 U3535 ( .A(n5728), .B(DATAIN[15]), .S(n6263), .Z(n3414) );
  MUX2_X1 U3536 ( .A(n5727), .B(DATAIN[16]), .S(n6263), .Z(n3415) );
  MUX2_X1 U3537 ( .A(n5726), .B(DATAIN[17]), .S(n6263), .Z(n3416) );
  MUX2_X1 U3538 ( .A(n5725), .B(DATAIN[18]), .S(n6263), .Z(n3417) );
  MUX2_X1 U3539 ( .A(n5724), .B(DATAIN[19]), .S(n6263), .Z(n3418) );
  MUX2_X1 U3540 ( .A(n5723), .B(DATAIN[20]), .S(n6263), .Z(n3419) );
  MUX2_X1 U3541 ( .A(n5722), .B(DATAIN[21]), .S(n6263), .Z(n3420) );
  MUX2_X1 U3542 ( .A(n5721), .B(DATAIN[22]), .S(n6263), .Z(n3421) );
  MUX2_X1 U3543 ( .A(n5720), .B(DATAIN[23]), .S(n6263), .Z(n3422) );
  MUX2_X1 U3544 ( .A(n5719), .B(DATAIN[24]), .S(n6264), .Z(n3423) );
  MUX2_X1 U3545 ( .A(n5718), .B(DATAIN[25]), .S(n6264), .Z(n3424) );
  MUX2_X1 U3546 ( .A(n5717), .B(DATAIN[26]), .S(n6264), .Z(n3425) );
  MUX2_X1 U3547 ( .A(n5716), .B(DATAIN[27]), .S(n6264), .Z(n3426) );
  MUX2_X1 U3548 ( .A(n5715), .B(DATAIN[28]), .S(n6264), .Z(n3427) );
  MUX2_X1 U3549 ( .A(n5714), .B(DATAIN[29]), .S(n6264), .Z(n3428) );
  MUX2_X1 U3550 ( .A(n5713), .B(DATAIN[30]), .S(n6264), .Z(n3429) );
  MUX2_X1 U3551 ( .A(n5712), .B(DATAIN[31]), .S(n6264), .Z(n3430) );
endmodule


module Decode ( CLK, RST, REG_LATCH_EN, RD1, RD2, RF_WE, ZERO_FLAG, PC_IN, 
        INS_IN, ADD_WR, DATA_WR_IN, PC_OUT, A_OUT, B_OUT, IMM_OUT, ADD_RS1_HDU, 
        ADD_RS2_HDU, ADD_WR_OUT, ADD_RS1_OUT, ADD_RS2_OUT );
  input [31:0] PC_IN;
  input [31:0] INS_IN;
  input [4:0] ADD_WR;
  input [31:0] DATA_WR_IN;
  output [31:0] PC_OUT;
  output [31:0] A_OUT;
  output [31:0] B_OUT;
  output [31:0] IMM_OUT;
  output [4:0] ADD_RS1_HDU;
  output [4:0] ADD_RS2_HDU;
  output [4:0] ADD_WR_OUT;
  output [4:0] ADD_RS1_OUT;
  output [4:0] ADD_RS2_OUT;
  input CLK, RST, REG_LATCH_EN, RD1, RD2, RF_WE, ZERO_FLAG;
  wire   sig_RST, sig_Rtype, sig_Itype, sig_Jtype, n2;
  wire   [4:0] sig_ADD_WR;
  wire   [31:0] sig_IMM;

  instruction_type ins_type ( .INST_IN(INS_IN), .Rtype(sig_Rtype), .Itype(
        sig_Itype), .Jtype(sig_Jtype) );
  instruction_decomposition ins_dec ( .INST_IN(INS_IN), .Rtype(sig_Rtype), 
        .Itype(sig_Itype), .Jtype(sig_Jtype), .ADD_RS1(ADD_RS1_HDU), .ADD_RS2(
        ADD_RS2_HDU), .ADD_WR(sig_ADD_WR), .IMM(sig_IMM) );
  regn_N32_8 regPC ( .DIN(PC_IN), .CLK(CLK), .EN(1'b1), .RST(sig_RST), .DOUT(
        PC_OUT) );
  regn_N32_7 regIMM ( .DIN(sig_IMM), .CLK(CLK), .EN(REG_LATCH_EN), .RST(
        sig_RST), .DOUT(IMM_OUT) );
  regn_N5_0 regWR ( .DIN(sig_ADD_WR), .CLK(CLK), .EN(REG_LATCH_EN), .RST(
        sig_RST), .DOUT(ADD_WR_OUT) );
  regn_N5_4 regRS1 ( .DIN(ADD_RS1_HDU), .CLK(CLK), .EN(REG_LATCH_EN), .RST(
        sig_RST), .DOUT(ADD_RS1_OUT) );
  regn_N5_3 regRS2 ( .DIN(ADD_RS2_HDU), .CLK(CLK), .EN(REG_LATCH_EN), .RST(
        sig_RST), .DOUT(ADD_RS2_OUT) );
  register_file_NBIT_ADD5_NBIT_DATA32 rf ( .CLK(CLK), .RST(RST), .ENABLE(
        REG_LATCH_EN), .RD1(RD1), .RD2(RD2), .WR(RF_WE), .ADD_WR(ADD_WR), 
        .ADD_RS1(ADD_RS1_HDU), .ADD_RS2(ADD_RS2_HDU), .DATAIN(DATA_WR_IN), 
        .OUT1(A_OUT), .OUT2(B_OUT) );
  NOR2_X1 U2 ( .A1(ZERO_FLAG), .A2(n2), .ZN(sig_RST) );
  INV_X1 U3 ( .A(RST), .ZN(n2) );
endmodule


module Branch_Cond_Unit_NBIT32 ( RST, A, .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , 
        \ALU_OPC[1] , \ALU_OPC[0] }), JUMP_TYPE, PC_SEL, ZERO );
  input [31:0] A;
  input [1:0] JUMP_TYPE;
  output [1:0] PC_SEL;
  input RST, \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] ;
  output ZERO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [3:0] ALU_OPC;

  NAND2_X1 U3 ( .A1(n2), .A2(n3), .ZN(ZERO) );
  NOR4_X1 U4 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n12) );
  NOR4_X1 U5 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n16) );
  NAND4_X1 U6 ( .A1(ALU_OPC[3]), .A2(RST), .A3(JUMP_TYPE[0]), .A4(n4), .ZN(n2)
         );
  NOR3_X1 U7 ( .A1(n5), .A2(ALU_OPC[2]), .A3(ALU_OPC[1]), .ZN(n4) );
  XNOR2_X1 U8 ( .A(ALU_OPC[0]), .B(n6), .ZN(n5) );
  NOR2_X1 U9 ( .A1(n7), .A2(n8), .ZN(n6) );
  NAND4_X1 U10 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n8) );
  NOR4_X1 U11 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n9) );
  NOR4_X1 U12 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n10) );
  NOR4_X1 U13 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n11) );
  NAND4_X1 U14 ( .A1(n13), .A2(n14), .A3(n15), .A4(n16), .ZN(n7) );
  NOR4_X1 U15 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n13) );
  NOR4_X1 U16 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n14) );
  NOR4_X1 U17 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n15) );
  NAND2_X1 U18 ( .A1(RST), .A2(JUMP_TYPE[1]), .ZN(n3) );
  OAI22_X1 U19 ( .A1(JUMP_TYPE[1]), .A2(n2), .B1(JUMP_TYPE[0]), .B2(n3), .ZN(
        PC_SEL[0]) );
  NOR2_X1 U20 ( .A1(n17), .A2(n3), .ZN(PC_SEL[1]) );
  INV_X1 U21 ( .A(JUMP_TYPE[0]), .ZN(n17) );
endmodule


module regn_N2 ( DIN, CLK, EN, RST, DOUT );
  input [1:0] DIN;
  output [1:0] DOUT;
  input CLK, EN, RST;
  wire   n3, n4, n5, n6, n1, n2;

  DFFR_X1 \DOUT_reg[1]  ( .D(n6), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n4) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n5), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n3) );
  OAI21_X1 U2 ( .B1(n3), .B2(EN), .A(n2), .ZN(n5) );
  NAND2_X1 U3 ( .A1(DIN[0]), .A2(EN), .ZN(n2) );
  OAI21_X1 U4 ( .B1(n4), .B2(EN), .A(n1), .ZN(n6) );
  NAND2_X1 U5 ( .A1(EN), .A2(DIN[1]), .ZN(n1) );
endmodule


module FWD_Unit ( RST, ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB, RF_WE_MEM, 
        RF_WE_WB, FWDA, FWDB );
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [4:0] ADD_WR_MEM;
  input [4:0] ADD_WR_WB;
  output [1:0] FWDA;
  output [1:0] FWDB;
  input RST, RF_WE_MEM, RF_WE_WB;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n43, n44, n45, n46;

  XOR2_X1 U38 ( .A(ADD_WR_WB[4]), .B(ADD_RS2[4]), .Z(n13) );
  XOR2_X1 U39 ( .A(ADD_WR_WB[0]), .B(ADD_RS2[0]), .Z(n12) );
  XOR2_X1 U40 ( .A(ADD_WR_MEM[4]), .B(ADD_RS2[4]), .Z(n19) );
  XOR2_X1 U41 ( .A(ADD_WR_MEM[3]), .B(ADD_RS2[3]), .Z(n18) );
  XOR2_X1 U42 ( .A(ADD_WR_WB[1]), .B(ADD_RS1[1]), .Z(n33) );
  XOR2_X1 U43 ( .A(ADD_WR_WB[0]), .B(ADD_RS1[0]), .Z(n32) );
  XOR2_X1 U44 ( .A(ADD_WR_MEM[4]), .B(ADD_RS1[4]), .Z(n39) );
  XOR2_X1 U45 ( .A(ADD_WR_MEM[3]), .B(ADD_RS1[3]), .Z(n38) );
  OAI22_X1 U3 ( .A1(n46), .A2(n6), .B1(n5), .B2(n7), .ZN(FWDB[0]) );
  INV_X1 U4 ( .A(n5), .ZN(n46) );
  OAI22_X1 U5 ( .A1(n45), .A2(n21), .B1(n20), .B2(n7), .ZN(FWDA[0]) );
  INV_X1 U6 ( .A(n20), .ZN(n45) );
  OAI22_X1 U7 ( .A1(n44), .A2(n5), .B1(n43), .B2(n6), .ZN(FWDB[1]) );
  OAI22_X1 U8 ( .A1(n44), .A2(n20), .B1(n43), .B2(n21), .ZN(FWDA[1]) );
  INV_X1 U9 ( .A(RST), .ZN(n44) );
  NOR3_X1 U10 ( .A1(n12), .A2(n44), .A3(n13), .ZN(n11) );
  NOR3_X1 U11 ( .A1(n32), .A2(n44), .A3(n33), .ZN(n31) );
  NAND4_X1 U12 ( .A1(n14), .A2(n15), .A3(n16), .A4(n17), .ZN(n5) );
  NOR2_X1 U13 ( .A1(n18), .A2(n19), .ZN(n17) );
  XNOR2_X1 U14 ( .A(ADD_RS2[0]), .B(ADD_WR_MEM[0]), .ZN(n14) );
  XNOR2_X1 U15 ( .A(ADD_RS2[1]), .B(ADD_WR_MEM[1]), .ZN(n15) );
  NAND4_X1 U16 ( .A1(n34), .A2(n35), .A3(n36), .A4(n37), .ZN(n20) );
  NOR2_X1 U17 ( .A1(n38), .A2(n39), .ZN(n37) );
  XNOR2_X1 U18 ( .A(ADD_RS1[0]), .B(ADD_WR_MEM[0]), .ZN(n34) );
  XNOR2_X1 U19 ( .A(ADD_RS1[1]), .B(ADD_WR_MEM[1]), .ZN(n35) );
  NAND4_X1 U20 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .ZN(n6) );
  XNOR2_X1 U21 ( .A(ADD_RS2[3]), .B(ADD_WR_WB[3]), .ZN(n8) );
  XNOR2_X1 U22 ( .A(ADD_RS2[1]), .B(ADD_WR_WB[1]), .ZN(n9) );
  XNOR2_X1 U23 ( .A(ADD_RS2[2]), .B(ADD_WR_WB[2]), .ZN(n10) );
  NAND4_X1 U24 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n21) );
  XNOR2_X1 U25 ( .A(ADD_RS1[4]), .B(ADD_WR_WB[4]), .ZN(n28) );
  XNOR2_X1 U26 ( .A(ADD_RS1[3]), .B(ADD_WR_WB[3]), .ZN(n29) );
  XNOR2_X1 U27 ( .A(ADD_RS1[2]), .B(ADD_WR_WB[2]), .ZN(n30) );
  XNOR2_X1 U28 ( .A(ADD_RS2[2]), .B(ADD_WR_MEM[2]), .ZN(n16) );
  XNOR2_X1 U29 ( .A(ADD_RS1[2]), .B(ADD_WR_MEM[2]), .ZN(n36) );
  NAND2_X1 U30 ( .A1(RST), .A2(n25), .ZN(n7) );
  OAI21_X1 U31 ( .B1(n26), .B2(n27), .A(RF_WE_MEM), .ZN(n25) );
  OR2_X1 U32 ( .A1(ADD_WR_MEM[0]), .A2(ADD_WR_MEM[1]), .ZN(n27) );
  OR3_X1 U33 ( .A1(ADD_WR_MEM[3]), .A2(ADD_WR_MEM[4]), .A3(ADD_WR_MEM[2]), 
        .ZN(n26) );
  INV_X1 U34 ( .A(n22), .ZN(n43) );
  OAI21_X1 U35 ( .B1(n23), .B2(n24), .A(RF_WE_WB), .ZN(n22) );
  OR2_X1 U36 ( .A1(ADD_WR_WB[0]), .A2(ADD_WR_WB[1]), .ZN(n24) );
  OR3_X1 U37 ( .A1(ADD_WR_WB[3]), .A2(ADD_WR_WB[4]), .A3(ADD_WR_WB[2]), .ZN(
        n23) );
endmodule


module comparator_NBIT32_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267;

  XOR2_X1 U103 ( .A(A[30]), .B(n208), .Z(n70) );
  NAND3_X1 U172 ( .A1(n197), .A2(n150), .A3(n147), .ZN(n196) );
  NAND3_X1 U176 ( .A1(n234), .A2(n199), .A3(n200), .ZN(n197) );
  INV_X1 U1 ( .A(n142), .ZN(n232) );
  INV_X1 U2 ( .A(n130), .ZN(n228) );
  INV_X1 U3 ( .A(n118), .ZN(n224) );
  INV_X1 U4 ( .A(n106), .ZN(n220) );
  INV_X1 U5 ( .A(n94), .ZN(n216) );
  INV_X1 U6 ( .A(n82), .ZN(n212) );
  NOR2_X1 U7 ( .A1(n193), .A2(n136), .ZN(n135) );
  NOR2_X1 U8 ( .A1(n187), .A2(n124), .ZN(n123) );
  NOR2_X1 U9 ( .A1(n181), .A2(n112), .ZN(n111) );
  NOR2_X1 U10 ( .A1(n175), .A2(n100), .ZN(n99) );
  NOR2_X1 U11 ( .A1(n169), .A2(n88), .ZN(n87) );
  NOR2_X1 U12 ( .A1(n163), .A2(n76), .ZN(n75) );
  OAI211_X1 U13 ( .C1(n161), .C2(n162), .A(n78), .B(n75), .ZN(n160) );
  NAND2_X1 U14 ( .A1(n210), .A2(n164), .ZN(n162) );
  AOI211_X1 U15 ( .C1(n165), .C2(n166), .A(n82), .B(n213), .ZN(n161) );
  INV_X1 U16 ( .A(n79), .ZN(n210) );
  OAI211_X1 U17 ( .C1(n191), .C2(n192), .A(n138), .B(n135), .ZN(n190) );
  NAND2_X1 U18 ( .A1(n230), .A2(n194), .ZN(n192) );
  AOI211_X1 U19 ( .C1(n195), .C2(n196), .A(n142), .B(n233), .ZN(n191) );
  INV_X1 U20 ( .A(n139), .ZN(n230) );
  OAI211_X1 U21 ( .C1(n185), .C2(n186), .A(n126), .B(n123), .ZN(n184) );
  NAND2_X1 U22 ( .A1(n226), .A2(n188), .ZN(n186) );
  AOI211_X1 U23 ( .C1(n189), .C2(n190), .A(n130), .B(n229), .ZN(n185) );
  INV_X1 U24 ( .A(n127), .ZN(n226) );
  OAI211_X1 U25 ( .C1(n179), .C2(n180), .A(n114), .B(n111), .ZN(n178) );
  NAND2_X1 U26 ( .A1(n222), .A2(n182), .ZN(n180) );
  AOI211_X1 U27 ( .C1(n183), .C2(n184), .A(n118), .B(n225), .ZN(n179) );
  INV_X1 U28 ( .A(n115), .ZN(n222) );
  OAI211_X1 U29 ( .C1(n173), .C2(n174), .A(n102), .B(n99), .ZN(n172) );
  NAND2_X1 U30 ( .A1(n218), .A2(n176), .ZN(n174) );
  AOI211_X1 U31 ( .C1(n177), .C2(n178), .A(n106), .B(n221), .ZN(n173) );
  INV_X1 U32 ( .A(n103), .ZN(n218) );
  OAI211_X1 U33 ( .C1(n167), .C2(n168), .A(n90), .B(n87), .ZN(n166) );
  NAND2_X1 U34 ( .A1(n214), .A2(n170), .ZN(n168) );
  AOI211_X1 U35 ( .C1(n171), .C2(n172), .A(n94), .B(n217), .ZN(n167) );
  INV_X1 U36 ( .A(n91), .ZN(n214) );
  AOI21_X1 U37 ( .B1(n143), .B2(n144), .A(n145), .ZN(n140) );
  AOI21_X1 U38 ( .B1(n146), .B2(n147), .A(n148), .ZN(n143) );
  AOI21_X1 U39 ( .B1(n149), .B2(n150), .A(n151), .ZN(n146) );
  AOI21_X1 U40 ( .B1(n152), .B2(n153), .A(n235), .ZN(n149) );
  AOI21_X1 U41 ( .B1(n131), .B2(n132), .A(n133), .ZN(n128) );
  AOI21_X1 U42 ( .B1(n134), .B2(n135), .A(n136), .ZN(n131) );
  AOI21_X1 U43 ( .B1(n137), .B2(n138), .A(n139), .ZN(n134) );
  AOI21_X1 U44 ( .B1(n140), .B2(n232), .A(n231), .ZN(n137) );
  AOI21_X1 U45 ( .B1(n119), .B2(n120), .A(n121), .ZN(n116) );
  AOI21_X1 U46 ( .B1(n122), .B2(n123), .A(n124), .ZN(n119) );
  AOI21_X1 U47 ( .B1(n125), .B2(n126), .A(n127), .ZN(n122) );
  AOI21_X1 U48 ( .B1(n128), .B2(n228), .A(n227), .ZN(n125) );
  AOI21_X1 U49 ( .B1(n107), .B2(n108), .A(n109), .ZN(n104) );
  AOI21_X1 U50 ( .B1(n110), .B2(n111), .A(n112), .ZN(n107) );
  AOI21_X1 U51 ( .B1(n113), .B2(n114), .A(n115), .ZN(n110) );
  AOI21_X1 U52 ( .B1(n116), .B2(n224), .A(n223), .ZN(n113) );
  AOI21_X1 U53 ( .B1(n95), .B2(n96), .A(n97), .ZN(n92) );
  AOI21_X1 U54 ( .B1(n98), .B2(n99), .A(n100), .ZN(n95) );
  AOI21_X1 U55 ( .B1(n101), .B2(n102), .A(n103), .ZN(n98) );
  AOI21_X1 U56 ( .B1(n104), .B2(n220), .A(n219), .ZN(n101) );
  AOI21_X1 U57 ( .B1(n83), .B2(n84), .A(n85), .ZN(n80) );
  AOI21_X1 U58 ( .B1(n86), .B2(n87), .A(n88), .ZN(n83) );
  AOI21_X1 U59 ( .B1(n89), .B2(n90), .A(n91), .ZN(n86) );
  AOI21_X1 U60 ( .B1(n92), .B2(n216), .A(n215), .ZN(n89) );
  AOI21_X1 U61 ( .B1(n71), .B2(n72), .A(n73), .ZN(n69) );
  AOI21_X1 U62 ( .B1(n74), .B2(n75), .A(n76), .ZN(n71) );
  AOI21_X1 U63 ( .B1(n77), .B2(n78), .A(n79), .ZN(n74) );
  AOI21_X1 U64 ( .B1(n80), .B2(n212), .A(n211), .ZN(n77) );
  NOR2_X1 U65 ( .A1(n198), .A2(n148), .ZN(n147) );
  NOR2_X1 U66 ( .A1(n198), .A2(n145), .ZN(n195) );
  NOR2_X1 U67 ( .A1(n193), .A2(n133), .ZN(n189) );
  NOR2_X1 U68 ( .A1(n187), .A2(n121), .ZN(n183) );
  NOR2_X1 U69 ( .A1(n181), .A2(n109), .ZN(n177) );
  NOR2_X1 U70 ( .A1(n175), .A2(n97), .ZN(n171) );
  NOR2_X1 U71 ( .A1(n169), .A2(n85), .ZN(n165) );
  NOR2_X1 U72 ( .A1(n163), .A2(n73), .ZN(n159) );
  NAND2_X1 U73 ( .A1(n194), .A2(n141), .ZN(n142) );
  NAND2_X1 U74 ( .A1(n188), .A2(n129), .ZN(n130) );
  NAND2_X1 U75 ( .A1(n182), .A2(n117), .ZN(n118) );
  NAND2_X1 U76 ( .A1(n176), .A2(n105), .ZN(n106) );
  NAND2_X1 U77 ( .A1(n170), .A2(n93), .ZN(n94) );
  NAND2_X1 U78 ( .A1(n164), .A2(n81), .ZN(n82) );
  AND2_X1 U79 ( .A1(n199), .A2(n154), .ZN(n153) );
  INV_X1 U80 ( .A(GT), .ZN(LE) );
  INV_X1 U81 ( .A(n108), .ZN(n221) );
  INV_X1 U82 ( .A(n96), .ZN(n217) );
  INV_X1 U83 ( .A(n84), .ZN(n213) );
  INV_X1 U84 ( .A(n144), .ZN(n233) );
  INV_X1 U85 ( .A(n132), .ZN(n229) );
  INV_X1 U86 ( .A(n120), .ZN(n225) );
  INV_X1 U87 ( .A(n141), .ZN(n231) );
  INV_X1 U88 ( .A(n129), .ZN(n227) );
  INV_X1 U89 ( .A(n117), .ZN(n223) );
  INV_X1 U90 ( .A(n105), .ZN(n219) );
  INV_X1 U91 ( .A(n93), .ZN(n215) );
  INV_X1 U92 ( .A(n81), .ZN(n211) );
  INV_X1 U93 ( .A(n154), .ZN(n235) );
  AOI21_X1 U94 ( .B1(n66), .B2(n207), .A(n67), .ZN(GE) );
  INV_X1 U95 ( .A(n68), .ZN(n207) );
  AOI22_X1 U96 ( .A1(B[30]), .A2(n238), .B1(n69), .B2(n70), .ZN(n68) );
  INV_X1 U97 ( .A(A[30]), .ZN(n238) );
  OAI21_X1 U98 ( .B1(n67), .B2(n157), .A(n66), .ZN(GT) );
  AOI22_X1 U99 ( .A1(A[30]), .A2(n208), .B1(n158), .B2(n70), .ZN(n157) );
  AOI21_X1 U100 ( .B1(n159), .B2(n160), .A(n209), .ZN(n158) );
  INV_X1 U101 ( .A(n72), .ZN(n209) );
  INV_X1 U102 ( .A(GE), .ZN(LT) );
  AOI22_X1 U104 ( .A1(n155), .A2(n237), .B1(A[1]), .B2(n156), .ZN(n152) );
  OR2_X1 U105 ( .A1(n156), .A2(A[1]), .ZN(n155) );
  NAND2_X1 U106 ( .A1(B[0]), .A2(n267), .ZN(n156) );
  NOR2_X1 U107 ( .A1(n267), .A2(B[0]), .ZN(n201) );
  NOR2_X1 U108 ( .A1(n264), .A2(B[4]), .ZN(n198) );
  NOR2_X1 U109 ( .A1(n260), .A2(B[8]), .ZN(n193) );
  NOR2_X1 U110 ( .A1(n256), .A2(B[12]), .ZN(n187) );
  NOR2_X1 U111 ( .A1(n252), .A2(B[16]), .ZN(n181) );
  NOR2_X1 U112 ( .A1(n248), .A2(B[20]), .ZN(n175) );
  NOR2_X1 U113 ( .A1(n244), .A2(B[24]), .ZN(n169) );
  NOR2_X1 U114 ( .A1(n240), .A2(B[28]), .ZN(n163) );
  NOR2_X1 U115 ( .A1(n263), .A2(B[5]), .ZN(n145) );
  NOR2_X1 U116 ( .A1(n259), .A2(B[9]), .ZN(n133) );
  NOR2_X1 U117 ( .A1(n255), .A2(B[13]), .ZN(n121) );
  NOR2_X1 U118 ( .A1(n251), .A2(B[17]), .ZN(n109) );
  NOR2_X1 U119 ( .A1(n247), .A2(B[21]), .ZN(n97) );
  NOR2_X1 U120 ( .A1(n243), .A2(B[25]), .ZN(n85) );
  NOR2_X1 U121 ( .A1(n239), .A2(B[29]), .ZN(n73) );
  NOR2_X1 U122 ( .A1(n265), .A2(B[3]), .ZN(n151) );
  NOR2_X1 U123 ( .A1(n261), .A2(B[7]), .ZN(n139) );
  NOR2_X1 U124 ( .A1(n257), .A2(B[11]), .ZN(n127) );
  NOR2_X1 U125 ( .A1(n253), .A2(B[15]), .ZN(n115) );
  NOR2_X1 U126 ( .A1(n249), .A2(B[19]), .ZN(n103) );
  NOR2_X1 U127 ( .A1(n245), .A2(B[23]), .ZN(n91) );
  NOR2_X1 U128 ( .A1(n241), .A2(B[27]), .ZN(n79) );
  NOR2_X1 U129 ( .A1(n206), .A2(A[31]), .ZN(n67) );
  INV_X1 U130 ( .A(NE), .ZN(EQ) );
  NAND2_X1 U131 ( .A1(LE), .A2(GE), .ZN(NE) );
  INV_X1 U132 ( .A(n151), .ZN(n234) );
  OAI211_X1 U133 ( .C1(A[1]), .C2(n201), .A(n236), .B(n153), .ZN(n200) );
  NAND2_X1 U134 ( .A1(B[7]), .A2(n261), .ZN(n138) );
  NAND2_X1 U135 ( .A1(B[11]), .A2(n257), .ZN(n126) );
  NAND2_X1 U136 ( .A1(B[15]), .A2(n253), .ZN(n114) );
  NAND2_X1 U137 ( .A1(B[19]), .A2(n249), .ZN(n102) );
  NAND2_X1 U138 ( .A1(B[23]), .A2(n245), .ZN(n90) );
  NAND2_X1 U139 ( .A1(B[27]), .A2(n241), .ZN(n78) );
  NAND2_X1 U140 ( .A1(B[5]), .A2(n263), .ZN(n144) );
  NAND2_X1 U141 ( .A1(B[9]), .A2(n259), .ZN(n132) );
  NAND2_X1 U142 ( .A1(B[13]), .A2(n255), .ZN(n120) );
  NAND2_X1 U143 ( .A1(B[17]), .A2(n251), .ZN(n108) );
  NAND2_X1 U144 ( .A1(B[21]), .A2(n247), .ZN(n96) );
  NAND2_X1 U145 ( .A1(B[25]), .A2(n243), .ZN(n84) );
  NAND2_X1 U146 ( .A1(B[29]), .A2(n239), .ZN(n72) );
  NAND2_X1 U147 ( .A1(B[6]), .A2(n262), .ZN(n141) );
  NAND2_X1 U148 ( .A1(B[10]), .A2(n258), .ZN(n129) );
  NAND2_X1 U149 ( .A1(B[14]), .A2(n254), .ZN(n117) );
  NAND2_X1 U150 ( .A1(B[18]), .A2(n250), .ZN(n105) );
  NAND2_X1 U151 ( .A1(B[22]), .A2(n246), .ZN(n93) );
  NAND2_X1 U152 ( .A1(B[26]), .A2(n242), .ZN(n81) );
  NAND2_X1 U153 ( .A1(A[31]), .A2(n206), .ZN(n66) );
  AND2_X1 U154 ( .A1(B[4]), .A2(n264), .ZN(n148) );
  AND2_X1 U155 ( .A1(B[8]), .A2(n260), .ZN(n136) );
  AND2_X1 U156 ( .A1(B[12]), .A2(n256), .ZN(n124) );
  AND2_X1 U157 ( .A1(B[16]), .A2(n252), .ZN(n112) );
  AND2_X1 U158 ( .A1(B[20]), .A2(n248), .ZN(n100) );
  AND2_X1 U159 ( .A1(B[24]), .A2(n244), .ZN(n88) );
  AND2_X1 U160 ( .A1(B[28]), .A2(n240), .ZN(n76) );
  NAND2_X1 U161 ( .A1(B[3]), .A2(n265), .ZN(n150) );
  NAND2_X1 U162 ( .A1(B[2]), .A2(n266), .ZN(n154) );
  INV_X1 U163 ( .A(A[0]), .ZN(n267) );
  INV_X1 U164 ( .A(A[3]), .ZN(n265) );
  INV_X1 U165 ( .A(A[5]), .ZN(n263) );
  INV_X1 U166 ( .A(A[7]), .ZN(n261) );
  INV_X1 U167 ( .A(A[9]), .ZN(n259) );
  INV_X1 U168 ( .A(A[11]), .ZN(n257) );
  INV_X1 U169 ( .A(A[13]), .ZN(n255) );
  INV_X1 U170 ( .A(A[15]), .ZN(n253) );
  INV_X1 U171 ( .A(A[17]), .ZN(n251) );
  INV_X1 U173 ( .A(A[19]), .ZN(n249) );
  INV_X1 U174 ( .A(A[21]), .ZN(n247) );
  INV_X1 U175 ( .A(A[23]), .ZN(n245) );
  INV_X1 U177 ( .A(A[25]), .ZN(n243) );
  INV_X1 U178 ( .A(A[29]), .ZN(n239) );
  INV_X1 U179 ( .A(A[27]), .ZN(n241) );
  INV_X1 U180 ( .A(B[31]), .ZN(n206) );
  INV_X1 U181 ( .A(B[1]), .ZN(n237) );
  OR2_X1 U182 ( .A1(n262), .A2(B[6]), .ZN(n194) );
  OR2_X1 U183 ( .A1(n258), .A2(B[10]), .ZN(n188) );
  OR2_X1 U184 ( .A1(n254), .A2(B[14]), .ZN(n182) );
  OR2_X1 U185 ( .A1(n250), .A2(B[18]), .ZN(n176) );
  OR2_X1 U186 ( .A1(n246), .A2(B[22]), .ZN(n170) );
  OR2_X1 U187 ( .A1(n242), .A2(B[26]), .ZN(n164) );
  INV_X1 U188 ( .A(B[30]), .ZN(n208) );
  INV_X1 U189 ( .A(A[2]), .ZN(n266) );
  INV_X1 U190 ( .A(A[6]), .ZN(n262) );
  INV_X1 U191 ( .A(A[10]), .ZN(n258) );
  INV_X1 U192 ( .A(A[14]), .ZN(n254) );
  INV_X1 U193 ( .A(A[18]), .ZN(n250) );
  INV_X1 U194 ( .A(A[22]), .ZN(n246) );
  INV_X1 U195 ( .A(A[26]), .ZN(n242) );
  INV_X1 U196 ( .A(A[4]), .ZN(n264) );
  INV_X1 U197 ( .A(A[8]), .ZN(n260) );
  INV_X1 U198 ( .A(A[12]), .ZN(n256) );
  INV_X1 U199 ( .A(A[16]), .ZN(n252) );
  INV_X1 U200 ( .A(A[20]), .ZN(n248) );
  INV_X1 U201 ( .A(A[24]), .ZN(n244) );
  INV_X1 U202 ( .A(A[28]), .ZN(n240) );
  OR2_X1 U203 ( .A1(n266), .A2(B[2]), .ZN(n199) );
  INV_X1 U204 ( .A(n202), .ZN(n236) );
  AOI21_X1 U205 ( .B1(A[1]), .B2(n201), .A(n237), .ZN(n202) );
endmodule


module comparator_NBIT32 ( A, B, .OPSel({\OPSel[2] , \OPSel[1] , \OPSel[0] }), 
        RES );
  input [31:0] A;
  input [31:0] B;
  output [31:0] RES;
  input \OPSel[2] , \OPSel[1] , \OPSel[0] ;
  wire   N26, N27, N28, N29, N30, N31, n6, n7, n8, n9, n11, n12, n10, n13, n14
;
  wire   [2:0] OPSel;
  assign RES[1] = 1'b0;
  assign RES[2] = 1'b0;
  assign RES[3] = 1'b0;
  assign RES[4] = 1'b0;
  assign RES[5] = 1'b0;
  assign RES[6] = 1'b0;
  assign RES[7] = 1'b0;
  assign RES[8] = 1'b0;
  assign RES[9] = 1'b0;
  assign RES[10] = 1'b0;
  assign RES[11] = 1'b0;
  assign RES[12] = 1'b0;
  assign RES[13] = 1'b0;
  assign RES[14] = 1'b0;
  assign RES[15] = 1'b0;
  assign RES[16] = 1'b0;
  assign RES[17] = 1'b0;
  assign RES[18] = 1'b0;
  assign RES[19] = 1'b0;
  assign RES[20] = 1'b0;
  assign RES[21] = 1'b0;
  assign RES[22] = 1'b0;
  assign RES[23] = 1'b0;
  assign RES[24] = 1'b0;
  assign RES[25] = 1'b0;
  assign RES[26] = 1'b0;
  assign RES[27] = 1'b0;
  assign RES[28] = 1'b0;
  assign RES[29] = 1'b0;
  assign RES[30] = 1'b0;
  assign RES[31] = 1'b0;

  comparator_NBIT32_DW01_cmp6_0 r57 ( .A(A), .B(B), .TC(1'b0), .LT(N30), .GT(
        N28), .EQ(N26), .LE(N31), .GE(N29), .NE(N27) );
  AOI22_X1 U2 ( .A1(N30), .A2(n14), .B1(OPSel[0]), .B2(N31), .ZN(n9) );
  AOI22_X1 U4 ( .A1(N26), .A2(n14), .B1(N27), .B2(OPSel[0]), .ZN(n12) );
  AOI22_X1 U5 ( .A1(N28), .A2(n14), .B1(N29), .B2(OPSel[0]), .ZN(n11) );
  INV_X1 U6 ( .A(OPSel[2]), .ZN(n10) );
  INV_X1 U7 ( .A(OPSel[1]), .ZN(n13) );
  INV_X1 U8 ( .A(n6), .ZN(RES[0]) );
  AOI21_X1 U9 ( .B1(n7), .B2(n10), .A(n8), .ZN(n6) );
  NOR3_X1 U10 ( .A1(n10), .A2(OPSel[1]), .A3(n9), .ZN(n8) );
  OAI22_X1 U11 ( .A1(n11), .A2(n13), .B1(OPSel[1]), .B2(n12), .ZN(n7) );
  INV_X1 U12 ( .A(OPSel[0]), .ZN(n14) );
endmodule


module carry_generator_NBIT32_NBIT_PER_BLOCK4 ( A, B, Cin, Co );
  input [32:1] A;
  input [32:1] B;
  output [7:0] Co;
  input Cin;
  wire   \G[1][1] , n3, \P[9][9] , \P[8][8] , \P[8][7] , \P[8][5] , \P[7][7] ,
         \P[6][6] , \P[6][5] , \P[5][5] , \P[4][4] , \P[4][3] , \P[3][3] ,
         \P[32][32] , \P[32][31] , \P[32][29] , \P[32][25] , \P[32][17] ,
         \P[31][31] , \P[30][30] , \P[30][29] , \P[2][2] , \P[29][29] ,
         \P[28][28] , \P[28][27] , \P[28][25] , \P[28][17] , \P[27][27] ,
         \P[26][26] , \P[26][25] , \P[25][25] , \P[24][24] , \P[24][23] ,
         \P[24][21] , \P[24][17] , \P[23][23] , \P[22][22] , \P[22][21] ,
         \P[21][21] , \P[20][20] , \P[20][19] , \P[20][17] , \P[19][19] ,
         \P[18][18] , \P[18][17] , \P[17][17] , \P[16][9] , \P[16][16] ,
         \P[16][15] , \P[16][13] , \P[15][15] , \P[14][14] , \P[14][13] ,
         \P[13][13] , \P[12][9] , \P[12][12] , \P[12][11] , \P[11][11] ,
         \P[10][9] , \P[10][10] , \G[9][9] , \G[8][8] , \G[8][7] , \G[8][5] ,
         \G[7][7] , \G[6][6] , \G[6][5] , \G[5][5] , \G[4][4] , \G[4][3] ,
         \G[3][3] , \G[32][32] , \G[32][31] , \G[32][29] , \G[32][25] ,
         \G[32][17] , \G[31][31] , \G[30][30] , \G[30][29] , \G[2][2] ,
         \G[2][1] , \G[29][29] , \G[28][28] , \G[28][27] , \G[28][25] ,
         \G[28][17] , \G[27][27] , \G[26][26] , \G[26][25] , \G[25][25] ,
         \G[24][24] , \G[24][23] , \G[24][21] , \G[24][17] , \G[23][23] ,
         \G[22][22] , \G[22][21] , \G[21][21] , \G[20][20] , \G[20][19] ,
         \G[20][17] , \G[19][19] , \G[18][18] , \G[18][17] , \G[17][17] ,
         \G[16][9] , \G[16][16] , \G[16][15] , \G[16][13] , \G[15][15] ,
         \G[14][14] , \G[14][13] , \G[13][13] , \G[12][9] , \G[12][12] ,
         \G[12][11] , \G[11][11] , \G[10][9] , \G[10][10] , n4, n5;

  PG_net_0 PGnetblock_2 ( .a(A[2]), .b(B[2]), .p(\P[2][2] ), .g(\G[2][2] ) );
  PG_net_30 PGnetblock_3 ( .a(A[3]), .b(B[3]), .p(\P[3][3] ), .g(\G[3][3] ) );
  PG_net_29 PGnetblock_4 ( .a(A[4]), .b(B[4]), .p(\P[4][4] ), .g(\G[4][4] ) );
  PG_net_28 PGnetblock_5 ( .a(A[5]), .b(B[5]), .p(\P[5][5] ), .g(\G[5][5] ) );
  PG_net_27 PGnetblock_6 ( .a(A[6]), .b(B[6]), .p(\P[6][6] ), .g(\G[6][6] ) );
  PG_net_26 PGnetblock_7 ( .a(A[7]), .b(B[7]), .p(\P[7][7] ), .g(\G[7][7] ) );
  PG_net_25 PGnetblock_8 ( .a(A[8]), .b(B[8]), .p(\P[8][8] ), .g(\G[8][8] ) );
  PG_net_24 PGnetblock_9 ( .a(A[9]), .b(B[9]), .p(\P[9][9] ), .g(\G[9][9] ) );
  PG_net_23 PGnetblock_10 ( .a(A[10]), .b(B[10]), .p(\P[10][10] ), .g(
        \G[10][10] ) );
  PG_net_22 PGnetblock_11 ( .a(A[11]), .b(B[11]), .p(\P[11][11] ), .g(
        \G[11][11] ) );
  PG_net_21 PGnetblock_12 ( .a(A[12]), .b(B[12]), .p(\P[12][12] ), .g(
        \G[12][12] ) );
  PG_net_20 PGnetblock_13 ( .a(A[13]), .b(B[13]), .p(\P[13][13] ), .g(
        \G[13][13] ) );
  PG_net_19 PGnetblock_14 ( .a(A[14]), .b(B[14]), .p(\P[14][14] ), .g(
        \G[14][14] ) );
  PG_net_18 PGnetblock_15 ( .a(A[15]), .b(B[15]), .p(\P[15][15] ), .g(
        \G[15][15] ) );
  PG_net_17 PGnetblock_16 ( .a(A[16]), .b(B[16]), .p(\P[16][16] ), .g(
        \G[16][16] ) );
  PG_net_16 PGnetblock_17 ( .a(A[17]), .b(B[17]), .p(\P[17][17] ), .g(
        \G[17][17] ) );
  PG_net_15 PGnetblock_18 ( .a(A[18]), .b(B[18]), .p(\P[18][18] ), .g(
        \G[18][18] ) );
  PG_net_14 PGnetblock_19 ( .a(A[19]), .b(B[19]), .p(\P[19][19] ), .g(
        \G[19][19] ) );
  PG_net_13 PGnetblock_20 ( .a(A[20]), .b(B[20]), .p(\P[20][20] ), .g(
        \G[20][20] ) );
  PG_net_12 PGnetblock_21 ( .a(A[21]), .b(B[21]), .p(\P[21][21] ), .g(
        \G[21][21] ) );
  PG_net_11 PGnetblock_22 ( .a(A[22]), .b(B[22]), .p(\P[22][22] ), .g(
        \G[22][22] ) );
  PG_net_10 PGnetblock_23 ( .a(A[23]), .b(B[23]), .p(\P[23][23] ), .g(
        \G[23][23] ) );
  PG_net_9 PGnetblock_24 ( .a(A[24]), .b(B[24]), .p(\P[24][24] ), .g(
        \G[24][24] ) );
  PG_net_8 PGnetblock_25 ( .a(A[25]), .b(B[25]), .p(\P[25][25] ), .g(
        \G[25][25] ) );
  PG_net_7 PGnetblock_26 ( .a(A[26]), .b(B[26]), .p(\P[26][26] ), .g(
        \G[26][26] ) );
  PG_net_6 PGnetblock_27 ( .a(A[27]), .b(B[27]), .p(\P[27][27] ), .g(
        \G[27][27] ) );
  PG_net_5 PGnetblock_28 ( .a(A[28]), .b(B[28]), .p(\P[28][28] ), .g(
        \G[28][28] ) );
  PG_net_4 PGnetblock_29 ( .a(A[29]), .b(B[29]), .p(\P[29][29] ), .g(
        \G[29][29] ) );
  PG_net_3 PGnetblock_30 ( .a(A[30]), .b(B[30]), .p(\P[30][30] ), .g(
        \G[30][30] ) );
  PG_net_2 PGnetblock_31 ( .a(A[31]), .b(B[31]), .p(\P[31][31] ), .g(
        \G[31][31] ) );
  PG_net_1 PGnetblock_32 ( .a(A[32]), .b(B[32]), .p(\P[32][32] ), .g(
        \G[32][32] ) );
  Gblock_0 GB_low_1_2 ( .Pik(\P[2][2] ), .Gik(\G[2][2] ), .Gk_1j(\G[1][1] ), 
        .Gij(\G[2][1] ) );
  Gblock_8 GB_low_2_4 ( .Pik(\P[4][3] ), .Gik(\G[4][3] ), .Gk_1j(\G[2][1] ), 
        .Gij(Co[0]) );
  Gblock_7 GB_low_3_8 ( .Pik(\P[8][5] ), .Gik(\G[8][5] ), .Gk_1j(Co[0]), .Gij(
        Co[1]) );
  Gblock_6 GB_high_4_16_0 ( .Pik(\P[16][9] ), .Gik(\G[16][9] ), .Gk_1j(Co[1]), 
        .Gij(Co[3]) );
  Gblock_5 GB_high_4_16_1 ( .Pik(\P[12][9] ), .Gik(\G[12][9] ), .Gk_1j(Co[1]), 
        .Gij(Co[2]) );
  Gblock_4 GB_high_5_32_0 ( .Pik(\P[32][17] ), .Gik(\G[32][17] ), .Gk_1j(Co[3]), .Gij(Co[7]) );
  Gblock_3 GB_high_5_32_1 ( .Pik(\P[28][17] ), .Gik(\G[28][17] ), .Gk_1j(Co[3]), .Gij(Co[6]) );
  Gblock_2 GB_high_5_32_2 ( .Pik(\P[24][17] ), .Gik(\G[24][17] ), .Gk_1j(Co[3]), .Gij(Co[5]) );
  Gblock_1 GB_high_5_32_3 ( .Pik(\P[20][17] ), .Gik(\G[20][17] ), .Gk_1j(Co[3]), .Gij(Co[4]) );
  PGblock_0 PGB_low_1_4 ( .Pik(\P[4][4] ), .Gik(\G[4][4] ), .Pk_1j(\P[3][3] ), 
        .Gk_1j(\G[3][3] ), .Pij(\P[4][3] ), .Gij(\G[4][3] ) );
  PGblock_26 PGB_low_1_6 ( .Pik(\P[6][6] ), .Gik(\G[6][6] ), .Pk_1j(\P[5][5] ), 
        .Gk_1j(\G[5][5] ), .Pij(\P[6][5] ), .Gij(\G[6][5] ) );
  PGblock_25 PGB_low_1_8 ( .Pik(\P[8][8] ), .Gik(\G[8][8] ), .Pk_1j(\P[7][7] ), 
        .Gk_1j(\G[7][7] ), .Pij(\P[8][7] ), .Gij(\G[8][7] ) );
  PGblock_24 PGB_low_1_10 ( .Pik(\P[10][10] ), .Gik(\G[10][10] ), .Pk_1j(
        \P[9][9] ), .Gk_1j(\G[9][9] ), .Pij(\P[10][9] ), .Gij(\G[10][9] ) );
  PGblock_23 PGB_low_1_12 ( .Pik(\P[12][12] ), .Gik(\G[12][12] ), .Pk_1j(
        \P[11][11] ), .Gk_1j(\G[11][11] ), .Pij(\P[12][11] ), .Gij(\G[12][11] ) );
  PGblock_22 PGB_low_1_14 ( .Pik(\P[14][14] ), .Gik(\G[14][14] ), .Pk_1j(
        \P[13][13] ), .Gk_1j(\G[13][13] ), .Pij(\P[14][13] ), .Gij(\G[14][13] ) );
  PGblock_21 PGB_low_1_16 ( .Pik(\P[16][16] ), .Gik(\G[16][16] ), .Pk_1j(
        \P[15][15] ), .Gk_1j(\G[15][15] ), .Pij(\P[16][15] ), .Gij(\G[16][15] ) );
  PGblock_20 PGB_low_1_18 ( .Pik(\P[18][18] ), .Gik(\G[18][18] ), .Pk_1j(
        \P[17][17] ), .Gk_1j(\G[17][17] ), .Pij(\P[18][17] ), .Gij(\G[18][17] ) );
  PGblock_19 PGB_low_1_20 ( .Pik(\P[20][20] ), .Gik(\G[20][20] ), .Pk_1j(
        \P[19][19] ), .Gk_1j(\G[19][19] ), .Pij(\P[20][19] ), .Gij(\G[20][19] ) );
  PGblock_18 PGB_low_1_22 ( .Pik(\P[22][22] ), .Gik(\G[22][22] ), .Pk_1j(
        \P[21][21] ), .Gk_1j(\G[21][21] ), .Pij(\P[22][21] ), .Gij(\G[22][21] ) );
  PGblock_17 PGB_low_1_24 ( .Pik(\P[24][24] ), .Gik(\G[24][24] ), .Pk_1j(
        \P[23][23] ), .Gk_1j(\G[23][23] ), .Pij(\P[24][23] ), .Gij(\G[24][23] ) );
  PGblock_16 PGB_low_1_26 ( .Pik(\P[26][26] ), .Gik(\G[26][26] ), .Pk_1j(
        \P[25][25] ), .Gk_1j(\G[25][25] ), .Pij(\P[26][25] ), .Gij(\G[26][25] ) );
  PGblock_15 PGB_low_1_28 ( .Pik(\P[28][28] ), .Gik(\G[28][28] ), .Pk_1j(
        \P[27][27] ), .Gk_1j(\G[27][27] ), .Pij(\P[28][27] ), .Gij(\G[28][27] ) );
  PGblock_14 PGB_low_1_30 ( .Pik(\P[30][30] ), .Gik(\G[30][30] ), .Pk_1j(
        \P[29][29] ), .Gk_1j(\G[29][29] ), .Pij(\P[30][29] ), .Gij(\G[30][29] ) );
  PGblock_13 PGB_low_1_32 ( .Pik(\P[32][32] ), .Gik(\G[32][32] ), .Pk_1j(
        \P[31][31] ), .Gk_1j(\G[31][31] ), .Pij(\P[32][31] ), .Gij(\G[32][31] ) );
  PGblock_12 PGB_low_2_8 ( .Pik(\P[8][7] ), .Gik(\G[8][7] ), .Pk_1j(\P[6][5] ), 
        .Gk_1j(\G[6][5] ), .Pij(\P[8][5] ), .Gij(\G[8][5] ) );
  PGblock_11 PGB_low_2_12 ( .Pik(\P[12][11] ), .Gik(\G[12][11] ), .Pk_1j(
        \P[10][9] ), .Gk_1j(\G[10][9] ), .Pij(\P[12][9] ), .Gij(\G[12][9] ) );
  PGblock_10 PGB_low_2_16 ( .Pik(\P[16][15] ), .Gik(\G[16][15] ), .Pk_1j(
        \P[14][13] ), .Gk_1j(\G[14][13] ), .Pij(\P[16][13] ), .Gij(\G[16][13] ) );
  PGblock_9 PGB_low_2_20 ( .Pik(\P[20][19] ), .Gik(\G[20][19] ), .Pk_1j(
        \P[18][17] ), .Gk_1j(\G[18][17] ), .Pij(\P[20][17] ), .Gij(\G[20][17] ) );
  PGblock_8 PGB_low_2_24 ( .Pik(\P[24][23] ), .Gik(\G[24][23] ), .Pk_1j(
        \P[22][21] ), .Gk_1j(\G[22][21] ), .Pij(\P[24][21] ), .Gij(\G[24][21] ) );
  PGblock_7 PGB_low_2_28 ( .Pik(\P[28][27] ), .Gik(\G[28][27] ), .Pk_1j(
        \P[26][25] ), .Gk_1j(\G[26][25] ), .Pij(\P[28][25] ), .Gij(\G[28][25] ) );
  PGblock_6 PGB_low_2_32 ( .Pik(\P[32][31] ), .Gik(\G[32][31] ), .Pk_1j(
        \P[30][29] ), .Gk_1j(\G[30][29] ), .Pij(\P[32][29] ), .Gij(\G[32][29] ) );
  PGblock_5 PGB_low_3_16 ( .Pik(\P[16][13] ), .Gik(\G[16][13] ), .Pk_1j(
        \P[12][9] ), .Gk_1j(\G[12][9] ), .Pij(\P[16][9] ), .Gij(\G[16][9] ) );
  PGblock_4 PGB_low_3_24 ( .Pik(\P[24][21] ), .Gik(\G[24][21] ), .Pk_1j(
        \P[20][17] ), .Gk_1j(\G[20][17] ), .Pij(\P[24][17] ), .Gij(\G[24][17] ) );
  PGblock_3 PGB_low_3_32 ( .Pik(\P[32][29] ), .Gik(\G[32][29] ), .Pk_1j(
        \P[28][25] ), .Gk_1j(\G[28][25] ), .Pij(\P[32][25] ), .Gij(\G[32][25] ) );
  PGblock_2 PGB_high_4_32_0 ( .Pik(\P[32][25] ), .Gik(\G[32][25] ), .Pk_1j(
        \P[24][17] ), .Gk_1j(\G[24][17] ), .Pij(\P[32][17] ), .Gij(\G[32][17] ) );
  PGblock_1 PGB_high_4_32_1 ( .Pik(\P[28][25] ), .Gik(\G[28][25] ), .Pk_1j(
        \P[24][17] ), .Gk_1j(\G[24][17] ), .Pij(\P[28][17] ), .Gij(\G[28][17] ) );
  OAI21_X1 U1 ( .B1(n4), .B2(n5), .A(n3), .ZN(\G[1][1] ) );
  INV_X1 U2 ( .A(A[1]), .ZN(n4) );
  INV_X1 U3 ( .A(B[1]), .ZN(n5) );
  OAI21_X1 U4 ( .B1(A[1]), .B2(B[1]), .A(Cin), .ZN(n3) );
endmodule


module SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_select_basic_N4_0 CSBI_1 ( .A(A[3:0]), .B(B[3:0]), .C_i(Ci[0]), .S(
        S[3:0]) );
  carry_select_basic_N4_7 CSBI_2 ( .A(A[7:4]), .B(B[7:4]), .C_i(Ci[1]), .S(
        S[7:4]) );
  carry_select_basic_N4_6 CSBI_3 ( .A(A[11:8]), .B(B[11:8]), .C_i(Ci[2]), .S(
        S[11:8]) );
  carry_select_basic_N4_5 CSBI_4 ( .A(A[15:12]), .B(B[15:12]), .C_i(Ci[3]), 
        .S(S[15:12]) );
  carry_select_basic_N4_4 CSBI_5 ( .A(A[19:16]), .B(B[19:16]), .C_i(Ci[4]), 
        .S(S[19:16]) );
  carry_select_basic_N4_3 CSBI_6 ( .A(A[23:20]), .B(B[23:20]), .C_i(Ci[5]), 
        .S(S[23:20]) );
  carry_select_basic_N4_2 CSBI_7 ( .A(A[27:24]), .B(B[27:24]), .C_i(Ci[6]), 
        .S(S[27:24]) );
  carry_select_basic_N4_1 CSBI_8 ( .A(A[31:28]), .B(B[31:28]), .C_i(Ci[7]), 
        .S(S[31:28]) );
endmodule


module P4Adder_NBIT32 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;

  wire   [7:1] Csum;

  carry_generator_NBIT32_NBIT_PER_BLOCK4 Carrygen0 ( .A(A), .B(B), .Cin(Cin), 
        .Co({Cout, Csum}) );
  SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 Sumgen0 ( .A(A), .B(B), .Ci({Csum, 
        Cin}), .S(S) );
endmodule


module ALU_NBIT32 ( OP1, OP2, .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , 
        \ALU_OPC[1] , \ALU_OPC[0] }), ALU_RES );
  input [31:0] OP1;
  input [31:0] OP2;
  output [31:0] ALU_RES;
  input \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] ;
  wire   select_zero_sig, ADD_SUB, LEFT_RIGHT, N176, N177, N178, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191,
         N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202,
         N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213,
         N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224,
         N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235,
         N236, N237, N238, N239, N240, N241, N242, N243, N244, N245,
         \COMP_RES[0] , n149, n71, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, \sig_intraMux[9] ,
         \sig_intraMux[8] , \sig_intraMux[7] , \sig_intraMux[6] ,
         \sig_intraMux[5] , \sig_intraMux[4] , \sig_intraMux[3] ,
         \sig_intraMux[31] , \sig_intraMux[30] , \sig_intraMux[2] ,
         \sig_intraMux[29] , \sig_intraMux[28] , \sig_intraMux[27] ,
         \sig_intraMux[26] , \sig_intraMux[25] , \sig_intraMux[24] ,
         \sig_intraMux[23] , \sig_intraMux[22] , \sig_intraMux[21] ,
         \sig_intraMux[20] , \sig_intraMux[1] , \sig_intraMux[19] ,
         \sig_intraMux[18] , \sig_intraMux[17] , \sig_intraMux[16] ,
         \sig_intraMux[15] , \sig_intraMux[14] , \sig_intraMux[13] ,
         \sig_intraMux[12] , \sig_intraMux[11] , \sig_intraMux[10] ,
         \sig_intraMux[0] , \SHIFT_RES[9] , \SHIFT_RES[8] , \SHIFT_RES[7] ,
         \SHIFT_RES[6] , \SHIFT_RES[5] , \SHIFT_RES[4] , \SHIFT_RES[3] ,
         \SHIFT_RES[31] , \SHIFT_RES[30] , \SHIFT_RES[2] , \SHIFT_RES[29] ,
         \SHIFT_RES[28] , \SHIFT_RES[27] , \SHIFT_RES[26] , \SHIFT_RES[25] ,
         \SHIFT_RES[24] , \SHIFT_RES[23] , \SHIFT_RES[22] , \SHIFT_RES[21] ,
         \SHIFT_RES[20] , \SHIFT_RES[1] , \SHIFT_RES[19] , \SHIFT_RES[18] ,
         \SHIFT_RES[17] , \SHIFT_RES[16] , \SHIFT_RES[15] , \SHIFT_RES[14] ,
         \SHIFT_RES[13] , \SHIFT_RES[12] , \SHIFT_RES[11] , \SHIFT_RES[10] ,
         \SHIFT_RES[0] , n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320;
  wire   [3:0] ALU_OPC;
  wire   [1:0] select_type_sig;
  wire   [31:0] A_ADD;
  wire   [31:0] B_ADD;
  wire   [31:0] LOGIC_RES;
  wire   [31:0] A_SHF;
  wire   [31:0] B_SHF;
  wire   [2:0] OPSel;
  wire   [31:0] A_CMP;
  wire   [31:0] B_CMP;
  wire   [31:0] ADD_SUB_RES;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  DLH_X1 \B_CMP_reg[31]  ( .G(n203), .D(OP2[31]), .Q(B_CMP[31]) );
  DLH_X1 \B_CMP_reg[30]  ( .G(n203), .D(OP2[30]), .Q(B_CMP[30]) );
  DLH_X1 \B_CMP_reg[29]  ( .G(n203), .D(OP2[29]), .Q(B_CMP[29]) );
  DLH_X1 \B_CMP_reg[28]  ( .G(n203), .D(OP2[28]), .Q(B_CMP[28]) );
  DLH_X1 \B_CMP_reg[27]  ( .G(n203), .D(OP2[27]), .Q(B_CMP[27]) );
  DLH_X1 \B_CMP_reg[26]  ( .G(n203), .D(OP2[26]), .Q(B_CMP[26]) );
  DLH_X1 \B_CMP_reg[25]  ( .G(n203), .D(OP2[25]), .Q(B_CMP[25]) );
  DLH_X1 \B_CMP_reg[24]  ( .G(n203), .D(OP2[24]), .Q(B_CMP[24]) );
  DLH_X1 \B_CMP_reg[23]  ( .G(n203), .D(OP2[23]), .Q(B_CMP[23]) );
  DLH_X1 \B_CMP_reg[22]  ( .G(n203), .D(OP2[22]), .Q(B_CMP[22]) );
  DLH_X1 \B_CMP_reg[21]  ( .G(n203), .D(OP2[21]), .Q(B_CMP[21]) );
  DLH_X1 \B_CMP_reg[20]  ( .G(n203), .D(OP2[20]), .Q(B_CMP[20]) );
  DLH_X1 \B_CMP_reg[19]  ( .G(n203), .D(OP2[19]), .Q(B_CMP[19]) );
  DLH_X1 \B_CMP_reg[18]  ( .G(n207), .D(OP2[18]), .Q(B_CMP[18]) );
  DLH_X1 \B_CMP_reg[17]  ( .G(n207), .D(OP2[17]), .Q(B_CMP[17]) );
  DLH_X1 \B_CMP_reg[16]  ( .G(n207), .D(OP2[16]), .Q(B_CMP[16]) );
  DLH_X1 \B_CMP_reg[15]  ( .G(n207), .D(OP2[15]), .Q(B_CMP[15]) );
  DLH_X1 \B_CMP_reg[14]  ( .G(n207), .D(OP2[14]), .Q(B_CMP[14]) );
  DLH_X1 \B_CMP_reg[13]  ( .G(n206), .D(OP2[13]), .Q(B_CMP[13]) );
  DLH_X1 \B_CMP_reg[12]  ( .G(n206), .D(OP2[12]), .Q(B_CMP[12]) );
  DLH_X1 \B_CMP_reg[11]  ( .G(n206), .D(OP2[11]), .Q(B_CMP[11]) );
  DLH_X1 \B_CMP_reg[10]  ( .G(n206), .D(OP2[10]), .Q(B_CMP[10]) );
  DLH_X1 \B_CMP_reg[9]  ( .G(n206), .D(OP2[9]), .Q(B_CMP[9]) );
  DLH_X1 \B_CMP_reg[8]  ( .G(n206), .D(OP2[8]), .Q(B_CMP[8]) );
  DLH_X1 \B_CMP_reg[7]  ( .G(n206), .D(OP2[7]), .Q(B_CMP[7]) );
  DLH_X1 \B_CMP_reg[6]  ( .G(n206), .D(OP2[6]), .Q(B_CMP[6]) );
  DLH_X1 \B_CMP_reg[5]  ( .G(n206), .D(OP2[5]), .Q(B_CMP[5]) );
  DLH_X1 \B_CMP_reg[4]  ( .G(n206), .D(OP2[4]), .Q(B_CMP[4]) );
  DLH_X1 \B_CMP_reg[3]  ( .G(n206), .D(OP2[3]), .Q(B_CMP[3]) );
  DLH_X1 \B_CMP_reg[2]  ( .G(n205), .D(OP2[2]), .Q(B_CMP[2]) );
  DLH_X1 \B_CMP_reg[1]  ( .G(n205), .D(OP2[1]), .Q(B_CMP[1]) );
  DLH_X1 \B_CMP_reg[0]  ( .G(n205), .D(OP2[0]), .Q(B_CMP[0]) );
  DLH_X1 select_zero_sig_reg ( .G(N176), .D(N177), .Q(select_zero_sig) );
  DLH_X1 ADD_SUB_reg ( .G(n215), .D(n184), .Q(ADD_SUB) );
  DLH_X1 \A_ADD_reg[31]  ( .G(n215), .D(OP1[31]), .Q(A_ADD[31]) );
  DLH_X1 \A_ADD_reg[30]  ( .G(n215), .D(OP1[30]), .Q(A_ADD[30]) );
  DLH_X1 \A_ADD_reg[29]  ( .G(n215), .D(OP1[29]), .Q(A_ADD[29]) );
  DLH_X1 \A_ADD_reg[28]  ( .G(n215), .D(OP1[28]), .Q(A_ADD[28]) );
  DLH_X1 \A_ADD_reg[27]  ( .G(n215), .D(OP1[27]), .Q(A_ADD[27]) );
  DLH_X1 \A_ADD_reg[26]  ( .G(n215), .D(OP1[26]), .Q(A_ADD[26]) );
  DLH_X1 \A_ADD_reg[25]  ( .G(n215), .D(OP1[25]), .Q(A_ADD[25]) );
  DLH_X1 \A_ADD_reg[24]  ( .G(n215), .D(OP1[24]), .Q(A_ADD[24]) );
  DLH_X1 \A_ADD_reg[23]  ( .G(n215), .D(OP1[23]), .Q(A_ADD[23]) );
  DLH_X1 \A_ADD_reg[22]  ( .G(n215), .D(OP1[22]), .Q(A_ADD[22]) );
  DLH_X1 \A_ADD_reg[21]  ( .G(n215), .D(OP1[21]), .Q(A_ADD[21]) );
  DLH_X1 \A_ADD_reg[20]  ( .G(n215), .D(OP1[20]), .Q(A_ADD[20]) );
  DLH_X1 \A_ADD_reg[19]  ( .G(n215), .D(OP1[19]), .Q(A_ADD[19]) );
  DLH_X1 \A_ADD_reg[18]  ( .G(n219), .D(OP1[18]), .Q(A_ADD[18]) );
  DLH_X1 \A_ADD_reg[17]  ( .G(n218), .D(OP1[17]), .Q(A_ADD[17]) );
  DLH_X1 \A_ADD_reg[16]  ( .G(n218), .D(OP1[16]), .Q(A_ADD[16]) );
  DLH_X1 \A_ADD_reg[15]  ( .G(n218), .D(OP1[15]), .Q(A_ADD[15]) );
  DLH_X1 \A_ADD_reg[14]  ( .G(n218), .D(OP1[14]), .Q(A_ADD[14]) );
  DLH_X1 \A_ADD_reg[13]  ( .G(n218), .D(OP1[13]), .Q(A_ADD[13]) );
  DLH_X1 \A_ADD_reg[12]  ( .G(n218), .D(OP1[12]), .Q(A_ADD[12]) );
  DLH_X1 \A_ADD_reg[11]  ( .G(n218), .D(OP1[11]), .Q(A_ADD[11]) );
  DLH_X1 \A_ADD_reg[10]  ( .G(n218), .D(OP1[10]), .Q(A_ADD[10]) );
  DLH_X1 \A_ADD_reg[9]  ( .G(n218), .D(OP1[9]), .Q(A_ADD[9]) );
  DLH_X1 \A_ADD_reg[8]  ( .G(n218), .D(OP1[8]), .Q(A_ADD[8]) );
  DLH_X1 \A_ADD_reg[7]  ( .G(n218), .D(OP1[7]), .Q(A_ADD[7]) );
  DLH_X1 \A_ADD_reg[6]  ( .G(n218), .D(OP1[6]), .Q(A_ADD[6]) );
  DLH_X1 \A_ADD_reg[5]  ( .G(n218), .D(OP1[5]), .Q(A_ADD[5]) );
  DLH_X1 \A_ADD_reg[4]  ( .G(n218), .D(OP1[4]), .Q(A_ADD[4]) );
  DLH_X1 \A_ADD_reg[3]  ( .G(n219), .D(OP1[3]), .Q(A_ADD[3]) );
  DLH_X1 \A_ADD_reg[2]  ( .G(n217), .D(OP1[2]), .Q(A_ADD[2]) );
  DLH_X1 \A_ADD_reg[1]  ( .G(n217), .D(OP1[1]), .Q(A_ADD[1]) );
  DLH_X1 \A_ADD_reg[0]  ( .G(n217), .D(OP1[0]), .Q(A_ADD[0]) );
  DLH_X1 \B_ADD_reg[31]  ( .G(n218), .D(N210), .Q(B_ADD[31]) );
  DLH_X1 \B_ADD_reg[30]  ( .G(n218), .D(N209), .Q(B_ADD[30]) );
  DLH_X1 \B_ADD_reg[29]  ( .G(n217), .D(N208), .Q(B_ADD[29]) );
  DLH_X1 \B_ADD_reg[28]  ( .G(n217), .D(N207), .Q(B_ADD[28]) );
  DLH_X1 \B_ADD_reg[27]  ( .G(n217), .D(N206), .Q(B_ADD[27]) );
  DLH_X1 \B_ADD_reg[26]  ( .G(n217), .D(N205), .Q(B_ADD[26]) );
  DLH_X1 \B_ADD_reg[25]  ( .G(n217), .D(N204), .Q(B_ADD[25]) );
  DLH_X1 \B_ADD_reg[24]  ( .G(n217), .D(N203), .Q(B_ADD[24]) );
  DLH_X1 \B_ADD_reg[23]  ( .G(n217), .D(N202), .Q(B_ADD[23]) );
  DLH_X1 \B_ADD_reg[22]  ( .G(n217), .D(N201), .Q(B_ADD[22]) );
  DLH_X1 \B_ADD_reg[21]  ( .G(n217), .D(N200), .Q(B_ADD[21]) );
  DLH_X1 \B_ADD_reg[20]  ( .G(n217), .D(N199), .Q(B_ADD[20]) );
  DLH_X1 \B_ADD_reg[19]  ( .G(n217), .D(N198), .Q(B_ADD[19]) );
  DLH_X1 \B_ADD_reg[18]  ( .G(n217), .D(N197), .Q(B_ADD[18]) );
  DLH_X1 \B_ADD_reg[17]  ( .G(n217), .D(N196), .Q(B_ADD[17]) );
  DLH_X1 \B_ADD_reg[16]  ( .G(n216), .D(N195), .Q(B_ADD[16]) );
  DLH_X1 \B_ADD_reg[15]  ( .G(n216), .D(N194), .Q(B_ADD[15]) );
  DLH_X1 \B_ADD_reg[14]  ( .G(n216), .D(N193), .Q(B_ADD[14]) );
  DLH_X1 \B_ADD_reg[13]  ( .G(n216), .D(N192), .Q(B_ADD[13]) );
  DLH_X1 \B_ADD_reg[12]  ( .G(n216), .D(N191), .Q(B_ADD[12]) );
  DLH_X1 \B_ADD_reg[11]  ( .G(n216), .D(N190), .Q(B_ADD[11]) );
  DLH_X1 \B_ADD_reg[10]  ( .G(n216), .D(N189), .Q(B_ADD[10]) );
  DLH_X1 \B_ADD_reg[9]  ( .G(n216), .D(N188), .Q(B_ADD[9]) );
  DLH_X1 \B_ADD_reg[8]  ( .G(n216), .D(N187), .Q(B_ADD[8]) );
  DLH_X1 \B_ADD_reg[7]  ( .G(n216), .D(N186), .Q(B_ADD[7]) );
  DLH_X1 \B_ADD_reg[6]  ( .G(n216), .D(N185), .Q(B_ADD[6]) );
  DLH_X1 \B_ADD_reg[5]  ( .G(n216), .D(N184), .Q(B_ADD[5]) );
  DLH_X1 \B_ADD_reg[4]  ( .G(n216), .D(N183), .Q(B_ADD[4]) );
  DLH_X1 \B_ADD_reg[3]  ( .G(n216), .D(N182), .Q(B_ADD[3]) );
  DLH_X1 \B_ADD_reg[2]  ( .G(n216), .D(N181), .Q(B_ADD[2]) );
  DLH_X1 \B_ADD_reg[1]  ( .G(n216), .D(N180), .Q(B_ADD[1]) );
  DLH_X1 \B_ADD_reg[0]  ( .G(n215), .D(N179), .Q(B_ADD[0]) );
  DLH_X1 \LOGIC_RES_reg[31]  ( .G(n213), .D(N243), .Q(LOGIC_RES[31]) );
  DLH_X1 \LOGIC_RES_reg[30]  ( .G(n213), .D(N242), .Q(LOGIC_RES[30]) );
  DLH_X1 \LOGIC_RES_reg[29]  ( .G(n213), .D(N241), .Q(LOGIC_RES[29]) );
  DLH_X1 \LOGIC_RES_reg[28]  ( .G(n213), .D(N240), .Q(LOGIC_RES[28]) );
  DLH_X1 \LOGIC_RES_reg[27]  ( .G(n213), .D(N239), .Q(LOGIC_RES[27]) );
  DLH_X1 \LOGIC_RES_reg[26]  ( .G(n213), .D(N238), .Q(LOGIC_RES[26]) );
  DLH_X1 \LOGIC_RES_reg[25]  ( .G(n213), .D(N237), .Q(LOGIC_RES[25]) );
  DLH_X1 \LOGIC_RES_reg[24]  ( .G(n213), .D(N236), .Q(LOGIC_RES[24]) );
  DLH_X1 \LOGIC_RES_reg[23]  ( .G(n213), .D(N235), .Q(LOGIC_RES[23]) );
  DLH_X1 \LOGIC_RES_reg[22]  ( .G(n213), .D(N234), .Q(LOGIC_RES[22]) );
  DLH_X1 \LOGIC_RES_reg[21]  ( .G(n213), .D(N233), .Q(LOGIC_RES[21]) );
  DLH_X1 \LOGIC_RES_reg[20]  ( .G(n213), .D(N232), .Q(LOGIC_RES[20]) );
  DLH_X1 \LOGIC_RES_reg[19]  ( .G(n213), .D(N231), .Q(LOGIC_RES[19]) );
  DLH_X1 \LOGIC_RES_reg[18]  ( .G(n213), .D(N230), .Q(LOGIC_RES[18]) );
  DLH_X1 \LOGIC_RES_reg[17]  ( .G(n213), .D(N229), .Q(LOGIC_RES[17]) );
  DLH_X1 \LOGIC_RES_reg[16]  ( .G(n214), .D(N228), .Q(LOGIC_RES[16]) );
  DLH_X1 \LOGIC_RES_reg[15]  ( .G(n214), .D(N227), .Q(LOGIC_RES[15]) );
  DLH_X1 \LOGIC_RES_reg[14]  ( .G(n214), .D(N226), .Q(LOGIC_RES[14]) );
  DLH_X1 \LOGIC_RES_reg[13]  ( .G(n214), .D(N225), .Q(LOGIC_RES[13]) );
  DLH_X1 \LOGIC_RES_reg[12]  ( .G(n214), .D(N224), .Q(LOGIC_RES[12]) );
  DLH_X1 \LOGIC_RES_reg[11]  ( .G(n214), .D(N223), .Q(LOGIC_RES[11]) );
  DLH_X1 \LOGIC_RES_reg[10]  ( .G(n214), .D(N222), .Q(LOGIC_RES[10]) );
  DLH_X1 \LOGIC_RES_reg[9]  ( .G(n214), .D(N221), .Q(LOGIC_RES[9]) );
  DLH_X1 \LOGIC_RES_reg[8]  ( .G(n214), .D(N220), .Q(LOGIC_RES[8]) );
  DLH_X1 \LOGIC_RES_reg[7]  ( .G(n214), .D(N219), .Q(LOGIC_RES[7]) );
  DLH_X1 \LOGIC_RES_reg[6]  ( .G(n214), .D(N218), .Q(LOGIC_RES[6]) );
  DLH_X1 \LOGIC_RES_reg[5]  ( .G(n214), .D(N217), .Q(LOGIC_RES[5]) );
  DLH_X1 \LOGIC_RES_reg[4]  ( .G(n214), .D(N216), .Q(LOGIC_RES[4]) );
  DLH_X1 \LOGIC_RES_reg[3]  ( .G(n214), .D(N215), .Q(LOGIC_RES[3]) );
  DLH_X1 \LOGIC_RES_reg[2]  ( .G(n214), .D(N214), .Q(LOGIC_RES[2]) );
  DLH_X1 \LOGIC_RES_reg[1]  ( .G(n214), .D(N213), .Q(LOGIC_RES[1]) );
  DLH_X1 \LOGIC_RES_reg[0]  ( .G(N211), .D(N212), .Q(LOGIC_RES[0]) );
  DLH_X1 LEFT_RIGHT_reg ( .G(n208), .D(n149), .Q(LEFT_RIGHT) );
  DLH_X1 \A_SHF_reg[31]  ( .G(n211), .D(OP1[31]), .Q(A_SHF[31]) );
  DLH_X1 \A_SHF_reg[30]  ( .G(n211), .D(OP1[30]), .Q(A_SHF[30]) );
  DLH_X1 \A_SHF_reg[29]  ( .G(n211), .D(OP1[29]), .Q(A_SHF[29]) );
  DLH_X1 \A_SHF_reg[28]  ( .G(n211), .D(OP1[28]), .Q(A_SHF[28]) );
  DLH_X1 \A_SHF_reg[27]  ( .G(n211), .D(OP1[27]), .Q(A_SHF[27]) );
  DLH_X1 \A_SHF_reg[26]  ( .G(n211), .D(OP1[26]), .Q(A_SHF[26]) );
  DLH_X1 \A_SHF_reg[25]  ( .G(n211), .D(OP1[25]), .Q(A_SHF[25]) );
  DLH_X1 \A_SHF_reg[24]  ( .G(n211), .D(OP1[24]), .Q(A_SHF[24]) );
  DLH_X1 \A_SHF_reg[23]  ( .G(n211), .D(OP1[23]), .Q(A_SHF[23]) );
  DLH_X1 \A_SHF_reg[22]  ( .G(n211), .D(OP1[22]), .Q(A_SHF[22]) );
  DLH_X1 \A_SHF_reg[21]  ( .G(n211), .D(OP1[21]), .Q(A_SHF[21]) );
  DLH_X1 \A_SHF_reg[20]  ( .G(n212), .D(OP1[20]), .Q(A_SHF[20]) );
  DLH_X1 \A_SHF_reg[19]  ( .G(n212), .D(OP1[19]), .Q(A_SHF[19]) );
  DLH_X1 \A_SHF_reg[18]  ( .G(n212), .D(OP1[18]), .Q(A_SHF[18]) );
  DLH_X1 \A_SHF_reg[17]  ( .G(n210), .D(OP1[17]), .Q(A_SHF[17]) );
  DLH_X1 \A_SHF_reg[16]  ( .G(n208), .D(OP1[16]), .Q(A_SHF[16]) );
  DLH_X1 \A_SHF_reg[15]  ( .G(n208), .D(OP1[15]), .Q(A_SHF[15]) );
  DLH_X1 \A_SHF_reg[14]  ( .G(n208), .D(OP1[14]), .Q(A_SHF[14]) );
  DLH_X1 \A_SHF_reg[13]  ( .G(n208), .D(OP1[13]), .Q(A_SHF[13]) );
  DLH_X1 \A_SHF_reg[12]  ( .G(n208), .D(OP1[12]), .Q(A_SHF[12]) );
  DLH_X1 \A_SHF_reg[11]  ( .G(n208), .D(OP1[11]), .Q(A_SHF[11]) );
  DLH_X1 \A_SHF_reg[10]  ( .G(n208), .D(OP1[10]), .Q(A_SHF[10]) );
  DLH_X1 \A_SHF_reg[9]  ( .G(n208), .D(OP1[9]), .Q(A_SHF[9]) );
  DLH_X1 \A_SHF_reg[8]  ( .G(n208), .D(OP1[8]), .Q(A_SHF[8]) );
  DLH_X1 \A_SHF_reg[7]  ( .G(n208), .D(OP1[7]), .Q(A_SHF[7]) );
  DLH_X1 \A_SHF_reg[6]  ( .G(n208), .D(OP1[6]), .Q(A_SHF[6]) );
  DLH_X1 \A_SHF_reg[5]  ( .G(n208), .D(OP1[5]), .Q(A_SHF[5]) );
  DLH_X1 \A_SHF_reg[4]  ( .G(n208), .D(OP1[4]), .Q(A_SHF[4]) );
  DLH_X1 \A_SHF_reg[3]  ( .G(n209), .D(OP1[3]), .Q(A_SHF[3]) );
  DLH_X1 \A_SHF_reg[2]  ( .G(n209), .D(OP1[2]), .Q(A_SHF[2]) );
  DLH_X1 \A_SHF_reg[1]  ( .G(n210), .D(OP1[1]), .Q(A_SHF[1]) );
  DLH_X1 \A_SHF_reg[0]  ( .G(n210), .D(OP1[0]), .Q(A_SHF[0]) );
  DLH_X1 \B_SHF_reg[31]  ( .G(n209), .D(OP2[31]), .Q(B_SHF[31]) );
  DLH_X1 \B_SHF_reg[30]  ( .G(n209), .D(OP2[30]), .Q(B_SHF[30]) );
  DLH_X1 \B_SHF_reg[29]  ( .G(n209), .D(OP2[29]), .Q(B_SHF[29]) );
  DLH_X1 \B_SHF_reg[28]  ( .G(n209), .D(OP2[28]), .Q(B_SHF[28]) );
  DLH_X1 \B_SHF_reg[27]  ( .G(n209), .D(OP2[27]), .Q(B_SHF[27]) );
  DLH_X1 \B_SHF_reg[26]  ( .G(n209), .D(OP2[26]), .Q(B_SHF[26]) );
  DLH_X1 \B_SHF_reg[25]  ( .G(n209), .D(OP2[25]), .Q(B_SHF[25]) );
  DLH_X1 \B_SHF_reg[24]  ( .G(n209), .D(OP2[24]), .Q(B_SHF[24]) );
  DLH_X1 \B_SHF_reg[23]  ( .G(n209), .D(OP2[23]), .Q(B_SHF[23]) );
  DLH_X1 \B_SHF_reg[22]  ( .G(n209), .D(OP2[22]), .Q(B_SHF[22]) );
  DLH_X1 \B_SHF_reg[21]  ( .G(n209), .D(OP2[21]), .Q(B_SHF[21]) );
  DLH_X1 \B_SHF_reg[20]  ( .G(n209), .D(OP2[20]), .Q(B_SHF[20]) );
  DLH_X1 \B_SHF_reg[19]  ( .G(n209), .D(OP2[19]), .Q(B_SHF[19]) );
  DLH_X1 \B_SHF_reg[18]  ( .G(n209), .D(OP2[18]), .Q(B_SHF[18]) );
  DLH_X1 \B_SHF_reg[17]  ( .G(n210), .D(OP2[17]), .Q(B_SHF[17]) );
  DLH_X1 \B_SHF_reg[16]  ( .G(n210), .D(OP2[16]), .Q(B_SHF[16]) );
  DLH_X1 \B_SHF_reg[15]  ( .G(n210), .D(OP2[15]), .Q(B_SHF[15]) );
  DLH_X1 \B_SHF_reg[14]  ( .G(n210), .D(OP2[14]), .Q(B_SHF[14]) );
  DLH_X1 \B_SHF_reg[13]  ( .G(n210), .D(OP2[13]), .Q(B_SHF[13]) );
  DLH_X1 \B_SHF_reg[12]  ( .G(n210), .D(OP2[12]), .Q(B_SHF[12]) );
  DLH_X1 \B_SHF_reg[11]  ( .G(n210), .D(OP2[11]), .Q(B_SHF[11]) );
  DLH_X1 \B_SHF_reg[10]  ( .G(n210), .D(OP2[10]), .Q(B_SHF[10]) );
  DLH_X1 \B_SHF_reg[9]  ( .G(n210), .D(OP2[9]), .Q(B_SHF[9]) );
  DLH_X1 \B_SHF_reg[8]  ( .G(n210), .D(OP2[8]), .Q(B_SHF[8]) );
  DLH_X1 \B_SHF_reg[7]  ( .G(n211), .D(OP2[7]), .Q(B_SHF[7]) );
  DLH_X1 \B_SHF_reg[6]  ( .G(n210), .D(OP2[6]), .Q(B_SHF[6]) );
  DLH_X1 \B_SHF_reg[5]  ( .G(n210), .D(OP2[5]), .Q(B_SHF[5]) );
  DLH_X1 \B_SHF_reg[4]  ( .G(n210), .D(OP2[4]), .Q(B_SHF[4]) );
  DLH_X1 \B_SHF_reg[3]  ( .G(n211), .D(OP2[3]), .Q(B_SHF[3]) );
  DLH_X1 \B_SHF_reg[2]  ( .G(n211), .D(OP2[2]), .Q(B_SHF[2]) );
  DLH_X1 \B_SHF_reg[1]  ( .G(n211), .D(OP2[1]), .Q(B_SHF[1]) );
  DLH_X1 \B_SHF_reg[0]  ( .G(n211), .D(OP2[0]), .Q(B_SHF[0]) );
  DLH_X1 \OPSel_reg[2]  ( .G(n205), .D(n146), .Q(OPSel[2]) );
  DLH_X1 \OPSel_reg[1]  ( .G(n205), .D(n145), .Q(OPSel[1]) );
  DLH_X1 \A_CMP_reg[31]  ( .G(n206), .D(OP1[31]), .Q(A_CMP[31]) );
  DLH_X1 \A_CMP_reg[30]  ( .G(n206), .D(OP1[30]), .Q(A_CMP[30]) );
  DLH_X1 \A_CMP_reg[29]  ( .G(n206), .D(OP1[29]), .Q(A_CMP[29]) );
  DLH_X1 \A_CMP_reg[28]  ( .G(n206), .D(OP1[28]), .Q(A_CMP[28]) );
  DLH_X1 \A_CMP_reg[27]  ( .G(n206), .D(OP1[27]), .Q(A_CMP[27]) );
  DLH_X1 \A_CMP_reg[26]  ( .G(n205), .D(OP1[26]), .Q(A_CMP[26]) );
  DLH_X1 \A_CMP_reg[25]  ( .G(n205), .D(OP1[25]), .Q(A_CMP[25]) );
  DLH_X1 \A_CMP_reg[24]  ( .G(n205), .D(OP1[24]), .Q(A_CMP[24]) );
  DLH_X1 \A_CMP_reg[23]  ( .G(n205), .D(OP1[23]), .Q(A_CMP[23]) );
  DLH_X1 \A_CMP_reg[22]  ( .G(n205), .D(OP1[22]), .Q(A_CMP[22]) );
  DLH_X1 \A_CMP_reg[21]  ( .G(n205), .D(OP1[21]), .Q(A_CMP[21]) );
  DLH_X1 \A_CMP_reg[20]  ( .G(n205), .D(OP1[20]), .Q(A_CMP[20]) );
  DLH_X1 \A_CMP_reg[19]  ( .G(n205), .D(OP1[19]), .Q(A_CMP[19]) );
  DLH_X1 \A_CMP_reg[18]  ( .G(n205), .D(OP1[18]), .Q(A_CMP[18]) );
  DLH_X1 \A_CMP_reg[17]  ( .G(n205), .D(OP1[17]), .Q(A_CMP[17]) );
  DLH_X1 \A_CMP_reg[16]  ( .G(n205), .D(OP1[16]), .Q(A_CMP[16]) );
  DLH_X1 \A_CMP_reg[15]  ( .G(n204), .D(OP1[15]), .Q(A_CMP[15]) );
  DLH_X1 \A_CMP_reg[14]  ( .G(n204), .D(OP1[14]), .Q(A_CMP[14]) );
  DLH_X1 \A_CMP_reg[13]  ( .G(n204), .D(OP1[13]), .Q(A_CMP[13]) );
  DLH_X1 \A_CMP_reg[12]  ( .G(n204), .D(OP1[12]), .Q(A_CMP[12]) );
  DLH_X1 \A_CMP_reg[11]  ( .G(n204), .D(OP1[11]), .Q(A_CMP[11]) );
  DLH_X1 \A_CMP_reg[10]  ( .G(n204), .D(OP1[10]), .Q(A_CMP[10]) );
  DLH_X1 \A_CMP_reg[9]  ( .G(n204), .D(OP1[9]), .Q(A_CMP[9]) );
  DLH_X1 \A_CMP_reg[8]  ( .G(n204), .D(OP1[8]), .Q(A_CMP[8]) );
  DLH_X1 \A_CMP_reg[7]  ( .G(n204), .D(OP1[7]), .Q(A_CMP[7]) );
  DLH_X1 \A_CMP_reg[6]  ( .G(n204), .D(OP1[6]), .Q(A_CMP[6]) );
  DLH_X1 \A_CMP_reg[5]  ( .G(n204), .D(OP1[5]), .Q(A_CMP[5]) );
  DLH_X1 \A_CMP_reg[4]  ( .G(n204), .D(OP1[4]), .Q(A_CMP[4]) );
  DLH_X1 \A_CMP_reg[3]  ( .G(n204), .D(OP1[3]), .Q(A_CMP[3]) );
  DLH_X1 \A_CMP_reg[2]  ( .G(n204), .D(OP1[2]), .Q(A_CMP[2]) );
  DLH_X1 \A_CMP_reg[1]  ( .G(n204), .D(OP1[1]), .Q(A_CMP[1]) );
  DLH_X1 \A_CMP_reg[0]  ( .G(n204), .D(OP1[0]), .Q(A_CMP[0]) );
  NAND3_X1 U188 ( .A1(n198), .A2(n284), .A3(OP2[31]), .ZN(n74) );
  NAND3_X1 U189 ( .A1(n200), .A2(n283), .A3(OP2[30]), .ZN(n79) );
  NAND3_X1 U190 ( .A1(n200), .A2(n282), .A3(OP2[29]), .ZN(n81) );
  NAND3_X1 U191 ( .A1(n200), .A2(n281), .A3(OP2[28]), .ZN(n83) );
  NAND3_X1 U192 ( .A1(n200), .A2(n280), .A3(OP2[27]), .ZN(n85) );
  NAND3_X1 U193 ( .A1(n200), .A2(n279), .A3(OP2[26]), .ZN(n87) );
  NAND3_X1 U194 ( .A1(n200), .A2(n278), .A3(OP2[25]), .ZN(n89) );
  NAND3_X1 U195 ( .A1(n200), .A2(n277), .A3(OP2[24]), .ZN(n91) );
  NAND3_X1 U196 ( .A1(n199), .A2(n276), .A3(OP2[23]), .ZN(n93) );
  NAND3_X1 U197 ( .A1(n199), .A2(n275), .A3(OP2[22]), .ZN(n95) );
  NAND3_X1 U198 ( .A1(n199), .A2(n274), .A3(OP2[21]), .ZN(n97) );
  NAND3_X1 U199 ( .A1(n199), .A2(n273), .A3(OP2[20]), .ZN(n99) );
  NAND3_X1 U200 ( .A1(n199), .A2(n272), .A3(OP2[19]), .ZN(n101) );
  NAND3_X1 U201 ( .A1(n199), .A2(n271), .A3(OP2[18]), .ZN(n103) );
  NAND3_X1 U202 ( .A1(n199), .A2(n270), .A3(OP2[17]), .ZN(n105) );
  NAND3_X1 U203 ( .A1(n199), .A2(n269), .A3(OP2[16]), .ZN(n107) );
  NAND3_X1 U204 ( .A1(n199), .A2(n268), .A3(OP2[15]), .ZN(n109) );
  NAND3_X1 U205 ( .A1(n199), .A2(n267), .A3(OP2[14]), .ZN(n111) );
  NAND3_X1 U206 ( .A1(n199), .A2(n266), .A3(OP2[13]), .ZN(n113) );
  NAND3_X1 U207 ( .A1(n199), .A2(n265), .A3(OP2[12]), .ZN(n115) );
  NAND3_X1 U208 ( .A1(n199), .A2(n264), .A3(OP2[11]), .ZN(n117) );
  NAND3_X1 U209 ( .A1(n200), .A2(n263), .A3(OP2[10]), .ZN(n119) );
  NAND3_X1 U210 ( .A1(n199), .A2(n262), .A3(OP2[9]), .ZN(n121) );
  NAND3_X1 U211 ( .A1(n199), .A2(n261), .A3(OP2[8]), .ZN(n123) );
  NAND3_X1 U212 ( .A1(n199), .A2(n260), .A3(OP2[7]), .ZN(n125) );
  NAND3_X1 U213 ( .A1(n199), .A2(n259), .A3(OP2[6]), .ZN(n127) );
  NAND3_X1 U214 ( .A1(n199), .A2(n258), .A3(OP2[5]), .ZN(n129) );
  NAND3_X1 U215 ( .A1(n199), .A2(n257), .A3(OP2[4]), .ZN(n131) );
  NAND3_X1 U216 ( .A1(n199), .A2(n256), .A3(OP2[3]), .ZN(n133) );
  NAND3_X1 U217 ( .A1(n198), .A2(n255), .A3(OP2[2]), .ZN(n135) );
  NAND3_X1 U218 ( .A1(n198), .A2(n254), .A3(OP2[1]), .ZN(n137) );
  NAND3_X1 U219 ( .A1(n198), .A2(n253), .A3(OP2[0]), .ZN(n139) );
  NAND3_X1 U220 ( .A1(ALU_OPC[1]), .A2(n318), .A3(ALU_OPC[3]), .ZN(n71) );
  NAND3_X1 U221 ( .A1(n319), .A2(n318), .A3(n320), .ZN(n144) );
  comparator_NBIT32 Comp ( .A(A_CMP), .B(B_CMP), .OPSel({OPSel[2:1], 1'b1}), 
        .RES({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, \COMP_RES[0] }) );
  shifter Shift ( .A(A_SHF), .B(B_SHF), .LOGIC_ARITH(1'b1), .LEFT_RIGHT(
        LEFT_RIGHT), .RES({\SHIFT_RES[31] , \SHIFT_RES[30] , \SHIFT_RES[29] , 
        \SHIFT_RES[28] , \SHIFT_RES[27] , \SHIFT_RES[26] , \SHIFT_RES[25] , 
        \SHIFT_RES[24] , \SHIFT_RES[23] , \SHIFT_RES[22] , \SHIFT_RES[21] , 
        \SHIFT_RES[20] , \SHIFT_RES[19] , \SHIFT_RES[18] , \SHIFT_RES[17] , 
        \SHIFT_RES[16] , \SHIFT_RES[15] , \SHIFT_RES[14] , \SHIFT_RES[13] , 
        \SHIFT_RES[12] , \SHIFT_RES[11] , \SHIFT_RES[10] , \SHIFT_RES[9] , 
        \SHIFT_RES[8] , \SHIFT_RES[7] , \SHIFT_RES[6] , \SHIFT_RES[5] , 
        \SHIFT_RES[4] , \SHIFT_RES[3] , \SHIFT_RES[2] , \SHIFT_RES[1] , 
        \SHIFT_RES[0] }) );
  P4Adder_NBIT32 Add_Sub_unit ( .A(A_ADD), .B(B_ADD), .Cin(ADD_SUB), .S(
        ADD_SUB_RES) );
  mux41_NBIT32_1 Res_mux ( .A(ADD_SUB_RES), .B(LOGIC_RES), .C({\SHIFT_RES[31] , 
        \SHIFT_RES[30] , \SHIFT_RES[29] , \SHIFT_RES[28] , \SHIFT_RES[27] , 
        \SHIFT_RES[26] , \SHIFT_RES[25] , \SHIFT_RES[24] , \SHIFT_RES[23] , 
        \SHIFT_RES[22] , \SHIFT_RES[21] , \SHIFT_RES[20] , \SHIFT_RES[19] , 
        \SHIFT_RES[18] , \SHIFT_RES[17] , \SHIFT_RES[16] , \SHIFT_RES[15] , 
        \SHIFT_RES[14] , \SHIFT_RES[13] , \SHIFT_RES[12] , \SHIFT_RES[11] , 
        \SHIFT_RES[10] , \SHIFT_RES[9] , \SHIFT_RES[8] , \SHIFT_RES[7] , 
        \SHIFT_RES[6] , \SHIFT_RES[5] , \SHIFT_RES[4] , \SHIFT_RES[3] , 
        \SHIFT_RES[2] , \SHIFT_RES[1] , \SHIFT_RES[0] }), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, \COMP_RES[0] }), .S(select_type_sig), .Z({
        \sig_intraMux[31] , \sig_intraMux[30] , \sig_intraMux[29] , 
        \sig_intraMux[28] , \sig_intraMux[27] , \sig_intraMux[26] , 
        \sig_intraMux[25] , \sig_intraMux[24] , \sig_intraMux[23] , 
        \sig_intraMux[22] , \sig_intraMux[21] , \sig_intraMux[20] , 
        \sig_intraMux[19] , \sig_intraMux[18] , \sig_intraMux[17] , 
        \sig_intraMux[16] , \sig_intraMux[15] , \sig_intraMux[14] , 
        \sig_intraMux[13] , \sig_intraMux[12] , \sig_intraMux[11] , 
        \sig_intraMux[10] , \sig_intraMux[9] , \sig_intraMux[8] , 
        \sig_intraMux[7] , \sig_intraMux[6] , \sig_intraMux[5] , 
        \sig_intraMux[4] , \sig_intraMux[3] , \sig_intraMux[2] , 
        \sig_intraMux[1] , \sig_intraMux[0] }) );
  mux21_NBIT32_1 Zeros_mux ( .A({\sig_intraMux[31] , \sig_intraMux[30] , 
        \sig_intraMux[29] , \sig_intraMux[28] , \sig_intraMux[27] , 
        \sig_intraMux[26] , \sig_intraMux[25] , \sig_intraMux[24] , 
        \sig_intraMux[23] , \sig_intraMux[22] , \sig_intraMux[21] , 
        \sig_intraMux[20] , \sig_intraMux[19] , \sig_intraMux[18] , 
        \sig_intraMux[17] , \sig_intraMux[16] , \sig_intraMux[15] , 
        \sig_intraMux[14] , \sig_intraMux[13] , \sig_intraMux[12] , 
        \sig_intraMux[11] , \sig_intraMux[10] , \sig_intraMux[9] , 
        \sig_intraMux[8] , \sig_intraMux[7] , \sig_intraMux[6] , 
        \sig_intraMux[5] , \sig_intraMux[4] , \sig_intraMux[3] , 
        \sig_intraMux[2] , \sig_intraMux[1] , \sig_intraMux[0] }), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(select_zero_sig), .Z(
        ALU_RES) );
  BUF_X1 U4 ( .A(N211), .Z(n213) );
  BUF_X1 U5 ( .A(N178), .Z(n215) );
  INV_X1 U6 ( .A(n184), .ZN(n201) );
  BUF_X1 U7 ( .A(n77), .Z(n188) );
  BUF_X1 U8 ( .A(n77), .Z(n189) );
  INV_X1 U9 ( .A(n184), .ZN(n202) );
  BUF_X1 U10 ( .A(n195), .Z(n199) );
  BUF_X1 U11 ( .A(n194), .Z(n197) );
  BUF_X1 U12 ( .A(n194), .Z(n196) );
  BUF_X1 U13 ( .A(n77), .Z(n190) );
  BUF_X1 U14 ( .A(n194), .Z(n198) );
  BUF_X1 U15 ( .A(n195), .Z(n200) );
  NAND2_X1 U16 ( .A1(n201), .A2(n185), .ZN(N178) );
  OR2_X1 U17 ( .A1(n198), .A2(n193), .ZN(N211) );
  OR2_X1 U18 ( .A1(n213), .A2(n203), .ZN(select_type_sig[0]) );
  OR2_X1 U19 ( .A1(n208), .A2(n203), .ZN(select_type_sig[1]) );
  BUF_X1 U20 ( .A(n76), .Z(n192) );
  BUF_X1 U21 ( .A(n76), .Z(n191) );
  BUF_X1 U22 ( .A(n140), .Z(n185) );
  BUF_X1 U23 ( .A(n76), .Z(n193) );
  BUF_X1 U24 ( .A(n140), .Z(n186) );
  BUF_X1 U25 ( .A(N244), .Z(n208) );
  BUF_X1 U26 ( .A(n140), .Z(n187) );
  BUF_X1 U27 ( .A(N245), .Z(n203) );
  AND2_X1 U28 ( .A1(n142), .A2(n320), .ZN(n184) );
  OR4_X1 U29 ( .A1(N177), .A2(n215), .A3(n149), .A4(select_type_sig[0]), .ZN(
        N176) );
  AND2_X1 U30 ( .A1(n198), .A2(n320), .ZN(n77) );
  NOR2_X1 U31 ( .A1(n320), .A2(n71), .ZN(n146) );
  BUF_X1 U32 ( .A(n75), .Z(n194) );
  BUF_X1 U33 ( .A(n75), .Z(n195) );
  AND2_X1 U34 ( .A1(n208), .A2(n320), .ZN(n149) );
  NOR3_X1 U35 ( .A1(n319), .A2(ALU_OPC[3]), .A3(n318), .ZN(N244) );
  NOR3_X1 U36 ( .A1(ALU_OPC[2]), .A2(ALU_OPC[3]), .A3(n319), .ZN(n142) );
  NAND4_X1 U37 ( .A1(ALU_OPC[0]), .A2(n319), .A3(n318), .A4(n317), .ZN(n140)
         );
  NOR3_X1 U38 ( .A1(ALU_OPC[1]), .A2(ALU_OPC[3]), .A3(n318), .ZN(n75) );
  INV_X1 U39 ( .A(ALU_OPC[1]), .ZN(n319) );
  OAI22_X1 U40 ( .A1(OP2[0]), .A2(n202), .B1(n285), .B2(n185), .ZN(N179) );
  OAI22_X1 U41 ( .A1(OP2[1]), .A2(n202), .B1(n286), .B2(n185), .ZN(N180) );
  OAI22_X1 U42 ( .A1(OP2[2]), .A2(n201), .B1(n287), .B2(n185), .ZN(N181) );
  OAI22_X1 U43 ( .A1(OP2[3]), .A2(n202), .B1(n288), .B2(n185), .ZN(N182) );
  OAI22_X1 U44 ( .A1(OP2[4]), .A2(n201), .B1(n289), .B2(n185), .ZN(N183) );
  OAI22_X1 U45 ( .A1(OP2[5]), .A2(n202), .B1(n290), .B2(n185), .ZN(N184) );
  OAI22_X1 U46 ( .A1(OP2[6]), .A2(n201), .B1(n291), .B2(n185), .ZN(N185) );
  OAI22_X1 U47 ( .A1(OP2[7]), .A2(n202), .B1(n292), .B2(n185), .ZN(N186) );
  OAI22_X1 U48 ( .A1(OP2[8]), .A2(n202), .B1(n293), .B2(n185), .ZN(N187) );
  OAI22_X1 U49 ( .A1(OP2[9]), .A2(n202), .B1(n294), .B2(n185), .ZN(N188) );
  OAI22_X1 U50 ( .A1(OP2[10]), .A2(n202), .B1(n295), .B2(n185), .ZN(N189) );
  OAI22_X1 U51 ( .A1(OP2[11]), .A2(n202), .B1(n296), .B2(n186), .ZN(N190) );
  OAI22_X1 U52 ( .A1(OP2[12]), .A2(n202), .B1(n297), .B2(n186), .ZN(N191) );
  OAI22_X1 U53 ( .A1(OP2[13]), .A2(n202), .B1(n298), .B2(n186), .ZN(N192) );
  OAI22_X1 U54 ( .A1(OP2[14]), .A2(n202), .B1(n299), .B2(n186), .ZN(N193) );
  OAI22_X1 U55 ( .A1(OP2[15]), .A2(n202), .B1(n300), .B2(n186), .ZN(N194) );
  OAI22_X1 U56 ( .A1(OP2[16]), .A2(n202), .B1(n301), .B2(n186), .ZN(N195) );
  OAI22_X1 U57 ( .A1(OP2[17]), .A2(n202), .B1(n302), .B2(n186), .ZN(N196) );
  OAI22_X1 U58 ( .A1(OP2[18]), .A2(n202), .B1(n303), .B2(n186), .ZN(N197) );
  OAI22_X1 U59 ( .A1(OP2[19]), .A2(n202), .B1(n304), .B2(n186), .ZN(N198) );
  OAI22_X1 U60 ( .A1(OP2[20]), .A2(n201), .B1(n305), .B2(n186), .ZN(N199) );
  OAI22_X1 U61 ( .A1(OP2[21]), .A2(n201), .B1(n306), .B2(n186), .ZN(N200) );
  OAI22_X1 U62 ( .A1(OP2[22]), .A2(n201), .B1(n307), .B2(n186), .ZN(N201) );
  OAI22_X1 U63 ( .A1(OP2[23]), .A2(n201), .B1(n308), .B2(n187), .ZN(N202) );
  OAI22_X1 U64 ( .A1(OP2[24]), .A2(n201), .B1(n309), .B2(n187), .ZN(N203) );
  OAI22_X1 U65 ( .A1(OP2[25]), .A2(n201), .B1(n310), .B2(n187), .ZN(N204) );
  OAI22_X1 U66 ( .A1(OP2[26]), .A2(n201), .B1(n311), .B2(n187), .ZN(N205) );
  OAI22_X1 U67 ( .A1(OP2[27]), .A2(n201), .B1(n312), .B2(n187), .ZN(N206) );
  OAI22_X1 U68 ( .A1(OP2[28]), .A2(n201), .B1(n313), .B2(n187), .ZN(N207) );
  OAI22_X1 U69 ( .A1(OP2[29]), .A2(n201), .B1(n314), .B2(n187), .ZN(N208) );
  OAI22_X1 U70 ( .A1(OP2[30]), .A2(n201), .B1(n315), .B2(n187), .ZN(N209) );
  OAI22_X1 U71 ( .A1(OP2[31]), .A2(n201), .B1(n316), .B2(n187), .ZN(N210) );
  INV_X1 U72 ( .A(ALU_OPC[0]), .ZN(n320) );
  INV_X1 U73 ( .A(ALU_OPC[2]), .ZN(n318) );
  OAI21_X1 U74 ( .B1(n143), .B2(n317), .A(n144), .ZN(N177) );
  AOI22_X1 U75 ( .A1(ALU_OPC[0]), .A2(n319), .B1(ALU_OPC[2]), .B2(ALU_OPC[1]), 
        .ZN(n143) );
  NAND2_X1 U76 ( .A1(n71), .A2(n141), .ZN(N245) );
  NAND4_X1 U77 ( .A1(ALU_OPC[3]), .A2(ALU_OPC[2]), .A3(n320), .A4(n319), .ZN(
        n141) );
  INV_X1 U78 ( .A(ALU_OPC[3]), .ZN(n317) );
  AND2_X1 U79 ( .A1(ALU_OPC[0]), .A2(n142), .ZN(n76) );
  OAI21_X1 U80 ( .B1(n122), .B2(n261), .A(n123), .ZN(N220) );
  AOI221_X1 U81 ( .B1(n197), .B2(n293), .C1(OP2[8]), .C2(n192), .A(n188), .ZN(
        n122) );
  INV_X1 U82 ( .A(OP1[8]), .ZN(n261) );
  OAI21_X1 U83 ( .B1(n120), .B2(n262), .A(n121), .ZN(N221) );
  AOI221_X1 U84 ( .B1(n197), .B2(n294), .C1(OP2[9]), .C2(n192), .A(n188), .ZN(
        n120) );
  INV_X1 U85 ( .A(OP1[9]), .ZN(n262) );
  OAI21_X1 U86 ( .B1(n118), .B2(n263), .A(n119), .ZN(N222) );
  AOI221_X1 U87 ( .B1(n197), .B2(n295), .C1(OP2[10]), .C2(n192), .A(n188), 
        .ZN(n118) );
  INV_X1 U88 ( .A(OP1[10]), .ZN(n263) );
  OAI21_X1 U89 ( .B1(n116), .B2(n264), .A(n117), .ZN(N223) );
  AOI221_X1 U90 ( .B1(n197), .B2(n296), .C1(OP2[11]), .C2(n192), .A(n188), 
        .ZN(n116) );
  INV_X1 U91 ( .A(OP1[11]), .ZN(n264) );
  OAI21_X1 U92 ( .B1(n114), .B2(n265), .A(n115), .ZN(N224) );
  AOI221_X1 U93 ( .B1(n197), .B2(n297), .C1(OP2[12]), .C2(n192), .A(n189), 
        .ZN(n114) );
  INV_X1 U94 ( .A(OP1[12]), .ZN(n265) );
  OAI21_X1 U95 ( .B1(n112), .B2(n266), .A(n113), .ZN(N225) );
  AOI221_X1 U96 ( .B1(n197), .B2(n298), .C1(OP2[13]), .C2(n192), .A(n189), 
        .ZN(n112) );
  INV_X1 U97 ( .A(OP1[13]), .ZN(n266) );
  OAI21_X1 U98 ( .B1(n110), .B2(n267), .A(n111), .ZN(N226) );
  AOI221_X1 U99 ( .B1(n197), .B2(n299), .C1(OP2[14]), .C2(n192), .A(n189), 
        .ZN(n110) );
  INV_X1 U100 ( .A(OP1[14]), .ZN(n267) );
  OAI21_X1 U101 ( .B1(n108), .B2(n268), .A(n109), .ZN(N227) );
  AOI221_X1 U102 ( .B1(n197), .B2(n300), .C1(OP2[15]), .C2(n192), .A(n189), 
        .ZN(n108) );
  INV_X1 U103 ( .A(OP1[15]), .ZN(n268) );
  OAI21_X1 U104 ( .B1(n106), .B2(n269), .A(n107), .ZN(N228) );
  AOI221_X1 U105 ( .B1(n197), .B2(n301), .C1(OP2[16]), .C2(n192), .A(n189), 
        .ZN(n106) );
  INV_X1 U106 ( .A(OP1[16]), .ZN(n269) );
  OAI21_X1 U107 ( .B1(n104), .B2(n270), .A(n105), .ZN(N229) );
  AOI221_X1 U108 ( .B1(n197), .B2(n302), .C1(OP2[17]), .C2(n192), .A(n189), 
        .ZN(n104) );
  INV_X1 U109 ( .A(OP1[17]), .ZN(n270) );
  OAI21_X1 U110 ( .B1(n102), .B2(n271), .A(n103), .ZN(N230) );
  AOI221_X1 U111 ( .B1(n197), .B2(n303), .C1(OP2[18]), .C2(n191), .A(n189), 
        .ZN(n102) );
  INV_X1 U112 ( .A(OP1[18]), .ZN(n271) );
  OAI21_X1 U113 ( .B1(n100), .B2(n272), .A(n101), .ZN(N231) );
  AOI221_X1 U114 ( .B1(n197), .B2(n304), .C1(OP2[19]), .C2(n191), .A(n189), 
        .ZN(n100) );
  INV_X1 U115 ( .A(OP1[19]), .ZN(n272) );
  OAI21_X1 U116 ( .B1(n98), .B2(n273), .A(n99), .ZN(N232) );
  AOI221_X1 U117 ( .B1(n196), .B2(n305), .C1(OP2[20]), .C2(n191), .A(n189), 
        .ZN(n98) );
  INV_X1 U118 ( .A(OP1[20]), .ZN(n273) );
  OAI21_X1 U119 ( .B1(n96), .B2(n274), .A(n97), .ZN(N233) );
  AOI221_X1 U120 ( .B1(n196), .B2(n306), .C1(OP2[21]), .C2(n191), .A(n189), 
        .ZN(n96) );
  INV_X1 U121 ( .A(OP1[21]), .ZN(n274) );
  OAI21_X1 U122 ( .B1(n94), .B2(n275), .A(n95), .ZN(N234) );
  AOI221_X1 U123 ( .B1(n196), .B2(n307), .C1(OP2[22]), .C2(n191), .A(n189), 
        .ZN(n94) );
  INV_X1 U124 ( .A(OP1[22]), .ZN(n275) );
  OAI21_X1 U125 ( .B1(n92), .B2(n276), .A(n93), .ZN(N235) );
  AOI221_X1 U126 ( .B1(n196), .B2(n308), .C1(OP2[23]), .C2(n192), .A(n189), 
        .ZN(n92) );
  INV_X1 U127 ( .A(OP1[23]), .ZN(n276) );
  OAI21_X1 U128 ( .B1(n90), .B2(n277), .A(n91), .ZN(N236) );
  AOI221_X1 U129 ( .B1(n196), .B2(n309), .C1(OP2[24]), .C2(n191), .A(n190), 
        .ZN(n90) );
  INV_X1 U130 ( .A(OP1[24]), .ZN(n277) );
  OAI21_X1 U131 ( .B1(n88), .B2(n278), .A(n89), .ZN(N237) );
  AOI221_X1 U132 ( .B1(n196), .B2(n310), .C1(OP2[25]), .C2(n191), .A(n190), 
        .ZN(n88) );
  INV_X1 U133 ( .A(OP1[25]), .ZN(n278) );
  OAI21_X1 U134 ( .B1(n86), .B2(n279), .A(n87), .ZN(N238) );
  AOI221_X1 U135 ( .B1(n196), .B2(n311), .C1(OP2[26]), .C2(n191), .A(n190), 
        .ZN(n86) );
  INV_X1 U136 ( .A(OP1[26]), .ZN(n279) );
  OAI21_X1 U137 ( .B1(n84), .B2(n280), .A(n85), .ZN(N239) );
  AOI221_X1 U138 ( .B1(n196), .B2(n312), .C1(OP2[27]), .C2(n191), .A(n190), 
        .ZN(n84) );
  INV_X1 U139 ( .A(OP1[27]), .ZN(n280) );
  OAI21_X1 U140 ( .B1(n82), .B2(n281), .A(n83), .ZN(N240) );
  AOI221_X1 U141 ( .B1(n196), .B2(n313), .C1(OP2[28]), .C2(n191), .A(n190), 
        .ZN(n82) );
  INV_X1 U142 ( .A(OP1[28]), .ZN(n281) );
  OAI21_X1 U143 ( .B1(n80), .B2(n282), .A(n81), .ZN(N241) );
  AOI221_X1 U144 ( .B1(n196), .B2(n314), .C1(OP2[29]), .C2(n191), .A(n190), 
        .ZN(n80) );
  INV_X1 U145 ( .A(OP1[29]), .ZN(n282) );
  OAI21_X1 U146 ( .B1(n78), .B2(n283), .A(n79), .ZN(N242) );
  AOI221_X1 U147 ( .B1(n196), .B2(n315), .C1(OP2[30]), .C2(n191), .A(n190), 
        .ZN(n78) );
  INV_X1 U148 ( .A(OP1[30]), .ZN(n283) );
  OAI21_X1 U149 ( .B1(n73), .B2(n284), .A(n74), .ZN(N243) );
  AOI221_X1 U150 ( .B1(n196), .B2(n316), .C1(n193), .C2(OP2[31]), .A(n190), 
        .ZN(n73) );
  INV_X1 U151 ( .A(OP1[31]), .ZN(n284) );
  OAI21_X1 U152 ( .B1(n138), .B2(n253), .A(n139), .ZN(N212) );
  AOI221_X1 U153 ( .B1(n198), .B2(n285), .C1(OP2[0]), .C2(n193), .A(n188), 
        .ZN(n138) );
  INV_X1 U154 ( .A(OP1[0]), .ZN(n253) );
  OAI21_X1 U155 ( .B1(n136), .B2(n254), .A(n137), .ZN(N213) );
  AOI221_X1 U156 ( .B1(n198), .B2(n286), .C1(OP2[1]), .C2(n193), .A(n188), 
        .ZN(n136) );
  INV_X1 U157 ( .A(OP1[1]), .ZN(n254) );
  OAI21_X1 U158 ( .B1(n134), .B2(n255), .A(n135), .ZN(N214) );
  AOI221_X1 U159 ( .B1(n198), .B2(n287), .C1(OP2[2]), .C2(n193), .A(n188), 
        .ZN(n134) );
  INV_X1 U160 ( .A(OP1[2]), .ZN(n255) );
  OAI21_X1 U161 ( .B1(n132), .B2(n256), .A(n133), .ZN(N215) );
  AOI221_X1 U162 ( .B1(n198), .B2(n288), .C1(OP2[3]), .C2(n193), .A(n188), 
        .ZN(n132) );
  INV_X1 U163 ( .A(OP1[3]), .ZN(n256) );
  OAI21_X1 U164 ( .B1(n130), .B2(n257), .A(n131), .ZN(N216) );
  AOI221_X1 U165 ( .B1(n198), .B2(n289), .C1(OP2[4]), .C2(n193), .A(n188), 
        .ZN(n130) );
  INV_X1 U166 ( .A(OP1[4]), .ZN(n257) );
  OAI21_X1 U167 ( .B1(n128), .B2(n258), .A(n129), .ZN(N217) );
  AOI221_X1 U168 ( .B1(n198), .B2(n290), .C1(OP2[5]), .C2(n193), .A(n188), 
        .ZN(n128) );
  INV_X1 U169 ( .A(OP1[5]), .ZN(n258) );
  OAI21_X1 U170 ( .B1(n126), .B2(n259), .A(n127), .ZN(N218) );
  AOI221_X1 U171 ( .B1(n198), .B2(n291), .C1(OP2[6]), .C2(n193), .A(n188), 
        .ZN(n126) );
  INV_X1 U172 ( .A(OP1[6]), .ZN(n259) );
  OAI21_X1 U173 ( .B1(n124), .B2(n260), .A(n125), .ZN(N219) );
  AOI221_X1 U174 ( .B1(n198), .B2(n292), .C1(OP2[7]), .C2(n192), .A(n188), 
        .ZN(n124) );
  INV_X1 U175 ( .A(OP1[7]), .ZN(n260) );
  NOR2_X1 U176 ( .A1(ALU_OPC[0]), .A2(n71), .ZN(n145) );
  INV_X1 U177 ( .A(OP2[0]), .ZN(n285) );
  INV_X1 U178 ( .A(OP2[1]), .ZN(n286) );
  INV_X1 U179 ( .A(OP2[2]), .ZN(n287) );
  INV_X1 U180 ( .A(OP2[3]), .ZN(n288) );
  INV_X1 U181 ( .A(OP2[4]), .ZN(n289) );
  INV_X1 U182 ( .A(OP2[5]), .ZN(n290) );
  INV_X1 U183 ( .A(OP2[6]), .ZN(n291) );
  INV_X1 U184 ( .A(OP2[7]), .ZN(n292) );
  INV_X1 U185 ( .A(OP2[8]), .ZN(n293) );
  INV_X1 U186 ( .A(OP2[9]), .ZN(n294) );
  INV_X1 U187 ( .A(OP2[10]), .ZN(n295) );
  INV_X1 U222 ( .A(OP2[11]), .ZN(n296) );
  INV_X1 U223 ( .A(OP2[12]), .ZN(n297) );
  INV_X1 U224 ( .A(OP2[13]), .ZN(n298) );
  INV_X1 U225 ( .A(OP2[14]), .ZN(n299) );
  INV_X1 U226 ( .A(OP2[15]), .ZN(n300) );
  INV_X1 U227 ( .A(OP2[16]), .ZN(n301) );
  INV_X1 U228 ( .A(OP2[17]), .ZN(n302) );
  INV_X1 U229 ( .A(OP2[18]), .ZN(n303) );
  INV_X1 U230 ( .A(OP2[19]), .ZN(n304) );
  INV_X1 U231 ( .A(OP2[20]), .ZN(n305) );
  INV_X1 U232 ( .A(OP2[21]), .ZN(n306) );
  INV_X1 U233 ( .A(OP2[22]), .ZN(n307) );
  INV_X1 U234 ( .A(OP2[23]), .ZN(n308) );
  INV_X1 U235 ( .A(OP2[24]), .ZN(n309) );
  INV_X1 U236 ( .A(OP2[25]), .ZN(n310) );
  INV_X1 U237 ( .A(OP2[26]), .ZN(n311) );
  INV_X1 U238 ( .A(OP2[27]), .ZN(n312) );
  INV_X1 U239 ( .A(OP2[28]), .ZN(n313) );
  INV_X1 U240 ( .A(OP2[29]), .ZN(n314) );
  INV_X1 U241 ( .A(OP2[30]), .ZN(n315) );
  INV_X1 U242 ( .A(OP2[31]), .ZN(n316) );
  CLKBUF_X1 U243 ( .A(N245), .Z(n204) );
  CLKBUF_X1 U244 ( .A(N245), .Z(n205) );
  CLKBUF_X1 U245 ( .A(N245), .Z(n206) );
  CLKBUF_X1 U246 ( .A(N245), .Z(n207) );
  CLKBUF_X1 U247 ( .A(N244), .Z(n209) );
  CLKBUF_X1 U248 ( .A(N244), .Z(n210) );
  CLKBUF_X1 U249 ( .A(N244), .Z(n211) );
  CLKBUF_X1 U250 ( .A(N244), .Z(n212) );
  CLKBUF_X1 U251 ( .A(N211), .Z(n214) );
  CLKBUF_X1 U252 ( .A(N178), .Z(n216) );
  CLKBUF_X1 U253 ( .A(N178), .Z(n217) );
  CLKBUF_X1 U254 ( .A(N178), .Z(n218) );
  CLKBUF_X1 U255 ( .A(N178), .Z(n219) );
endmodule


module Execute_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \B[0] , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57;
  assign SUM[1] = B[1];
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U4 ( .A(B[3]), .B(B[2]), .Z(SUM[3]) );
  XOR2_X1 U5 ( .A(B[4]), .B(n30), .Z(SUM[4]) );
  XOR2_X1 U6 ( .A(B[5]), .B(n31), .Z(SUM[5]) );
  XOR2_X1 U7 ( .A(B[6]), .B(n32), .Z(SUM[6]) );
  XOR2_X1 U8 ( .A(B[7]), .B(n33), .Z(SUM[7]) );
  XOR2_X1 U9 ( .A(B[8]), .B(n34), .Z(SUM[8]) );
  XOR2_X1 U10 ( .A(B[9]), .B(n35), .Z(SUM[9]) );
  XOR2_X1 U11 ( .A(B[10]), .B(n36), .Z(SUM[10]) );
  XOR2_X1 U12 ( .A(B[11]), .B(n37), .Z(SUM[11]) );
  XOR2_X1 U13 ( .A(B[12]), .B(n38), .Z(SUM[12]) );
  XOR2_X1 U14 ( .A(B[13]), .B(n39), .Z(SUM[13]) );
  XOR2_X1 U15 ( .A(B[14]), .B(n40), .Z(SUM[14]) );
  XOR2_X1 U16 ( .A(B[15]), .B(n41), .Z(SUM[15]) );
  XOR2_X1 U17 ( .A(B[16]), .B(n42), .Z(SUM[16]) );
  XOR2_X1 U18 ( .A(B[17]), .B(n43), .Z(SUM[17]) );
  XOR2_X1 U19 ( .A(B[18]), .B(n44), .Z(SUM[18]) );
  XOR2_X1 U20 ( .A(B[19]), .B(n45), .Z(SUM[19]) );
  XOR2_X1 U21 ( .A(B[20]), .B(n46), .Z(SUM[20]) );
  XOR2_X1 U22 ( .A(B[21]), .B(n47), .Z(SUM[21]) );
  XOR2_X1 U23 ( .A(B[22]), .B(n48), .Z(SUM[22]) );
  XOR2_X1 U24 ( .A(B[23]), .B(n49), .Z(SUM[23]) );
  XOR2_X1 U25 ( .A(B[24]), .B(n50), .Z(SUM[24]) );
  XOR2_X1 U26 ( .A(B[25]), .B(n51), .Z(SUM[25]) );
  XOR2_X1 U27 ( .A(B[26]), .B(n52), .Z(SUM[26]) );
  XOR2_X1 U28 ( .A(B[27]), .B(n53), .Z(SUM[27]) );
  XOR2_X1 U29 ( .A(B[28]), .B(n54), .Z(SUM[28]) );
  XOR2_X1 U30 ( .A(B[29]), .B(n55), .Z(SUM[29]) );
  XOR2_X1 U31 ( .A(B[30]), .B(n56), .Z(SUM[30]) );
  INV_X1 U1 ( .A(B[2]), .ZN(SUM[2]) );
  AND2_X1 U2 ( .A1(B[29]), .A2(n55), .ZN(n56) );
  AND2_X1 U3 ( .A1(B[4]), .A2(n30), .ZN(n31) );
  AND2_X1 U32 ( .A1(B[5]), .A2(n31), .ZN(n32) );
  AND2_X1 U33 ( .A1(B[6]), .A2(n32), .ZN(n33) );
  AND2_X1 U34 ( .A1(B[7]), .A2(n33), .ZN(n34) );
  AND2_X1 U35 ( .A1(B[8]), .A2(n34), .ZN(n35) );
  AND2_X1 U36 ( .A1(B[9]), .A2(n35), .ZN(n36) );
  AND2_X1 U37 ( .A1(B[10]), .A2(n36), .ZN(n37) );
  AND2_X1 U38 ( .A1(B[11]), .A2(n37), .ZN(n38) );
  AND2_X1 U39 ( .A1(B[12]), .A2(n38), .ZN(n39) );
  AND2_X1 U40 ( .A1(B[13]), .A2(n39), .ZN(n40) );
  AND2_X1 U41 ( .A1(B[14]), .A2(n40), .ZN(n41) );
  AND2_X1 U42 ( .A1(B[15]), .A2(n41), .ZN(n42) );
  AND2_X1 U43 ( .A1(B[16]), .A2(n42), .ZN(n43) );
  AND2_X1 U44 ( .A1(B[17]), .A2(n43), .ZN(n44) );
  AND2_X1 U45 ( .A1(B[18]), .A2(n44), .ZN(n45) );
  AND2_X1 U46 ( .A1(B[19]), .A2(n45), .ZN(n46) );
  AND2_X1 U47 ( .A1(B[20]), .A2(n46), .ZN(n47) );
  AND2_X1 U48 ( .A1(B[21]), .A2(n47), .ZN(n48) );
  AND2_X1 U49 ( .A1(B[22]), .A2(n48), .ZN(n49) );
  AND2_X1 U50 ( .A1(B[23]), .A2(n49), .ZN(n50) );
  AND2_X1 U51 ( .A1(B[24]), .A2(n50), .ZN(n51) );
  AND2_X1 U52 ( .A1(B[25]), .A2(n51), .ZN(n52) );
  AND2_X1 U53 ( .A1(B[26]), .A2(n52), .ZN(n53) );
  AND2_X1 U54 ( .A1(B[27]), .A2(n53), .ZN(n54) );
  AND2_X1 U55 ( .A1(B[28]), .A2(n54), .ZN(n55) );
  AND2_X1 U56 ( .A1(B[3]), .A2(B[2]), .ZN(n30) );
  XNOR2_X1 U57 ( .A(B[31]), .B(n57), .ZN(SUM[31]) );
  NAND2_X1 U58 ( .A1(B[30]), .A2(n56), .ZN(n57) );
endmodule


module Execute_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module Execute ( CLK, RST, MUX_A_SEL, MUX_B_SEL, .ALU_OPC({\ALU_OPC[3] , 
        \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), ALU_OUTREG_EN, JUMP_TYPE, 
        PC_IN, A_IN, B_IN, IMM_IN, ADD_WR_IN, ADD_RS1_IN, ADD_RS2_IN, 
        ADD_WR_MEM, ADD_WR_WB, RF_WE_MEM, RF_WE_WB, OP_MEM, OP_WB, PC_SEL, 
        ZERO_FLAG, NPC_ABS, NPC_REL, ALU_RES, B_OUT, ADD_WR_OUT );
  input [1:0] MUX_B_SEL;
  input [1:0] JUMP_TYPE;
  input [31:0] PC_IN;
  input [31:0] A_IN;
  input [31:0] B_IN;
  input [31:0] IMM_IN;
  input [4:0] ADD_WR_IN;
  input [4:0] ADD_RS1_IN;
  input [4:0] ADD_RS2_IN;
  input [4:0] ADD_WR_MEM;
  input [4:0] ADD_WR_WB;
  input [31:0] OP_MEM;
  input [31:0] OP_WB;
  output [1:0] PC_SEL;
  output [31:0] NPC_ABS;
  output [31:0] NPC_REL;
  output [31:0] ALU_RES;
  output [31:0] B_OUT;
  output [4:0] ADD_WR_OUT;
  input CLK, RST, MUX_A_SEL, \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] ,
         \ALU_OPC[0] , ALU_OUTREG_EN, RF_WE_MEM, RF_WE_WB;
  output ZERO_FLAG;
  wire   sig_RST, sig_ZERO_FLAG, N9, N8, N7, N6, N5, N4, N31, N30, N3, N29,
         N28, N27, N26, N25, N24, N23, N22, N21, N20, N2, N19, N18, N17, N16,
         N15, N14, N13, N12, N11, N10, N1, N0, \OP2_FW[9] , \OP2_FW[8] ,
         \OP2_FW[7] , \OP2_FW[6] , \OP2_FW[5] , \OP2_FW[4] , \OP2_FW[3] ,
         \OP2_FW[31] , \OP2_FW[30] , \OP2_FW[2] , \OP2_FW[29] , \OP2_FW[28] ,
         \OP2_FW[27] , \OP2_FW[26] , \OP2_FW[25] , \OP2_FW[24] , \OP2_FW[23] ,
         \OP2_FW[22] , \OP2_FW[21] , \OP2_FW[20] , \OP2_FW[1] , \OP2_FW[19] ,
         \OP2_FW[18] , \OP2_FW[17] , \OP2_FW[16] , \OP2_FW[15] , \OP2_FW[14] ,
         \OP2_FW[13] , \OP2_FW[12] , \OP2_FW[11] , \OP2_FW[10] , \OP2_FW[0] ,
         n11;
  wire   [3:0] ALU_OPC;
  wire   [31:0] sig_NPC_ABS;
  wire   [31:0] sig_NPC_REL;
  wire   [1:0] sig_PC_SEL;
  wire   [1:0] FWDA;
  wire   [1:0] FWDB;
  wire   [31:0] sig_OP1;
  wire   [31:0] sig_OP2;
  wire   [31:0] sig_ALU_RES;

  Branch_Cond_Unit_NBIT32 Branch_Cond ( .RST(sig_RST), .A(sig_NPC_ABS), 
        .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), 
        .JUMP_TYPE(JUMP_TYPE), .PC_SEL(sig_PC_SEL), .ZERO(sig_ZERO_FLAG) );
  ff_1 ff0 ( .D(sig_ZERO_FLAG), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(ZERO_FLAG)
         );
  regn_N2 reg0 ( .DIN(sig_PC_SEL), .CLK(CLK), .EN(1'b1), .RST(RST), .DOUT(
        PC_SEL) );
  FWD_Unit FWD ( .RST(sig_RST), .ADD_RS1(ADD_RS1_IN), .ADD_RS2(ADD_RS2_IN), 
        .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_WB(ADD_WR_WB), .RF_WE_MEM(RF_WE_MEM), 
        .RF_WE_WB(RF_WE_WB), .FWDA(FWDA), .FWDB(FWDB) );
  mux41_NBIT32_0 FW1 ( .A(A_IN), .B(OP_WB), .C(OP_MEM), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(FWDA), .Z(sig_NPC_ABS) );
  mux41_NBIT32_4 FW2 ( .A(B_IN), .B(OP_WB), .C(OP_MEM), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(FWDB), .Z({\OP2_FW[31] , 
        \OP2_FW[30] , \OP2_FW[29] , \OP2_FW[28] , \OP2_FW[27] , \OP2_FW[26] , 
        \OP2_FW[25] , \OP2_FW[24] , \OP2_FW[23] , \OP2_FW[22] , \OP2_FW[21] , 
        \OP2_FW[20] , \OP2_FW[19] , \OP2_FW[18] , \OP2_FW[17] , \OP2_FW[16] , 
        \OP2_FW[15] , \OP2_FW[14] , \OP2_FW[13] , \OP2_FW[12] , \OP2_FW[11] , 
        \OP2_FW[10] , \OP2_FW[9] , \OP2_FW[8] , \OP2_FW[7] , \OP2_FW[6] , 
        \OP2_FW[5] , \OP2_FW[4] , \OP2_FW[3] , \OP2_FW[2] , \OP2_FW[1] , 
        \OP2_FW[0] }) );
  mux21_NBIT32_3 muxA ( .A(sig_NPC_ABS), .B(PC_IN), .S(MUX_A_SEL), .Z(sig_OP1)
         );
  mux41_NBIT32_3 muxB ( .A({\OP2_FW[31] , \OP2_FW[30] , \OP2_FW[29] , 
        \OP2_FW[28] , \OP2_FW[27] , \OP2_FW[26] , \OP2_FW[25] , \OP2_FW[24] , 
        \OP2_FW[23] , \OP2_FW[22] , \OP2_FW[21] , \OP2_FW[20] , \OP2_FW[19] , 
        \OP2_FW[18] , \OP2_FW[17] , \OP2_FW[16] , \OP2_FW[15] , \OP2_FW[14] , 
        \OP2_FW[13] , \OP2_FW[12] , \OP2_FW[11] , \OP2_FW[10] , \OP2_FW[9] , 
        \OP2_FW[8] , \OP2_FW[7] , \OP2_FW[6] , \OP2_FW[5] , \OP2_FW[4] , 
        \OP2_FW[3] , \OP2_FW[2] , \OP2_FW[1] , \OP2_FW[0] }), .B(IMM_IN), .C({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(MUX_B_SEL), .Z(sig_OP2) );
  ALU_NBIT32 alu0 ( .OP1(sig_OP1), .OP2(sig_OP2), .ALU_OPC({\ALU_OPC[3] , 
        \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), .ALU_RES(sig_ALU_RES) );
  regn_N32_6 alureg ( .DIN(sig_ALU_RES), .CLK(CLK), .EN(ALU_OUTREG_EN), .RST(
        RST), .DOUT(ALU_RES) );
  regn_N32_5 B_reg ( .DIN({\OP2_FW[31] , \OP2_FW[30] , \OP2_FW[29] , 
        \OP2_FW[28] , \OP2_FW[27] , \OP2_FW[26] , \OP2_FW[25] , \OP2_FW[24] , 
        \OP2_FW[23] , \OP2_FW[22] , \OP2_FW[21] , \OP2_FW[20] , \OP2_FW[19] , 
        \OP2_FW[18] , \OP2_FW[17] , \OP2_FW[16] , \OP2_FW[15] , \OP2_FW[14] , 
        \OP2_FW[13] , \OP2_FW[12] , \OP2_FW[11] , \OP2_FW[10] , \OP2_FW[9] , 
        \OP2_FW[8] , \OP2_FW[7] , \OP2_FW[6] , \OP2_FW[5] , \OP2_FW[4] , 
        \OP2_FW[3] , \OP2_FW[2] , \OP2_FW[1] , \OP2_FW[0] }), .CLK(CLK), .EN(
        ALU_OUTREG_EN), .RST(RST), .DOUT(B_OUT) );
  regn_N5_2 ADD_WR_reg ( .DIN(ADD_WR_IN), .CLK(CLK), .EN(ALU_OUTREG_EN), .RST(
        RST), .DOUT(ADD_WR_OUT) );
  regn_N32_4 NPC_ABS_reg ( .DIN(sig_NPC_ABS), .CLK(CLK), .EN(ALU_OUTREG_EN), 
        .RST(RST), .DOUT(NPC_ABS) );
  regn_N32_3 NPC_REL_reg ( .DIN(sig_NPC_REL), .CLK(CLK), .EN(ALU_OUTREG_EN), 
        .RST(RST), .DOUT(NPC_REL) );
  Execute_DW01_add_1 add_1_root_add_0_root_add_118_2 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .B(IMM_IN), .CI(1'b0), .SUM({N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0})
         );
  Execute_DW01_add_0 add_0_root_add_0_root_add_118_2 ( .A(PC_IN), .B({N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}), 
        .CI(1'b0), .SUM(sig_NPC_REL) );
  NOR2_X1 U5 ( .A1(ZERO_FLAG), .A2(n11), .ZN(sig_RST) );
  INV_X1 U6 ( .A(RST), .ZN(n11) );
endmodule


module Memory ( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, DRAM_EN_IN, PC_SEL, 
        NPC_IN, NPC_ABS, NPC_REL, ALU_RES_IN, B_IN, ADD_WR_IN, DRAM_DATA_IN, 
        PC_OUT, DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, DRAM_ADDR_OUT, 
        DRAM_DATA_OUT, DATA_OUT, ALU_RES_OUT, OP_MEM, ADD_WR_MEM, ADD_WR_OUT
 );
  input [1:0] PC_SEL;
  input [31:0] NPC_IN;
  input [31:0] NPC_ABS;
  input [31:0] NPC_REL;
  input [31:0] ALU_RES_IN;
  input [31:0] B_IN;
  input [4:0] ADD_WR_IN;
  input [31:0] DRAM_DATA_IN;
  output [31:0] PC_OUT;
  output [31:0] DRAM_ADDR_OUT;
  output [31:0] DRAM_DATA_OUT;
  output [31:0] DATA_OUT;
  output [31:0] ALU_RES_OUT;
  output [31:0] OP_MEM;
  output [4:0] ADD_WR_MEM;
  output [4:0] ADD_WR_OUT;
  input CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, DRAM_EN_IN;
  output DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT;
  wire   DRAM_EN_IN, DRAM_R_IN, DRAM_W_IN;
  assign DRAM_EN_OUT = DRAM_EN_IN;
  assign DRAM_R_OUT = DRAM_R_IN;
  assign DRAM_W_OUT = DRAM_W_IN;
  assign OP_MEM[31] = ALU_RES_IN[31];
  assign DRAM_ADDR_OUT[31] = ALU_RES_IN[31];
  assign OP_MEM[30] = ALU_RES_IN[30];
  assign DRAM_ADDR_OUT[30] = ALU_RES_IN[30];
  assign OP_MEM[29] = ALU_RES_IN[29];
  assign DRAM_ADDR_OUT[29] = ALU_RES_IN[29];
  assign OP_MEM[28] = ALU_RES_IN[28];
  assign DRAM_ADDR_OUT[28] = ALU_RES_IN[28];
  assign OP_MEM[27] = ALU_RES_IN[27];
  assign DRAM_ADDR_OUT[27] = ALU_RES_IN[27];
  assign OP_MEM[26] = ALU_RES_IN[26];
  assign DRAM_ADDR_OUT[26] = ALU_RES_IN[26];
  assign OP_MEM[25] = ALU_RES_IN[25];
  assign DRAM_ADDR_OUT[25] = ALU_RES_IN[25];
  assign OP_MEM[24] = ALU_RES_IN[24];
  assign DRAM_ADDR_OUT[24] = ALU_RES_IN[24];
  assign OP_MEM[23] = ALU_RES_IN[23];
  assign DRAM_ADDR_OUT[23] = ALU_RES_IN[23];
  assign OP_MEM[22] = ALU_RES_IN[22];
  assign DRAM_ADDR_OUT[22] = ALU_RES_IN[22];
  assign OP_MEM[21] = ALU_RES_IN[21];
  assign DRAM_ADDR_OUT[21] = ALU_RES_IN[21];
  assign OP_MEM[20] = ALU_RES_IN[20];
  assign DRAM_ADDR_OUT[20] = ALU_RES_IN[20];
  assign OP_MEM[19] = ALU_RES_IN[19];
  assign DRAM_ADDR_OUT[19] = ALU_RES_IN[19];
  assign OP_MEM[18] = ALU_RES_IN[18];
  assign DRAM_ADDR_OUT[18] = ALU_RES_IN[18];
  assign OP_MEM[17] = ALU_RES_IN[17];
  assign DRAM_ADDR_OUT[17] = ALU_RES_IN[17];
  assign OP_MEM[16] = ALU_RES_IN[16];
  assign DRAM_ADDR_OUT[16] = ALU_RES_IN[16];
  assign OP_MEM[15] = ALU_RES_IN[15];
  assign DRAM_ADDR_OUT[15] = ALU_RES_IN[15];
  assign OP_MEM[14] = ALU_RES_IN[14];
  assign DRAM_ADDR_OUT[14] = ALU_RES_IN[14];
  assign OP_MEM[13] = ALU_RES_IN[13];
  assign DRAM_ADDR_OUT[13] = ALU_RES_IN[13];
  assign OP_MEM[12] = ALU_RES_IN[12];
  assign DRAM_ADDR_OUT[12] = ALU_RES_IN[12];
  assign OP_MEM[11] = ALU_RES_IN[11];
  assign DRAM_ADDR_OUT[11] = ALU_RES_IN[11];
  assign OP_MEM[10] = ALU_RES_IN[10];
  assign DRAM_ADDR_OUT[10] = ALU_RES_IN[10];
  assign OP_MEM[9] = ALU_RES_IN[9];
  assign DRAM_ADDR_OUT[9] = ALU_RES_IN[9];
  assign OP_MEM[8] = ALU_RES_IN[8];
  assign DRAM_ADDR_OUT[8] = ALU_RES_IN[8];
  assign OP_MEM[7] = ALU_RES_IN[7];
  assign DRAM_ADDR_OUT[7] = ALU_RES_IN[7];
  assign OP_MEM[6] = ALU_RES_IN[6];
  assign DRAM_ADDR_OUT[6] = ALU_RES_IN[6];
  assign OP_MEM[5] = ALU_RES_IN[5];
  assign DRAM_ADDR_OUT[5] = ALU_RES_IN[5];
  assign OP_MEM[4] = ALU_RES_IN[4];
  assign DRAM_ADDR_OUT[4] = ALU_RES_IN[4];
  assign OP_MEM[3] = ALU_RES_IN[3];
  assign DRAM_ADDR_OUT[3] = ALU_RES_IN[3];
  assign OP_MEM[2] = ALU_RES_IN[2];
  assign DRAM_ADDR_OUT[2] = ALU_RES_IN[2];
  assign OP_MEM[1] = ALU_RES_IN[1];
  assign DRAM_ADDR_OUT[1] = ALU_RES_IN[1];
  assign OP_MEM[0] = ALU_RES_IN[0];
  assign DRAM_ADDR_OUT[0] = ALU_RES_IN[0];
  assign DRAM_DATA_OUT[31] = B_IN[31];
  assign DRAM_DATA_OUT[30] = B_IN[30];
  assign DRAM_DATA_OUT[29] = B_IN[29];
  assign DRAM_DATA_OUT[28] = B_IN[28];
  assign DRAM_DATA_OUT[27] = B_IN[27];
  assign DRAM_DATA_OUT[26] = B_IN[26];
  assign DRAM_DATA_OUT[25] = B_IN[25];
  assign DRAM_DATA_OUT[24] = B_IN[24];
  assign DRAM_DATA_OUT[23] = B_IN[23];
  assign DRAM_DATA_OUT[22] = B_IN[22];
  assign DRAM_DATA_OUT[21] = B_IN[21];
  assign DRAM_DATA_OUT[20] = B_IN[20];
  assign DRAM_DATA_OUT[19] = B_IN[19];
  assign DRAM_DATA_OUT[18] = B_IN[18];
  assign DRAM_DATA_OUT[17] = B_IN[17];
  assign DRAM_DATA_OUT[16] = B_IN[16];
  assign DRAM_DATA_OUT[15] = B_IN[15];
  assign DRAM_DATA_OUT[14] = B_IN[14];
  assign DRAM_DATA_OUT[13] = B_IN[13];
  assign DRAM_DATA_OUT[12] = B_IN[12];
  assign DRAM_DATA_OUT[11] = B_IN[11];
  assign DRAM_DATA_OUT[10] = B_IN[10];
  assign DRAM_DATA_OUT[9] = B_IN[9];
  assign DRAM_DATA_OUT[8] = B_IN[8];
  assign DRAM_DATA_OUT[7] = B_IN[7];
  assign DRAM_DATA_OUT[6] = B_IN[6];
  assign DRAM_DATA_OUT[5] = B_IN[5];
  assign DRAM_DATA_OUT[4] = B_IN[4];
  assign DRAM_DATA_OUT[3] = B_IN[3];
  assign DRAM_DATA_OUT[2] = B_IN[2];
  assign DRAM_DATA_OUT[1] = B_IN[1];
  assign DRAM_DATA_OUT[0] = B_IN[0];
  assign ADD_WR_MEM[4] = ADD_WR_IN[4];
  assign ADD_WR_MEM[3] = ADD_WR_IN[3];
  assign ADD_WR_MEM[2] = ADD_WR_IN[2];
  assign ADD_WR_MEM[1] = ADD_WR_IN[1];
  assign ADD_WR_MEM[0] = ADD_WR_IN[0];

  regn_N32_2 LMD ( .DIN(DRAM_DATA_IN), .CLK(CLK), .EN(MEM_EN_IN), .RST(RST), 
        .DOUT(DATA_OUT) );
  regn_N5_1 reg0 ( .DIN(ADD_WR_IN), .CLK(CLK), .EN(MEM_EN_IN), .RST(RST), 
        .DOUT(ADD_WR_OUT) );
  regn_N32_1 reg1 ( .DIN(ALU_RES_IN), .CLK(CLK), .EN(MEM_EN_IN), .RST(RST), 
        .DOUT(ALU_RES_OUT) );
  mux41_NBIT32_2 PCsel ( .A(NPC_IN), .B(NPC_REL), .C(NPC_ABS), .D({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(PC_SEL), .Z(PC_OUT) );
endmodule


module Writeback ( WB_MUX_SEL, DATA_IN, ALU_RES_IN, ADD_WR_IN, DATA_OUT, 
        ADD_WR_OUT );
  input [31:0] DATA_IN;
  input [31:0] ALU_RES_IN;
  input [4:0] ADD_WR_IN;
  output [31:0] DATA_OUT;
  output [4:0] ADD_WR_OUT;
  input WB_MUX_SEL;

  assign ADD_WR_OUT[4] = ADD_WR_IN[4];
  assign ADD_WR_OUT[3] = ADD_WR_IN[3];
  assign ADD_WR_OUT[2] = ADD_WR_IN[2];
  assign ADD_WR_OUT[1] = ADD_WR_IN[1];
  assign ADD_WR_OUT[0] = ADD_WR_IN[0];

  mux21_NBIT32_2 WBmux ( .A(DATA_IN), .B(ALU_RES_IN), .S(WB_MUX_SEL), .Z(
        DATA_OUT) );
endmodule


module HazardDetection_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \A[0] , n2;
  wire   [32:0] carry;
  assign DIFF[1] = A[1];
  assign DIFF[0] = \A[0] ;
  assign \A[0]  = A[0];

  OR2_X1 U1 ( .A1(A[4]), .A2(carry[4]), .ZN(carry[5]) );
  OR2_X1 U2 ( .A1(A[5]), .A2(carry[5]), .ZN(carry[6]) );
  OR2_X1 U3 ( .A1(A[6]), .A2(carry[6]), .ZN(carry[7]) );
  OR2_X1 U4 ( .A1(A[7]), .A2(carry[7]), .ZN(carry[8]) );
  OR2_X1 U5 ( .A1(A[8]), .A2(carry[8]), .ZN(carry[9]) );
  OR2_X1 U6 ( .A1(A[9]), .A2(carry[9]), .ZN(carry[10]) );
  OR2_X1 U7 ( .A1(A[10]), .A2(carry[10]), .ZN(carry[11]) );
  OR2_X1 U8 ( .A1(A[11]), .A2(carry[11]), .ZN(carry[12]) );
  OR2_X1 U9 ( .A1(A[12]), .A2(carry[12]), .ZN(carry[13]) );
  OR2_X1 U10 ( .A1(A[13]), .A2(carry[13]), .ZN(carry[14]) );
  OR2_X1 U11 ( .A1(A[14]), .A2(carry[14]), .ZN(carry[15]) );
  OR2_X1 U12 ( .A1(A[15]), .A2(carry[15]), .ZN(carry[16]) );
  OR2_X1 U13 ( .A1(A[16]), .A2(carry[16]), .ZN(carry[17]) );
  OR2_X1 U14 ( .A1(A[17]), .A2(carry[17]), .ZN(carry[18]) );
  OR2_X1 U15 ( .A1(A[18]), .A2(carry[18]), .ZN(carry[19]) );
  OR2_X1 U16 ( .A1(A[19]), .A2(carry[19]), .ZN(carry[20]) );
  OR2_X1 U17 ( .A1(A[20]), .A2(carry[20]), .ZN(carry[21]) );
  OR2_X1 U18 ( .A1(A[21]), .A2(carry[21]), .ZN(carry[22]) );
  OR2_X1 U19 ( .A1(A[22]), .A2(carry[22]), .ZN(carry[23]) );
  OR2_X1 U20 ( .A1(A[23]), .A2(carry[23]), .ZN(carry[24]) );
  OR2_X1 U21 ( .A1(A[24]), .A2(carry[24]), .ZN(carry[25]) );
  OR2_X1 U22 ( .A1(A[25]), .A2(carry[25]), .ZN(carry[26]) );
  OR2_X1 U23 ( .A1(A[26]), .A2(carry[26]), .ZN(carry[27]) );
  OR2_X1 U24 ( .A1(A[27]), .A2(carry[27]), .ZN(carry[28]) );
  OR2_X1 U25 ( .A1(A[28]), .A2(carry[28]), .ZN(carry[29]) );
  OR2_X1 U26 ( .A1(A[29]), .A2(carry[29]), .ZN(carry[30]) );
  OR2_X1 U27 ( .A1(A[3]), .A2(A[2]), .ZN(carry[4]) );
  XNOR2_X1 U28 ( .A(A[4]), .B(carry[4]), .ZN(DIFF[4]) );
  XNOR2_X1 U29 ( .A(A[5]), .B(carry[5]), .ZN(DIFF[5]) );
  XNOR2_X1 U30 ( .A(A[6]), .B(carry[6]), .ZN(DIFF[6]) );
  XNOR2_X1 U31 ( .A(A[7]), .B(carry[7]), .ZN(DIFF[7]) );
  XNOR2_X1 U32 ( .A(A[8]), .B(carry[8]), .ZN(DIFF[8]) );
  XNOR2_X1 U33 ( .A(A[9]), .B(carry[9]), .ZN(DIFF[9]) );
  XNOR2_X1 U34 ( .A(A[10]), .B(carry[10]), .ZN(DIFF[10]) );
  XNOR2_X1 U35 ( .A(A[11]), .B(carry[11]), .ZN(DIFF[11]) );
  XNOR2_X1 U36 ( .A(A[12]), .B(carry[12]), .ZN(DIFF[12]) );
  XNOR2_X1 U37 ( .A(A[13]), .B(carry[13]), .ZN(DIFF[13]) );
  XNOR2_X1 U38 ( .A(A[14]), .B(carry[14]), .ZN(DIFF[14]) );
  XNOR2_X1 U39 ( .A(A[15]), .B(carry[15]), .ZN(DIFF[15]) );
  XNOR2_X1 U40 ( .A(A[16]), .B(carry[16]), .ZN(DIFF[16]) );
  XNOR2_X1 U41 ( .A(A[17]), .B(carry[17]), .ZN(DIFF[17]) );
  XNOR2_X1 U42 ( .A(A[18]), .B(carry[18]), .ZN(DIFF[18]) );
  XNOR2_X1 U43 ( .A(A[19]), .B(carry[19]), .ZN(DIFF[19]) );
  XNOR2_X1 U44 ( .A(A[20]), .B(carry[20]), .ZN(DIFF[20]) );
  XNOR2_X1 U45 ( .A(A[21]), .B(carry[21]), .ZN(DIFF[21]) );
  XNOR2_X1 U46 ( .A(A[22]), .B(carry[22]), .ZN(DIFF[22]) );
  XNOR2_X1 U47 ( .A(A[23]), .B(carry[23]), .ZN(DIFF[23]) );
  XNOR2_X1 U48 ( .A(A[24]), .B(carry[24]), .ZN(DIFF[24]) );
  XNOR2_X1 U49 ( .A(A[25]), .B(carry[25]), .ZN(DIFF[25]) );
  XNOR2_X1 U50 ( .A(A[26]), .B(carry[26]), .ZN(DIFF[26]) );
  XNOR2_X1 U51 ( .A(A[27]), .B(carry[27]), .ZN(DIFF[27]) );
  XNOR2_X1 U52 ( .A(A[28]), .B(carry[28]), .ZN(DIFF[28]) );
  XNOR2_X1 U53 ( .A(A[29]), .B(carry[29]), .ZN(DIFF[29]) );
  XNOR2_X1 U54 ( .A(A[30]), .B(carry[30]), .ZN(DIFF[30]) );
  XOR2_X1 U55 ( .A(A[31]), .B(n2), .Z(DIFF[31]) );
  NOR2_X1 U56 ( .A1(A[30]), .A2(carry[30]), .ZN(n2) );
  XNOR2_X1 U57 ( .A(A[3]), .B(A[2]), .ZN(DIFF[3]) );
  INV_X1 U58 ( .A(A[2]), .ZN(DIFF[2]) );
endmodule


module HazardDetection ( RST, ADD_RS1, ADD_RS2, ADD_WR, DRAM_R, INS_IN, PC_IN, 
        Bubble, HDU_INS_OUT, HDU_PC_OUT, HDU_NPC_OUT );
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [4:0] ADD_WR;
  input [31:0] INS_IN;
  input [31:0] PC_IN;
  output [31:0] HDU_INS_OUT;
  output [31:0] HDU_PC_OUT;
  output [31:0] HDU_NPC_OUT;
  input RST, DRAM_R;
  output Bubble;
  wire   n4, n5, n6, n9, n10, n12, n13, n14, n15, n16, n17, n18, n19;
  assign HDU_INS_OUT[31] = INS_IN[31];
  assign HDU_INS_OUT[30] = INS_IN[30];
  assign HDU_INS_OUT[29] = INS_IN[29];
  assign HDU_INS_OUT[28] = INS_IN[28];
  assign HDU_INS_OUT[27] = INS_IN[27];
  assign HDU_INS_OUT[26] = INS_IN[26];
  assign HDU_INS_OUT[25] = INS_IN[25];
  assign HDU_INS_OUT[24] = INS_IN[24];
  assign HDU_INS_OUT[23] = INS_IN[23];
  assign HDU_INS_OUT[22] = INS_IN[22];
  assign HDU_INS_OUT[21] = INS_IN[21];
  assign HDU_INS_OUT[20] = INS_IN[20];
  assign HDU_INS_OUT[19] = INS_IN[19];
  assign HDU_INS_OUT[18] = INS_IN[18];
  assign HDU_INS_OUT[17] = INS_IN[17];
  assign HDU_INS_OUT[16] = INS_IN[16];
  assign HDU_INS_OUT[15] = INS_IN[15];
  assign HDU_INS_OUT[14] = INS_IN[14];
  assign HDU_INS_OUT[13] = INS_IN[13];
  assign HDU_INS_OUT[12] = INS_IN[12];
  assign HDU_INS_OUT[11] = INS_IN[11];
  assign HDU_INS_OUT[10] = INS_IN[10];
  assign HDU_INS_OUT[9] = INS_IN[9];
  assign HDU_INS_OUT[8] = INS_IN[8];
  assign HDU_INS_OUT[7] = INS_IN[7];
  assign HDU_INS_OUT[6] = INS_IN[6];
  assign HDU_INS_OUT[5] = INS_IN[5];
  assign HDU_INS_OUT[4] = INS_IN[4];
  assign HDU_INS_OUT[3] = INS_IN[3];
  assign HDU_INS_OUT[2] = INS_IN[2];
  assign HDU_INS_OUT[1] = INS_IN[1];
  assign HDU_INS_OUT[0] = INS_IN[0];
  assign HDU_NPC_OUT[31] = PC_IN[31];
  assign HDU_NPC_OUT[30] = PC_IN[30];
  assign HDU_NPC_OUT[29] = PC_IN[29];
  assign HDU_NPC_OUT[28] = PC_IN[28];
  assign HDU_NPC_OUT[27] = PC_IN[27];
  assign HDU_NPC_OUT[26] = PC_IN[26];
  assign HDU_NPC_OUT[25] = PC_IN[25];
  assign HDU_NPC_OUT[24] = PC_IN[24];
  assign HDU_NPC_OUT[23] = PC_IN[23];
  assign HDU_NPC_OUT[22] = PC_IN[22];
  assign HDU_NPC_OUT[21] = PC_IN[21];
  assign HDU_NPC_OUT[20] = PC_IN[20];
  assign HDU_NPC_OUT[19] = PC_IN[19];
  assign HDU_NPC_OUT[18] = PC_IN[18];
  assign HDU_NPC_OUT[17] = PC_IN[17];
  assign HDU_NPC_OUT[16] = PC_IN[16];
  assign HDU_NPC_OUT[15] = PC_IN[15];
  assign HDU_NPC_OUT[14] = PC_IN[14];
  assign HDU_NPC_OUT[13] = PC_IN[13];
  assign HDU_NPC_OUT[12] = PC_IN[12];
  assign HDU_NPC_OUT[11] = PC_IN[11];
  assign HDU_NPC_OUT[10] = PC_IN[10];
  assign HDU_NPC_OUT[9] = PC_IN[9];
  assign HDU_NPC_OUT[8] = PC_IN[8];
  assign HDU_NPC_OUT[7] = PC_IN[7];
  assign HDU_NPC_OUT[6] = PC_IN[6];
  assign HDU_NPC_OUT[5] = PC_IN[5];
  assign HDU_NPC_OUT[4] = PC_IN[4];
  assign HDU_NPC_OUT[3] = PC_IN[3];
  assign HDU_NPC_OUT[2] = PC_IN[2];
  assign HDU_NPC_OUT[1] = PC_IN[1];
  assign HDU_NPC_OUT[0] = PC_IN[0];

  OAI33_X1 U16 ( .A1(n5), .A2(n6), .A3(n9), .B1(n10), .B2(n12), .B3(n13), .ZN(
        n4) );
  XOR2_X1 U17 ( .A(ADD_WR[4]), .B(ADD_RS2[4]), .Z(n13) );
  XOR2_X1 U18 ( .A(ADD_WR[2]), .B(ADD_RS2[2]), .Z(n12) );
  NAND3_X1 U19 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n10) );
  XOR2_X1 U20 ( .A(ADD_WR[4]), .B(ADD_RS1[4]), .Z(n9) );
  XOR2_X1 U21 ( .A(ADD_WR[2]), .B(ADD_RS1[2]), .Z(n6) );
  NAND3_X1 U22 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n5) );
  HazardDetection_DW01_sub_0 sub_25 ( .A(PC_IN), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .DIFF(HDU_PC_OUT) );
  AND3_X1 U3 ( .A1(DRAM_R), .A2(n4), .A3(RST), .ZN(Bubble) );
  XNOR2_X1 U7 ( .A(ADD_WR[3]), .B(ADD_RS1[3]), .ZN(n17) );
  XNOR2_X1 U8 ( .A(ADD_WR[3]), .B(ADD_RS2[3]), .ZN(n14) );
  XNOR2_X1 U9 ( .A(ADD_WR[0]), .B(ADD_RS1[0]), .ZN(n18) );
  XNOR2_X1 U10 ( .A(ADD_WR[0]), .B(ADD_RS2[0]), .ZN(n15) );
  XNOR2_X1 U11 ( .A(ADD_WR[1]), .B(ADD_RS1[1]), .ZN(n19) );
  XNOR2_X1 U12 ( .A(ADD_WR[1]), .B(ADD_RS2[1]), .ZN(n16) );
endmodule


module Datapath ( CLK, RST, INS_IN, DATA_IN, REG_LATCH_EN, RD1, RD2, MUX_A_SEL, 
        MUX_B_SEL, .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , 
        \ALU_OPC[0] }), ALU_OUTREG_EN, JUMP_TYPE, DRAM_R_IN, MEM_EN_IN, 
        DRAM_W_IN, RF_WE, DRAM_EN_IN, WB_MUX_SEL, INS_OUT, IRAM_ADDR_OUT, 
        DRAM_ADDR_OUT, DATA_OUT, DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, 
        Bubble_out );
  input [31:0] INS_IN;
  input [31:0] DATA_IN;
  input [1:0] MUX_B_SEL;
  input [1:0] JUMP_TYPE;
  output [31:0] INS_OUT;
  output [31:0] IRAM_ADDR_OUT;
  output [31:0] DRAM_ADDR_OUT;
  output [31:0] DATA_OUT;
  input CLK, RST, REG_LATCH_EN, RD1, RD2, MUX_A_SEL, \ALU_OPC[3] ,
         \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] , ALU_OUTREG_EN, DRAM_R_IN,
         MEM_EN_IN, DRAM_W_IN, RF_WE, DRAM_EN_IN, WB_MUX_SEL;
  output DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble_out;
  wire   ZERO_FLAG_EX, RF_WE_WB, DRAM_R_MEM;
  wire   [3:0] ALU_OPC;
  wire   [31:0] PC_MEM_OUT;
  wire   [31:0] sig_HDU_INS_OUT;
  wire   [31:0] sig_HDU_PC_OUT;
  wire   [31:0] sig_HDU_NPC_OUT;
  wire   [31:0] PC_FETCH_OUT;
  wire   [31:0] NPC_FETCH_OUT;
  wire   [4:0] ADD_WR_WB;
  wire   [31:0] OP_WB;
  wire   [31:0] PC_DECODE_OUT;
  wire   [31:0] A_DECODE_OUT;
  wire   [31:0] B_DECODE_OUT;
  wire   [31:0] IMM_DECODE_OUT;
  wire   [4:0] ADD_RS1_HDU;
  wire   [4:0] ADD_RS2_HDU;
  wire   [4:0] ADD_WR_DECODE_OUT;
  wire   [4:0] ADD_RS1_DECODE_OUT;
  wire   [4:0] ADD_RS2_DECODE_OUT;
  wire   [4:0] ADD_WR_MEM;
  wire   [31:0] OP_MEM;
  wire   [1:0] PC_SEL_EX;
  wire   [31:0] NPC_ABS_EX;
  wire   [31:0] NPC_REL_EX;
  wire   [31:0] ALU_RES_EX;
  wire   [31:0] B_EX_OUT;
  wire   [4:0] ADD_WR_EX_OUT;
  wire   [31:0] DATA_MEM_OUT;
  wire   [31:0] ALU_RES_MEM;
  wire   [4:0] ADD_WR_MEM_OUT;

  Fetch FetchStage ( .CLK(CLK), .RST(RST), .ZERO_FLAG(ZERO_FLAG_EX), .PC_EXT(
        PC_MEM_OUT), .INS_IN(INS_IN), .Bubble_in(Bubble_out), .HDU_INS_IN(
        sig_HDU_INS_OUT), .HDU_PC_IN(sig_HDU_PC_OUT), .HDU_NPC_IN(
        sig_HDU_NPC_OUT), .PC_OUT(PC_FETCH_OUT), .ADDR_OUT(IRAM_ADDR_OUT), 
        .NPC_OUT(NPC_FETCH_OUT), .INS_OUT(INS_OUT) );
  Decode DecodeStage ( .CLK(CLK), .RST(RST), .REG_LATCH_EN(REG_LATCH_EN), 
        .RD1(RD1), .RD2(RD2), .RF_WE(RF_WE_WB), .ZERO_FLAG(ZERO_FLAG_EX), 
        .PC_IN(PC_FETCH_OUT), .INS_IN(INS_OUT), .ADD_WR(ADD_WR_WB), 
        .DATA_WR_IN(OP_WB), .PC_OUT(PC_DECODE_OUT), .A_OUT(A_DECODE_OUT), 
        .B_OUT(B_DECODE_OUT), .IMM_OUT(IMM_DECODE_OUT), .ADD_RS1_HDU(
        ADD_RS1_HDU), .ADD_RS2_HDU(ADD_RS2_HDU), .ADD_WR_OUT(ADD_WR_DECODE_OUT), .ADD_RS1_OUT(ADD_RS1_DECODE_OUT), .ADD_RS2_OUT(ADD_RS2_DECODE_OUT) );
  Execute ExecuteStage ( .CLK(CLK), .RST(RST), .MUX_A_SEL(MUX_A_SEL), 
        .MUX_B_SEL(MUX_B_SEL), .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , 
        \ALU_OPC[1] , \ALU_OPC[0] }), .ALU_OUTREG_EN(ALU_OUTREG_EN), 
        .JUMP_TYPE(JUMP_TYPE), .PC_IN(PC_DECODE_OUT), .A_IN(A_DECODE_OUT), 
        .B_IN(B_DECODE_OUT), .IMM_IN(IMM_DECODE_OUT), .ADD_WR_IN(
        ADD_WR_DECODE_OUT), .ADD_RS1_IN(ADD_RS1_DECODE_OUT), .ADD_RS2_IN(
        ADD_RS2_DECODE_OUT), .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_WB(ADD_WR_WB), 
        .RF_WE_MEM(RF_WE), .RF_WE_WB(RF_WE_WB), .OP_MEM(OP_MEM), .OP_WB(OP_WB), 
        .PC_SEL(PC_SEL_EX), .ZERO_FLAG(ZERO_FLAG_EX), .NPC_ABS(NPC_ABS_EX), 
        .NPC_REL(NPC_REL_EX), .ALU_RES(ALU_RES_EX), .B_OUT(B_EX_OUT), 
        .ADD_WR_OUT(ADD_WR_EX_OUT) );
  ff_0 DRAM_R_ff ( .D(DRAM_R_IN), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(
        DRAM_R_MEM) );
  Memory MemoryStage ( .CLK(CLK), .RST(RST), .MEM_EN_IN(MEM_EN_IN), 
        .DRAM_R_IN(DRAM_R_MEM), .DRAM_W_IN(DRAM_W_IN), .DRAM_EN_IN(DRAM_EN_IN), 
        .PC_SEL(PC_SEL_EX), .NPC_IN(NPC_FETCH_OUT), .NPC_ABS(NPC_ABS_EX), 
        .NPC_REL(NPC_REL_EX), .ALU_RES_IN(ALU_RES_EX), .B_IN(B_EX_OUT), 
        .ADD_WR_IN(ADD_WR_EX_OUT), .DRAM_DATA_IN(DATA_IN), .PC_OUT(PC_MEM_OUT), 
        .DRAM_EN_OUT(DRAM_EN_OUT), .DRAM_R_OUT(DRAM_R_OUT), .DRAM_W_OUT(
        DRAM_W_OUT), .DRAM_ADDR_OUT(DRAM_ADDR_OUT), .DRAM_DATA_OUT(DATA_OUT), 
        .DATA_OUT(DATA_MEM_OUT), .ALU_RES_OUT(ALU_RES_MEM), .OP_MEM(OP_MEM), 
        .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_OUT(ADD_WR_MEM_OUT) );
  ff_2 RF_WE_ff ( .D(RF_WE), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(RF_WE_WB) );
  Writeback WritebackStage ( .WB_MUX_SEL(WB_MUX_SEL), .DATA_IN(DATA_MEM_OUT), 
        .ALU_RES_IN(ALU_RES_MEM), .ADD_WR_IN(ADD_WR_MEM_OUT), .DATA_OUT(OP_WB), 
        .ADD_WR_OUT(ADD_WR_WB) );
  HazardDetection HDU ( .RST(RST), .ADD_RS1(ADD_RS1_HDU), .ADD_RS2(ADD_RS2_HDU), .ADD_WR(ADD_WR_DECODE_OUT), .DRAM_R(DRAM_R_IN), .INS_IN(INS_OUT), .PC_IN(
        PC_FETCH_OUT), .Bubble(Bubble_out), .HDU_INS_OUT(sig_HDU_INS_OUT), 
        .HDU_PC_OUT(sig_HDU_PC_OUT), .HDU_NPC_OUT(sig_HDU_NPC_OUT) );
endmodule


module hardwired_cu_NBIT32 ( REG_LATCH_EN, RD1, RD2, MUX_A_SEL, MUX_B_SEL, 
    .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), 
        ALU_OUTREG_EN, DRAM_R_IN, JUMP_TYPE, MEM_EN_IN, DRAM_W_IN, RF_WE, 
        DRAM_EN_IN, WB_MUX_SEL, INS_IN, Bubble, Clk, Rst );
  output [1:0] MUX_B_SEL;
  output [1:0] JUMP_TYPE;
  input [31:0] INS_IN;
  input Bubble, Clk, Rst;
  output REG_LATCH_EN, RD1, RD2, MUX_A_SEL, \ALU_OPC[3] , \ALU_OPC[2] ,
         \ALU_OPC[1] , \ALU_OPC[0] , ALU_OUTREG_EN, DRAM_R_IN, MEM_EN_IN,
         DRAM_W_IN, RF_WE, DRAM_EN_IN, WB_MUX_SEL;
  wire   INS_IN_31, INS_IN_30, INS_IN_29, INS_IN_28, INS_IN_27, INS_IN_26, N24,
         N25, N26, N27, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76;
  wire   [3:0] ALU_OPC;
  wire   [3:0] AluOP_E;
  assign REG_LATCH_EN = 1'b0;
  assign RD1 = 1'b0;
  assign RD2 = 1'b0;
  assign MUX_A_SEL = 1'b0;
  assign MUX_B_SEL[1] = 1'b0;
  assign MUX_B_SEL[0] = 1'b0;
  assign ALU_OUTREG_EN = 1'b0;
  assign DRAM_R_IN = 1'b0;
  assign JUMP_TYPE[1] = 1'b0;
  assign JUMP_TYPE[0] = 1'b0;
  assign MEM_EN_IN = 1'b0;
  assign DRAM_W_IN = 1'b0;
  assign RF_WE = 1'b0;
  assign DRAM_EN_IN = 1'b0;
  assign WB_MUX_SEL = 1'b0;
  assign INS_IN_31 = INS_IN[31];
  assign INS_IN_30 = INS_IN[30];
  assign INS_IN_29 = INS_IN[29];
  assign INS_IN_28 = INS_IN[28];
  assign INS_IN_27 = INS_IN[27];
  assign INS_IN_26 = INS_IN[26];

  DFFR_X1 \AluOP_E_reg[3]  ( .D(N27), .CK(Clk), .RN(Rst), .Q(AluOP_E[3]) );
  DFFR_X1 \ALU_OPC_reg[3]  ( .D(AluOP_E[3]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[3]) );
  DFFR_X1 \AluOP_E_reg[2]  ( .D(N26), .CK(Clk), .RN(Rst), .Q(AluOP_E[2]) );
  DFFR_X1 \ALU_OPC_reg[2]  ( .D(AluOP_E[2]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[2]) );
  DFFR_X1 \AluOP_E_reg[1]  ( .D(N25), .CK(Clk), .RN(Rst), .Q(AluOP_E[1]) );
  DFFR_X1 \ALU_OPC_reg[1]  ( .D(AluOP_E[1]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[1]) );
  DFFR_X1 \AluOP_E_reg[0]  ( .D(N24), .CK(Clk), .RN(Rst), .Q(AluOP_E[0]) );
  DFFR_X1 \ALU_OPC_reg[0]  ( .D(AluOP_E[0]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[0]) );
  XOR2_X1 U73 ( .A(INS_IN[1]), .B(INS_IN[0]), .Z(n25) );
  NAND3_X1 U74 ( .A1(n37), .A2(n38), .A3(n61), .ZN(n27) );
  NAND3_X1 U75 ( .A1(n39), .A2(INS_IN_30), .A3(n40), .ZN(n37) );
  NAND3_X1 U76 ( .A1(n43), .A2(n26), .A3(INS_IN_30), .ZN(n30) );
  NAND3_X1 U77 ( .A1(n63), .A2(n66), .A3(n24), .ZN(n31) );
  OAI33_X1 U78 ( .A1(n53), .A2(n71), .A3(n73), .B1(n54), .B2(INS_IN[1]), .B3(
        n55), .ZN(n20) );
  NAND3_X1 U79 ( .A1(n43), .A2(n75), .A3(INS_IN_28), .ZN(n52) );
  NAND3_X1 U80 ( .A1(n73), .A2(n75), .A3(n43), .ZN(n42) );
  INV_X1 U18 ( .A(n36), .ZN(n62) );
  OAI22_X1 U19 ( .A1(n73), .A2(n30), .B1(n41), .B2(n42), .ZN(n35) );
  AOI21_X1 U20 ( .B1(n39), .B2(n74), .A(n20), .ZN(n36) );
  NOR2_X1 U21 ( .A1(n41), .A2(n52), .ZN(n29) );
  INV_X1 U22 ( .A(n40), .ZN(n72) );
  INV_X1 U23 ( .A(n30), .ZN(n69) );
  INV_X1 U24 ( .A(n52), .ZN(n74) );
  INV_X1 U25 ( .A(n39), .ZN(n71) );
  INV_X1 U26 ( .A(n26), .ZN(n67) );
  INV_X1 U27 ( .A(n56), .ZN(n61) );
  OAI21_X1 U28 ( .B1(n65), .B2(n38), .A(n57), .ZN(n56) );
  OR3_X1 U29 ( .A1(n72), .A2(n75), .A3(n41), .ZN(n57) );
  INV_X1 U30 ( .A(n28), .ZN(n68) );
  AOI21_X1 U31 ( .B1(n73), .B2(n69), .A(n29), .ZN(n28) );
  NAND2_X1 U32 ( .A1(INS_IN[5]), .A2(INS_IN[3]), .ZN(n54) );
  NAND2_X1 U33 ( .A1(INS_IN_30), .A2(n43), .ZN(n53) );
  NOR4_X1 U34 ( .A1(INS_IN[6]), .A2(INS_IN[4]), .A3(INS_IN[10]), .A4(n59), 
        .ZN(n46) );
  OR3_X1 U35 ( .A1(INS_IN[9]), .A2(INS_IN[8]), .A3(INS_IN[7]), .ZN(n59) );
  NOR3_X1 U36 ( .A1(INS_IN_29), .A2(INS_IN_31), .A3(n73), .ZN(n40) );
  NOR2_X1 U37 ( .A1(INS_IN_27), .A2(INS_IN_26), .ZN(n39) );
  OAI221_X1 U38 ( .B1(n64), .B2(n31), .C1(Bubble), .C2(n32), .A(n33), .ZN(N25)
         );
  INV_X1 U39 ( .A(n44), .ZN(n64) );
  OAI211_X1 U40 ( .C1(INS_IN[3]), .C2(n63), .A(n65), .B(n34), .ZN(n33) );
  NOR3_X1 U41 ( .A1(n35), .A2(n27), .A3(n62), .ZN(n32) );
  OAI221_X1 U42 ( .B1(INS_IN[2]), .B2(n19), .C1(Bubble), .C2(n22), .A(n23), 
        .ZN(N26) );
  NAND4_X1 U43 ( .A1(n24), .A2(INS_IN[2]), .A3(n25), .A4(n66), .ZN(n23) );
  AOI211_X1 U44 ( .C1(n74), .C2(n26), .A(n68), .B(n27), .ZN(n22) );
  OAI22_X1 U45 ( .A1(INS_IN_29), .A2(INS_IN_31), .B1(n76), .B2(INS_IN_30), 
        .ZN(n51) );
  NOR2_X1 U46 ( .A1(n70), .A2(INS_IN_27), .ZN(n26) );
  NOR3_X1 U47 ( .A1(n72), .A2(INS_IN_30), .A3(n67), .ZN(n49) );
  INV_X1 U48 ( .A(INS_IN_28), .ZN(n73) );
  NAND4_X1 U49 ( .A1(INS_IN[2]), .A2(n46), .A3(n47), .A4(n63), .ZN(n55) );
  OAI22_X1 U50 ( .A1(Bubble), .A2(n45), .B1(n44), .B2(n31), .ZN(N24) );
  NOR4_X1 U51 ( .A1(n48), .A2(n49), .A3(n29), .A4(n50), .ZN(n45) );
  AND4_X1 U52 ( .A1(n73), .A2(n51), .A3(INS_IN_26), .A4(INS_IN_27), .ZN(n50)
         );
  OAI211_X1 U53 ( .C1(n71), .C2(n42), .A(n61), .B(n36), .ZN(n48) );
  NOR2_X1 U54 ( .A1(n65), .A2(INS_IN[2]), .ZN(n44) );
  NAND4_X1 U55 ( .A1(INS_IN[0]), .A2(n24), .A3(INS_IN[3]), .A4(n65), .ZN(n19)
         );
  INV_X1 U56 ( .A(INS_IN[1]), .ZN(n65) );
  NAND2_X1 U57 ( .A1(INS_IN_27), .A2(n70), .ZN(n41) );
  AND2_X1 U58 ( .A1(INS_IN_29), .A2(n76), .ZN(n43) );
  AND3_X1 U59 ( .A1(n39), .A2(n73), .A3(n58), .ZN(n47) );
  NOR3_X1 U60 ( .A1(INS_IN_29), .A2(INS_IN_31), .A3(INS_IN_30), .ZN(n58) );
  AND4_X1 U61 ( .A1(INS_IN[5]), .A2(n46), .A3(n47), .A4(n60), .ZN(n24) );
  INV_X1 U62 ( .A(Bubble), .ZN(n60) );
  OAI21_X1 U63 ( .B1(Bubble), .B2(n18), .A(n19), .ZN(N27) );
  NOR3_X1 U64 ( .A1(n20), .A2(n69), .A3(n21), .ZN(n18) );
  AOI211_X1 U65 ( .C1(n71), .C2(n67), .A(n72), .B(INS_IN_30), .ZN(n21) );
  INV_X1 U66 ( .A(INS_IN[0]), .ZN(n63) );
  OR3_X1 U67 ( .A1(INS_IN[3]), .A2(INS_IN[5]), .A3(n55), .ZN(n38) );
  INV_X1 U68 ( .A(INS_IN_30), .ZN(n75) );
  INV_X1 U69 ( .A(INS_IN_26), .ZN(n70) );
  INV_X1 U70 ( .A(INS_IN[3]), .ZN(n66) );
  INV_X1 U71 ( .A(INS_IN_31), .ZN(n76) );
  AND2_X1 U72 ( .A1(INS_IN[2]), .A2(n24), .ZN(n34) );
endmodule


module DLX ( Clk, Rst );
  input Clk, Rst;
  wire   DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble;
  wire   [31:0] INS_IN;
  wire   [31:0] DATA_IN;
  wire   [1:0] MUX_B_SEL;
  wire   [3:0] ALU_OPC;
  wire   [1:0] JUMP_TYPE;
  wire   [31:0] IRAM_ADDR_OUT;
  wire   [31:0] DRAM_ADDR_OUT;
  wire   [31:0] DATA_OUT;

  Datapath DP ( .CLK(Clk), .RST(Rst), .INS_IN(INS_IN), .DATA_IN(DATA_IN), 
        .REG_LATCH_EN(1'b0), .RD1(1'b0), .RD2(1'b0), .MUX_A_SEL(1'b0), 
        .MUX_B_SEL({1'b0, 1'b0}), .ALU_OPC(ALU_OPC), .ALU_OUTREG_EN(1'b0), 
        .JUMP_TYPE({1'b0, 1'b0}), .DRAM_R_IN(1'b0), .MEM_EN_IN(1'b0), 
        .DRAM_W_IN(1'b0), .RF_WE(1'b0), .DRAM_EN_IN(1'b0), .WB_MUX_SEL(1'b0), 
        .IRAM_ADDR_OUT(IRAM_ADDR_OUT), .DRAM_ADDR_OUT(DRAM_ADDR_OUT), 
        .DATA_OUT(DATA_OUT), .DRAM_EN_OUT(DRAM_EN_OUT), .DRAM_R_OUT(DRAM_R_OUT), .DRAM_W_OUT(DRAM_W_OUT), .Bubble_out(Bubble) );
  hardwired_cu_NBIT32 CU ( .ALU_OPC(ALU_OPC), .INS_IN(INS_IN), .Bubble(Bubble), 
        .Clk(Clk), .Rst(Rst) );
  IRAM IRAM_I ( .Rst(Rst), .Addr(IRAM_ADDR_OUT), .Iout(INS_IN) );
  DRAM DRAM_I ( .En(DRAM_EN_OUT), .Rst(Rst), .ADDR_IN(DRAM_ADDR_OUT), 
        .DATA_IN(DATA_OUT), .DRAM_W(DRAM_W_OUT), .DRAM_R(DRAM_R_OUT), 
        .DATA_OUT(DATA_IN) );
endmodule

