library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;
use work.constants.all;

entity tb_RF is
end entity;

architecture test of tb_RF is

component register_file is
 generic( NBIT_ADD: integer;
		  NBIT_DATA: integer);
 port ( CLK: 		IN std_logic;
        RESET:  	IN std_logic;
	ENABLE: 	IN std_logic;
        RD1:            IN std_logic;
        RD2:            IN std_logic; 
        WR: 		IN std_logic;
        ADD_WR: 	IN std_logic_vector(NBIT_ADD-1 downto 0);
        ADD_RD1: 	IN std_logic_vector(NBIT_ADD-1 downto 0);
        ADD_RD2: 	IN std_logic_vector(NBIT_ADD-1 downto 0);
        DATAIN: 	IN std_logic_vector(NBIT_DATA-1 downto 0);
        OUT1: 		OUT std_logic_vector(NBIT_DATA-1 downto 0);
        OUT2: 		OUT std_logic_vector(NBIT_DATA-1 downto 0));
end component;

  constant tb_period : time := 30ns;
  constant tb_clk    : time := 10ns;

  signal      CLK: 	std_logic;

  signal      RESET:  	std_logic;
  signal      ENABLE:   std_logic;
  signal      RD1:      std_logic;
  signal      RD2:      std_logic;
  signal      WR:       std_logic;
  signal      ADD_WR: 	std_logic_vector(NBIT_ADD-1 downto 0);
  signal      ADD_RD1: 	std_logic_vector(NBIT_ADD-1 downto 0);
  signal      ADD_RD2: 	std_logic_vector(NBIT_ADD-1 downto 0);
  signal      DATAIN: 	std_logic_vector(NBIT_DATA-1 downto 0);

  signal      OUT1:     std_logic_vector(NBIT_DATA-1 downto 0);
  signal      OUT2:     std_logic_vector(NBIT_DATA-1 downto 0);

begin

  DUT : register_file
    generic map (NBIT_ADD => 5,
                 NBIT_DATA => 32)
    port map(
                 CLK => CLK,
                 RESET => RESET,
                 ENABLE => ENABLE,
                 RD1 => RD1,
                 RD2 => RD2,
                 WR => WR,
                 ADD_WR => ADD_WR,
                 ADD_RD1 => ADD_RD1,
                 ADD_RD2 => ADD_RD2,
                 DATAIN => DATAIN,
                 OUT1 => OUT1,
                 OUT2 => OUT2
                );

  

  stimuli : process

                procedure apply_stimuli (
                         constant      RESET_val:    in std_logic;
                         constant      ENABLE_val:   in std_logic;
                         constant      RD1_val:          in std_logic;
                         constant      RD2_val:          in std_logic;
                         constant      WR_val:       in std_logic;
                         constant      ADD_WR_val:   in integer;
                         constant      ADD_RD1_val:  in integer;
                         constant      ADD_RD2_val:  in integer;
                         constant      DATAIN_val:   in integer;

                         signal      RESET:    out std_logic;
                         signal      ENABLE:   out std_logic;
                         signal      RD1:      out std_logic;
                         signal      RD2:      out std_logic;
                         signal      WR:       out std_logic;
                         signal      ADD_WR:   out std_logic_vector(NBIT_ADD-1 downto 0);
                         signal      ADD_RD1:  out std_logic_vector(NBIT_ADD-1 downto 0);
                         signal      ADD_RD2:  out std_logic_vector(NBIT_ADD-1 downto 0);
                         signal      DATAIN:   out std_logic_vector(NBIT_DATA-1 downto 0)) is
                begin

                        RESET <= RESET_val;
                        ENABLE <= ENABLE_val;
                        RD1 <= RD1_val;
                        RD2 <= RD2_val;
                        WR <= WR_val;
                        ADD_WR <= conv_std_logic_vector(ADD_WR_val, NBIT_ADD);
                        ADD_RD1 <= conv_std_logic_vector(ADD_RD1_val, NBIT_ADD);
                        ADD_RD2 <= conv_std_logic_vector(ADD_RD2_val, NBIT_ADD);
                        DATAIN <= conv_std_logic_vector(DATAIN_val, NBIT_DATA);

                        wait for tb_period;
                       
                end apply_stimuli;

                
  begin

   --apply_stimuli(input values, signals);

    -- perform RESET (active low)
    apply_stimuli('0','1','1','1','1',0,0,0,0, RESET, ENABLE, RD1, RD2, WR, ADD_WR, ADD_RD1, ADD_RD2, DATAIN);
    
    -- apply stimuli
    apply_stimuli('1','1','1','1','1',2,0,0,7, RESET, ENABLE, RD1, RD2, WR, ADD_WR, ADD_RD1, ADD_RD2, DATAIN);
    apply_stimuli('1','1','1','1','0',2,2,0,9, RESET, ENABLE, RD1, RD2, WR, ADD_WR, ADD_RD1, ADD_RD2, DATAIN);
    
    apply_stimuli('1','1','1','1','1',5,9,0,23, RESET, ENABLE, RD1, RD2, WR, ADD_WR, ADD_RD1, ADD_RD2, DATAIN);
  
  end process;

  CLK_process : process

    begin

      CLK <= '0';

      wait for tb_clk;

      CLK <= '1';

      wait for tb_clk;
      
  end process;

end test;
