
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type VHDLOUT_TYPE is range 0 to 5;
type aluOp is (NOP, ADDS, SUBS, ANDS, ORS, XORS, SLLS, SRLS, BEQZS, BNEZS, 
   SGES, SLES, NEQS);
attribute ENUM_ENCODING of aluOp : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010 1011 1100";
   
   -- Declarations for conversion functions.
   function integer_to_unsigned(arg, size : in INTEGER) return std_logic_vector
               ;
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 4 )) 
               return aluOp;
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX;

package body CONV_PACK_DLX is
   
   -- integer type to std_logic_vector function
   function integer_to_unsigned(arg, size : in INTEGER) return std_logic_vector
   is 
      variable result: std_logic_vector(size-1 downto 0);
      variable temp: INTEGER;
      -- synopsys built_in SYN_INTEGER_TO_UNSIGNED
   begin
      temp := arg;
      for i in 0 to size-1 loop
         if (temp mod 2) = 1 then
            result(i) := '1';
         else
            result(i) := '0';
         end if;
         temp := temp / 2;
      end loop;
      return result;
   end;
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 4 )) 
   return aluOp is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "0000" => return NOP;
         when "0001" => return ADDS;
         when "0010" => return SUBS;
         when "0011" => return ANDS;
         when "0100" => return ORS;
         when "0101" => return XORS;
         when "0110" => return SLLS;
         when "0111" => return SRLS;
         when "1000" => return BEQZS;
         when "1001" => return BNEZS;
         when "1010" => return SGES;
         when "1011" => return SLES;
         when "1100" => return NEQS;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "0000";
         when ADDS => return "0001";
         when SUBS => return "0010";
         when ANDS => return "0011";
         when ORS => return "0100";
         when XORS => return "0101";
         when SLLS => return "0110";
         when SRLS => return "0111";
         when BEQZS => return "1000";
         when BNEZS => return "1001";
         when SGES => return "1010";
         when SLES => return "1011";
         when NEQS => return "1100";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Fetch_DW01_add_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Fetch_DW01_add_1;

architecture SYN_cla of Fetch_DW01_add_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
      n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53
      , n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
      SUM_2_port, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, 
      n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95
      , n96, n97, n98, n99 : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U2 : AND2_X1 port map( A1 => n11, A2 => n42, ZN => n36);
   U3 : AND2_X1 port map( A1 => n54, A2 => n92, ZN => n49);
   U4 : AND3_X1 port map( A1 => A(11), A2 => A(13), A3 => A(12), ZN => n1);
   U5 : AND2_X1 port map( A1 => A(25), A2 => A(24), ZN => n2);
   U6 : AND3_X1 port map( A1 => n12, A2 => A(14), A3 => A(15), ZN => n3);
   U7 : NOR2_X1 port map( A1 => n27, A2 => n70, ZN => n4);
   U8 : AND2_X1 port map( A1 => n10, A2 => n42, ZN => n5);
   U9 : AND4_X1 port map( A1 => A(25), A2 => A(24), A3 => n10, A4 => n42, ZN =>
                           n73);
   U10 : AND3_X1 port map( A1 => n37, A2 => n14, A3 => n4, ZN => n30);
   U11 : NOR2_X1 port map( A1 => n95, A2 => n94, ZN => n52);
   U12 : AND4_X1 port map( A1 => A(26), A2 => n22, A3 => n5, A4 => n2, ZN => 
                           n72);
   U13 : AND4_X1 port map( A1 => n83, A2 => n84, A3 => A(16), A4 => A(17), ZN 
                           => n47);
   U14 : AND4_X1 port map( A1 => n67, A2 => n34, A3 => n36, A4 => A(30), ZN => 
                           n15);
   U15 : AND3_X1 port map( A1 => n54, A2 => n92, A3 => A(13), ZN => n90);
   U16 : AND3_X2 port map( A1 => n23, A2 => n3, A3 => n1, ZN => n22);
   U17 : XOR2_X1 port map( A => A(25), B => n51, Z => SUM_25_port);
   U18 : AND3_X1 port map( A1 => n14, A2 => n36, A3 => n6, ZN => n41);
   U19 : INV_X1 port map( A => n27, ZN => n6);
   U20 : NAND4_X1 port map( A1 => A(10), A2 => A(6), A3 => A(8), A4 => A(9), ZN
                           => n87);
   U21 : BUF_X1 port map( A => A(6), Z => n7);
   U22 : AND2_X1 port map( A1 => A(22), A2 => A(23), ZN => n8);
   U23 : AND2_X1 port map( A1 => A(22), A2 => A(23), ZN => n24);
   U24 : AND2_X2 port map( A1 => n61, A2 => n9, ZN => n56);
   U25 : AND4_X1 port map( A1 => n32, A2 => A(5), A3 => n7, A4 => A(4), ZN => 
                           n9);
   U26 : XNOR2_X1 port map( A => n44, B => n98, ZN => SUM_10_port);
   U27 : AND2_X1 port map( A1 => n8, A2 => n25, ZN => n10);
   U28 : AND2_X1 port map( A1 => n24, A2 => n25, ZN => n11);
   U29 : AND2_X1 port map( A1 => n8, A2 => n25, ZN => n74);
   U30 : AND2_X1 port map( A1 => A(3), A2 => A(7), ZN => n12);
   U31 : CLKBUF_X1 port map( A => n7, Z => n13);
   U32 : AND2_X1 port map( A1 => n84, A2 => n83, ZN => n14);
   U33 : AND2_X1 port map( A1 => n83, A2 => n84, ZN => n34);
   U34 : XOR2_X1 port map( A => A(31), B => n15, Z => SUM_31_port);
   U35 : XOR2_X1 port map( A => n16, B => A(21), Z => SUM_21_port);
   U36 : AND2_X1 port map( A1 => n78, A2 => n22, ZN => n16);
   U37 : CLKBUF_X1 port map( A => n22, Z => n17);
   U38 : AND3_X1 port map( A1 => n34, A2 => n67, A3 => n36, ZN => n48);
   U39 : XNOR2_X1 port map( A => A(23), B => n18, ZN => SUM_23_port);
   U40 : NAND2_X1 port map( A1 => n22, A2 => n31, ZN => n18);
   U41 : AND3_X1 port map( A1 => A(5), A2 => A(6), A3 => A(4), ZN => n19);
   U42 : AND2_X1 port map( A1 => n32, A2 => n19, ZN => n28);
   U43 : CLKBUF_X1 port map( A => A(7), Z => n32);
   U44 : AND2_X1 port map( A1 => A(22), A2 => n20, ZN => n21);
   U45 : INV_X1 port map( A => n76, ZN => n20);
   U46 : NOR2_X1 port map( A1 => n87, A2 => n88, ZN => n23);
   U47 : AND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n25);
   U48 : OR2_X1 port map( A1 => n69, A2 => n70, ZN => n26);
   U49 : NAND4_X1 port map( A1 => A(24), A2 => A(25), A3 => A(26), A4 => A(27),
                           ZN => n27);
   U50 : AND2_X1 port map( A1 => n37, A2 => A(24), ZN => n29);
   U51 : XOR2_X1 port map( A => A(29), B => n30, Z => SUM_29_port);
   U52 : AND2_X1 port map( A1 => n42, A2 => n21, ZN => n31);
   U53 : AND2_X1 port map( A1 => n22, A2 => n75, ZN => n33);
   U54 : AND2_X1 port map( A1 => n56, A2 => n35, ZN => n99);
   U55 : NOR2_X1 port map( A1 => n96, A2 => n97, ZN => n35);
   U56 : AND2_X1 port map( A1 => n74, A2 => n42, ZN => n37);
   U57 : NOR2_X1 port map( A1 => n66, A2 => SUM_2_port, ZN => n38);
   U58 : NOR2_X1 port map( A1 => n66, A2 => SUM_2_port, ZN => n61);
   U59 : AND2_X1 port map( A1 => n37, A2 => n22, ZN => n39);
   U60 : AND2_X1 port map( A1 => A(3), A2 => A(7), ZN => n40);
   U61 : AND4_X2 port map( A1 => A(16), A2 => A(17), A3 => A(18), A4 => A(19), 
                           ZN => n42);
   U62 : NOR2_X1 port map( A1 => n26, A2 => n27, ZN => n67);
   U63 : NAND3_X1 port map( A1 => n40, A2 => A(14), A3 => A(15), ZN => n85);
   U64 : AND2_X1 port map( A1 => n47, A2 => A(18), ZN => n81);
   U65 : XOR2_X1 port map( A => A(19), B => n81, Z => SUM_19_port);
   U66 : XNOR2_X1 port map( A => n41, B => n70, ZN => SUM_28_port);
   U67 : XOR2_X1 port map( A => n43, B => A(11), Z => SUM_11_port);
   U68 : AND2_X1 port map( A1 => A(10), A2 => n99, ZN => n43);
   U69 : NOR2_X1 port map( A1 => n55, A2 => n97, ZN => n44);
   U70 : AND2_X1 port map( A1 => n45, A2 => A(5), ZN => n59);
   U71 : NAND4_X1 port map( A1 => A(16), A2 => A(17), A3 => A(18), A4 => A(19),
                           ZN => n77);
   U72 : AND2_X1 port map( A1 => n61, A2 => n62, ZN => n45);
   U73 : AND2_X1 port map( A1 => n73, A2 => n22, ZN => n46);
   U74 : INV_X1 port map( A => n66, ZN => n65);
   U75 : AND2_X1 port map( A1 => n28, A2 => n38, ZN => n54);
   U76 : INV_X1 port map( A => n64, ZN => n62);
   U77 : INV_X1 port map( A => n96, ZN => n57);
   U78 : NAND2_X1 port map( A1 => A(21), A2 => A(20), ZN => n76);
   U79 : AND2_X1 port map( A1 => n13, A2 => n59, ZN => n50);
   U80 : AND2_X1 port map( A1 => n22, A2 => n29, ZN => n51);
   U81 : INV_X1 port map( A => A(27), ZN => n71);
   U82 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U83 : INV_X1 port map( A => A(14), ZN => n91);
   U84 : XOR2_X1 port map( A => A(22), B => n33, Z => SUM_22_port);
   U85 : XNOR2_X1 port map( A => n52, B => n93, ZN => SUM_12_port);
   U86 : XOR2_X1 port map( A => n55, B => n97, Z => SUM_9_port);
   U87 : XOR2_X1 port map( A => A(13), B => n49, Z => SUM_13_port);
   U88 : XOR2_X1 port map( A => n46, B => A(26), Z => SUM_26_port);
   U89 : XOR2_X1 port map( A => n48, B => A(30), Z => SUM_30_port);
   U90 : XOR2_X1 port map( A => n47, B => A(18), Z => SUM_18_port);
   U91 : XNOR2_X1 port map( A => n53, B => n89, ZN => SUM_15_port);
   U92 : AND2_X1 port map( A1 => A(14), A2 => n90, ZN => n53);
   U93 : XOR2_X1 port map( A => n39, B => A(24), Z => SUM_24_port);
   U94 : XOR2_X1 port map( A => n17, B => A(16), Z => SUM_16_port);
   U95 : XOR2_X1 port map( A => n56, B => n57, Z => SUM_8_port);
   U96 : XNOR2_X1 port map( A => n80, B => A(20), ZN => SUM_20_port);
   U97 : XNOR2_X1 port map( A => n82, B => A(17), ZN => SUM_17_port);
   U98 : INV_X1 port map( A => A(28), ZN => n70);
   U99 : XNOR2_X1 port map( A => n63, B => n45, ZN => SUM_5_port);
   U100 : XNOR2_X1 port map( A => SUM_2_port, B => n65, ZN => SUM_3_port);
   U101 : INV_X1 port map( A => A(29), ZN => n69);
   U102 : INV_X1 port map( A => n32, ZN => n58);
   U103 : NOR2_X1 port map( A1 => n93, A2 => n94, ZN => n92);
   U104 : INV_X1 port map( A => n54, ZN => n95);
   U105 : INV_X1 port map( A => A(4), ZN => n64);
   U106 : NOR2_X1 port map( A1 => n87, A2 => n88, ZN => n83);
   U107 : XNOR2_X1 port map( A => n58, B => n50, ZN => SUM_7_port);
   U108 : NOR2_X1 port map( A1 => n77, A2 => n76, ZN => n75);
   U109 : NOR2_X1 port map( A1 => n79, A2 => n77, ZN => n78);
   U110 : NOR2_X1 port map( A1 => n85, A2 => n86, ZN => n84);
   U111 : NAND4_X1 port map( A1 => A(10), A2 => A(9), A3 => A(8), A4 => A(11), 
                           ZN => n94);
   U112 : INV_X1 port map( A => A(5), ZN => n63);
   U113 : INV_X1 port map( A => A(10), ZN => n98);
   U114 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => n55);
   U115 : INV_X1 port map( A => n13, ZN => n60);
   U116 : XNOR2_X1 port map( A => n60, B => n59, ZN => SUM_6_port);
   U117 : XNOR2_X1 port map( A => n64, B => n38, ZN => SUM_4_port);
   U118 : INV_X1 port map( A => A(8), ZN => n96);
   U119 : NAND2_X1 port map( A1 => n22, A2 => n42, ZN => n80);
   U120 : NAND2_X1 port map( A1 => n22, A2 => A(16), ZN => n82);
   U121 : INV_X1 port map( A => A(9), ZN => n97);
   U122 : XNOR2_X1 port map( A => n72, B => n71, ZN => SUM_27_port);
   U123 : INV_X1 port map( A => A(20), ZN => n79);
   U124 : NAND3_X1 port map( A1 => A(11), A2 => A(13), A3 => A(12), ZN => n86);
   U125 : NAND3_X1 port map( A1 => A(5), A2 => A(2), A3 => A(4), ZN => n88);
   U126 : INV_X1 port map( A => A(15), ZN => n89);
   U127 : XNOR2_X1 port map( A => n91, B => n90, ZN => SUM_14_port);
   U128 : INV_X1 port map( A => A(12), ZN => n93);
   U129 : INV_X1 port map( A => A(3), ZN => n66);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute_DW01_add_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Execute_DW01_add_1;

architecture SYN_rpl of Execute_DW01_add_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_3_port, SUM_4_port, SUM_5_port, SUM_6_port, 
      SUM_7_port, SUM_8_port, SUM_9_port, SUM_10_port, SUM_11_port, SUM_12_port
      , SUM_13_port, SUM_14_port, SUM_15_port, SUM_16_port, SUM_17_port, 
      SUM_18_port, SUM_19_port, SUM_20_port, SUM_21_port, SUM_22_port, 
      SUM_23_port, SUM_24_port, SUM_25_port, SUM_26_port, SUM_27_port, 
      SUM_28_port, SUM_29_port, SUM_30_port, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n54, n55, n56, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, B(1), B(0) );
   
   U1 : XNOR2_X1 port map( A => B(31), B => n57, ZN => SUM_31_port);
   U2 : NAND2_X1 port map( A1 => B(30), A2 => n56, ZN => n57);
   U3 : INV_X1 port map( A => B(2), ZN => SUM_2_port);
   U4 : XOR2_X1 port map( A => B(3), B => B(2), Z => SUM_3_port);
   U5 : XOR2_X1 port map( A => B(4), B => n30, Z => SUM_4_port);
   U6 : XOR2_X1 port map( A => B(5), B => n31, Z => SUM_5_port);
   U7 : XOR2_X1 port map( A => B(6), B => n32, Z => SUM_6_port);
   U8 : XOR2_X1 port map( A => B(7), B => n33, Z => SUM_7_port);
   U9 : XOR2_X1 port map( A => B(8), B => n34, Z => SUM_8_port);
   U10 : XOR2_X1 port map( A => B(9), B => n35, Z => SUM_9_port);
   U11 : XOR2_X1 port map( A => B(10), B => n36, Z => SUM_10_port);
   U12 : XOR2_X1 port map( A => B(11), B => n37, Z => SUM_11_port);
   U13 : XOR2_X1 port map( A => B(12), B => n38, Z => SUM_12_port);
   U14 : XOR2_X1 port map( A => B(13), B => n39, Z => SUM_13_port);
   U15 : XOR2_X1 port map( A => B(14), B => n40, Z => SUM_14_port);
   U16 : XOR2_X1 port map( A => B(15), B => n41, Z => SUM_15_port);
   U17 : XOR2_X1 port map( A => B(16), B => n42, Z => SUM_16_port);
   U18 : XOR2_X1 port map( A => B(17), B => n43, Z => SUM_17_port);
   U19 : XOR2_X1 port map( A => B(18), B => n44, Z => SUM_18_port);
   U20 : XOR2_X1 port map( A => B(19), B => n45, Z => SUM_19_port);
   U21 : XOR2_X1 port map( A => B(20), B => n46, Z => SUM_20_port);
   U22 : XOR2_X1 port map( A => B(21), B => n47, Z => SUM_21_port);
   U23 : XOR2_X1 port map( A => B(22), B => n48, Z => SUM_22_port);
   U24 : XOR2_X1 port map( A => B(23), B => n49, Z => SUM_23_port);
   U25 : XOR2_X1 port map( A => B(24), B => n50, Z => SUM_24_port);
   U26 : XOR2_X1 port map( A => B(25), B => n51, Z => SUM_25_port);
   U27 : XOR2_X1 port map( A => B(26), B => n52, Z => SUM_26_port);
   U28 : XOR2_X1 port map( A => B(27), B => n53, Z => SUM_27_port);
   U29 : XOR2_X1 port map( A => B(28), B => n54, Z => SUM_28_port);
   U30 : XOR2_X1 port map( A => B(29), B => n55, Z => SUM_29_port);
   U31 : XOR2_X1 port map( A => B(30), B => n56, Z => SUM_30_port);
   U32 : AND2_X1 port map( A1 => B(3), A2 => B(2), ZN => n30);
   U33 : AND2_X1 port map( A1 => B(4), A2 => n30, ZN => n31);
   U34 : AND2_X1 port map( A1 => B(5), A2 => n31, ZN => n32);
   U35 : AND2_X1 port map( A1 => B(6), A2 => n32, ZN => n33);
   U36 : AND2_X1 port map( A1 => B(7), A2 => n33, ZN => n34);
   U37 : AND2_X1 port map( A1 => B(8), A2 => n34, ZN => n35);
   U38 : AND2_X1 port map( A1 => B(9), A2 => n35, ZN => n36);
   U39 : AND2_X1 port map( A1 => B(10), A2 => n36, ZN => n37);
   U40 : AND2_X1 port map( A1 => B(11), A2 => n37, ZN => n38);
   U41 : AND2_X1 port map( A1 => B(12), A2 => n38, ZN => n39);
   U42 : AND2_X1 port map( A1 => B(13), A2 => n39, ZN => n40);
   U43 : AND2_X1 port map( A1 => B(14), A2 => n40, ZN => n41);
   U44 : AND2_X1 port map( A1 => B(15), A2 => n41, ZN => n42);
   U45 : AND2_X1 port map( A1 => B(16), A2 => n42, ZN => n43);
   U46 : AND2_X1 port map( A1 => B(17), A2 => n43, ZN => n44);
   U47 : AND2_X1 port map( A1 => B(18), A2 => n44, ZN => n45);
   U48 : AND2_X1 port map( A1 => B(19), A2 => n45, ZN => n46);
   U49 : AND2_X1 port map( A1 => B(20), A2 => n46, ZN => n47);
   U50 : AND2_X1 port map( A1 => B(21), A2 => n47, ZN => n48);
   U51 : AND2_X1 port map( A1 => B(22), A2 => n48, ZN => n49);
   U52 : AND2_X1 port map( A1 => B(23), A2 => n49, ZN => n50);
   U53 : AND2_X1 port map( A1 => B(24), A2 => n50, ZN => n51);
   U54 : AND2_X1 port map( A1 => B(25), A2 => n51, ZN => n52);
   U55 : AND2_X1 port map( A1 => B(26), A2 => n52, ZN => n53);
   U56 : AND2_X1 port map( A1 => B(27), A2 => n53, ZN => n54);
   U57 : AND2_X1 port map( A1 => B(28), A2 => n54, ZN => n55);
   U58 : AND2_X1 port map( A1 => B(29), A2 => n55, ZN => n56);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Execute_DW01_add_0;

architecture SYN_rpl of Execute_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n2, n_1070 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1070, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n2, CO => carry_2_port, S
                           => SUM(1));
   U1 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U2 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n2);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity comparator_NBIT32_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end comparator_NBIT32_DW01_cmp6_0;

architecture SYN_rpl of comparator_NBIT32_DW01_cmp6_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal GT_port, GE_port, NE_port, n3, LE_port, n5, n6, n7, n8, n9, n10, n11,
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55
      , n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, 
      n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84
      , n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, 
      n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202 : std_logic;

begin
   GT <= GT_port;
   LE <= LE_port;
   GE <= GE_port;
   NE <= NE_port;
   
   U1 : INV_X1 port map( A => n142, ZN => n10);
   U2 : INV_X1 port map( A => n130, ZN => n14);
   U3 : INV_X1 port map( A => n118, ZN => n18);
   U4 : INV_X1 port map( A => n106, ZN => n22);
   U5 : INV_X1 port map( A => n94, ZN => n26);
   U6 : INV_X1 port map( A => n82, ZN => n30);
   U7 : INV_X1 port map( A => GE_port, ZN => LT);
   U8 : INV_X1 port map( A => NE_port, ZN => EQ);
   U9 : INV_X1 port map( A => n139, ZN => n12);
   U10 : INV_X1 port map( A => n127, ZN => n16);
   U11 : INV_X1 port map( A => n115, ZN => n20);
   U12 : INV_X1 port map( A => n103, ZN => n24);
   U13 : INV_X1 port map( A => n91, ZN => n28);
   U14 : INV_X1 port map( A => n79, ZN => n32);
   U15 : INV_X1 port map( A => GT_port, ZN => LE_port);
   U16 : INV_X1 port map( A => n144, ZN => n9);
   U17 : INV_X1 port map( A => n132, ZN => n13);
   U18 : INV_X1 port map( A => n120, ZN => n17);
   U19 : INV_X1 port map( A => n108, ZN => n21);
   U20 : INV_X1 port map( A => n96, ZN => n25);
   U21 : INV_X1 port map( A => n84, ZN => n29);
   U22 : INV_X1 port map( A => n154, ZN => n7);
   U23 : INV_X1 port map( A => n141, ZN => n11);
   U24 : INV_X1 port map( A => n129, ZN => n15);
   U25 : INV_X1 port map( A => n117, ZN => n19);
   U26 : INV_X1 port map( A => n105, ZN => n23);
   U27 : INV_X1 port map( A => n93, ZN => n27);
   U28 : INV_X1 port map( A => n81, ZN => n31);
   U29 : INV_X1 port map( A => n68, ZN => n3);
   U30 : INV_X1 port map( A => A(30), ZN => n65);
   U31 : INV_X1 port map( A => n72, ZN => n33);
   U32 : INV_X1 port map( A => n151, ZN => n8);
   U33 : INV_X1 port map( A => n202, ZN => n5);
   U34 : INV_X1 port map( A => B(30), ZN => n34);
   U35 : INV_X1 port map( A => A(0), ZN => n36);
   U36 : INV_X1 port map( A => A(3), ZN => n38);
   U37 : INV_X1 port map( A => A(5), ZN => n40);
   U38 : INV_X1 port map( A => A(7), ZN => n42);
   U39 : INV_X1 port map( A => A(9), ZN => n44);
   U40 : INV_X1 port map( A => A(11), ZN => n46);
   U41 : INV_X1 port map( A => A(13), ZN => n48);
   U42 : INV_X1 port map( A => A(15), ZN => n50);
   U43 : INV_X1 port map( A => A(17), ZN => n52);
   U44 : INV_X1 port map( A => A(19), ZN => n54);
   U45 : INV_X1 port map( A => A(21), ZN => n56);
   U46 : INV_X1 port map( A => A(23), ZN => n58);
   U47 : INV_X1 port map( A => A(25), ZN => n60);
   U48 : INV_X1 port map( A => A(27), ZN => n62);
   U49 : INV_X1 port map( A => A(29), ZN => n64);
   U50 : INV_X1 port map( A => B(31), ZN => n35);
   U51 : INV_X1 port map( A => B(1), ZN => n6);
   U52 : INV_X1 port map( A => A(4), ZN => n39);
   U53 : INV_X1 port map( A => A(8), ZN => n43);
   U54 : INV_X1 port map( A => A(12), ZN => n47);
   U55 : INV_X1 port map( A => A(16), ZN => n51);
   U56 : INV_X1 port map( A => A(20), ZN => n55);
   U57 : INV_X1 port map( A => A(24), ZN => n59);
   U58 : INV_X1 port map( A => A(28), ZN => n63);
   U59 : INV_X1 port map( A => A(2), ZN => n37);
   U60 : INV_X1 port map( A => A(6), ZN => n41);
   U61 : INV_X1 port map( A => A(10), ZN => n45);
   U62 : INV_X1 port map( A => A(14), ZN => n49);
   U63 : INV_X1 port map( A => A(18), ZN => n53);
   U64 : INV_X1 port map( A => A(22), ZN => n57);
   U65 : INV_X1 port map( A => A(26), ZN => n61);
   U66 : NAND2_X1 port map( A1 => LE_port, A2 => GE_port, ZN => NE_port);
   U67 : AOI21_X1 port map( B1 => n66, B2 => n3, A => n67, ZN => GE_port);
   U68 : AOI22_X1 port map( A1 => B(30), A2 => n65, B1 => n69, B2 => n70, ZN =>
                           n68);
   U69 : AOI21_X1 port map( B1 => n71, B2 => n72, A => n73, ZN => n69);
   U70 : AOI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => n71);
   U71 : AOI21_X1 port map( B1 => n77, B2 => n78, A => n79, ZN => n74);
   U72 : AOI21_X1 port map( B1 => n80, B2 => n30, A => n31, ZN => n77);
   U73 : AOI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n80);
   U74 : AOI21_X1 port map( B1 => n86, B2 => n87, A => n88, ZN => n83);
   U75 : AOI21_X1 port map( B1 => n89, B2 => n90, A => n91, ZN => n86);
   U76 : AOI21_X1 port map( B1 => n92, B2 => n26, A => n27, ZN => n89);
   U77 : AOI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n92);
   U78 : AOI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => n95);
   U79 : AOI21_X1 port map( B1 => n101, B2 => n102, A => n103, ZN => n98);
   U80 : AOI21_X1 port map( B1 => n104, B2 => n22, A => n23, ZN => n101);
   U81 : AOI21_X1 port map( B1 => n107, B2 => n108, A => n109, ZN => n104);
   U82 : AOI21_X1 port map( B1 => n110, B2 => n111, A => n112, ZN => n107);
   U83 : AOI21_X1 port map( B1 => n113, B2 => n114, A => n115, ZN => n110);
   U84 : AOI21_X1 port map( B1 => n116, B2 => n18, A => n19, ZN => n113);
   U85 : AOI21_X1 port map( B1 => n119, B2 => n120, A => n121, ZN => n116);
   U86 : AOI21_X1 port map( B1 => n122, B2 => n123, A => n124, ZN => n119);
   U87 : AOI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n122);
   U88 : AOI21_X1 port map( B1 => n128, B2 => n14, A => n15, ZN => n125);
   U89 : AOI21_X1 port map( B1 => n131, B2 => n132, A => n133, ZN => n128);
   U90 : AOI21_X1 port map( B1 => n134, B2 => n135, A => n136, ZN => n131);
   U91 : AOI21_X1 port map( B1 => n137, B2 => n138, A => n139, ZN => n134);
   U92 : AOI21_X1 port map( B1 => n140, B2 => n10, A => n11, ZN => n137);
   U93 : AOI21_X1 port map( B1 => n143, B2 => n144, A => n145, ZN => n140);
   U94 : AOI21_X1 port map( B1 => n146, B2 => n147, A => n148, ZN => n143);
   U95 : AOI21_X1 port map( B1 => n149, B2 => n150, A => n151, ZN => n146);
   U96 : AOI21_X1 port map( B1 => n152, B2 => n153, A => n7, ZN => n149);
   U97 : AOI22_X1 port map( A1 => n155, A2 => n6, B1 => A(1), B2 => n156, ZN =>
                           n152);
   U98 : OR2_X1 port map( A1 => n156, A2 => A(1), ZN => n155);
   U99 : NAND2_X1 port map( A1 => B(0), A2 => n36, ZN => n156);
   U100 : OAI21_X1 port map( B1 => n67, B2 => n157, A => n66, ZN => GT_port);
   U101 : NAND2_X1 port map( A1 => A(31), A2 => n35, ZN => n66);
   U102 : AOI22_X1 port map( A1 => A(30), A2 => n34, B1 => n158, B2 => n70, ZN 
                           => n157);
   U103 : XOR2_X1 port map( A => A(30), B => n34, Z => n70);
   U104 : AOI21_X1 port map( B1 => n159, B2 => n160, A => n33, ZN => n158);
   U105 : NAND2_X1 port map( A1 => B(29), A2 => n64, ZN => n72);
   U106 : OAI211_X1 port map( C1 => n161, C2 => n162, A => n78, B => n75, ZN =>
                           n160);
   U107 : NOR2_X1 port map( A1 => n163, A2 => n76, ZN => n75);
   U108 : AND2_X1 port map( A1 => B(28), A2 => n63, ZN => n76);
   U109 : NAND2_X1 port map( A1 => B(27), A2 => n62, ZN => n78);
   U110 : NAND2_X1 port map( A1 => n32, A2 => n164, ZN => n162);
   U111 : NOR2_X1 port map( A1 => n62, A2 => B(27), ZN => n79);
   U112 : AOI211_X1 port map( C1 => n165, C2 => n166, A => n82, B => n29, ZN =>
                           n161);
   U113 : NAND2_X1 port map( A1 => B(25), A2 => n60, ZN => n84);
   U114 : NAND2_X1 port map( A1 => n164, A2 => n81, ZN => n82);
   U115 : NAND2_X1 port map( A1 => B(26), A2 => n61, ZN => n81);
   U116 : OR2_X1 port map( A1 => n61, A2 => B(26), ZN => n164);
   U117 : OAI211_X1 port map( C1 => n167, C2 => n168, A => n90, B => n87, ZN =>
                           n166);
   U118 : NOR2_X1 port map( A1 => n169, A2 => n88, ZN => n87);
   U119 : AND2_X1 port map( A1 => B(24), A2 => n59, ZN => n88);
   U120 : NAND2_X1 port map( A1 => B(23), A2 => n58, ZN => n90);
   U121 : NAND2_X1 port map( A1 => n28, A2 => n170, ZN => n168);
   U122 : NOR2_X1 port map( A1 => n58, A2 => B(23), ZN => n91);
   U123 : AOI211_X1 port map( C1 => n171, C2 => n172, A => n94, B => n25, ZN =>
                           n167);
   U124 : NAND2_X1 port map( A1 => B(21), A2 => n56, ZN => n96);
   U125 : NAND2_X1 port map( A1 => n170, A2 => n93, ZN => n94);
   U126 : NAND2_X1 port map( A1 => B(22), A2 => n57, ZN => n93);
   U127 : OR2_X1 port map( A1 => n57, A2 => B(22), ZN => n170);
   U128 : OAI211_X1 port map( C1 => n173, C2 => n174, A => n102, B => n99, ZN 
                           => n172);
   U129 : NOR2_X1 port map( A1 => n175, A2 => n100, ZN => n99);
   U130 : AND2_X1 port map( A1 => B(20), A2 => n55, ZN => n100);
   U131 : NAND2_X1 port map( A1 => B(19), A2 => n54, ZN => n102);
   U132 : NAND2_X1 port map( A1 => n24, A2 => n176, ZN => n174);
   U133 : NOR2_X1 port map( A1 => n54, A2 => B(19), ZN => n103);
   U134 : AOI211_X1 port map( C1 => n177, C2 => n178, A => n106, B => n21, ZN 
                           => n173);
   U135 : NAND2_X1 port map( A1 => B(17), A2 => n52, ZN => n108);
   U136 : NAND2_X1 port map( A1 => n176, A2 => n105, ZN => n106);
   U137 : NAND2_X1 port map( A1 => B(18), A2 => n53, ZN => n105);
   U138 : OR2_X1 port map( A1 => n53, A2 => B(18), ZN => n176);
   U139 : OAI211_X1 port map( C1 => n179, C2 => n180, A => n114, B => n111, ZN 
                           => n178);
   U140 : NOR2_X1 port map( A1 => n181, A2 => n112, ZN => n111);
   U141 : AND2_X1 port map( A1 => B(16), A2 => n51, ZN => n112);
   U142 : NAND2_X1 port map( A1 => B(15), A2 => n50, ZN => n114);
   U143 : NAND2_X1 port map( A1 => n20, A2 => n182, ZN => n180);
   U144 : NOR2_X1 port map( A1 => n50, A2 => B(15), ZN => n115);
   U145 : AOI211_X1 port map( C1 => n183, C2 => n184, A => n118, B => n17, ZN 
                           => n179);
   U146 : NAND2_X1 port map( A1 => B(13), A2 => n48, ZN => n120);
   U147 : NAND2_X1 port map( A1 => n182, A2 => n117, ZN => n118);
   U148 : NAND2_X1 port map( A1 => B(14), A2 => n49, ZN => n117);
   U149 : OR2_X1 port map( A1 => n49, A2 => B(14), ZN => n182);
   U150 : OAI211_X1 port map( C1 => n185, C2 => n186, A => n126, B => n123, ZN 
                           => n184);
   U151 : NOR2_X1 port map( A1 => n187, A2 => n124, ZN => n123);
   U152 : AND2_X1 port map( A1 => B(12), A2 => n47, ZN => n124);
   U153 : NAND2_X1 port map( A1 => B(11), A2 => n46, ZN => n126);
   U154 : NAND2_X1 port map( A1 => n16, A2 => n188, ZN => n186);
   U155 : NOR2_X1 port map( A1 => n46, A2 => B(11), ZN => n127);
   U156 : AOI211_X1 port map( C1 => n189, C2 => n190, A => n130, B => n13, ZN 
                           => n185);
   U157 : NAND2_X1 port map( A1 => B(9), A2 => n44, ZN => n132);
   U158 : NAND2_X1 port map( A1 => n188, A2 => n129, ZN => n130);
   U159 : NAND2_X1 port map( A1 => B(10), A2 => n45, ZN => n129);
   U160 : OR2_X1 port map( A1 => n45, A2 => B(10), ZN => n188);
   U161 : OAI211_X1 port map( C1 => n191, C2 => n192, A => n138, B => n135, ZN 
                           => n190);
   U162 : NOR2_X1 port map( A1 => n193, A2 => n136, ZN => n135);
   U163 : AND2_X1 port map( A1 => B(8), A2 => n43, ZN => n136);
   U164 : NAND2_X1 port map( A1 => B(7), A2 => n42, ZN => n138);
   U165 : NAND2_X1 port map( A1 => n12, A2 => n194, ZN => n192);
   U166 : NOR2_X1 port map( A1 => n42, A2 => B(7), ZN => n139);
   U167 : AOI211_X1 port map( C1 => n195, C2 => n196, A => n142, B => n9, ZN =>
                           n191);
   U168 : NAND2_X1 port map( A1 => B(5), A2 => n40, ZN => n144);
   U169 : NAND2_X1 port map( A1 => n194, A2 => n141, ZN => n142);
   U170 : NAND2_X1 port map( A1 => B(6), A2 => n41, ZN => n141);
   U171 : OR2_X1 port map( A1 => n41, A2 => B(6), ZN => n194);
   U172 : NAND3_X1 port map( A1 => n197, A2 => n150, A3 => n147, ZN => n196);
   U173 : NOR2_X1 port map( A1 => n198, A2 => n148, ZN => n147);
   U174 : AND2_X1 port map( A1 => B(4), A2 => n39, ZN => n148);
   U175 : NAND2_X1 port map( A1 => B(3), A2 => n38, ZN => n150);
   U176 : NAND3_X1 port map( A1 => n8, A2 => n199, A3 => n200, ZN => n197);
   U177 : OAI211_X1 port map( C1 => A(1), C2 => n201, A => n5, B => n153, ZN =>
                           n200);
   U178 : AND2_X1 port map( A1 => n199, A2 => n154, ZN => n153);
   U179 : NAND2_X1 port map( A1 => B(2), A2 => n37, ZN => n154);
   U180 : AOI21_X1 port map( B1 => A(1), B2 => n201, A => n6, ZN => n202);
   U181 : NOR2_X1 port map( A1 => n36, A2 => B(0), ZN => n201);
   U182 : OR2_X1 port map( A1 => n37, A2 => B(2), ZN => n199);
   U183 : NOR2_X1 port map( A1 => n38, A2 => B(3), ZN => n151);
   U184 : NOR2_X1 port map( A1 => n198, A2 => n145, ZN => n195);
   U185 : NOR2_X1 port map( A1 => n40, A2 => B(5), ZN => n145);
   U186 : NOR2_X1 port map( A1 => n39, A2 => B(4), ZN => n198);
   U187 : NOR2_X1 port map( A1 => n193, A2 => n133, ZN => n189);
   U188 : NOR2_X1 port map( A1 => n44, A2 => B(9), ZN => n133);
   U189 : NOR2_X1 port map( A1 => n43, A2 => B(8), ZN => n193);
   U190 : NOR2_X1 port map( A1 => n187, A2 => n121, ZN => n183);
   U191 : NOR2_X1 port map( A1 => n48, A2 => B(13), ZN => n121);
   U192 : NOR2_X1 port map( A1 => n47, A2 => B(12), ZN => n187);
   U193 : NOR2_X1 port map( A1 => n181, A2 => n109, ZN => n177);
   U194 : NOR2_X1 port map( A1 => n52, A2 => B(17), ZN => n109);
   U195 : NOR2_X1 port map( A1 => n51, A2 => B(16), ZN => n181);
   U196 : NOR2_X1 port map( A1 => n175, A2 => n97, ZN => n171);
   U197 : NOR2_X1 port map( A1 => n56, A2 => B(21), ZN => n97);
   U198 : NOR2_X1 port map( A1 => n55, A2 => B(20), ZN => n175);
   U199 : NOR2_X1 port map( A1 => n169, A2 => n85, ZN => n165);
   U200 : NOR2_X1 port map( A1 => n60, A2 => B(25), ZN => n85);
   U201 : NOR2_X1 port map( A1 => n59, A2 => B(24), ZN => n169);
   U202 : NOR2_X1 port map( A1 => n163, A2 => n73, ZN => n159);
   U203 : NOR2_X1 port map( A1 => n64, A2 => B(29), ZN => n73);
   U204 : NOR2_X1 port map( A1 => n63, A2 => B(28), ZN => n163);
   U205 : NOR2_X1 port map( A1 => n35, A2 => A(31), ZN => n67);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HazardDetection_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end HazardDetection_DW01_sub_0;

architecture SYN_rpl of HazardDetection_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port,
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, carry_31_port, 
      carry_30_port, carry_29_port, carry_28_port, carry_27_port, carry_26_port
      , carry_25_port, carry_24_port, carry_23_port, carry_22_port, 
      carry_21_port, carry_20_port, carry_19_port, carry_18_port, carry_17_port
      , carry_16_port, carry_15_port, carry_14_port, carry_13_port, 
      carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, n1, n2, 
      DIFF_2_port : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, A(1), A(0) );
   
   U1 : XNOR2_X1 port map( A => A(4), B => carry_4_port, ZN => DIFF_4_port);
   U2 : XNOR2_X1 port map( A => A(21), B => carry_21_port, ZN => DIFF_21_port);
   U3 : XNOR2_X1 port map( A => A(22), B => carry_22_port, ZN => DIFF_22_port);
   U4 : XNOR2_X1 port map( A => A(23), B => carry_23_port, ZN => DIFF_23_port);
   U5 : XNOR2_X1 port map( A => A(28), B => carry_28_port, ZN => DIFF_28_port);
   U6 : XNOR2_X1 port map( A => A(29), B => carry_29_port, ZN => DIFF_29_port);
   U7 : XNOR2_X1 port map( A => A(30), B => carry_30_port, ZN => DIFF_30_port);
   U8 : XNOR2_X1 port map( A => A(31), B => carry_31_port, ZN => DIFF_31_port);
   U9 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => carry_31_port);
   U10 : INV_X1 port map( A => carry_30_port, ZN => n2);
   U11 : INV_X1 port map( A => A(30), ZN => n1);
   U12 : XNOR2_X1 port map( A => A(3), B => A(2), ZN => DIFF_3_port);
   U13 : XNOR2_X1 port map( A => A(5), B => carry_5_port, ZN => DIFF_5_port);
   U14 : XNOR2_X1 port map( A => A(6), B => carry_6_port, ZN => DIFF_6_port);
   U15 : XNOR2_X1 port map( A => A(7), B => carry_7_port, ZN => DIFF_7_port);
   U16 : OR2_X1 port map( A1 => A(3), A2 => A(2), ZN => carry_4_port);
   U17 : XNOR2_X1 port map( A => A(25), B => carry_25_port, ZN => DIFF_25_port)
                           ;
   U18 : XNOR2_X1 port map( A => A(9), B => carry_9_port, ZN => DIFF_9_port);
   U19 : OR2_X1 port map( A1 => A(4), A2 => carry_4_port, ZN => carry_5_port);
   U20 : OR2_X1 port map( A1 => A(5), A2 => carry_5_port, ZN => carry_6_port);
   U21 : OR2_X1 port map( A1 => A(6), A2 => carry_6_port, ZN => carry_7_port);
   U22 : OR2_X1 port map( A1 => A(7), A2 => carry_7_port, ZN => carry_8_port);
   U23 : OR2_X1 port map( A1 => A(8), A2 => carry_8_port, ZN => carry_9_port);
   U24 : OR2_X1 port map( A1 => A(9), A2 => carry_9_port, ZN => carry_10_port);
   U25 : OR2_X1 port map( A1 => A(10), A2 => carry_10_port, ZN => carry_11_port
                           );
   U26 : OR2_X1 port map( A1 => A(11), A2 => carry_11_port, ZN => carry_12_port
                           );
   U27 : OR2_X1 port map( A1 => A(12), A2 => carry_12_port, ZN => carry_13_port
                           );
   U28 : OR2_X1 port map( A1 => A(13), A2 => carry_13_port, ZN => carry_14_port
                           );
   U29 : OR2_X1 port map( A1 => A(14), A2 => carry_14_port, ZN => carry_15_port
                           );
   U30 : OR2_X1 port map( A1 => A(15), A2 => carry_15_port, ZN => carry_16_port
                           );
   U31 : OR2_X1 port map( A1 => A(16), A2 => carry_16_port, ZN => carry_17_port
                           );
   U32 : OR2_X1 port map( A1 => A(17), A2 => carry_17_port, ZN => carry_18_port
                           );
   U33 : OR2_X1 port map( A1 => A(18), A2 => carry_18_port, ZN => carry_19_port
                           );
   U34 : OR2_X1 port map( A1 => A(19), A2 => carry_19_port, ZN => carry_20_port
                           );
   U35 : OR2_X1 port map( A1 => A(20), A2 => carry_20_port, ZN => carry_21_port
                           );
   U36 : OR2_X1 port map( A1 => A(21), A2 => carry_21_port, ZN => carry_22_port
                           );
   U37 : OR2_X1 port map( A1 => A(22), A2 => carry_22_port, ZN => carry_23_port
                           );
   U38 : OR2_X1 port map( A1 => A(23), A2 => carry_23_port, ZN => carry_24_port
                           );
   U39 : OR2_X1 port map( A1 => A(24), A2 => carry_24_port, ZN => carry_25_port
                           );
   U40 : OR2_X1 port map( A1 => A(25), A2 => carry_25_port, ZN => carry_26_port
                           );
   U41 : OR2_X1 port map( A1 => A(26), A2 => carry_26_port, ZN => carry_27_port
                           );
   U42 : OR2_X1 port map( A1 => A(27), A2 => carry_27_port, ZN => carry_28_port
                           );
   U43 : OR2_X1 port map( A1 => A(28), A2 => carry_28_port, ZN => carry_29_port
                           );
   U44 : OR2_X1 port map( A1 => A(29), A2 => carry_29_port, ZN => carry_30_port
                           );
   U45 : XNOR2_X1 port map( A => A(8), B => carry_8_port, ZN => DIFF_8_port);
   U46 : XNOR2_X1 port map( A => A(10), B => carry_10_port, ZN => DIFF_10_port)
                           ;
   U47 : XNOR2_X1 port map( A => A(11), B => carry_11_port, ZN => DIFF_11_port)
                           ;
   U48 : XNOR2_X1 port map( A => A(12), B => carry_12_port, ZN => DIFF_12_port)
                           ;
   U49 : XNOR2_X1 port map( A => A(13), B => carry_13_port, ZN => DIFF_13_port)
                           ;
   U50 : XNOR2_X1 port map( A => A(14), B => carry_14_port, ZN => DIFF_14_port)
                           ;
   U51 : XNOR2_X1 port map( A => A(15), B => carry_15_port, ZN => DIFF_15_port)
                           ;
   U52 : XNOR2_X1 port map( A => A(16), B => carry_16_port, ZN => DIFF_16_port)
                           ;
   U53 : XNOR2_X1 port map( A => A(17), B => carry_17_port, ZN => DIFF_17_port)
                           ;
   U54 : XNOR2_X1 port map( A => A(18), B => carry_18_port, ZN => DIFF_18_port)
                           ;
   U55 : XNOR2_X1 port map( A => A(19), B => carry_19_port, ZN => DIFF_19_port)
                           ;
   U56 : XNOR2_X1 port map( A => A(20), B => carry_20_port, ZN => DIFF_20_port)
                           ;
   U57 : XNOR2_X1 port map( A => A(24), B => carry_24_port, ZN => DIFF_24_port)
                           ;
   U58 : XNOR2_X1 port map( A => A(26), B => carry_26_port, ZN => DIFF_26_port)
                           ;
   U59 : XNOR2_X1 port map( A => A(27), B => carry_27_port, ZN => DIFF_27_port)
                           ;
   U60 : INV_X1 port map( A => A(2), ZN => DIFF_2_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_15;

architecture SYN_STRUCTURAL of RCA_N4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_14;

architecture SYN_STRUCTURAL of RCA_N4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_13;

architecture SYN_STRUCTURAL of RCA_N4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_12;

architecture SYN_STRUCTURAL of RCA_N4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_11;

architecture SYN_STRUCTURAL of RCA_N4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_10;

architecture SYN_STRUCTURAL of RCA_N4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_9;

architecture SYN_STRUCTURAL of RCA_N4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_8;

architecture SYN_STRUCTURAL of RCA_N4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_7;

architecture SYN_STRUCTURAL of RCA_N4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_6;

architecture SYN_STRUCTURAL of RCA_N4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_5;

architecture SYN_STRUCTURAL of RCA_N4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_4;

architecture SYN_STRUCTURAL of RCA_N4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_3;

architecture SYN_STRUCTURAL of RCA_N4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_2;

architecture SYN_STRUCTURAL of RCA_N4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_1;

architecture SYN_STRUCTURAL of RCA_N4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_7;

architecture SYN_struct of carry_select_basic_N4_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1106, n_1107 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1106);
   RCA1 : RCA_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1107);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n11, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_6;

architecture SYN_struct of carry_select_basic_N4_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1108, n_1109 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1108);
   RCA1 : RCA_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1109);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n11, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_5;

architecture SYN_struct of carry_select_basic_N4_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1110, n_1111 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1110);
   RCA1 : RCA_N4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1111);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n11, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_4;

architecture SYN_struct of carry_select_basic_N4_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1112, n_1113 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1112);
   RCA1 : RCA_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1113);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n11, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_3;

architecture SYN_struct of carry_select_basic_N4_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1114, n_1115 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1114);
   RCA1 : RCA_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1115);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n11, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_2;

architecture SYN_struct of carry_select_basic_N4_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1116, n_1117 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1116);
   RCA1 : RCA_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1117);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n11, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_1;

architecture SYN_struct of carry_select_basic_N4_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1118, n_1119 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1118);
   RCA1 : RCA_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1119);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n11, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_26 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_26;

architecture SYN_bhv of PGblock_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_25 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_25;

architecture SYN_bhv of PGblock_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_24 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_24;

architecture SYN_bhv of PGblock_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_23 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_23;

architecture SYN_bhv of PGblock_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_22 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_22;

architecture SYN_bhv of PGblock_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_21 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_21;

architecture SYN_bhv of PGblock_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_20 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_20;

architecture SYN_bhv of PGblock_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_19 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_19;

architecture SYN_bhv of PGblock_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_18 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_18;

architecture SYN_bhv of PGblock_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_17 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_17;

architecture SYN_bhv of PGblock_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_16 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_16;

architecture SYN_bhv of PGblock_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_15 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_15;

architecture SYN_bhv of PGblock_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_14 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_14;

architecture SYN_bhv of PGblock_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_13 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_13;

architecture SYN_bhv of PGblock_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_12 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_12;

architecture SYN_bhv of PGblock_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_11 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_11;

architecture SYN_bhv of PGblock_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_10 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_10;

architecture SYN_bhv of PGblock_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_9 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_9;

architecture SYN_bhv of PGblock_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_8 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_8;

architecture SYN_bhv of PGblock_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_7 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_7;

architecture SYN_bhv of PGblock_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_6 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_6;

architecture SYN_bhv of PGblock_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_5 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_5;

architecture SYN_bhv of PGblock_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_4 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_4;

architecture SYN_bhv of PGblock_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_3 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_3;

architecture SYN_bhv of PGblock_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_2 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_2;

architecture SYN_bhv of PGblock_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_1 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_1;

architecture SYN_bhv of PGblock_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_8 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_8;

architecture SYN_bhv of Gblock_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_7 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_7;

architecture SYN_bhv of Gblock_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_6 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_6;

architecture SYN_bhv of Gblock_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_5 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_5;

architecture SYN_bhv of Gblock_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_4 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_4;

architecture SYN_bhv of Gblock_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_3 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_3;

architecture SYN_bhv of Gblock_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_2 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_2;

architecture SYN_bhv of Gblock_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_1 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_1;

architecture SYN_bhv of Gblock_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_30 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_30;

architecture SYN_bhv of PG_net_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_29 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_29;

architecture SYN_bhv of PG_net_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_28 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_28;

architecture SYN_bhv of PG_net_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_27 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_27;

architecture SYN_bhv of PG_net_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_26 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_26;

architecture SYN_bhv of PG_net_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_25 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_25;

architecture SYN_bhv of PG_net_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_24 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_24;

architecture SYN_bhv of PG_net_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_23 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_23;

architecture SYN_bhv of PG_net_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_22 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_22;

architecture SYN_bhv of PG_net_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_21 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_21;

architecture SYN_bhv of PG_net_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_20 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_20;

architecture SYN_bhv of PG_net_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_19 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_19;

architecture SYN_bhv of PG_net_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_18 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_18;

architecture SYN_bhv of PG_net_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_17 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_17;

architecture SYN_bhv of PG_net_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_16 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_16;

architecture SYN_bhv of PG_net_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_15 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_15;

architecture SYN_bhv of PG_net_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_14 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_14;

architecture SYN_bhv of PG_net_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_13 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_13;

architecture SYN_bhv of PG_net_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_12 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_12;

architecture SYN_bhv of PG_net_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_11 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_11;

architecture SYN_bhv of PG_net_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_10 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_10;

architecture SYN_bhv of PG_net_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_9 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_9;

architecture SYN_bhv of PG_net_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_8 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_8;

architecture SYN_bhv of PG_net_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_7 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_7;

architecture SYN_bhv of PG_net_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_6 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_6;

architecture SYN_bhv of PG_net_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_5 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_5;

architecture SYN_bhv of PG_net_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_4 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_4;

architecture SYN_bhv of PG_net_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_3 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_3;

architecture SYN_bhv of PG_net_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_2 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_2;

architecture SYN_bhv of PG_net_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_1 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_1;

architecture SYN_bhv of PG_net_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_4 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_4;

architecture SYN_bhv of mux41_NBIT32_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n145, Z => n72);
   U2 : BUF_X1 port map( A => n145, Z => n73);
   U3 : BUF_X1 port map( A => n147, Z => n78);
   U4 : BUF_X1 port map( A => n147, Z => n79);
   U5 : BUF_X1 port map( A => n144, Z => n1);
   U6 : BUF_X1 port map( A => n144, Z => n70);
   U7 : BUF_X1 port map( A => n146, Z => n75);
   U8 : BUF_X1 port map( A => n146, Z => n76);
   U9 : BUF_X1 port map( A => n145, Z => n74);
   U10 : BUF_X1 port map( A => n147, Z => n80);
   U11 : BUF_X1 port map( A => n144, Z => n71);
   U12 : BUF_X1 port map( A => n146, Z => n77);
   U13 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n145);
   U14 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n144);
   U15 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n147);
   U16 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n146);
   U17 : INV_X1 port map( A => S(0), ZN => n81);
   U18 : NAND2_X1 port map( A1 => n83, A2 => n82, ZN => Z(0));
   U19 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n82);
   U20 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n83);
   U21 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(1));
   U22 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN =>
                           n104);
   U23 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN => 
                           n105);
   U24 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(2));
   U25 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN =>
                           n126);
   U26 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN =>
                           n127);
   U27 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(6));
   U28 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n138);
   U29 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n139);
   U30 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(5));
   U31 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN =>
                           n136);
   U32 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN =>
                           n137);
   U33 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(4));
   U34 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN =>
                           n134);
   U35 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN =>
                           n135);
   U36 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => Z(13));
   U37 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN 
                           => n90);
   U38 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n91);
   U39 : NAND2_X1 port map( A1 => n93, A2 => n92, ZN => Z(14));
   U40 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN 
                           => n92);
   U41 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n93);
   U42 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => Z(12));
   U43 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN 
                           => n88);
   U44 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n89);
   U45 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(16));
   U46 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n96);
   U47 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n97);
   U48 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(17));
   U49 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n98);
   U50 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n99);
   U51 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(8));
   U52 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n142);
   U53 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n143);
   U54 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(9));
   U55 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN =>
                           n148);
   U56 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN =>
                           n149);
   U57 : NAND2_X1 port map( A1 => n85, A2 => n84, ZN => Z(10));
   U58 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN 
                           => n84);
   U59 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n85);
   U60 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(18));
   U61 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n100);
   U62 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n101);
   U63 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(21));
   U64 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n108);
   U65 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n109);
   U66 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(20));
   U67 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN 
                           => n106);
   U68 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN 
                           => n107);
   U69 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(30));
   U70 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN 
                           => n128);
   U71 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN 
                           => n129);
   U72 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(29));
   U73 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n124);
   U74 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n125);
   U75 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(24));
   U76 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN 
                           => n114);
   U77 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN 
                           => n115);
   U78 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(22));
   U79 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n110);
   U80 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n111);
   U81 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(25));
   U82 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n116);
   U83 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n117);
   U84 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(26));
   U85 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n118);
   U86 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n119);
   U87 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(28));
   U88 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n122);
   U89 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n123);
   U90 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(3));
   U91 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN =>
                           n132);
   U92 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN =>
                           n133);
   U93 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(7));
   U94 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n140);
   U95 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n141);
   U96 : NAND2_X1 port map( A1 => n87, A2 => n86, ZN => Z(11));
   U97 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN 
                           => n86);
   U98 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n87);
   U99 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => Z(15));
   U100 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN
                           => n94);
   U101 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n95);
   U102 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(19));
   U103 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN
                           => n102);
   U104 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n103);
   U105 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(23));
   U106 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN
                           => n112);
   U107 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN
                           => n113);
   U108 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(27));
   U109 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN
                           => n120);
   U110 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN
                           => n121);
   U111 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(31));
   U112 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN
                           => n130);
   U113 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN
                           => n131);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_3 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_3;

architecture SYN_bhv of mux41_NBIT32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n145, Z => n72);
   U2 : BUF_X1 port map( A => n147, Z => n78);
   U3 : BUF_X1 port map( A => n145, Z => n73);
   U4 : BUF_X1 port map( A => n147, Z => n79);
   U5 : BUF_X1 port map( A => n144, Z => n1);
   U6 : BUF_X1 port map( A => n146, Z => n75);
   U7 : BUF_X1 port map( A => n144, Z => n70);
   U8 : BUF_X1 port map( A => n146, Z => n76);
   U9 : BUF_X1 port map( A => n145, Z => n74);
   U10 : BUF_X1 port map( A => n147, Z => n80);
   U11 : BUF_X1 port map( A => n144, Z => n71);
   U12 : BUF_X1 port map( A => n146, Z => n77);
   U13 : NAND2_X1 port map( A1 => n83, A2 => n82, ZN => Z(0));
   U14 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n82);
   U15 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n83);
   U16 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(1));
   U17 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN =>
                           n104);
   U18 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN => 
                           n105);
   U19 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(2));
   U20 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN =>
                           n126);
   U21 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN =>
                           n127);
   U22 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(6));
   U23 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n138);
   U24 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n139);
   U25 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(5));
   U26 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN =>
                           n136);
   U27 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN =>
                           n137);
   U28 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(4));
   U29 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN =>
                           n134);
   U30 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN =>
                           n135);
   U31 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => Z(13));
   U32 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN 
                           => n90);
   U33 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n91);
   U34 : NAND2_X1 port map( A1 => n93, A2 => n92, ZN => Z(14));
   U35 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN 
                           => n92);
   U36 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n93);
   U37 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => Z(12));
   U38 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN 
                           => n88);
   U39 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n89);
   U40 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(16));
   U41 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n96);
   U42 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n97);
   U43 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(17));
   U44 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n98);
   U45 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n99);
   U46 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(8));
   U47 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n142);
   U48 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n143);
   U49 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(9));
   U50 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN =>
                           n148);
   U51 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN =>
                           n149);
   U52 : NAND2_X1 port map( A1 => n85, A2 => n84, ZN => Z(10));
   U53 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN 
                           => n84);
   U54 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n85);
   U55 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(18));
   U56 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n100);
   U57 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n101);
   U58 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(21));
   U59 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n108);
   U60 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n109);
   U61 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(20));
   U62 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN 
                           => n106);
   U63 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN 
                           => n107);
   U64 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(30));
   U65 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN 
                           => n128);
   U66 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN 
                           => n129);
   U67 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(29));
   U68 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n124);
   U69 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n125);
   U70 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(24));
   U71 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN 
                           => n114);
   U72 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN 
                           => n115);
   U73 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(22));
   U74 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n110);
   U75 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n111);
   U76 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(25));
   U77 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n116);
   U78 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n117);
   U79 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(26));
   U80 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n118);
   U81 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n119);
   U82 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(28));
   U83 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n122);
   U84 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n123);
   U85 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(3));
   U86 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN =>
                           n132);
   U87 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN =>
                           n133);
   U88 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(7));
   U89 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n140);
   U90 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n141);
   U91 : NAND2_X1 port map( A1 => n87, A2 => n86, ZN => Z(11));
   U92 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN 
                           => n86);
   U93 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n87);
   U94 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => Z(15));
   U95 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN 
                           => n94);
   U96 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n95);
   U97 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(19));
   U98 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN 
                           => n102);
   U99 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n103);
   U100 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(23));
   U101 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN
                           => n112);
   U102 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN
                           => n113);
   U103 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(27));
   U104 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN
                           => n120);
   U105 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN
                           => n121);
   U106 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(31));
   U107 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN
                           => n130);
   U108 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN
                           => n131);
   U109 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n145);
   U110 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n144);
   U111 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n147);
   U112 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n146);
   U113 : INV_X1 port map( A => S(0), ZN => n81);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_2 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_2;

architecture SYN_bhv of mux41_NBIT32_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n20, n21, n22, n23, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n71, n72, n73, n74, 
      n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105 : std_logic;

begin
   
   U1 : OAI221_X1 port map( B1 => n1, B2 => n9, C1 => n2, C2 => n3, A => n105, 
                           ZN => Z(7));
   U2 : INV_X1 port map( A => B(7), ZN => n1);
   U3 : INV_X1 port map( A => A(7), ZN => n2);
   U4 : INV_X1 port map( A => n32, ZN => n3);
   U5 : OAI221_X1 port map( B1 => n4, B2 => n5, C1 => n6, C2 => n7, A => n50, 
                           ZN => Z(9));
   U6 : INV_X1 port map( A => B(9), ZN => n4);
   U7 : INV_X1 port map( A => n34, ZN => n5);
   U8 : INV_X1 port map( A => A(9), ZN => n6);
   U9 : INV_X1 port map( A => n32, ZN => n7);
   U10 : AOI22_X1 port map( A1 => B(27), A2 => n34, B1 => A(27), B2 => n32, ZN 
                           => n82);
   U11 : OAI221_X1 port map( B1 => n8, B2 => n9, C1 => n10, C2 => n7, A => n78,
                           ZN => Z(25));
   U12 : INV_X1 port map( A => B(25), ZN => n8);
   U13 : INV_X1 port map( A => n34, ZN => n9);
   U14 : INV_X1 port map( A => A(25), ZN => n10);
   U15 : OAI221_X1 port map( B1 => n20, B2 => n5, C1 => n21, C2 => n3, A => n63
                           , ZN => Z(17));
   U16 : INV_X1 port map( A => B(17), ZN => n20);
   U17 : INV_X1 port map( A => A(17), ZN => n21);
   U18 : OAI221_X1 port map( B1 => n22, B2 => n5, C1 => n23, C2 => n7, A => n51
                           , ZN => Z(10));
   U19 : INV_X1 port map( A => B(10), ZN => n22);
   U20 : INV_X1 port map( A => A(10), ZN => n23);
   U21 : OAI221_X1 port map( B1 => n26, B2 => n9, C1 => n27, C2 => n7, A => n52
                           , ZN => Z(11));
   U22 : INV_X1 port map( A => B(11), ZN => n26);
   U23 : INV_X1 port map( A => A(11), ZN => n27);
   U24 : AOI221_X1 port map( B1 => B(19), B2 => n34, C1 => A(19), C2 => n32, A 
                           => n28, ZN => n29);
   U25 : INV_X1 port map( A => n66, ZN => n28);
   U26 : INV_X1 port map( A => n29, ZN => Z(19));
   U27 : OAI221_X1 port map( B1 => n30, B2 => n5, C1 => n31, C2 => n3, A => n67
                           , ZN => Z(20));
   U28 : INV_X1 port map( A => B(20), ZN => n30);
   U29 : INV_X1 port map( A => A(20), ZN => n31);
   U30 : AOI22_X1 port map( A1 => B(28), A2 => n34, B1 => A(28), B2 => n32, ZN 
                           => n84);
   U31 : AOI22_X1 port map( A1 => B(31), A2 => n34, B1 => A(31), B2 => n32, ZN 
                           => n90);
   U32 : AOI22_X1 port map( A1 => B(15), A2 => n34, B1 => A(15), B2 => n32, ZN 
                           => n60);
   U33 : BUF_X1 port map( A => n32, Z => n41);
   U34 : BUF_X1 port map( A => n32, Z => n40);
   U35 : BUF_X1 port map( A => n34, Z => n43);
   U36 : BUF_X1 port map( A => n33, Z => n37);
   U37 : BUF_X1 port map( A => n33, Z => n36);
   U38 : BUF_X1 port map( A => n34, Z => n42);
   U39 : AND2_X1 port map( A1 => n44, A2 => n45, ZN => n32);
   U40 : BUF_X1 port map( A => n35, Z => n39);
   U41 : BUF_X1 port map( A => n35, Z => n38);
   U42 : NAND2_X1 port map( A1 => n92, A2 => n91, ZN => Z(0));
   U43 : AOI22_X1 port map( A1 => D(0), A2 => n38, B1 => C(0), B2 => n36, ZN =>
                           n91);
   U44 : AOI22_X1 port map( A1 => B(0), A2 => n42, B1 => A(0), B2 => n40, ZN =>
                           n92);
   U45 : AND2_X1 port map( A1 => S(1), A2 => n45, ZN => n33);
   U46 : AND2_X1 port map( A1 => S(0), A2 => n44, ZN => n34);
   U47 : AOI22_X1 port map( A1 => D(7), A2 => n38, B1 => C(7), B2 => n36, ZN =>
                           n105);
   U48 : NAND2_X1 port map( A1 => n96, A2 => n95, ZN => Z(2));
   U49 : AOI22_X1 port map( A1 => D(2), A2 => n38, B1 => C(2), B2 => n36, ZN =>
                           n95);
   U50 : AOI22_X1 port map( A1 => B(2), A2 => n42, B1 => A(2), B2 => n40, ZN =>
                           n96);
   U51 : NAND2_X1 port map( A1 => n104, A2 => n103, ZN => Z(6));
   U52 : AOI22_X1 port map( A1 => D(6), A2 => n38, B1 => C(6), B2 => n36, ZN =>
                           n103);
   U53 : AOI22_X1 port map( A1 => B(6), A2 => n42, B1 => A(6), B2 => n40, ZN =>
                           n104);
   U54 : NAND2_X1 port map( A1 => n102, A2 => n101, ZN => Z(5));
   U55 : AOI22_X1 port map( A1 => D(5), A2 => n38, B1 => C(5), B2 => n36, ZN =>
                           n101);
   U56 : AOI22_X1 port map( A1 => B(5), A2 => n42, B1 => A(5), B2 => n40, ZN =>
                           n102);
   U57 : NAND2_X1 port map( A1 => n94, A2 => n93, ZN => Z(1));
   U58 : AOI22_X1 port map( A1 => D(1), A2 => n38, B1 => C(1), B2 => n36, ZN =>
                           n93);
   U59 : AOI22_X1 port map( A1 => B(1), A2 => n42, B1 => A(1), B2 => n40, ZN =>
                           n94);
   U60 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => Z(3));
   U61 : AOI22_X1 port map( A1 => D(3), A2 => n38, B1 => C(3), B2 => n36, ZN =>
                           n97);
   U62 : AOI22_X1 port map( A1 => B(3), A2 => n42, B1 => A(3), B2 => n40, ZN =>
                           n98);
   U63 : NAND2_X1 port map( A1 => n100, A2 => n99, ZN => Z(4));
   U64 : AOI22_X1 port map( A1 => D(4), A2 => n38, B1 => C(4), B2 => n36, ZN =>
                           n99);
   U65 : AOI22_X1 port map( A1 => B(4), A2 => n42, B1 => A(4), B2 => n40, ZN =>
                           n100);
   U66 : AND2_X1 port map( A1 => S(0), A2 => S(1), ZN => n35);
   U67 : INV_X1 port map( A => S(1), ZN => n44);
   U68 : INV_X1 port map( A => S(0), ZN => n45);
   U69 : AOI22_X1 port map( A1 => B(8), A2 => n43, B1 => A(8), B2 => n41, ZN =>
                           n49);
   U70 : AOI22_X1 port map( A1 => D(8), A2 => n39, B1 => C(8), B2 => n37, ZN =>
                           n48);
   U71 : NAND2_X1 port map( A1 => n49, A2 => n48, ZN => Z(8));
   U72 : AOI22_X1 port map( A1 => D(9), A2 => n39, B1 => C(9), B2 => n37, ZN =>
                           n50);
   U73 : AOI22_X1 port map( A1 => D(10), A2 => n39, B1 => C(10), B2 => n37, ZN 
                           => n51);
   U74 : AOI22_X1 port map( A1 => D(11), A2 => n39, B1 => C(11), B2 => n37, ZN 
                           => n52);
   U75 : AOI22_X1 port map( A1 => B(12), A2 => n43, B1 => A(12), B2 => n41, ZN 
                           => n54);
   U76 : AOI22_X1 port map( A1 => D(12), A2 => n39, B1 => C(12), B2 => n37, ZN 
                           => n53);
   U77 : NAND2_X1 port map( A1 => n54, A2 => n53, ZN => Z(12));
   U78 : AOI22_X1 port map( A1 => B(13), A2 => n43, B1 => A(13), B2 => n41, ZN 
                           => n56);
   U79 : AOI22_X1 port map( A1 => D(13), A2 => n39, B1 => C(13), B2 => n37, ZN 
                           => n55);
   U80 : NAND2_X1 port map( A1 => n56, A2 => n55, ZN => Z(13));
   U81 : AOI22_X1 port map( A1 => B(14), A2 => n43, B1 => A(14), B2 => n41, ZN 
                           => n58);
   U82 : AOI22_X1 port map( A1 => D(14), A2 => n39, B1 => C(14), B2 => n37, ZN 
                           => n57);
   U83 : NAND2_X1 port map( A1 => n58, A2 => n57, ZN => Z(14));
   U84 : AOI22_X1 port map( A1 => D(15), A2 => n39, B1 => C(15), B2 => n37, ZN 
                           => n59);
   U85 : NAND2_X1 port map( A1 => n60, A2 => n59, ZN => Z(15));
   U86 : AOI22_X1 port map( A1 => B(16), A2 => n43, B1 => A(16), B2 => n41, ZN 
                           => n62);
   U87 : AOI22_X1 port map( A1 => D(16), A2 => n39, B1 => C(16), B2 => n37, ZN 
                           => n61);
   U88 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => Z(16));
   U89 : AOI22_X1 port map( A1 => D(17), A2 => n39, B1 => C(17), B2 => n37, ZN 
                           => n63);
   U90 : AOI22_X1 port map( A1 => B(18), A2 => n43, B1 => A(18), B2 => n41, ZN 
                           => n65);
   U91 : AOI22_X1 port map( A1 => D(18), A2 => n39, B1 => C(18), B2 => n37, ZN 
                           => n64);
   U92 : NAND2_X1 port map( A1 => n65, A2 => n64, ZN => Z(18));
   U93 : AOI22_X1 port map( A1 => D(19), A2 => n39, B1 => C(19), B2 => n37, ZN 
                           => n66);
   U94 : AOI22_X1 port map( A1 => D(20), A2 => n39, B1 => C(20), B2 => n37, ZN 
                           => n67);
   U95 : AOI22_X1 port map( A1 => B(21), A2 => n43, B1 => A(21), B2 => n41, ZN 
                           => n71);
   U96 : AOI22_X1 port map( A1 => D(21), A2 => n39, B1 => C(21), B2 => n37, ZN 
                           => n70);
   U97 : NAND2_X1 port map( A1 => n71, A2 => n70, ZN => Z(21));
   U98 : AOI22_X1 port map( A1 => B(22), A2 => n43, B1 => A(22), B2 => n41, ZN 
                           => n73);
   U99 : AOI22_X1 port map( A1 => D(22), A2 => n39, B1 => C(22), B2 => n37, ZN 
                           => n72);
   U100 : NAND2_X1 port map( A1 => n73, A2 => n72, ZN => Z(22));
   U101 : AOI22_X1 port map( A1 => B(23), A2 => n43, B1 => A(23), B2 => n41, ZN
                           => n75);
   U102 : AOI22_X1 port map( A1 => D(23), A2 => n39, B1 => C(23), B2 => n37, ZN
                           => n74);
   U103 : NAND2_X1 port map( A1 => n75, A2 => n74, ZN => Z(23));
   U104 : AOI22_X1 port map( A1 => B(24), A2 => n43, B1 => A(24), B2 => n41, ZN
                           => n77);
   U105 : AOI22_X1 port map( A1 => D(24), A2 => n39, B1 => C(24), B2 => n37, ZN
                           => n76);
   U106 : NAND2_X1 port map( A1 => n77, A2 => n76, ZN => Z(24));
   U107 : AOI22_X1 port map( A1 => D(25), A2 => n38, B1 => C(25), B2 => n36, ZN
                           => n78);
   U108 : AOI22_X1 port map( A1 => B(26), A2 => n42, B1 => A(26), B2 => n40, ZN
                           => n80);
   U109 : AOI22_X1 port map( A1 => D(26), A2 => n38, B1 => C(26), B2 => n36, ZN
                           => n79);
   U110 : NAND2_X1 port map( A1 => n80, A2 => n79, ZN => Z(26));
   U111 : AOI22_X1 port map( A1 => D(27), A2 => n38, B1 => C(27), B2 => n36, ZN
                           => n81);
   U112 : NAND2_X1 port map( A1 => n82, A2 => n81, ZN => Z(27));
   U113 : AOI22_X1 port map( A1 => D(28), A2 => n38, B1 => C(28), B2 => n36, ZN
                           => n83);
   U114 : NAND2_X1 port map( A1 => n84, A2 => n83, ZN => Z(28));
   U115 : AOI22_X1 port map( A1 => B(29), A2 => n42, B1 => A(29), B2 => n40, ZN
                           => n86);
   U116 : AOI22_X1 port map( A1 => D(29), A2 => n38, B1 => C(29), B2 => n36, ZN
                           => n85);
   U117 : NAND2_X1 port map( A1 => n86, A2 => n85, ZN => Z(29));
   U118 : AOI22_X1 port map( A1 => B(30), A2 => n42, B1 => A(30), B2 => n40, ZN
                           => n88);
   U119 : AOI22_X1 port map( A1 => D(30), A2 => n38, B1 => C(30), B2 => n36, ZN
                           => n87);
   U120 : NAND2_X1 port map( A1 => n88, A2 => n87, ZN => Z(30));
   U121 : AOI22_X1 port map( A1 => D(31), A2 => n38, B1 => C(31), B2 => n36, ZN
                           => n89);
   U122 : NAND2_X1 port map( A1 => n90, A2 => n89, ZN => Z(31));

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_1 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_1;

architecture SYN_bhv of mux41_NBIT32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n145, Z => n72);
   U2 : BUF_X1 port map( A => n145, Z => n73);
   U3 : BUF_X1 port map( A => n147, Z => n78);
   U4 : BUF_X1 port map( A => n147, Z => n79);
   U5 : BUF_X1 port map( A => n144, Z => n1);
   U6 : BUF_X1 port map( A => n144, Z => n70);
   U7 : BUF_X1 port map( A => n146, Z => n75);
   U8 : BUF_X1 port map( A => n146, Z => n76);
   U9 : BUF_X1 port map( A => n145, Z => n74);
   U10 : BUF_X1 port map( A => n147, Z => n80);
   U11 : BUF_X1 port map( A => n144, Z => n71);
   U12 : BUF_X1 port map( A => n146, Z => n77);
   U13 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n144);
   U14 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n145);
   U15 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n147);
   U16 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n146);
   U17 : INV_X1 port map( A => S(0), ZN => n81);
   U18 : NAND2_X1 port map( A1 => n83, A2 => n82, ZN => Z(0));
   U19 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n83);
   U20 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n82);
   U21 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(31));
   U22 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN 
                           => n130);
   U23 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN 
                           => n131);
   U24 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(7));
   U25 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n140);
   U26 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n141);
   U27 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(8));
   U28 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n142);
   U29 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n143);
   U30 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(9));
   U31 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN =>
                           n148);
   U32 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN =>
                           n149);
   U33 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => Z(12));
   U34 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN 
                           => n88);
   U35 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n89);
   U36 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => Z(13));
   U37 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN 
                           => n90);
   U38 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n91);
   U39 : NAND2_X1 port map( A1 => n93, A2 => n92, ZN => Z(14));
   U40 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN 
                           => n92);
   U41 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n93);
   U42 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(17));
   U43 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n98);
   U44 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n99);
   U45 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => Z(15));
   U46 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN 
                           => n94);
   U47 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n95);
   U48 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(18));
   U49 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n100);
   U50 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n101);
   U51 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(16));
   U52 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n96);
   U53 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n97);
   U54 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(19));
   U55 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN 
                           => n102);
   U56 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n103);
   U57 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(20));
   U58 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN 
                           => n106);
   U59 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN 
                           => n107);
   U60 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(21));
   U61 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n108);
   U62 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n109);
   U63 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(22));
   U64 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n110);
   U65 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n111);
   U66 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(23));
   U67 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN 
                           => n112);
   U68 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN 
                           => n113);
   U69 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(24));
   U70 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN 
                           => n114);
   U71 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN 
                           => n115);
   U72 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(25));
   U73 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n116);
   U74 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n117);
   U75 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(6));
   U76 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n138);
   U77 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n139);
   U78 : NAND2_X1 port map( A1 => n85, A2 => n84, ZN => Z(10));
   U79 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN 
                           => n84);
   U80 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n85);
   U81 : NAND2_X1 port map( A1 => n87, A2 => n86, ZN => Z(11));
   U82 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN 
                           => n86);
   U83 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n87);
   U84 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(26));
   U85 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n118);
   U86 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n119);
   U87 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(27));
   U88 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN 
                           => n120);
   U89 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN 
                           => n121);
   U90 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(5));
   U91 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN =>
                           n136);
   U92 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN =>
                           n137);
   U93 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(28));
   U94 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n122);
   U95 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n123);
   U96 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(29));
   U97 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n124);
   U98 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n125);
   U99 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(30));
   U100 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN
                           => n128);
   U101 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN
                           => n129);
   U102 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(2));
   U103 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN 
                           => n126);
   U104 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN 
                           => n127);
   U105 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(1));
   U106 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN 
                           => n104);
   U107 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN =>
                           n105);
   U108 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(3));
   U109 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN 
                           => n132);
   U110 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN 
                           => n133);
   U111 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(4));
   U112 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN 
                           => n134);
   U113 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN 
                           => n135);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_4 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_4;

architecture SYN_bhv of regn_N5_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n16, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n21);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n17, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n22);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n18, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n23);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n19, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n24);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n20, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n25);
   U2 : OAI21_X1 port map( B1 => n25, B2 => EN, A => n30, ZN => n20);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n30);
   U4 : OAI21_X1 port map( B1 => n24, B2 => EN, A => n29, ZN => n19);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n29);
   U6 : OAI21_X1 port map( B1 => n23, B2 => EN, A => n28, ZN => n18);
   U7 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n28);
   U8 : OAI21_X1 port map( B1 => n22, B2 => EN, A => n27, ZN => n17);
   U9 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n27);
   U10 : OAI21_X1 port map( B1 => n21, B2 => EN, A => n26, ZN => n16);
   U11 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n26);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_3 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_3;

architecture SYN_bhv of regn_N5_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n16, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n21);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n17, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n22);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n18, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n23);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n19, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n24);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n20, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n25);
   U2 : OAI21_X1 port map( B1 => n25, B2 => EN, A => n30, ZN => n20);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n30);
   U4 : OAI21_X1 port map( B1 => n24, B2 => EN, A => n29, ZN => n19);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n29);
   U6 : OAI21_X1 port map( B1 => n23, B2 => EN, A => n28, ZN => n18);
   U7 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n28);
   U8 : OAI21_X1 port map( B1 => n22, B2 => EN, A => n27, ZN => n17);
   U9 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n27);
   U10 : OAI21_X1 port map( B1 => n21, B2 => EN, A => n26, ZN => n16);
   U11 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n26);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_2 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_2;

architecture SYN_bhv of regn_N5_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n16, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n21);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n17, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n22);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n18, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n23);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n19, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n24);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n20, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n25);
   U2 : OAI21_X1 port map( B1 => n25, B2 => EN, A => n30, ZN => n20);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n30);
   U4 : OAI21_X1 port map( B1 => n24, B2 => EN, A => n29, ZN => n19);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n29);
   U6 : OAI21_X1 port map( B1 => n23, B2 => EN, A => n28, ZN => n18);
   U7 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n28);
   U8 : OAI21_X1 port map( B1 => n22, B2 => EN, A => n27, ZN => n17);
   U9 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n27);
   U10 : OAI21_X1 port map( B1 => n21, B2 => EN, A => n26, ZN => n16);
   U11 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n26);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_1 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_1;

architecture SYN_bhv of regn_N5_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n16, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n21);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n17, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n22);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n18, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n23);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n19, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n24);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n20, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n25);
   U2 : OAI21_X1 port map( B1 => n25, B2 => EN, A => n30, ZN => n20);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n30);
   U4 : OAI21_X1 port map( B1 => n24, B2 => EN, A => n29, ZN => n19);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n29);
   U6 : OAI21_X1 port map( B1 => n23, B2 => EN, A => n28, ZN => n18);
   U7 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n28);
   U8 : OAI21_X1 port map( B1 => n22, B2 => EN, A => n27, ZN => n17);
   U9 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n27);
   U10 : OAI21_X1 port map( B1 => n21, B2 => EN, A => n26, ZN => n16);
   U11 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n26);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_10 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_10;

architecture SYN_bhv of regn_N32_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U6 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U7 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U8 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U9 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U10 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U11 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U12 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U13 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U14 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U15 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U16 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U17 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U18 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U19 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U20 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U21 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U22 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U23 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U24 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U25 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U26 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U27 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U28 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U29 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U30 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U31 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U32 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U33 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U34 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U35 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U36 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U37 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U38 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U39 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U40 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U41 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U42 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U43 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U44 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U45 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U46 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U47 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U48 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U49 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U50 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U51 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U52 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U53 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U54 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U55 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U56 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U57 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U58 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U59 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U60 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U61 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_9 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_9;

architecture SYN_bhv of regn_N32_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U6 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U7 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U8 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U9 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U10 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U11 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U12 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U13 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U14 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U15 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U16 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U17 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U18 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U19 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U20 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U21 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U22 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U23 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U24 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U25 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U26 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U27 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U28 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U29 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U30 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U31 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U32 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U33 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U34 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U35 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U36 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U37 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U38 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U39 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U40 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U41 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U42 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U43 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U44 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U45 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U46 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U47 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U48 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U49 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U50 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U51 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U52 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U53 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U54 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U55 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U56 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U57 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U58 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U59 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U60 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U61 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U62 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U63 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U64 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);
   U65 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U66 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U67 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U68 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_8 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_8;

architecture SYN_bhv of regn_N32_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U6 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U7 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U8 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U9 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U10 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U11 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U12 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U13 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U14 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U15 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U16 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U17 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U18 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U19 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U20 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U21 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U22 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U23 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U24 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U25 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U26 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U27 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U28 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U29 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U30 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U31 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U32 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U33 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U34 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U35 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U36 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U37 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U38 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U39 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U40 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U41 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U42 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U43 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U44 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U45 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U46 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U47 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U48 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U49 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U50 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U51 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U52 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U53 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U54 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U55 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U56 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U57 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U58 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U59 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U60 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U61 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U62 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U63 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U64 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);
   U65 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U66 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U67 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U68 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_7 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_7;

architecture SYN_bhv of regn_N32_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_6 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_6;

architecture SYN_bhv of regn_N32_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_5 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_5;

architecture SYN_bhv of regn_N32_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_4 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_4;

architecture SYN_bhv of regn_N32_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_3 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_3;

architecture SYN_bhv of regn_N32_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_2 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_2;

architecture SYN_bhv of regn_N32_2 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U4 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U6 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U7 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U8 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U9 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U10 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U11 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U12 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U13 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U14 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U15 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U16 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U17 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U18 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U19 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U20 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U21 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U22 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U23 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U24 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U25 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U26 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U27 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U28 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U29 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U30 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U31 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U32 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U33 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U34 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U35 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U36 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U37 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U38 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U39 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U40 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U41 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U42 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U43 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U44 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U45 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U46 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U47 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U48 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U49 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U50 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U51 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U52 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U53 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U54 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U55 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U56 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U57 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U58 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U59 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U60 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U61 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U62 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U63 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U64 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U65 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);
   U66 : BUF_X1 port map( A => RST, Z => n97);
   U67 : BUF_X1 port map( A => RST, Z => n98);
   U68 : BUF_X1 port map( A => RST, Z => n99);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_1 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_1;

architecture SYN_bhv of regn_N32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U4 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U6 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U7 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U8 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U9 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U10 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U11 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U12 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U13 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U14 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U15 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U16 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U17 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U18 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U19 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U20 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U21 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U22 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U23 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U24 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U25 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U26 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U27 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U28 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U29 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U30 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U31 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U32 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U33 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U34 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U35 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U36 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U37 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U38 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U39 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U40 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U41 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U42 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U43 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U44 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U45 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U46 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U47 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U48 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U49 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U50 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U51 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U52 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U53 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U54 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U55 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U56 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U57 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U58 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U59 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U60 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U61 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U62 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U63 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U64 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U65 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);
   U66 : BUF_X1 port map( A => RST, Z => n97);
   U67 : BUF_X1 port map( A => RST, Z => n98);
   U68 : BUF_X1 port map( A => RST, Z => n99);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_5;

architecture SYN_bhv of mux21_NBIT32_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n15, ZN => n5);
   U2 : INV_X1 port map( A => n15, ZN => n4);
   U3 : BUF_X1 port map( A => n3, Z => n15);
   U4 : BUF_X1 port map( A => n2, Z => n11);
   U5 : BUF_X1 port map( A => n1, Z => n8);
   U6 : BUF_X1 port map( A => n2, Z => n10);
   U7 : BUF_X1 port map( A => n1, Z => n9);
   U8 : BUF_X1 port map( A => n3, Z => n14);
   U9 : BUF_X1 port map( A => n1, Z => n7);
   U10 : BUF_X1 port map( A => n3, Z => n13);
   U11 : BUF_X1 port map( A => n2, Z => n12);
   U12 : BUF_X1 port map( A => S, Z => n3);
   U13 : BUF_X1 port map( A => S, Z => n2);
   U14 : BUF_X1 port map( A => S, Z => n1);
   U15 : INV_X1 port map( A => n107, ZN => Z(5));
   U16 : INV_X1 port map( A => n99, ZN => Z(27));
   U17 : INV_X1 port map( A => n82, ZN => Z(11));
   U18 : INV_X1 port map( A => n83, ZN => Z(12));
   U19 : INV_X1 port map( A => n84, ZN => Z(13));
   U20 : INV_X1 port map( A => n87, ZN => Z(16));
   U21 : INV_X1 port map( A => n88, ZN => Z(17));
   U22 : INV_X1 port map( A => n89, ZN => Z(18));
   U23 : INV_X1 port map( A => n92, ZN => Z(20));
   U24 : INV_X1 port map( A => n96, ZN => Z(24));
   U25 : INV_X1 port map( A => n98, ZN => Z(26));
   U26 : INV_X1 port map( A => n108, ZN => Z(6));
   U27 : INV_X1 port map( A => n81, ZN => Z(10));
   U28 : INV_X1 port map( A => n102, ZN => Z(2));
   U29 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => n8, ZN => 
                           n102);
   U30 : INV_X1 port map( A => n110, ZN => Z(8));
   U31 : INV_X1 port map( A => n91, ZN => Z(1));
   U32 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n11, ZN => 
                           n91);
   U33 : INV_X1 port map( A => n80, ZN => Z(0));
   U34 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => n14, ZN => 
                           n80);
   U35 : INV_X1 port map( A => n85, ZN => Z(14));
   U36 : INV_X1 port map( A => n90, ZN => Z(19));
   U37 : INV_X1 port map( A => n105, ZN => Z(3));
   U38 : INV_X1 port map( A => n109, ZN => Z(7));
   U39 : INV_X1 port map( A => n111, ZN => Z(9));
   U40 : INV_X1 port map( A => n86, ZN => Z(15));
   U41 : INV_X1 port map( A => n97, ZN => Z(25));
   U42 : INV_X1 port map( A => n106, ZN => Z(4));
   U43 : AOI22_X1 port map( A1 => A(4), A2 => n6, B1 => B(4), B2 => n8, ZN => 
                           n106);
   U44 : INV_X1 port map( A => n93, ZN => Z(21));
   U45 : AOI22_X1 port map( A1 => A(21), A2 => n5, B1 => B(21), B2 => n11, ZN 
                           => n93);
   U46 : INV_X1 port map( A => n94, ZN => Z(22));
   U47 : AOI22_X1 port map( A1 => A(22), A2 => n5, B1 => B(22), B2 => n10, ZN 
                           => n94);
   U48 : INV_X1 port map( A => n95, ZN => Z(23));
   U49 : AOI22_X1 port map( A1 => A(23), A2 => n5, B1 => B(23), B2 => n10, ZN 
                           => n95);
   U50 : INV_X1 port map( A => n100, ZN => Z(28));
   U51 : AOI22_X1 port map( A1 => A(28), A2 => n5, B1 => B(28), B2 => n9, ZN =>
                           n100);
   U52 : INV_X1 port map( A => n101, ZN => Z(29));
   U53 : AOI22_X1 port map( A1 => A(29), A2 => n5, B1 => B(29), B2 => n9, ZN =>
                           n101);
   U54 : INV_X1 port map( A => n103, ZN => Z(30));
   U55 : AOI22_X1 port map( A1 => A(30), A2 => n5, B1 => B(30), B2 => n11, ZN 
                           => n103);
   U56 : INV_X1 port map( A => n104, ZN => Z(31));
   U57 : AOI22_X1 port map( A1 => A(31), A2 => n6, B1 => B(31), B2 => n8, ZN =>
                           n104);
   U58 : AOI22_X1 port map( A1 => A(20), A2 => n5, B1 => B(20), B2 => n11, ZN 
                           => n92);
   U59 : AOI22_X1 port map( A1 => A(27), A2 => n5, B1 => B(27), B2 => n9, ZN =>
                           n99);
   U60 : AOI22_X1 port map( A1 => A(24), A2 => n5, B1 => B(24), B2 => n10, ZN 
                           => n96);
   U61 : AOI22_X1 port map( A1 => A(25), A2 => n5, B1 => B(25), B2 => n10, ZN 
                           => n97);
   U62 : AOI22_X1 port map( A1 => A(26), A2 => n5, B1 => B(26), B2 => n9, ZN =>
                           n98);
   U63 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n13, ZN 
                           => n86);
   U64 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => B(11), B2 => n14, ZN 
                           => n82);
   U65 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n13, ZN 
                           => n84);
   U66 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => B(12), B2 => n13, ZN 
                           => n83);
   U67 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => B(19), B2 => n12, ZN 
                           => n90);
   U68 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n12, ZN 
                           => n88);
   U69 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => B(18), B2 => n12, ZN 
                           => n89);
   U70 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => B(16), B2 => n12, ZN 
                           => n87);
   U71 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n13, ZN 
                           => n85);
   U72 : AOI22_X1 port map( A1 => A(5), A2 => n6, B1 => B(5), B2 => n7, ZN => 
                           n107);
   U73 : AOI22_X1 port map( A1 => A(7), A2 => n6, B1 => B(7), B2 => n7, ZN => 
                           n109);
   U74 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => B(10), B2 => n14, ZN 
                           => n81);
   U75 : AOI22_X1 port map( A1 => A(3), A2 => n6, B1 => B(3), B2 => n8, ZN => 
                           n105);
   U76 : AOI22_X1 port map( A1 => A(6), A2 => n6, B1 => B(6), B2 => n7, ZN => 
                           n108);
   U77 : AOI22_X1 port map( A1 => A(8), A2 => n6, B1 => B(8), B2 => n7, ZN => 
                           n110);
   U78 : AOI22_X1 port map( A1 => A(9), A2 => n6, B1 => n14, B2 => B(9), ZN => 
                           n111);
   U79 : INV_X1 port map( A => n15, ZN => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_4;

architecture SYN_bhv of mux21_NBIT32_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => n4);
   U2 : INV_X1 port map( A => n14, ZN => n5);
   U3 : BUF_X1 port map( A => n1, Z => n6);
   U4 : BUF_X1 port map( A => n3, Z => n12);
   U5 : BUF_X1 port map( A => n2, Z => n11);
   U6 : BUF_X1 port map( A => n2, Z => n9);
   U7 : BUF_X1 port map( A => n1, Z => n8);
   U8 : BUF_X1 port map( A => n2, Z => n10);
   U9 : BUF_X1 port map( A => n1, Z => n7);
   U10 : BUF_X1 port map( A => n3, Z => n14);
   U11 : BUF_X1 port map( A => n3, Z => n13);
   U12 : BUF_X1 port map( A => S, Z => n3);
   U13 : BUF_X1 port map( A => S, Z => n2);
   U14 : BUF_X1 port map( A => S, Z => n1);
   U15 : INV_X1 port map( A => n90, ZN => Z(1));
   U16 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n10, ZN => 
                           n90);
   U17 : INV_X1 port map( A => n101, ZN => Z(2));
   U18 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           n101);
   U19 : INV_X1 port map( A => n104, ZN => Z(3));
   U20 : AOI22_X1 port map( A1 => A(3), A2 => n4, B1 => B(3), B2 => n7, ZN => 
                           n104);
   U21 : INV_X1 port map( A => n105, ZN => Z(4));
   U22 : AOI22_X1 port map( A1 => A(4), A2 => n5, B1 => B(4), B2 => n7, ZN => 
                           n105);
   U23 : INV_X1 port map( A => n106, ZN => Z(5));
   U24 : AOI22_X1 port map( A1 => A(5), A2 => n4, B1 => B(5), B2 => n6, ZN => 
                           n106);
   U25 : INV_X1 port map( A => n107, ZN => Z(6));
   U26 : AOI22_X1 port map( A1 => A(6), A2 => n5, B1 => B(6), B2 => n6, ZN => 
                           n107);
   U27 : INV_X1 port map( A => n108, ZN => Z(7));
   U28 : AOI22_X1 port map( A1 => A(7), A2 => n4, B1 => B(7), B2 => n6, ZN => 
                           n108);
   U29 : INV_X1 port map( A => n109, ZN => Z(8));
   U30 : AOI22_X1 port map( A1 => A(8), A2 => n5, B1 => B(8), B2 => n6, ZN => 
                           n109);
   U31 : INV_X1 port map( A => n80, ZN => Z(10));
   U32 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => B(10), B2 => n13, ZN 
                           => n80);
   U33 : INV_X1 port map( A => n81, ZN => Z(11));
   U34 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => B(11), B2 => n13, ZN 
                           => n81);
   U35 : INV_X1 port map( A => n82, ZN => Z(12));
   U36 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => B(12), B2 => n12, ZN 
                           => n82);
   U37 : INV_X1 port map( A => n83, ZN => Z(13));
   U38 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n12, ZN 
                           => n83);
   U39 : INV_X1 port map( A => n84, ZN => Z(14));
   U40 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n12, ZN 
                           => n84);
   U41 : INV_X1 port map( A => n85, ZN => Z(15));
   U42 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n12, ZN 
                           => n85);
   U43 : INV_X1 port map( A => n86, ZN => Z(16));
   U44 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => B(16), B2 => n11, ZN 
                           => n86);
   U45 : INV_X1 port map( A => n87, ZN => Z(17));
   U46 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n11, ZN 
                           => n87);
   U47 : INV_X1 port map( A => n88, ZN => Z(18));
   U48 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => B(18), B2 => n11, ZN 
                           => n88);
   U49 : INV_X1 port map( A => n89, ZN => Z(19));
   U50 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => B(19), B2 => n11, ZN 
                           => n89);
   U51 : INV_X1 port map( A => n91, ZN => Z(20));
   U52 : AOI22_X1 port map( A1 => A(20), A2 => n5, B1 => B(20), B2 => n10, ZN 
                           => n91);
   U53 : INV_X1 port map( A => n92, ZN => Z(21));
   U54 : AOI22_X1 port map( A1 => A(21), A2 => n5, B1 => B(21), B2 => n10, ZN 
                           => n92);
   U55 : INV_X1 port map( A => n93, ZN => Z(22));
   U56 : AOI22_X1 port map( A1 => A(22), A2 => n5, B1 => B(22), B2 => n9, ZN =>
                           n93);
   U57 : INV_X1 port map( A => n94, ZN => Z(23));
   U58 : AOI22_X1 port map( A1 => A(23), A2 => n5, B1 => B(23), B2 => n9, ZN =>
                           n94);
   U59 : INV_X1 port map( A => n95, ZN => Z(24));
   U60 : AOI22_X1 port map( A1 => A(24), A2 => n5, B1 => B(24), B2 => n9, ZN =>
                           n95);
   U61 : INV_X1 port map( A => n96, ZN => Z(25));
   U62 : AOI22_X1 port map( A1 => A(25), A2 => n5, B1 => B(25), B2 => n9, ZN =>
                           n96);
   U63 : INV_X1 port map( A => n97, ZN => Z(26));
   U64 : AOI22_X1 port map( A1 => A(26), A2 => n5, B1 => B(26), B2 => n8, ZN =>
                           n97);
   U65 : INV_X1 port map( A => n98, ZN => Z(27));
   U66 : AOI22_X1 port map( A1 => A(27), A2 => n5, B1 => B(27), B2 => n8, ZN =>
                           n98);
   U67 : INV_X1 port map( A => n99, ZN => Z(28));
   U68 : AOI22_X1 port map( A1 => A(28), A2 => n5, B1 => B(28), B2 => n8, ZN =>
                           n99);
   U69 : INV_X1 port map( A => n100, ZN => Z(29));
   U70 : AOI22_X1 port map( A1 => A(29), A2 => n5, B1 => B(29), B2 => n8, ZN =>
                           n100);
   U71 : INV_X1 port map( A => n102, ZN => Z(30));
   U72 : AOI22_X1 port map( A1 => A(30), A2 => n5, B1 => B(30), B2 => n10, ZN 
                           => n102);
   U73 : INV_X1 port map( A => n103, ZN => Z(31));
   U74 : AOI22_X1 port map( A1 => A(31), A2 => n4, B1 => B(31), B2 => n7, ZN =>
                           n103);
   U75 : INV_X1 port map( A => n110, ZN => Z(9));
   U76 : AOI22_X1 port map( A1 => A(9), A2 => n5, B1 => n13, B2 => B(9), ZN => 
                           n110);
   U77 : INV_X1 port map( A => n79, ZN => Z(0));
   U78 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => n13, ZN => 
                           n79);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_3;

architecture SYN_bhv of mux21_NBIT32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n68, Z => n1);
   U2 : BUF_X1 port map( A => n68, Z => n2);
   U3 : BUF_X1 port map( A => n68, Z => n3);
   U4 : INV_X1 port map( A => n69, ZN => Z(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => S, ZN => n69
                           );
   U6 : INV_X1 port map( A => n81, ZN => Z(20));
   U7 : AOI22_X1 port map( A1 => A(20), A2 => n2, B1 => B(20), B2 => S, ZN => 
                           n81);
   U8 : INV_X1 port map( A => n73, ZN => Z(13));
   U9 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => S, ZN => 
                           n73);
   U10 : INV_X1 port map( A => n77, ZN => Z(17));
   U11 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => S, ZN => 
                           n77);
   U12 : INV_X1 port map( A => n97, ZN => Z(6));
   U13 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => S, ZN => 
                           n97);
   U14 : INV_X1 port map( A => n85, ZN => Z(24));
   U15 : AOI22_X1 port map( A1 => A(24), A2 => n2, B1 => B(24), B2 => S, ZN => 
                           n85);
   U16 : INV_X1 port map( A => n89, ZN => Z(28));
   U17 : AOI22_X1 port map( A1 => A(28), A2 => n2, B1 => B(28), B2 => S, ZN => 
                           n89);
   U18 : INV_X1 port map( A => n93, ZN => Z(31));
   U19 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => S, ZN => 
                           n93);
   U20 : INV_X1 port map( A => n70, ZN => Z(10));
   U21 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => S, ZN => 
                           n70);
   U22 : INV_X1 port map( A => n82, ZN => Z(21));
   U23 : AOI22_X1 port map( A1 => A(21), A2 => n2, B1 => B(21), B2 => S, ZN => 
                           n82);
   U24 : INV_X1 port map( A => n74, ZN => Z(14));
   U25 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => S, ZN => 
                           n74);
   U26 : INV_X1 port map( A => n78, ZN => Z(18));
   U27 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => S, ZN => 
                           n78);
   U28 : INV_X1 port map( A => n86, ZN => Z(25));
   U29 : AOI22_X1 port map( A1 => A(25), A2 => n2, B1 => B(25), B2 => S, ZN => 
                           n86);
   U30 : INV_X1 port map( A => n90, ZN => Z(29));
   U31 : AOI22_X1 port map( A1 => A(29), A2 => n2, B1 => B(29), B2 => S, ZN => 
                           n90);
   U32 : INV_X1 port map( A => n94, ZN => Z(3));
   U33 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => S, ZN => 
                           n94);
   U34 : INV_X1 port map( A => n98, ZN => Z(7));
   U35 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => S, ZN => 
                           n98);
   U36 : INV_X1 port map( A => n95, ZN => Z(4));
   U37 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => S, ZN => 
                           n95);
   U38 : INV_X1 port map( A => n83, ZN => Z(22));
   U39 : AOI22_X1 port map( A1 => A(22), A2 => n2, B1 => B(22), B2 => S, ZN => 
                           n83);
   U40 : INV_X1 port map( A => n91, ZN => Z(2));
   U41 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => S, ZN => 
                           n91);
   U42 : INV_X1 port map( A => n99, ZN => Z(8));
   U43 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => S, ZN => 
                           n99);
   U44 : INV_X1 port map( A => n87, ZN => Z(26));
   U45 : AOI22_X1 port map( A1 => A(26), A2 => n2, B1 => B(26), B2 => S, ZN => 
                           n87);
   U46 : INV_X1 port map( A => n71, ZN => Z(11));
   U47 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => S, ZN => 
                           n71);
   U48 : INV_X1 port map( A => n75, ZN => Z(15));
   U49 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => S, ZN => 
                           n75);
   U50 : INV_X1 port map( A => n79, ZN => Z(19));
   U51 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => S, ZN => 
                           n79);
   U52 : INV_X1 port map( A => n76, ZN => Z(16));
   U53 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => S, ZN => 
                           n76);
   U54 : INV_X1 port map( A => n72, ZN => Z(12));
   U55 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => S, ZN => 
                           n72);
   U56 : INV_X1 port map( A => n80, ZN => Z(1));
   U57 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => S, ZN => 
                           n80);
   U58 : INV_X1 port map( A => n96, ZN => Z(5));
   U59 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => S, ZN => 
                           n96);
   U60 : INV_X1 port map( A => n92, ZN => Z(30));
   U61 : AOI22_X1 port map( A1 => A(30), A2 => n2, B1 => B(30), B2 => S, ZN => 
                           n92);
   U62 : INV_X1 port map( A => n84, ZN => Z(23));
   U63 : AOI22_X1 port map( A1 => A(23), A2 => n2, B1 => B(23), B2 => S, ZN => 
                           n84);
   U64 : INV_X1 port map( A => n88, ZN => Z(27));
   U65 : AOI22_X1 port map( A1 => A(27), A2 => n2, B1 => B(27), B2 => S, ZN => 
                           n88);
   U66 : INV_X1 port map( A => n100, ZN => Z(9));
   U67 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => S, B2 => B(9), ZN => 
                           n100);
   U68 : INV_X1 port map( A => S, ZN => n68);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_2;

architecture SYN_bhv of mux21_NBIT32_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n68, Z => n1);
   U2 : BUF_X1 port map( A => n68, Z => n2);
   U3 : BUF_X1 port map( A => n68, Z => n3);
   U4 : INV_X1 port map( A => n81, ZN => Z(20));
   U5 : AOI22_X1 port map( A1 => A(20), A2 => n2, B1 => B(20), B2 => S, ZN => 
                           n81);
   U6 : INV_X1 port map( A => n82, ZN => Z(21));
   U7 : AOI22_X1 port map( A1 => A(21), A2 => n2, B1 => B(21), B2 => S, ZN => 
                           n82);
   U8 : INV_X1 port map( A => n83, ZN => Z(22));
   U9 : AOI22_X1 port map( A1 => A(22), A2 => n2, B1 => B(22), B2 => S, ZN => 
                           n83);
   U10 : INV_X1 port map( A => n84, ZN => Z(23));
   U11 : AOI22_X1 port map( A1 => A(23), A2 => n2, B1 => B(23), B2 => S, ZN => 
                           n84);
   U12 : INV_X1 port map( A => n77, ZN => Z(17));
   U13 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => S, ZN => 
                           n77);
   U14 : INV_X1 port map( A => n78, ZN => Z(18));
   U15 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => S, ZN => 
                           n78);
   U16 : INV_X1 port map( A => n79, ZN => Z(19));
   U17 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => S, ZN => 
                           n79);
   U18 : INV_X1 port map( A => n80, ZN => Z(1));
   U19 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => S, ZN => 
                           n80);
   U20 : INV_X1 port map( A => n73, ZN => Z(13));
   U21 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => S, ZN => 
                           n73);
   U22 : INV_X1 port map( A => n74, ZN => Z(14));
   U23 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => S, ZN => 
                           n74);
   U24 : INV_X1 port map( A => n75, ZN => Z(15));
   U25 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => S, ZN => 
                           n75);
   U26 : INV_X1 port map( A => n76, ZN => Z(16));
   U27 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => S, ZN => 
                           n76);
   U28 : INV_X1 port map( A => n69, ZN => Z(0));
   U29 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => S, ZN => 
                           n69);
   U30 : INV_X1 port map( A => n70, ZN => Z(10));
   U31 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => S, ZN => 
                           n70);
   U32 : INV_X1 port map( A => n71, ZN => Z(11));
   U33 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => S, ZN => 
                           n71);
   U34 : INV_X1 port map( A => n72, ZN => Z(12));
   U35 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => S, ZN => 
                           n72);
   U36 : INV_X1 port map( A => n97, ZN => Z(6));
   U37 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => S, ZN => 
                           n97);
   U38 : INV_X1 port map( A => n98, ZN => Z(7));
   U39 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => S, ZN => 
                           n98);
   U40 : INV_X1 port map( A => n99, ZN => Z(8));
   U41 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => S, ZN => 
                           n99);
   U42 : INV_X1 port map( A => n94, ZN => Z(3));
   U43 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => S, ZN => 
                           n94);
   U44 : INV_X1 port map( A => n95, ZN => Z(4));
   U45 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => S, ZN => 
                           n95);
   U46 : INV_X1 port map( A => n96, ZN => Z(5));
   U47 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => S, ZN => 
                           n96);
   U48 : INV_X1 port map( A => n89, ZN => Z(28));
   U49 : AOI22_X1 port map( A1 => A(28), A2 => n2, B1 => B(28), B2 => S, ZN => 
                           n89);
   U50 : INV_X1 port map( A => n90, ZN => Z(29));
   U51 : AOI22_X1 port map( A1 => A(29), A2 => n2, B1 => B(29), B2 => S, ZN => 
                           n90);
   U52 : INV_X1 port map( A => n91, ZN => Z(2));
   U53 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => S, ZN => 
                           n91);
   U54 : INV_X1 port map( A => n92, ZN => Z(30));
   U55 : AOI22_X1 port map( A1 => A(30), A2 => n2, B1 => B(30), B2 => S, ZN => 
                           n92);
   U56 : INV_X1 port map( A => n85, ZN => Z(24));
   U57 : AOI22_X1 port map( A1 => A(24), A2 => n2, B1 => B(24), B2 => S, ZN => 
                           n85);
   U58 : INV_X1 port map( A => n86, ZN => Z(25));
   U59 : AOI22_X1 port map( A1 => A(25), A2 => n2, B1 => B(25), B2 => S, ZN => 
                           n86);
   U60 : INV_X1 port map( A => n87, ZN => Z(26));
   U61 : AOI22_X1 port map( A1 => A(26), A2 => n2, B1 => B(26), B2 => S, ZN => 
                           n87);
   U62 : INV_X1 port map( A => n88, ZN => Z(27));
   U63 : AOI22_X1 port map( A1 => A(27), A2 => n2, B1 => B(27), B2 => S, ZN => 
                           n88);
   U64 : INV_X1 port map( A => n93, ZN => Z(31));
   U65 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => S, ZN => 
                           n93);
   U66 : INV_X1 port map( A => n100, ZN => Z(9));
   U67 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => S, B2 => B(9), ZN => 
                           n100);
   U68 : INV_X1 port map( A => S, ZN => n68);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_1;

architecture SYN_bhv of mux21_NBIT32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => n4);
   U2 : INV_X1 port map( A => n14, ZN => n5);
   U3 : BUF_X1 port map( A => n1, Z => n6);
   U4 : BUF_X1 port map( A => n3, Z => n12);
   U5 : BUF_X1 port map( A => n2, Z => n11);
   U6 : BUF_X1 port map( A => n2, Z => n9);
   U7 : BUF_X1 port map( A => n1, Z => n8);
   U8 : BUF_X1 port map( A => n2, Z => n10);
   U9 : BUF_X1 port map( A => n1, Z => n7);
   U10 : BUF_X1 port map( A => n3, Z => n14);
   U11 : BUF_X1 port map( A => n3, Z => n13);
   U12 : BUF_X1 port map( A => S, Z => n3);
   U13 : BUF_X1 port map( A => S, Z => n2);
   U14 : BUF_X1 port map( A => S, Z => n1);
   U15 : INV_X1 port map( A => n79, ZN => Z(0));
   U16 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => n13, ZN => 
                           n79);
   U17 : INV_X1 port map( A => n90, ZN => Z(1));
   U18 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n10, ZN => 
                           n90);
   U19 : INV_X1 port map( A => n101, ZN => Z(2));
   U20 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           n101);
   U21 : INV_X1 port map( A => n104, ZN => Z(3));
   U22 : AOI22_X1 port map( A1 => A(3), A2 => n4, B1 => B(3), B2 => n7, ZN => 
                           n104);
   U23 : INV_X1 port map( A => n105, ZN => Z(4));
   U24 : AOI22_X1 port map( A1 => A(4), A2 => n5, B1 => B(4), B2 => n7, ZN => 
                           n105);
   U25 : INV_X1 port map( A => n106, ZN => Z(5));
   U26 : AOI22_X1 port map( A1 => A(5), A2 => n4, B1 => B(5), B2 => n6, ZN => 
                           n106);
   U27 : INV_X1 port map( A => n107, ZN => Z(6));
   U28 : AOI22_X1 port map( A1 => A(6), A2 => n5, B1 => B(6), B2 => n6, ZN => 
                           n107);
   U29 : INV_X1 port map( A => n108, ZN => Z(7));
   U30 : AOI22_X1 port map( A1 => A(7), A2 => n4, B1 => B(7), B2 => n6, ZN => 
                           n108);
   U31 : INV_X1 port map( A => n109, ZN => Z(8));
   U32 : AOI22_X1 port map( A1 => A(8), A2 => n5, B1 => B(8), B2 => n6, ZN => 
                           n109);
   U33 : INV_X1 port map( A => n110, ZN => Z(9));
   U34 : AOI22_X1 port map( A1 => A(9), A2 => n4, B1 => n13, B2 => B(9), ZN => 
                           n110);
   U35 : INV_X1 port map( A => n80, ZN => Z(10));
   U36 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => B(10), B2 => n13, ZN 
                           => n80);
   U37 : INV_X1 port map( A => n81, ZN => Z(11));
   U38 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => B(11), B2 => n13, ZN 
                           => n81);
   U39 : INV_X1 port map( A => n82, ZN => Z(12));
   U40 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => B(12), B2 => n12, ZN 
                           => n82);
   U41 : INV_X1 port map( A => n83, ZN => Z(13));
   U42 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n12, ZN 
                           => n83);
   U43 : INV_X1 port map( A => n84, ZN => Z(14));
   U44 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n12, ZN 
                           => n84);
   U45 : INV_X1 port map( A => n85, ZN => Z(15));
   U46 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n12, ZN 
                           => n85);
   U47 : INV_X1 port map( A => n86, ZN => Z(16));
   U48 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => B(16), B2 => n11, ZN 
                           => n86);
   U49 : INV_X1 port map( A => n87, ZN => Z(17));
   U50 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n11, ZN 
                           => n87);
   U51 : INV_X1 port map( A => n88, ZN => Z(18));
   U52 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => B(18), B2 => n11, ZN 
                           => n88);
   U53 : INV_X1 port map( A => n89, ZN => Z(19));
   U54 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => B(19), B2 => n11, ZN 
                           => n89);
   U55 : INV_X1 port map( A => n91, ZN => Z(20));
   U56 : AOI22_X1 port map( A1 => A(20), A2 => n5, B1 => B(20), B2 => n10, ZN 
                           => n91);
   U57 : INV_X1 port map( A => n92, ZN => Z(21));
   U58 : AOI22_X1 port map( A1 => A(21), A2 => n5, B1 => B(21), B2 => n10, ZN 
                           => n92);
   U59 : INV_X1 port map( A => n93, ZN => Z(22));
   U60 : AOI22_X1 port map( A1 => A(22), A2 => n5, B1 => B(22), B2 => n9, ZN =>
                           n93);
   U61 : INV_X1 port map( A => n94, ZN => Z(23));
   U62 : AOI22_X1 port map( A1 => A(23), A2 => n5, B1 => B(23), B2 => n9, ZN =>
                           n94);
   U63 : INV_X1 port map( A => n95, ZN => Z(24));
   U64 : AOI22_X1 port map( A1 => A(24), A2 => n5, B1 => B(24), B2 => n9, ZN =>
                           n95);
   U65 : INV_X1 port map( A => n96, ZN => Z(25));
   U66 : AOI22_X1 port map( A1 => A(25), A2 => n5, B1 => B(25), B2 => n9, ZN =>
                           n96);
   U67 : INV_X1 port map( A => n97, ZN => Z(26));
   U68 : AOI22_X1 port map( A1 => A(26), A2 => n5, B1 => B(26), B2 => n8, ZN =>
                           n97);
   U69 : INV_X1 port map( A => n98, ZN => Z(27));
   U70 : AOI22_X1 port map( A1 => A(27), A2 => n5, B1 => B(27), B2 => n8, ZN =>
                           n98);
   U71 : INV_X1 port map( A => n99, ZN => Z(28));
   U72 : AOI22_X1 port map( A1 => A(28), A2 => n5, B1 => B(28), B2 => n8, ZN =>
                           n99);
   U73 : INV_X1 port map( A => n100, ZN => Z(29));
   U74 : AOI22_X1 port map( A1 => A(29), A2 => n5, B1 => B(29), B2 => n8, ZN =>
                           n100);
   U75 : INV_X1 port map( A => n102, ZN => Z(30));
   U76 : AOI22_X1 port map( A1 => A(30), A2 => n5, B1 => B(30), B2 => n10, ZN 
                           => n102);
   U77 : INV_X1 port map( A => n103, ZN => Z(31));
   U78 : AOI22_X1 port map( A1 => A(31), A2 => n5, B1 => B(31), B2 => n7, ZN =>
                           n103);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ff_2 is

   port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);

end ff_2;

architecture SYN_bhv of ff_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CLK, RN => RST, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => EN, A => n6, ZN => n4);
   U3 : NAND2_X1 port map( A1 => EN, A2 => D, ZN => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ff_1 is

   port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);

end ff_1;

architecture SYN_bhv of ff_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CLK, RN => RST, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => EN, A => n6, ZN => n4);
   U3 : NAND2_X1 port map( A1 => EN, A2 => D, ZN => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_0;

architecture SYN_STRUCTURAL of RCA_N4_0 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_0;

architecture SYN_struct of carry_select_basic_N4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n6, n7, n8, n9, n1
      , n_1120, n_1121 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1120);
   RCA1 : RCA_N4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1121);
   U3 : INV_X1 port map( A => n7, ZN => S(2));
   U4 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n1, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n7);
   U5 : INV_X1 port map( A => n6, ZN => S(3));
   U6 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n1, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n6);
   U7 : INV_X1 port map( A => n9, ZN => S(0));
   U8 : INV_X1 port map( A => n8, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n1, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n8);
   U10 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n1, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n9);
   U11 : INV_X1 port map( A => C_i, ZN => n1);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_0 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_0;

architecture SYN_bhv of PGblock_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n2);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_0 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_0;

architecture SYN_bhv of Gblock_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_0 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_0;

architecture SYN_bhv of PG_net_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8;

architecture SYN_structural of SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   component carry_select_basic_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CSBI_1 : carry_select_basic_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) 
                           => A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), 
                           B(1) => B(1), B(0) => B(0), C_i => Ci(0), S(3) => 
                           S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CSBI_2 : carry_select_basic_N4_7 port map( A(3) => A(7), A(2) => A(6), A(1) 
                           => A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), 
                           B(1) => B(5), B(0) => B(4), C_i => Ci(1), S(3) => 
                           S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   CSBI_3 : carry_select_basic_N4_6 port map( A(3) => A(11), A(2) => A(10), 
                           A(1) => A(9), A(0) => A(8), B(3) => B(11), B(2) => 
                           B(10), B(1) => B(9), B(0) => B(8), C_i => Ci(2), 
                           S(3) => S(11), S(2) => S(10), S(1) => S(9), S(0) => 
                           S(8));
   CSBI_4 : carry_select_basic_N4_5 port map( A(3) => A(15), A(2) => A(14), 
                           A(1) => A(13), A(0) => A(12), B(3) => B(15), B(2) =>
                           B(14), B(1) => B(13), B(0) => B(12), C_i => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   CSBI_5 : carry_select_basic_N4_4 port map( A(3) => A(19), A(2) => A(18), 
                           A(1) => A(17), A(0) => A(16), B(3) => B(19), B(2) =>
                           B(18), B(1) => B(17), B(0) => B(16), C_i => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   CSBI_6 : carry_select_basic_N4_3 port map( A(3) => A(23), A(2) => A(22), 
                           A(1) => A(21), A(0) => A(20), B(3) => B(23), B(2) =>
                           B(22), B(1) => B(21), B(0) => B(20), C_i => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   CSBI_7 : carry_select_basic_N4_2 port map( A(3) => A(27), A(2) => A(26), 
                           A(1) => A(25), A(0) => A(24), B(3) => B(27), B(2) =>
                           B(26), B(1) => B(25), B(0) => B(24), C_i => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   CSBI_8 : carry_select_basic_N4_1 port map( A(3) => A(31), A(2) => A(30), 
                           A(1) => A(29), A(0) => A(28), B(3) => B(31), B(2) =>
                           B(30), B(1) => B(29), B(0) => B(28), C_i => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_generator_NBIT32_NBIT_PER_BLOCK4 is

   port( A, B : in std_logic_vector (32 downto 1);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end carry_generator_NBIT32_NBIT_PER_BLOCK4;

architecture SYN_struct of carry_generator_NBIT32_NBIT_PER_BLOCK4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component PGblock_1
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_2
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_3
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_4
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_5
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_6
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_7
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_8
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_9
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_10
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_11
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_12
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_13
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_14
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_15
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_16
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_17
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_18
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_19
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_20
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_21
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_22
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_23
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_24
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_25
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_26
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_0
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component Gblock_1
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_2
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_3
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_4
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_5
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_6
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_7
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_8
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_0
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_net_1
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_2
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_3
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_4
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_5
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_6
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_7
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_8
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_9
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_10
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_11
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_12
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_13
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_14
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_15
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_16
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_17
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_18
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_19
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_20
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_21
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_22
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_23
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_24
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_25
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_26
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_27
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_28
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_29
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_30
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_0
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   signal Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port, G_16_16_port, G_16_15_port, G_16_13_port, 
      G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, G_13_13_port, 
      G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, G_10_10_port, 
      G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port, G_7_7_port, 
      G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port, G_3_3_port, 
      G_2_2_port, G_2_1_port, G_1_1_port, P_16_16_port, P_16_15_port, 
      P_16_13_port, P_16_9_port, P_15_15_port, P_14_14_port, P_14_13_port, 
      P_13_13_port, P_12_12_port, P_12_11_port, P_12_9_port, P_11_11_port, 
      P_10_10_port, P_10_9_port, P_9_9_port, P_8_8_port, P_8_7_port, P_8_5_port
      , P_7_7_port, P_6_6_port, P_6_5_port, P_5_5_port, P_4_4_port, P_4_3_port,
      P_3_3_port, P_2_2_port, G_32_32_port, G_32_31_port, G_32_29_port, 
      G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, G_30_29_port, 
      G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, G_28_17_port, 
      G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, G_24_24_port, 
      G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, G_22_22_port, 
      G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, G_20_17_port, 
      G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, P_32_32_port, 
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n3, n1, n2 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port );
   
   PGnetblock_2 : PG_net_0 port map( a => A(2), b => B(2), p => P_2_2_port, g 
                           => G_2_2_port);
   PGnetblock_3 : PG_net_30 port map( a => A(3), b => B(3), p => P_3_3_port, g 
                           => G_3_3_port);
   PGnetblock_4 : PG_net_29 port map( a => A(4), b => B(4), p => P_4_4_port, g 
                           => G_4_4_port);
   PGnetblock_5 : PG_net_28 port map( a => A(5), b => B(5), p => P_5_5_port, g 
                           => G_5_5_port);
   PGnetblock_6 : PG_net_27 port map( a => A(6), b => B(6), p => P_6_6_port, g 
                           => G_6_6_port);
   PGnetblock_7 : PG_net_26 port map( a => A(7), b => B(7), p => P_7_7_port, g 
                           => G_7_7_port);
   PGnetblock_8 : PG_net_25 port map( a => A(8), b => B(8), p => P_8_8_port, g 
                           => G_8_8_port);
   PGnetblock_9 : PG_net_24 port map( a => A(9), b => B(9), p => P_9_9_port, g 
                           => G_9_9_port);
   PGnetblock_10 : PG_net_23 port map( a => A(10), b => B(10), p => 
                           P_10_10_port, g => G_10_10_port);
   PGnetblock_11 : PG_net_22 port map( a => A(11), b => B(11), p => 
                           P_11_11_port, g => G_11_11_port);
   PGnetblock_12 : PG_net_21 port map( a => A(12), b => B(12), p => 
                           P_12_12_port, g => G_12_12_port);
   PGnetblock_13 : PG_net_20 port map( a => A(13), b => B(13), p => 
                           P_13_13_port, g => G_13_13_port);
   PGnetblock_14 : PG_net_19 port map( a => A(14), b => B(14), p => 
                           P_14_14_port, g => G_14_14_port);
   PGnetblock_15 : PG_net_18 port map( a => A(15), b => B(15), p => 
                           P_15_15_port, g => G_15_15_port);
   PGnetblock_16 : PG_net_17 port map( a => A(16), b => B(16), p => 
                           P_16_16_port, g => G_16_16_port);
   PGnetblock_17 : PG_net_16 port map( a => A(17), b => B(17), p => 
                           P_17_17_port, g => G_17_17_port);
   PGnetblock_18 : PG_net_15 port map( a => A(18), b => B(18), p => 
                           P_18_18_port, g => G_18_18_port);
   PGnetblock_19 : PG_net_14 port map( a => A(19), b => B(19), p => 
                           P_19_19_port, g => G_19_19_port);
   PGnetblock_20 : PG_net_13 port map( a => A(20), b => B(20), p => 
                           P_20_20_port, g => G_20_20_port);
   PGnetblock_21 : PG_net_12 port map( a => A(21), b => B(21), p => 
                           P_21_21_port, g => G_21_21_port);
   PGnetblock_22 : PG_net_11 port map( a => A(22), b => B(22), p => 
                           P_22_22_port, g => G_22_22_port);
   PGnetblock_23 : PG_net_10 port map( a => A(23), b => B(23), p => 
                           P_23_23_port, g => G_23_23_port);
   PGnetblock_24 : PG_net_9 port map( a => A(24), b => B(24), p => P_24_24_port
                           , g => G_24_24_port);
   PGnetblock_25 : PG_net_8 port map( a => A(25), b => B(25), p => P_25_25_port
                           , g => G_25_25_port);
   PGnetblock_26 : PG_net_7 port map( a => A(26), b => B(26), p => P_26_26_port
                           , g => G_26_26_port);
   PGnetblock_27 : PG_net_6 port map( a => A(27), b => B(27), p => P_27_27_port
                           , g => G_27_27_port);
   PGnetblock_28 : PG_net_5 port map( a => A(28), b => B(28), p => P_28_28_port
                           , g => G_28_28_port);
   PGnetblock_29 : PG_net_4 port map( a => A(29), b => B(29), p => P_29_29_port
                           , g => G_29_29_port);
   PGnetblock_30 : PG_net_3 port map( a => A(30), b => B(30), p => P_30_30_port
                           , g => G_30_30_port);
   PGnetblock_31 : PG_net_2 port map( a => A(31), b => B(31), p => P_31_31_port
                           , g => G_31_31_port);
   PGnetblock_32 : PG_net_1 port map( a => A(32), b => B(32), p => P_32_32_port
                           , g => G_32_32_port);
   GB_low_1_2 : Gblock_0 port map( Pik => P_2_2_port, Gik => G_2_2_port, Gk_1j 
                           => G_1_1_port, Gij => G_2_1_port);
   GB_low_2_4 : Gblock_8 port map( Pik => P_4_3_port, Gik => G_4_3_port, Gk_1j 
                           => G_2_1_port, Gij => Co_0_port);
   GB_low_3_8 : Gblock_7 port map( Pik => P_8_5_port, Gik => G_8_5_port, Gk_1j 
                           => Co_0_port, Gij => Co_1_port);
   GB_high_4_16_0 : Gblock_6 port map( Pik => P_16_9_port, Gik => G_16_9_port, 
                           Gk_1j => Co_1_port, Gij => Co_3_port);
   GB_high_4_16_1 : Gblock_5 port map( Pik => P_12_9_port, Gik => G_12_9_port, 
                           Gk_1j => Co_1_port, Gij => Co_2_port);
   GB_high_5_32_0 : Gblock_4 port map( Pik => P_32_17_port, Gik => G_32_17_port
                           , Gk_1j => Co_3_port, Gij => Co_7_port);
   GB_high_5_32_1 : Gblock_3 port map( Pik => P_28_17_port, Gik => G_28_17_port
                           , Gk_1j => Co_3_port, Gij => Co_6_port);
   GB_high_5_32_2 : Gblock_2 port map( Pik => P_24_17_port, Gik => G_24_17_port
                           , Gk_1j => Co_3_port, Gij => Co_5_port);
   GB_high_5_32_3 : Gblock_1 port map( Pik => P_20_17_port, Gik => G_20_17_port
                           , Gk_1j => Co_3_port, Gij => Co_4_port);
   PGB_low_1_4 : PGblock_0 port map( Pik => P_4_4_port, Gik => G_4_4_port, 
                           Pk_1j => P_3_3_port, Gk_1j => G_3_3_port, Pij => 
                           P_4_3_port, Gij => G_4_3_port);
   PGB_low_1_6 : PGblock_26 port map( Pik => P_6_6_port, Gik => G_6_6_port, 
                           Pk_1j => P_5_5_port, Gk_1j => G_5_5_port, Pij => 
                           P_6_5_port, Gij => G_6_5_port);
   PGB_low_1_8 : PGblock_25 port map( Pik => P_8_8_port, Gik => G_8_8_port, 
                           Pk_1j => P_7_7_port, Gk_1j => G_7_7_port, Pij => 
                           P_8_7_port, Gij => G_8_7_port);
   PGB_low_1_10 : PGblock_24 port map( Pik => P_10_10_port, Gik => G_10_10_port
                           , Pk_1j => P_9_9_port, Gk_1j => G_9_9_port, Pij => 
                           P_10_9_port, Gij => G_10_9_port);
   PGB_low_1_12 : PGblock_23 port map( Pik => P_12_12_port, Gik => G_12_12_port
                           , Pk_1j => P_11_11_port, Gk_1j => G_11_11_port, Pij 
                           => P_12_11_port, Gij => G_12_11_port);
   PGB_low_1_14 : PGblock_22 port map( Pik => P_14_14_port, Gik => G_14_14_port
                           , Pk_1j => P_13_13_port, Gk_1j => G_13_13_port, Pij 
                           => P_14_13_port, Gij => G_14_13_port);
   PGB_low_1_16 : PGblock_21 port map( Pik => P_16_16_port, Gik => G_16_16_port
                           , Pk_1j => P_15_15_port, Gk_1j => G_15_15_port, Pij 
                           => P_16_15_port, Gij => G_16_15_port);
   PGB_low_1_18 : PGblock_20 port map( Pik => P_18_18_port, Gik => G_18_18_port
                           , Pk_1j => P_17_17_port, Gk_1j => G_17_17_port, Pij 
                           => P_18_17_port, Gij => G_18_17_port);
   PGB_low_1_20 : PGblock_19 port map( Pik => P_20_20_port, Gik => G_20_20_port
                           , Pk_1j => P_19_19_port, Gk_1j => G_19_19_port, Pij 
                           => P_20_19_port, Gij => G_20_19_port);
   PGB_low_1_22 : PGblock_18 port map( Pik => P_22_22_port, Gik => G_22_22_port
                           , Pk_1j => P_21_21_port, Gk_1j => G_21_21_port, Pij 
                           => P_22_21_port, Gij => G_22_21_port);
   PGB_low_1_24 : PGblock_17 port map( Pik => P_24_24_port, Gik => G_24_24_port
                           , Pk_1j => P_23_23_port, Gk_1j => G_23_23_port, Pij 
                           => P_24_23_port, Gij => G_24_23_port);
   PGB_low_1_26 : PGblock_16 port map( Pik => P_26_26_port, Gik => G_26_26_port
                           , Pk_1j => P_25_25_port, Gk_1j => G_25_25_port, Pij 
                           => P_26_25_port, Gij => G_26_25_port);
   PGB_low_1_28 : PGblock_15 port map( Pik => P_28_28_port, Gik => G_28_28_port
                           , Pk_1j => P_27_27_port, Gk_1j => G_27_27_port, Pij 
                           => P_28_27_port, Gij => G_28_27_port);
   PGB_low_1_30 : PGblock_14 port map( Pik => P_30_30_port, Gik => G_30_30_port
                           , Pk_1j => P_29_29_port, Gk_1j => G_29_29_port, Pij 
                           => P_30_29_port, Gij => G_30_29_port);
   PGB_low_1_32 : PGblock_13 port map( Pik => P_32_32_port, Gik => G_32_32_port
                           , Pk_1j => P_31_31_port, Gk_1j => G_31_31_port, Pij 
                           => P_32_31_port, Gij => G_32_31_port);
   PGB_low_2_8 : PGblock_12 port map( Pik => P_8_7_port, Gik => G_8_7_port, 
                           Pk_1j => P_6_5_port, Gk_1j => G_6_5_port, Pij => 
                           P_8_5_port, Gij => G_8_5_port);
   PGB_low_2_12 : PGblock_11 port map( Pik => P_12_11_port, Gik => G_12_11_port
                           , Pk_1j => P_10_9_port, Gk_1j => G_10_9_port, Pij =>
                           P_12_9_port, Gij => G_12_9_port);
   PGB_low_2_16 : PGblock_10 port map( Pik => P_16_15_port, Gik => G_16_15_port
                           , Pk_1j => P_14_13_port, Gk_1j => G_14_13_port, Pij 
                           => P_16_13_port, Gij => G_16_13_port);
   PGB_low_2_20 : PGblock_9 port map( Pik => P_20_19_port, Gik => G_20_19_port,
                           Pk_1j => P_18_17_port, Gk_1j => G_18_17_port, Pij =>
                           P_20_17_port, Gij => G_20_17_port);
   PGB_low_2_24 : PGblock_8 port map( Pik => P_24_23_port, Gik => G_24_23_port,
                           Pk_1j => P_22_21_port, Gk_1j => G_22_21_port, Pij =>
                           P_24_21_port, Gij => G_24_21_port);
   PGB_low_2_28 : PGblock_7 port map( Pik => P_28_27_port, Gik => G_28_27_port,
                           Pk_1j => P_26_25_port, Gk_1j => G_26_25_port, Pij =>
                           P_28_25_port, Gij => G_28_25_port);
   PGB_low_2_32 : PGblock_6 port map( Pik => P_32_31_port, Gik => G_32_31_port,
                           Pk_1j => P_30_29_port, Gk_1j => G_30_29_port, Pij =>
                           P_32_29_port, Gij => G_32_29_port);
   PGB_low_3_16 : PGblock_5 port map( Pik => P_16_13_port, Gik => G_16_13_port,
                           Pk_1j => P_12_9_port, Gk_1j => G_12_9_port, Pij => 
                           P_16_9_port, Gij => G_16_9_port);
   PGB_low_3_24 : PGblock_4 port map( Pik => P_24_21_port, Gik => G_24_21_port,
                           Pk_1j => P_20_17_port, Gk_1j => G_20_17_port, Pij =>
                           P_24_17_port, Gij => G_24_17_port);
   PGB_low_3_32 : PGblock_3 port map( Pik => P_32_29_port, Gik => G_32_29_port,
                           Pk_1j => P_28_25_port, Gk_1j => G_28_25_port, Pij =>
                           P_32_25_port, Gij => G_32_25_port);
   PGB_high_4_32_0 : PGblock_2 port map( Pik => P_32_25_port, Gik => 
                           G_32_25_port, Pk_1j => P_24_17_port, Gk_1j => 
                           G_24_17_port, Pij => P_32_17_port, Gij => 
                           G_32_17_port);
   PGB_high_4_32_1 : PGblock_1 port map( Pik => P_28_25_port, Gik => 
                           G_28_25_port, Pk_1j => P_24_17_port, Gk_1j => 
                           G_24_17_port, Pij => P_28_17_port, Gij => 
                           G_28_17_port);
   U1 : INV_X1 port map( A => A(1), ZN => n1);
   U2 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => G_1_1_port);
   U3 : OAI21_X1 port map( B1 => A(1), B2 => B(1), A => Cin, ZN => n3);
   U4 : INV_X1 port map( A => B(1), ZN => n2);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity P4Adder_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (31 downto 0);  Cout : out std_logic);

end P4Adder_NBIT32;

architecture SYN_struct of P4Adder_NBIT32 is

   component SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component carry_generator_NBIT32_NBIT_PER_BLOCK4
      port( A, B : in std_logic_vector (32 downto 1);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal Csum_7_port, Csum_6_port, Csum_5_port, Csum_4_port, Csum_3_port, 
      Csum_2_port, Csum_1_port : std_logic;

begin
   
   Carrygen0 : carry_generator_NBIT32_NBIT_PER_BLOCK4 port map( A(32) => A(31),
                           A(31) => A(30), A(30) => A(29), A(29) => A(28), 
                           A(28) => A(27), A(27) => A(26), A(26) => A(25), 
                           A(25) => A(24), A(24) => A(23), A(23) => A(22), 
                           A(22) => A(21), A(21) => A(20), A(20) => A(19), 
                           A(19) => A(18), A(18) => A(17), A(17) => A(16), 
                           A(16) => A(15), A(15) => A(14), A(14) => A(13), 
                           A(13) => A(12), A(12) => A(11), A(11) => A(10), 
                           A(10) => A(9), A(9) => A(8), A(8) => A(7), A(7) => 
                           A(6), A(6) => A(5), A(5) => A(4), A(4) => A(3), A(3)
                           => A(2), A(2) => A(1), A(1) => A(0), B(32) => B(31),
                           B(31) => B(30), B(30) => B(29), B(29) => B(28), 
                           B(28) => B(27), B(27) => B(26), B(26) => B(25), 
                           B(25) => B(24), B(24) => B(23), B(23) => B(22), 
                           B(22) => B(21), B(21) => B(20), B(20) => B(19), 
                           B(19) => B(18), B(18) => B(17), B(17) => B(16), 
                           B(16) => B(15), B(15) => B(14), B(14) => B(13), 
                           B(13) => B(12), B(12) => B(11), B(11) => B(10), 
                           B(10) => B(9), B(9) => B(8), B(8) => B(7), B(7) => 
                           B(6), B(6) => B(5), B(5) => B(4), B(4) => B(3), B(3)
                           => B(2), B(2) => B(1), B(1) => B(0), Cin => Cin, 
                           Co(7) => Cout, Co(6) => Csum_7_port, Co(5) => 
                           Csum_6_port, Co(4) => Csum_5_port, Co(3) => 
                           Csum_4_port, Co(2) => Csum_3_port, Co(1) => 
                           Csum_2_port, Co(0) => Csum_1_port);
   Sumgen0 : SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), Ci(7) => 
                           Csum_7_port, Ci(6) => Csum_6_port, Ci(5) => 
                           Csum_5_port, Ci(4) => Csum_4_port, Ci(3) => 
                           Csum_3_port, Ci(2) => Csum_2_port, Ci(1) => 
                           Csum_1_port, Ci(0) => Cin, S(31) => S(31), S(30) => 
                           S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           S(21), S(20) => S(20), S(19) => S(19), S(18) => 
                           S(18), S(17) => S(17), S(16) => S(16), S(15) => 
                           S(15), S(14) => S(14), S(13) => S(13), S(12) => 
                           S(12), S(11) => S(11), S(10) => S(10), S(9) => S(9),
                           S(8) => S(8), S(7) => S(7), S(6) => S(6), S(5) => 
                           S(5), S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1)
                           => S(1), S(0) => S(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity shifter_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  LOGIC_ARITH, LEFT_RIGHT : 
         in std_logic;  RES : out std_logic_vector (31 downto 0));

end shifter_NBIT32;

architecture SYN_bhv of shifter_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X4
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X2
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, 
      n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
      n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, 
      n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, 
      n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n1, n2, n3, n4, n5, n6, 
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n266, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648 : std_logic;

begin
   
   U264 : AOI21_X2 port map( B1 => A(31), B2 => B(18), A => n483, ZN => n282);
   U267 : OAI21_X2 port map( B1 => n612, B2 => n628, A => n486, ZN => n285);
   U269 : AOI21_X2 port map( B1 => A(31), B2 => n38, A => n487, ZN => n288);
   U388 : AOI221_X2 port map( B1 => n30, B2 => A(18), C1 => n21, C2 => A(17), A
                           => n568, ZN => n196);
   U428 : NOR2_X2 port map( A1 => n638, A2 => n38, ZN => n165);
   U461 : NOR2_X2 port map( A1 => n642, A2 => n38, ZN => n199);
   U637 : NAND3_X1 port map( A1 => n227, A2 => n646, A3 => n228, ZN => n226);
   U638 : NAND3_X1 port map( A1 => n227, A2 => n646, A3 => B(4), ZN => n428);
   U639 : NAND3_X1 port map( A1 => n445, A2 => n199, A3 => LEFT_RIGHT, ZN => 
                           n240);
   U641 : NAND3_X1 port map( A1 => n489, A2 => n628, A3 => n579, ZN => n255);
   U642 : NAND3_X1 port map( A1 => n7, A2 => n199, A3 => n445, ZN => n138);
   U2 : NOR4_X1 port map( A1 => B(20), A2 => B(21), A3 => B(19), A4 => n594, ZN
                           => n484);
   U3 : NOR2_X2 port map( A1 => n639, A2 => B(3), ZN => n262);
   U4 : AOI221_X1 port map( B1 => n29, B2 => A(6), C1 => n19, C2 => A(7), A => 
                           n525, ZN => n363);
   U5 : AOI221_X1 port map( B1 => n30, B2 => A(7), C1 => n20, C2 => A(8), A => 
                           n570, ZN => n405);
   U6 : AOI221_X1 port map( B1 => n29, B2 => A(8), C1 => n21, C2 => A(9), A => 
                           n552, ZN => n387);
   U7 : OAI21_X2 port map( B1 => n266, B2 => n632, A => n481, ZN => n279);
   U8 : AOI222_X1 port map( A1 => n11, A2 => A(1), B1 => A(0), B2 => n18, C1 =>
                           n7, C2 => A(2), ZN => n293);
   U9 : INV_X1 port map( A => n167, ZN => n635);
   U10 : NOR2_X1 port map( A1 => n636, A2 => B(4), ZN => n167);
   U11 : INV_X1 port map( A => n169, ZN => n644);
   U12 : INV_X1 port map( A => n165, ZN => n637);
   U13 : INV_X1 port map( A => n199, ZN => n641);
   U14 : INV_X1 port map( A => n28, ZN => n26);
   U15 : INV_X1 port map( A => n31, ZN => n24);
   U16 : INV_X1 port map( A => n31, ZN => n25);
   U17 : INV_X1 port map( A => n21, ZN => n14);
   U18 : INV_X1 port map( A => n19, ZN => n16);
   U19 : INV_X1 port map( A => n19, ZN => n15);
   U20 : INV_X1 port map( A => n505, ZN => n643);
   U21 : INV_X1 port map( A => n29, ZN => n27);
   U22 : INV_X1 port map( A => n493, ZN => n640);
   U23 : NOR2_X1 port map( A1 => n645, A2 => n38, ZN => n169);
   U24 : NAND2_X1 port map( A1 => n488, A2 => n454, ZN => n161);
   U25 : INV_X1 port map( A => n41, ZN => n38);
   U26 : OAI222_X1 port map( A1 => n637, A2 => n70, B1 => n635, B2 => n92, C1 
                           => n644, C2 => n80, ZN => n224);
   U27 : OAI222_X1 port map( A1 => n637, A2 => n67, B1 => n635, B2 => n96, C1 
                           => n644, C2 => n83, ZN => n212);
   U28 : NOR2_X1 port map( A1 => n40, A2 => n642, ZN => n493);
   U29 : OAI22_X1 port map( A1 => n115, A2 => n642, B1 => n126, B2 => n638, ZN 
                           => n383);
   U30 : INV_X1 port map( A => n454, ZN => n636);
   U31 : AOI21_X1 port map( B1 => n134, B2 => n2, A => n519, ZN => n286);
   U32 : AOI21_X1 port map( B1 => n129, B2 => n3, A => n519, ZN => n312);
   U33 : BUF_X1 port map( A => n138, Z => n33);
   U34 : BUF_X1 port map( A => n138, Z => n32);
   U35 : NOR2_X1 port map( A1 => n383, A2 => n359, ZN => n197);
   U36 : NOR2_X1 port map( A1 => n118, A2 => n359, ZN => n181);
   U37 : BUF_X1 port map( A => n138, Z => n34);
   U38 : NAND2_X1 port map( A1 => n488, A2 => n5, ZN => n505);
   U39 : INV_X1 port map( A => n182, ZN => n118);
   U40 : INV_X1 port map( A => n172, ZN => n54);
   U41 : INV_X1 port map( A => n139, ZN => n58);
   U42 : INV_X1 port map( A => n348, ZN => n52);
   U43 : INV_X1 port map( A => n337, ZN => n44);
   U44 : INV_X1 port map( A => n480, ZN => n88);
   U45 : INV_X1 port map( A => n314, ZN => n56);
   U46 : INV_X1 port map( A => n290, ZN => n50);
   U47 : INV_X1 port map( A => n271, ZN => n46);
   U48 : INV_X1 port map( A => n257, ZN => n101);
   U49 : INV_X1 port map( A => n440, ZN => n93);
   U50 : INV_X1 port map( A => n302, ZN => n97);
   U51 : NOR2_X1 port map( A1 => n612, A2 => n148, ZN => n150);
   U52 : NOR2_X1 port map( A1 => n639, A2 => n646, ZN => n454);
   U53 : NAND2_X1 port map( A1 => n484, A2 => n630, ZN => n281);
   U54 : AOI222_X1 port map( A1 => n370, A2 => n262, B1 => n320, B2 => n260, C1
                           => n185, C2 => n3, ZN => n238);
   U55 : INV_X1 port map( A => n356, ZN => n642);
   U56 : AOI222_X1 port map( A1 => n168, A2 => n262, B1 => n355, B2 => n260, C1
                           => n170, C2 => n3, ZN => n471);
   U57 : AOI222_X1 port map( A1 => n402, A2 => n262, B1 => n403, B2 => n260, C1
                           => n464, C2 => n2, ZN => n461);
   U58 : NAND2_X1 port map( A1 => n488, A2 => n262, ZN => n157);
   U59 : NAND2_X1 port map( A1 => n488, A2 => n260, ZN => n158);
   U60 : OAI222_X1 port map( A1 => n374, A2 => n638, B1 => n645, B2 => n375, C1
                           => n376, C2 => n642, ZN => n172);
   U61 : OAI222_X1 port map( A1 => n131, A2 => n638, B1 => n362, B2 => n645, C1
                           => n363, C2 => n642, ZN => n139);
   U62 : OAI222_X1 port map( A1 => n613, A2 => n638, B1 => n293, B2 => n645, C1
                           => n405, C2 => n642, ZN => n348);
   U63 : OAI222_X1 port map( A1 => n615, A2 => n638, B1 => n45, B2 => n645, C1 
                           => n387, C2 => n642, ZN => n337);
   U64 : AOI221_X1 port map( B1 => n129, B2 => n262, C1 => n355, C2 => n2, A =>
                           n359, ZN => n159);
   U65 : AOI221_X1 port map( B1 => n134, B2 => n262, C1 => n403, C2 => n3, A =>
                           n359, ZN => n347);
   U66 : OAI221_X1 port map( B1 => n105, B2 => n638, C1 => n89, C2 => n642, A 
                           => n607, ZN => n480);
   U67 : AOI22_X1 port map( A1 => n454, A2 => n320, B1 => n260, B2 => n370, ZN 
                           => n607);
   U68 : AOI222_X1 port map( A1 => n169, A2 => n185, B1 => n493, B2 => n320, C1
                           => n167, C2 => n370, ZN => n550);
   U69 : AOI222_X1 port map( A1 => n165, A2 => n166, B1 => n167, B2 => n168, C1
                           => n169, C2 => n170, ZN => n164);
   U70 : AOI222_X1 port map( A1 => n165, A2 => n516, B1 => n167, B2 => n402, C1
                           => n169, C2 => n464, ZN => n581);
   U71 : AOI222_X1 port map( A1 => n165, A2 => n184, B1 => n167, B2 => n185, C1
                           => n169, C2 => n186, ZN => n183);
   U72 : AOI222_X1 port map( A1 => n165, A2 => n178, B1 => n167, B2 => n186, C1
                           => n169, C2 => n184, ZN => n239);
   U73 : AOI222_X1 port map( A1 => n169, A2 => n168, B1 => n493, B2 => n128, C1
                           => n167, C2 => n355, ZN => n534);
   U74 : AOI222_X1 port map( A1 => n169, A2 => n402, B1 => n493, B2 => n133, C1
                           => n167, C2 => n403, ZN => n520);
   U75 : AOI222_X1 port map( A1 => n169, A2 => n453, B1 => n493, B2 => n382, C1
                           => n167, C2 => n506, ZN => n507);
   U76 : OAI222_X1 port map( A1 => n637, A2 => n74, B1 => n635, B2 => n100, C1 
                           => n644, C2 => n196, ZN => n200);
   U77 : INV_X1 port map( A => n260, ZN => n645);
   U78 : NOR2_X1 port map( A1 => n647, A2 => B(4), ZN => n488);
   U79 : INV_X1 port map( A => n262, ZN => n638);
   U80 : OAI222_X1 port map( A1 => n132, A2 => n14, B1 => n27, B2 => n614, C1 
                           => n1, C2 => n102, ZN => n602);
   U81 : OAI221_X1 port map( B1 => n363, B2 => n638, C1 => n61, C2 => n642, A 
                           => n522, ZN => n314);
   U82 : AOI22_X1 port map( A1 => n454, A2 => n57, B1 => n260, B2 => n420, ZN 
                           => n522);
   U83 : OAI221_X1 port map( B1 => n405, B2 => n638, C1 => n72, C2 => n642, A 
                           => n509, ZN => n290);
   U84 : AOI22_X1 port map( A1 => n454, A2 => n51, B1 => n260, B2 => n407, ZN 
                           => n509);
   U85 : OAI221_X1 port map( B1 => n387, B2 => n638, C1 => n75, C2 => n642, A 
                           => n496, ZN => n271);
   U86 : AOI22_X1 port map( A1 => n454, A2 => n390, B1 => n260, B2 => n389, ZN 
                           => n496);
   U87 : INV_X1 port map( A => n228, ZN => n625);
   U88 : OAI21_X1 port map( B1 => n612, B2 => n630, A => n486, ZN => n253);
   U89 : AOI221_X1 port map( B1 => n199, B2 => n361, C1 => B(4), C2 => n55, A 
                           => n418, ZN => n409);
   U90 : INV_X1 port map( A => n214, ZN => n55);
   U91 : OAI222_X1 port map( A1 => n61, A2 => n644, B1 => n363, B2 => n635, C1 
                           => n81, C2 => n637, ZN => n418);
   U92 : AOI221_X1 port map( B1 => n199, B2 => n350, C1 => B(4), C2 => n49, A 
                           => n404, ZN => n392);
   U93 : INV_X1 port map( A => n202, ZN => n49);
   U94 : OAI222_X1 port map( A1 => n72, A2 => n644, B1 => n405, B2 => n635, C1 
                           => n84, C2 => n637, ZN => n404);
   U95 : AOI221_X1 port map( B1 => n199, B2 => n339, C1 => B(4), C2 => n47, A 
                           => n386, ZN => n378);
   U96 : INV_X1 port map( A => n188, ZN => n47);
   U97 : OAI222_X1 port map( A1 => n75, A2 => n644, B1 => n387, B2 => n635, C1 
                           => n86, C2 => n637, ZN => n386);
   U98 : AOI221_X1 port map( B1 => n199, B2 => n324, C1 => n38, C2 => n172, A 
                           => n371, ZN => n365);
   U99 : OAI222_X1 port map( A1 => n78, A2 => n644, B1 => n62, B2 => n635, C1 
                           => n90, C2 => n637, ZN => n371);
   U100 : AOI221_X1 port map( B1 => n199, B2 => n313, C1 => n38, C2 => n139, A 
                           => n360, ZN => n352);
   U101 : OAI222_X1 port map( A1 => n81, A2 => n644, B1 => n61, B2 => n635, C1 
                           => n94, C2 => n637, ZN => n360);
   U102 : AOI221_X1 port map( B1 => n199, B2 => n289, C1 => n38, C2 => n348, A 
                           => n349, ZN => n341);
   U103 : OAI222_X1 port map( A1 => n84, A2 => n644, B1 => n72, B2 => n635, C1 
                           => n98, C2 => n637, ZN => n349);
   U104 : AOI221_X1 port map( B1 => n199, B2 => n270, C1 => n38, C2 => n337, A 
                           => n338, ZN => n328);
   U105 : OAI222_X1 port map( A1 => n86, A2 => n644, B1 => n75, B2 => n635, C1 
                           => n103, C2 => n637, ZN => n338);
   U106 : NOR2_X1 port map( A1 => n612, A2 => n646, ZN => n359);
   U107 : AOI221_X1 port map( B1 => n276, B2 => n479, C1 => n627, C2 => n480, A
                           => n279, ZN => n478);
   U108 : OAI21_X1 port map( B1 => n482, B2 => n281, A => n282, ZN => n479);
   U109 : AOI21_X1 port map( B1 => n283, B2 => n485, A => n285, ZN => n482);
   U110 : OAI21_X1 port map( B1 => n88, B2 => n287, A => n288, ZN => n485);
   U111 : AOI221_X1 port map( B1 => n276, B2 => n470, C1 => n627, C2 => n434, A
                           => n279, ZN => n469);
   U112 : OAI21_X1 port map( B1 => n472, B2 => n281, A => n282, ZN => n470);
   U113 : AOI21_X1 port map( B1 => n283, B2 => n473, A => n285, ZN => n472);
   U114 : OAI21_X1 port map( B1 => n93, B2 => n287, A => n288, ZN => n473);
   U115 : AOI221_X1 port map( B1 => n276, B2 => n460, C1 => n627, C2 => n297, A
                           => n279, ZN => n459);
   U116 : OAI21_X1 port map( B1 => n462, B2 => n281, A => n282, ZN => n460);
   U117 : AOI21_X1 port map( B1 => n283, B2 => n463, A => n285, ZN => n462);
   U118 : OAI21_X1 port map( B1 => n97, B2 => n287, A => n288, ZN => n463);
   U119 : AOI221_X1 port map( B1 => n276, B2 => n448, C1 => n627, C2 => n246, A
                           => n279, ZN => n447);
   U120 : OAI21_X1 port map( B1 => n450, B2 => n281, A => n282, ZN => n448);
   U121 : AOI21_X1 port map( B1 => n283, B2 => n451, A => n285, ZN => n450);
   U122 : OAI21_X1 port map( B1 => n101, B2 => n287, A => n288, ZN => n451);
   U123 : AOI221_X1 port map( B1 => n276, B2 => n424, C1 => n627, C2 => n106, A
                           => n279, ZN => n423);
   U124 : INV_X1 port map( A => n238, ZN => n106);
   U125 : OAI21_X1 port map( B1 => n425, B2 => n281, A => n282, ZN => n424);
   U126 : AOI21_X1 port map( B1 => n283, B2 => n426, A => n285, ZN => n425);
   U127 : AOI221_X1 port map( B1 => n276, B2 => n411, C1 => n627, C2 => n223, A
                           => n279, ZN => n410);
   U128 : OAI21_X1 port map( B1 => n414, B2 => n281, A => n282, ZN => n411);
   U129 : AOI21_X1 port map( B1 => n283, B2 => n415, A => n285, ZN => n414);
   U130 : OAI21_X1 port map( B1 => n109, B2 => n287, A => n288, ZN => n415);
   U131 : AOI221_X1 port map( B1 => n276, B2 => n394, C1 => n627, C2 => n211, A
                           => n279, ZN => n393);
   U132 : OAI21_X1 port map( B1 => n397, B2 => n281, A => n282, ZN => n394);
   U133 : AOI21_X1 port map( B1 => n283, B2 => n398, A => n285, ZN => n397);
   U134 : OAI21_X1 port map( B1 => n112, B2 => n287, A => n288, ZN => n398);
   U135 : AOI221_X1 port map( B1 => n276, B2 => n380, C1 => n627, C2 => n114, A
                           => n279, ZN => n379);
   U136 : OAI21_X1 port map( B1 => n384, B2 => n281, A => n282, ZN => n380);
   U137 : AOI21_X1 port map( B1 => n283, B2 => n385, A => n285, ZN => n384);
   U138 : OAI21_X1 port map( B1 => n197, B2 => n287, A => n288, ZN => n385);
   U139 : AOI221_X1 port map( B1 => n276, B2 => n367, C1 => n627, C2 => n118, A
                           => n279, ZN => n366);
   U140 : OAI21_X1 port map( B1 => n368, B2 => n281, A => n282, ZN => n367);
   U141 : AOI21_X1 port map( B1 => n283, B2 => n369, A => n285, ZN => n368);
   U142 : OAI21_X1 port map( B1 => n181, B2 => n287, A => n288, ZN => n369);
   U143 : AOI221_X1 port map( B1 => n276, B2 => n354, C1 => n627, C2 => n121, A
                           => n279, ZN => n353);
   U144 : INV_X1 port map( A => n163, ZN => n121);
   U145 : OAI21_X1 port map( B1 => n357, B2 => n281, A => n282, ZN => n354);
   U146 : AOI21_X1 port map( B1 => n283, B2 => n358, A => n285, ZN => n357);
   U147 : AOI221_X1 port map( B1 => n276, B2 => n343, C1 => n627, C2 => n124, A
                           => n279, ZN => n342);
   U148 : INV_X1 port map( A => n344, ZN => n124);
   U149 : OAI21_X1 port map( B1 => n345, B2 => n281, A => n282, ZN => n343);
   U150 : AOI21_X1 port map( B1 => n283, B2 => n346, A => n285, ZN => n345);
   U151 : NOR2_X1 port map( A1 => n612, A2 => n2, ZN => n519);
   U152 : AOI221_X1 port map( B1 => n165, B2 => n429, C1 => n199, C2 => n373, A
                           => n492, ZN => n477);
   U153 : OAI222_X1 port map( A1 => n374, A2 => n635, B1 => n375, B2 => n640, 
                           C1 => n376, C2 => n644, ZN => n492);
   U154 : AOI221_X1 port map( B1 => n165, B2 => n474, C1 => n199, C2 => n419, A
                           => n475, ZN => n468);
   U155 : OAI222_X1 port map( A1 => n131, A2 => n635, B1 => n362, B2 => n640, 
                           C1 => n363, C2 => n644, ZN => n475);
   U156 : AOI221_X1 port map( B1 => n165, B2 => n465, C1 => n199, C2 => n406, A
                           => n466, ZN => n458);
   U157 : OAI222_X1 port map( A1 => n613, A2 => n635, B1 => n293, B2 => n640, 
                           C1 => n405, C2 => n644, ZN => n466);
   U158 : AOI221_X1 port map( B1 => n165, B2 => n455, C1 => n199, C2 => n388, A
                           => n456, ZN => n446);
   U159 : OAI222_X1 port map( A1 => n615, A2 => n635, B1 => n45, B2 => n640, C1
                           => n387, C2 => n644, ZN => n456);
   U160 : AOI221_X1 port map( B1 => n165, B2 => n373, C1 => n199, C2 => n372, A
                           => n427, ZN => n422);
   U161 : OAI221_X1 port map( B1 => n376, B2 => n635, C1 => n62, C2 => n644, A 
                           => n428, ZN => n427);
   U162 : OAI22_X1 port map( A1 => n8, A2 => n130, B1 => n1, B2 => n135, ZN => 
                           n533);
   U163 : NOR2_X1 port map( A1 => n612, A2 => n8, ZN => n382);
   U164 : OAI221_X1 port map( B1 => n109, B2 => n160, C1 => n92, C2 => n161, A 
                           => n162, ZN => n220);
   U165 : OAI221_X1 port map( B1 => n112, B2 => n160, C1 => n96, C2 => n161, A 
                           => n162, ZN => n208);
   U166 : OAI221_X1 port map( B1 => n197, B2 => n160, C1 => n100, C2 => n161, A
                           => n162, ZN => n194);
   U167 : AOI22_X1 port map( A1 => n480, A2 => n38, B1 => n42, B2 => n63, ZN =>
                           n587);
   U168 : INV_X1 port map( A => n601, ZN => n63);
   U169 : AOI221_X1 port map( B1 => n4, B2 => n602, C1 => n454, C2 => n184, A 
                           => n603, ZN => n601);
   U170 : OAI22_X1 port map( A1 => n617, A2 => n638, B1 => n64, B2 => n645, ZN 
                           => n603);
   U171 : AOI22_X1 port map( A1 => n420, A2 => n2, B1 => n57, B2 => n262, ZN =>
                           n214);
   U172 : AOI22_X1 port map( A1 => n407, A2 => n5, B1 => n51, B2 => n262, ZN =>
                           n202);
   U173 : AOI22_X1 port map( A1 => n389, A2 => n3, B1 => n390, B2 => n262, ZN 
                           => n188);
   U174 : AOI22_X1 port map( A1 => n452, A2 => n4, B1 => n453, B2 => n262, ZN 
                           => n449);
   U175 : AOI22_X1 port map( A1 => n168, A2 => n3, B1 => n355, B2 => n262, ZN 
                           => n413);
   U176 : AOI22_X1 port map( A1 => n402, A2 => n5, B1 => n403, B2 => n262, ZN 
                           => n396);
   U177 : AOI22_X1 port map( A1 => n370, A2 => n4, B1 => n320, B2 => n262, ZN 
                           => n182);
   U178 : AOI22_X1 port map( A1 => n355, A2 => n2, B1 => n128, B2 => n262, ZN 
                           => n163);
   U179 : AOI22_X1 port map( A1 => n403, A2 => n4, B1 => n133, B2 => n262, ZN 
                           => n344);
   U180 : AOI21_X1 port map( B1 => n148, B2 => n217, A => n150, ZN => n216);
   U181 : OAI21_X1 port map( B1 => n218, B2 => n152, A => n153, ZN => n217);
   U182 : AOI211_X1 port map( C1 => n643, C2 => n219, A => n220, B => n221, ZN 
                           => n218);
   U183 : OAI22_X1 port map( A1 => n70, A2 => n157, B1 => n80, B2 => n158, ZN 
                           => n221);
   U184 : AOI21_X1 port map( B1 => n148, B2 => n205, A => n150, ZN => n204);
   U185 : OAI21_X1 port map( B1 => n206, B2 => n152, A => n153, ZN => n205);
   U186 : AOI211_X1 port map( C1 => n643, C2 => n207, A => n208, B => n209, ZN 
                           => n206);
   U187 : OAI22_X1 port map( A1 => n67, A2 => n157, B1 => n83, B2 => n158, ZN 
                           => n209);
   U188 : AOI21_X1 port map( B1 => n148, B2 => n191, A => n150, ZN => n190);
   U189 : OAI21_X1 port map( B1 => n192, B2 => n152, A => n153, ZN => n191);
   U190 : AOI211_X1 port map( C1 => n643, C2 => n193, A => n194, B => n195, ZN 
                           => n192);
   U191 : OAI22_X1 port map( A1 => n74, A2 => n157, B1 => n196, B2 => n158, ZN 
                           => n195);
   U192 : OAI211_X1 port map( C1 => n126, C2 => n645, A => n401, B => n449, ZN 
                           => n257);
   U193 : AOI21_X1 port map( B1 => n320, B2 => n4, A => n519, ZN => n323);
   U194 : AOI21_X1 port map( B1 => n506, B2 => n5, A => n519, ZN => n336);
   U195 : NAND2_X1 port map( A1 => n484, A2 => n632, ZN => n249);
   U196 : OAI21_X1 port map( B1 => n417, B2 => n636, A => n471, ZN => n440);
   U197 : OAI21_X1 port map( B1 => n400, B2 => n636, A => n461, ZN => n302);
   U198 : OAI21_X1 port map( B1 => n412, B2 => n636, A => n471, ZN => n434);
   U199 : OAI21_X1 port map( B1 => n395, B2 => n636, A => n461, ZN => n297);
   U200 : OAI21_X1 port map( B1 => n412, B2 => n645, A => n413, ZN => n223);
   U201 : OAI21_X1 port map( B1 => n395, B2 => n645, A => n396, ZN => n211);
   U202 : OAI21_X1 port map( B1 => n333, B2 => n646, A => n449, ZN => n246);
   U203 : NOR2_X1 port map( A1 => n612, A2 => n484, ZN => n483);
   U204 : OAI21_X1 port map( B1 => n237, B2 => n287, A => n288, ZN => n426);
   U205 : OAI21_X1 port map( B1 => n159, B2 => n287, A => n288, ZN => n358);
   U206 : OAI21_X1 port map( B1 => n347, B2 => n287, A => n288, ZN => n346);
   U207 : OAI21_X1 port map( B1 => n336, B2 => n287, A => n288, ZN => n335);
   U208 : BUF_X1 port map( A => n137, Z => n35);
   U209 : BUF_X1 port map( A => n137, Z => n36);
   U210 : OAI21_X1 port map( B1 => n233, B2 => n152, A => n153, ZN => n232);
   U211 : AOI211_X1 port map( C1 => n643, C2 => n234, A => n235, B => n236, ZN 
                           => n233);
   U212 : OAI22_X1 port map( A1 => n64, A2 => n157, B1 => n77, B2 => n158, ZN 
                           => n236);
   U213 : OAI221_X1 port map( B1 => n237, B2 => n160, C1 => n89, C2 => n161, A 
                           => n162, ZN => n235);
   U214 : OAI21_X1 port map( B1 => n177, B2 => n152, A => n153, ZN => n176);
   U215 : AOI211_X1 port map( C1 => n643, C2 => n178, A => n179, B => n180, ZN 
                           => n177);
   U216 : OAI22_X1 port map( A1 => n77, A2 => n157, B1 => n89, B2 => n158, ZN 
                           => n180);
   U217 : OAI221_X1 port map( B1 => n181, B2 => n160, C1 => n105, C2 => n161, A
                           => n162, ZN => n179);
   U218 : OAI21_X1 port map( B1 => n151, B2 => n152, A => n153, ZN => n149);
   U219 : AOI211_X1 port map( C1 => n643, C2 => n154, A => n155, B => n156, ZN 
                           => n151);
   U220 : OAI22_X1 port map( A1 => n80, A2 => n157, B1 => n92, B2 => n158, ZN 
                           => n156);
   U221 : OAI221_X1 port map( B1 => n159, B2 => n160, C1 => n108, C2 => n161, A
                           => n162, ZN => n155);
   U222 : OAI21_X1 port map( B1 => n576, B2 => n152, A => n153, ZN => n575);
   U223 : AOI211_X1 port map( C1 => n643, C2 => n305, A => n577, B => n578, ZN 
                           => n576);
   U224 : OAI22_X1 port map( A1 => n83, A2 => n157, B1 => n96, B2 => n158, ZN 
                           => n578);
   U225 : OAI221_X1 port map( B1 => n347, B2 => n160, C1 => n111, C2 => n161, A
                           => n162, ZN => n577);
   U226 : OAI21_X1 port map( B1 => n559, B2 => n152, A => n153, ZN => n558);
   U227 : AOI211_X1 port map( C1 => n643, C2 => n261, A => n560, B => n561, ZN 
                           => n559);
   U228 : OAI22_X1 port map( A1 => n196, A2 => n157, B1 => n100, B2 => n158, ZN
                           => n561);
   U229 : OAI221_X1 port map( B1 => n336, B2 => n160, C1 => n115, C2 => n161, A
                           => n162, ZN => n560);
   U230 : OAI21_X1 port map( B1 => n547, B2 => n152, A => n153, ZN => n546);
   U231 : AOI211_X1 port map( C1 => n643, C2 => n184, A => n548, B => n549, ZN 
                           => n547);
   U232 : OAI22_X1 port map( A1 => n89, A2 => n157, B1 => n105, B2 => n158, ZN 
                           => n549);
   U233 : OAI221_X1 port map( B1 => n323, B2 => n160, C1 => n117, C2 => n161, A
                           => n162, ZN => n548);
   U234 : OAI21_X1 port map( B1 => n530, B2 => n152, A => n153, ZN => n529);
   U235 : AOI211_X1 port map( C1 => n643, C2 => n166, A => n531, B => n532, ZN 
                           => n530);
   U236 : OAI22_X1 port map( A1 => n92, A2 => n157, B1 => n108, B2 => n158, ZN 
                           => n532);
   U237 : OAI221_X1 port map( B1 => n312, B2 => n160, C1 => n120, C2 => n161, A
                           => n162, ZN => n531);
   U238 : OAI21_X1 port map( B1 => n515, B2 => n152, A => n153, ZN => n514);
   U239 : AOI211_X1 port map( C1 => n643, C2 => n516, A => n517, B => n518, ZN 
                           => n515);
   U240 : OAI22_X1 port map( A1 => n96, A2 => n157, B1 => n111, B2 => n158, ZN 
                           => n518);
   U241 : OAI221_X1 port map( B1 => n286, B2 => n160, C1 => n123, C2 => n161, A
                           => n162, ZN => n517);
   U242 : INV_X1 port map( A => n452, ZN => n100);
   U243 : INV_X1 port map( A => n170, ZN => n92);
   U244 : INV_X1 port map( A => n464, ZN => n96);
   U245 : INV_X1 port map( A => n186, ZN => n89);
   U246 : INV_X1 port map( A => n166, ZN => n80);
   U247 : INV_X1 port map( A => n516, ZN => n83);
   U248 : NOR2_X1 port map( A1 => n135, A2 => n8, ZN => n580);
   U249 : OAI21_X1 port map( B1 => n587, B2 => n255, A => n256, ZN => n595);
   U250 : AOI21_X1 port map( B1 => n251, B2 => n438, A => n253, ZN => n437);
   U251 : OAI21_X1 port map( B1 => n439, B2 => n255, A => n256, ZN => n438);
   U252 : AOI22_X1 port map( A1 => n435, A2 => n39, B1 => B(4), B2 => n440, ZN 
                           => n439);
   U253 : AOI21_X1 port map( B1 => n251, B2 => n300, A => n253, ZN => n299);
   U254 : OAI21_X1 port map( B1 => n301, B2 => n255, A => n256, ZN => n300);
   U255 : AOI22_X1 port map( A1 => n298, A2 => n39, B1 => B(4), B2 => n302, ZN 
                           => n301);
   U256 : AOI21_X1 port map( B1 => n251, B2 => n252, A => n253, ZN => n248);
   U257 : OAI21_X1 port map( B1 => n254, B2 => n255, A => n256, ZN => n252);
   U258 : AOI22_X1 port map( A1 => n247, A2 => n39, B1 => B(4), B2 => n257, ZN 
                           => n254);
   U259 : BUF_X1 port map( A => n356, Z => n2);
   U260 : BUF_X1 port map( A => n356, Z => n3);
   U261 : INV_X1 port map( A => n293, ZN => n51);
   U262 : INV_X1 port map( A => n184, ZN => n77);
   U263 : INV_X1 port map( A => n506, ZN => n126);
   U265 : INV_X1 port map( A => n185, ZN => n105);
   U266 : INV_X1 port map( A => n390, ZN => n45);
   U268 : BUF_X1 port map( A => n356, Z => n4);
   U270 : BUF_X1 port map( A => n356, Z => n5);
   U271 : INV_X1 port map( A => n453, ZN => n115);
   U272 : INV_X1 port map( A => n412, ZN => n128);
   U273 : INV_X1 port map( A => n395, ZN => n133);
   U274 : INV_X1 port map( A => n154, ZN => n70);
   U275 : INV_X1 port map( A => n305, ZN => n67);
   U276 : INV_X1 port map( A => n178, ZN => n64);
   U277 : INV_X1 port map( A => n168, ZN => n108);
   U278 : INV_X1 port map( A => n402, ZN => n111);
   U279 : INV_X1 port map( A => n261, ZN => n74);
   U280 : INV_X1 port map( A => n419, ZN => n81);
   U281 : INV_X1 port map( A => n406, ZN => n84);
   U282 : INV_X1 port map( A => n388, ZN => n86);
   U283 : BUF_X1 port map( A => n43, Z => n41);
   U284 : INV_X1 port map( A => n362, ZN => n57);
   U285 : INV_X1 port map( A => n474, ZN => n61);
   U286 : INV_X1 port map( A => n465, ZN => n72);
   U287 : INV_X1 port map( A => n455, ZN => n75);
   U288 : INV_X1 port map( A => n267, ZN => n8);
   U289 : INV_X1 port map( A => n355, ZN => n120);
   U290 : INV_X1 port map( A => n403, ZN => n123);
   U291 : BUF_X1 port map( A => n43, Z => n42);
   U292 : BUF_X1 port map( A => n43, Z => n39);
   U293 : BUF_X1 port map( A => n43, Z => n40);
   U294 : INV_X1 port map( A => n370, ZN => n117);
   U295 : INV_X1 port map( A => n373, ZN => n78);
   U296 : INV_X1 port map( A => n420, ZN => n131);
   U297 : INV_X1 port map( A => n407, ZN => n613);
   U298 : INV_X1 port map( A => n389, ZN => n615);
   U299 : INV_X1 port map( A => n417, ZN => n129);
   U300 : INV_X1 port map( A => n400, ZN => n134);
   U301 : INV_X1 port map( A => n429, ZN => n62);
   U302 : INV_X1 port map( A => n372, ZN => n90);
   U303 : INV_X1 port map( A => n361, ZN => n94);
   U304 : INV_X1 port map( A => n350, ZN => n98);
   U305 : INV_X1 port map( A => n339, ZN => n103);
   U306 : AND2_X1 port map( A1 => n238, A2 => n401, ZN => n237);
   U307 : INV_X1 port map( A => n234, ZN => n617);
   U308 : INV_X1 port map( A => n416, ZN => n109);
   U309 : OAI211_X1 port map( C1 => n417, C2 => n645, A => n401, B => n413, ZN 
                           => n416);
   U310 : INV_X1 port map( A => n399, ZN => n112);
   U311 : OAI211_X1 port map( C1 => n400, C2 => n645, A => n401, B => n396, ZN 
                           => n399);
   U312 : INV_X1 port map( A => n381, ZN => n114);
   U313 : AOI21_X1 port map( B1 => n260, B2 => n382, A => n383, ZN => n381);
   U314 : BUF_X1 port map( A => n137, Z => n37);
   U315 : OR4_X1 port map( A1 => B(21), A2 => B(20), A3 => B(19), A4 => B(18), 
                           ZN => n598);
   U316 : OAI22_X1 port map( A1 => n87, A2 => n1, B1 => n85, B2 => n8, ZN => 
                           n568);
   U317 : OAI22_X1 port map( A1 => n622, A2 => n1, B1 => n623, B2 => n8, ZN => 
                           n525);
   U318 : OAI22_X1 port map( A1 => n623, A2 => n1, B1 => n65, B2 => n8, ZN => 
                           n570);
   U319 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n73, B2 => n8, ZN => 
                           n552);
   U320 : AOI221_X1 port map( B1 => n31, B2 => A(5), C1 => n20, C2 => A(6), A 
                           => n541, ZN => n376);
   U321 : OAI22_X1 port map( A1 => n621, A2 => n1, B1 => n622, B2 => n8, ZN => 
                           n541);
   U322 : OAI221_X1 port map( B1 => n27, B2 => n612, C1 => n17, C2 => n135, A 
                           => n609, ZN => n320);
   U323 : AOI22_X1 port map( A1 => A(29), A2 => n10, B1 => A(28), B2 => n7, ZN 
                           => n609);
   U324 : OAI221_X1 port map( B1 => n25, B2 => n127, C1 => n15, C2 => n125, A 
                           => n535, ZN => n355);
   U325 : AOI22_X1 port map( A1 => A(26), A2 => n9, B1 => A(25), B2 => n267, ZN
                           => n535);
   U326 : OAI221_X1 port map( B1 => n26, B2 => n130, C1 => n16, C2 => n127, A 
                           => n585, ZN => n403);
   U327 : AOI22_X1 port map( A1 => A(27), A2 => n10, B1 => A(26), B2 => n7, ZN 
                           => n585);
   U328 : OR3_X1 port map( A1 => B(22), A2 => B(24), A3 => B(23), ZN => n594);
   U329 : NAND3_X1 port map( A1 => n489, A2 => n628, A3 => n600, ZN => n152);
   U330 : NOR3_X1 port map( A1 => B(12), A2 => B(14), A3 => B(13), ZN => n600);
   U331 : NAND3_X1 port map( A1 => n592, A2 => n631, A3 => n599, ZN => n146);
   U332 : INV_X1 port map( A => B(22), ZN => n631);
   U333 : NOR3_X1 port map( A1 => B(23), A2 => B(25), A3 => B(24), ZN => n599);
   U334 : OAI221_X1 port map( B1 => n27, B2 => n85, C1 => n17, C2 => n82, A => 
                           n606, ZN => n184);
   U335 : AOI22_X1 port map( A1 => A(13), A2 => n11, B1 => A(12), B2 => n7, ZN 
                           => n606);
   U336 : OAI221_X1 port map( B1 => n27, B2 => n125, C1 => n17, C2 => n122, A 
                           => n608, ZN => n370);
   U337 : AOI22_X1 port map( A1 => A(25), A2 => n9, B1 => A(24), B2 => n7, ZN 
                           => n608);
   U338 : NAND2_X1 port map( A1 => n488, A2 => n489, ZN => n287);
   U339 : OAI221_X1 port map( B1 => n25, B2 => n116, C1 => n15, C2 => n113, A 
                           => n536, ZN => n168);
   U340 : AOI22_X1 port map( A1 => A(22), A2 => n9, B1 => A(21), B2 => n267, ZN
                           => n536);
   U341 : OAI221_X1 port map( B1 => n26, B2 => n119, C1 => n16, C2 => n116, A 
                           => n583, ZN => n402);
   U342 : AOI22_X1 port map( A1 => A(23), A2 => n10, B1 => A(22), B2 => n7, ZN 
                           => n583);
   U343 : NOR2_X2 port map( A1 => n490, A2 => B(11), ZN => n283);
   U344 : NAND2_X1 port map( A1 => A(31), A2 => n647, ZN => n162);
   U345 : AOI221_X1 port map( B1 => A(1), B2 => n31, C1 => A(2), C2 => n21, A 
                           => n540, ZN => n374);
   U346 : OAI22_X1 port map( A1 => n614, A2 => n1, B1 => n616, B2 => n8, ZN => 
                           n540);
   U347 : NOR2_X2 port map( A1 => n266, A2 => n591, ZN => n144);
   U348 : NAND2_X1 port map( A1 => A(31), A2 => n152, ZN => n153);
   U349 : NAND2_X1 port map( A1 => A(31), A2 => n146, ZN => n147);
   U350 : OAI221_X1 port map( B1 => n26, B2 => n135, C1 => n16, C2 => n130, A 
                           => n564, ZN => n506);
   U351 : AOI22_X1 port map( A1 => A(28), A2 => n10, B1 => A(27), B2 => n6, ZN 
                           => n564);
   U352 : OAI221_X1 port map( B1 => n26, B2 => n122, C1 => n16, C2 => n119, A 
                           => n565, ZN => n453);
   U353 : AOI22_X1 port map( A1 => A(24), A2 => n10, B1 => A(23), B2 => n6, ZN 
                           => n565);
   U354 : NOR2_X2 port map( A1 => n646, A2 => B(2), ZN => n260);
   U355 : OAI221_X1 port map( B1 => n24, B2 => n113, C1 => n14, C2 => n110, A 
                           => n611, ZN => n185);
   U356 : AOI22_X1 port map( A1 => A(21), A2 => n11, B1 => A(20), B2 => n6, ZN 
                           => n611);
   U357 : AOI222_X1 port map( A1 => n429, A2 => n5, B1 => n619, B2 => n262, C1 
                           => n227, C2 => B(3), ZN => n327);
   U358 : INV_X1 port map( A => n376, ZN => n619);
   U359 : OAI221_X1 port map( B1 => n24, B2 => n76, C1 => n15, C2 => n73, A => 
                           n444, ZN => n154);
   U360 : AOI22_X1 port map( A1 => A(10), A2 => n11, B1 => A(9), B2 => n267, ZN
                           => n444);
   U361 : OAI221_X1 port map( B1 => n27, B2 => n79, C1 => n16, C2 => n76, A => 
                           n586, ZN => n305);
   U362 : AOI22_X1 port map( A1 => A(11), A2 => n10, B1 => A(10), B2 => n7, ZN 
                           => n586);
   U363 : OAI221_X1 port map( B1 => n26, B2 => n82, C1 => n16, C2 => n79, A => 
                           n567, ZN => n261);
   U364 : AOI22_X1 port map( A1 => A(12), A2 => n10, B1 => A(11), B2 => n6, ZN 
                           => n567);
   U365 : OAI221_X1 port map( B1 => n24, B2 => n622, C1 => n14, C2 => n621, A 
                           => n443, ZN => n219);
   U366 : AOI22_X1 port map( A1 => A(6), A2 => n11, B1 => A(5), B2 => n267, ZN 
                           => n443);
   U367 : OAI221_X1 port map( B1 => n24, B2 => n623, C1 => n14, C2 => n622, A 
                           => n306, ZN => n207);
   U368 : AOI22_X1 port map( A1 => A(7), A2 => n11, B1 => A(6), B2 => n7, ZN =>
                           n306);
   U369 : OAI221_X1 port map( B1 => n25, B2 => n65, C1 => n15, C2 => n623, A =>
                           n265, ZN => n193);
   U370 : AOI22_X1 port map( A1 => A(8), A2 => n9, B1 => A(7), B2 => n6, ZN => 
                           n265);
   U371 : OAI221_X1 port map( B1 => n27, B2 => n99, C1 => n17, C2 => n95, A => 
                           n610, ZN => n186);
   U372 : AOI22_X1 port map( A1 => A(17), A2 => n11, B1 => A(16), B2 => n7, ZN 
                           => n610);
   U373 : OAI221_X1 port map( B1 => n27, B2 => n73, C1 => n17, C2 => n65, A => 
                           n604, ZN => n178);
   U374 : AOI22_X1 port map( A1 => A(9), A2 => n9, B1 => A(8), B2 => n7, ZN => 
                           n604);
   U375 : OAI221_X1 port map( B1 => n25, B2 => n87, C1 => n15, C2 => n85, A => 
                           n537, ZN => n166);
   U376 : AOI22_X1 port map( A1 => A(14), A2 => n9, B1 => A(13), B2 => n6, ZN 
                           => n537);
   U377 : OAI221_X1 port map( B1 => n26, B2 => n91, C1 => n16, C2 => n87, A => 
                           n584, ZN => n516);
   U378 : AOI22_X1 port map( A1 => A(15), A2 => n10, B1 => A(14), B2 => n6, ZN 
                           => n584);
   U379 : OAI221_X1 port map( B1 => n25, B2 => n79, C1 => n15, C2 => n82, A => 
                           n494, ZN => n373);
   U380 : AOI22_X1 port map( A1 => A(15), A2 => n9, B1 => A(16), B2 => n267, ZN
                           => n494);
   U381 : OAI221_X1 port map( B1 => n25, B2 => n132, C1 => n15, C2 => n614, A 
                           => n523, ZN => n420);
   U382 : AOI22_X1 port map( A1 => A(4), A2 => n9, B1 => A(5), B2 => n267, ZN 
                           => n523);
   U383 : OAI221_X1 port map( B1 => n26, B2 => n614, C1 => n16, C2 => n616, A 
                           => n571, ZN => n407);
   U384 : AOI22_X1 port map( A1 => A(5), A2 => n10, B1 => A(6), B2 => n6, ZN =>
                           n571);
   U385 : OAI221_X1 port map( B1 => n26, B2 => n616, C1 => n16, C2 => n618, A 
                           => n554, ZN => n389);
   U386 : AOI22_X1 port map( A1 => A(6), A2 => n10, B1 => A(7), B2 => n6, ZN =>
                           n554);
   U387 : OAI221_X1 port map( B1 => n48, B2 => n27, C1 => n102, C2 => n14, A =>
                           n553, ZN => n390);
   U389 : AOI22_X1 port map( A1 => A(2), A2 => n10, B1 => A(3), B2 => n6, ZN =>
                           n553);
   U390 : OAI221_X1 port map( B1 => n26, B2 => n623, C1 => n16, C2 => n65, A =>
                           n542, ZN => n429);
   U391 : AOI22_X1 port map( A1 => A(11), A2 => n10, B1 => A(12), B2 => n6, ZN 
                           => n542);
   U392 : OAI221_X1 port map( B1 => n26, B2 => n110, C1 => n16, C2 => n107, A 
                           => n566, ZN => n452);
   U393 : AOI22_X1 port map( A1 => A(20), A2 => n10, B1 => A(19), B2 => n6, ZN 
                           => n566);
   U394 : OAI221_X1 port map( B1 => n26, B2 => n104, C1 => n16, C2 => n99, A =>
                           n538, ZN => n170);
   U395 : AOI22_X1 port map( A1 => A(18), A2 => n10, B1 => A(17), B2 => n6, ZN 
                           => n538);
   U396 : OAI221_X1 port map( B1 => n26, B2 => n107, C1 => n16, C2 => n104, A 
                           => n582, ZN => n464);
   U397 : AOI22_X1 port map( A1 => A(19), A2 => n10, B1 => A(18), B2 => n6, ZN 
                           => n582);
   U398 : AOI22_X1 port map( A1 => n7, A2 => A(1), B1 => n11, B2 => A(0), ZN =>
                           n362);
   U399 : NAND2_X1 port map( A1 => B(4), A2 => n579, ZN => n160);
   U400 : INV_X1 port map( A => A(31), ZN => n612);
   U401 : INV_X1 port map( A => n332, ZN => n627);
   U402 : AOI21_X1 port map( B1 => A(31), B2 => B(11), A => n487, ZN => n256);
   U403 : AOI21_X1 port map( B1 => A(31), B2 => B(25), A => n483, ZN => n250);
   U404 : OAI221_X1 port map( B1 => n24, B2 => n91, C1 => n14, C2 => n95, A => 
                           n430, ZN => n372);
   U405 : AOI22_X1 port map( A1 => A(19), A2 => n11, B1 => A(20), B2 => n7, ZN 
                           => n430);
   U406 : OAI221_X1 port map( B1 => n25, B2 => n82, C1 => n15, C2 => n85, A => 
                           n476, ZN => n419);
   U407 : AOI22_X1 port map( A1 => A(16), A2 => n9, B1 => A(17), B2 => n267, ZN
                           => n476);
   U408 : OAI221_X1 port map( B1 => n25, B2 => n85, C1 => n15, C2 => n87, A => 
                           n467, ZN => n406);
   U409 : AOI22_X1 port map( A1 => A(17), A2 => n9, B1 => A(18), B2 => n267, ZN
                           => n467);
   U410 : OAI221_X1 port map( B1 => n25, B2 => n87, C1 => n15, C2 => n91, A => 
                           n457, ZN => n388);
   U411 : AOI22_X1 port map( A1 => A(18), A2 => n9, B1 => A(19), B2 => n267, ZN
                           => n457);
   U412 : OAI221_X1 port map( B1 => n27, B2 => n621, C1 => n17, C2 => n620, A 
                           => n605, ZN => n234);
   U413 : AOI22_X1 port map( A1 => A(5), A2 => n11, B1 => A(4), B2 => n7, ZN =>
                           n605);
   U414 : OAI221_X1 port map( B1 => n258, B2 => n642, C1 => n196, C2 => n636, A
                           => n259, ZN => n247);
   U415 : AOI22_X1 port map( A1 => n260, A2 => n261, B1 => n262, B2 => n193, ZN
                           => n259);
   U416 : AOI222_X1 port map( A1 => A(4), A2 => n11, B1 => A(6), B2 => n29, C1 
                           => A(5), C2 => n18, ZN => n258);
   U417 : OAI221_X1 port map( B1 => n303, B2 => n642, C1 => n83, C2 => n636, A 
                           => n304, ZN => n298);
   U418 : AOI22_X1 port map( A1 => n260, A2 => n305, B1 => n262, B2 => n207, ZN
                           => n304);
   U419 : AOI222_X1 port map( A1 => A(3), A2 => n11, B1 => A(5), B2 => n28, C1 
                           => A(4), C2 => n19, ZN => n303);
   U420 : OAI221_X1 port map( B1 => n441, B2 => n642, C1 => n80, C2 => n636, A 
                           => n442, ZN => n435);
   U421 : AOI22_X1 port map( A1 => n260, A2 => n154, B1 => n262, B2 => n219, ZN
                           => n442);
   U422 : AOI222_X1 port map( A1 => A(2), A2 => n9, B1 => A(4), B2 => n28, C1 
                           => A(3), C2 => n18, ZN => n441);
   U423 : OAI221_X1 port map( B1 => n24, B2 => n95, C1 => n14, C2 => n99, A => 
                           n421, ZN => n361);
   U424 : AOI22_X1 port map( A1 => A(20), A2 => n11, B1 => A(21), B2 => n6, ZN 
                           => n421);
   U425 : OAI221_X1 port map( B1 => n25, B2 => n65, C1 => n15, C2 => n73, A => 
                           n524, ZN => n474);
   U426 : AOI22_X1 port map( A1 => A(12), A2 => n9, B1 => A(13), B2 => n267, ZN
                           => n524);
   U427 : OAI221_X1 port map( B1 => n24, B2 => n99, C1 => n14, C2 => n104, A =>
                           n408, ZN => n350);
   U429 : AOI22_X1 port map( A1 => A(21), A2 => n9, B1 => A(22), B2 => n7, ZN 
                           => n408);
   U430 : OAI221_X1 port map( B1 => n25, B2 => n73, C1 => n15, C2 => n76, A => 
                           n510, ZN => n465);
   U431 : AOI22_X1 port map( A1 => A(13), A2 => n9, B1 => A(14), B2 => n267, ZN
                           => n510);
   U432 : OAI221_X1 port map( B1 => n24, B2 => n104, C1 => n14, C2 => n107, A 
                           => n391, ZN => n339);
   U433 : AOI22_X1 port map( A1 => A(22), A2 => n10, B1 => A(23), B2 => n6, ZN 
                           => n391);
   U434 : OAI221_X1 port map( B1 => n25, B2 => n76, C1 => n15, C2 => n79, A => 
                           n497, ZN => n455);
   U435 : AOI22_X1 port map( A1 => A(14), A2 => n9, B1 => A(15), B2 => n6, ZN 
                           => n497);
   U436 : OAI221_X1 port map( B1 => n24, B2 => n107, C1 => n14, C2 => n110, A 
                           => n377, ZN => n324);
   U437 : AOI22_X1 port map( A1 => A(23), A2 => n9, B1 => A(24), B2 => n7, ZN 
                           => n377);
   U438 : OAI221_X1 port map( B1 => n24, B2 => n110, C1 => n14, C2 => n113, A 
                           => n364, ZN => n313);
   U439 : AOI22_X1 port map( A1 => A(24), A2 => n11, B1 => A(25), B2 => n6, ZN 
                           => n364);
   U440 : OAI221_X1 port map( B1 => n24, B2 => n113, C1 => n14, C2 => n116, A 
                           => n351, ZN => n289);
   U441 : AOI22_X1 port map( A1 => A(25), A2 => n9, B1 => A(26), B2 => n7, ZN 
                           => n351);
   U442 : OAI221_X1 port map( B1 => n24, B2 => n116, C1 => n14, C2 => n119, A 
                           => n340, ZN => n270);
   U443 : AOI22_X1 port map( A1 => A(26), A2 => n10, B1 => A(27), B2 => n6, ZN 
                           => n340);
   U444 : AOI221_X1 port map( B1 => n169, B2 => n452, C1 => n167, C2 => n453, A
                           => n563, ZN => n562);
   U445 : NOR3_X1 port map( A1 => n40, A2 => B(3), A3 => n333, ZN => n563);
   U446 : AOI221_X1 port map( B1 => n242, B2 => n432, C1 => n626, C2 => n71, A 
                           => n244, ZN => n431);
   U447 : INV_X1 port map( A => n433, ZN => n71);
   U448 : OAI21_X1 port map( B1 => n437, B2 => n249, A => n250, ZN => n432);
   U449 : AOI22_X1 port map( A1 => n434, A2 => n38, B1 => n41, B2 => n435, ZN 
                           => n433);
   U450 : AOI221_X1 port map( B1 => n242, B2 => n295, C1 => n626, C2 => n68, A 
                           => n244, ZN => n294);
   U451 : INV_X1 port map( A => n296, ZN => n68);
   U452 : OAI21_X1 port map( B1 => n299, B2 => n249, A => n250, ZN => n295);
   U453 : AOI22_X1 port map( A1 => n297, A2 => n38, B1 => n41, B2 => n298, ZN 
                           => n296);
   U454 : AOI221_X1 port map( B1 => n242, B2 => n243, C1 => n626, C2 => n59, A 
                           => n244, ZN => n241);
   U455 : INV_X1 port map( A => n245, ZN => n59);
   U456 : OAI21_X1 port map( B1 => n248, B2 => n249, A => n250, ZN => n243);
   U457 : AOI22_X1 port map( A1 => n246, A2 => n38, B1 => n42, B2 => n247, ZN 
                           => n245);
   U458 : AOI22_X1 port map( A1 => n639, A2 => n506, B1 => B(2), B2 => n382, ZN
                           => n333);
   U459 : AOI221_X1 port map( B1 => n276, B2 => n319, C1 => n278, C2 => n320, A
                           => n279, ZN => n318);
   U460 : OAI21_X1 port map( B1 => n321, B2 => n281, A => n282, ZN => n319);
   U462 : AOI21_X1 port map( B1 => n283, B2 => n322, A => n285, ZN => n321);
   U463 : OAI21_X1 port map( B1 => n323, B2 => n287, A => n288, ZN => n322);
   U464 : AOI221_X1 port map( B1 => n276, B2 => n309, C1 => n278, C2 => n128, A
                           => n279, ZN => n308);
   U465 : OAI21_X1 port map( B1 => n310, B2 => n281, A => n282, ZN => n309);
   U466 : AOI21_X1 port map( B1 => n283, B2 => n311, A => n285, ZN => n310);
   U467 : OAI21_X1 port map( B1 => n312, B2 => n287, A => n288, ZN => n311);
   U468 : AOI221_X1 port map( B1 => n276, B2 => n277, C1 => n278, C2 => n133, A
                           => n279, ZN => n275);
   U469 : OAI21_X1 port map( B1 => n280, B2 => n281, A => n282, ZN => n277);
   U470 : AOI21_X1 port map( B1 => n283, B2 => n284, A => n285, ZN => n280);
   U471 : OAI21_X1 port map( B1 => n286, B2 => n287, A => n288, ZN => n284);
   U472 : AOI221_X1 port map( B1 => n165, B2 => n324, C1 => n38, C2 => n53, A 
                           => n325, ZN => n317);
   U473 : INV_X1 port map( A => n327, ZN => n53);
   U474 : OAI222_X1 port map( A1 => n78, A2 => n635, B1 => n326, B2 => n641, C1
                           => n90, C2 => n644, ZN => n325);
   U475 : AOI222_X1 port map( A1 => A(27), A2 => n10, B1 => A(25), B2 => n28, 
                           C1 => A(26), C2 => n19, ZN => n326);
   U476 : AOI221_X1 port map( B1 => n165, B2 => n313, C1 => n38, C2 => n314, A 
                           => n315, ZN => n307);
   U477 : OAI222_X1 port map( A1 => n81, A2 => n635, B1 => n316, B2 => n641, C1
                           => n94, C2 => n644, ZN => n315);
   U478 : AOI222_X1 port map( A1 => A(28), A2 => n11, B1 => A(26), B2 => n28, 
                           C1 => A(27), C2 => n18, ZN => n316);
   U479 : AOI221_X1 port map( B1 => n165, B2 => n289, C1 => n38, C2 => n290, A 
                           => n291, ZN => n274);
   U480 : OAI222_X1 port map( A1 => n84, A2 => n635, B1 => n292, B2 => n641, C1
                           => n98, C2 => n644, ZN => n291);
   U481 : AOI222_X1 port map( A1 => A(29), A2 => n11, B1 => A(27), B2 => n31, 
                           C1 => A(28), C2 => n18, ZN => n292);
   U482 : AOI221_X1 port map( B1 => n165, B2 => n270, C1 => n38, C2 => n271, A 
                           => n272, ZN => n268);
   U483 : OAI222_X1 port map( A1 => n86, A2 => n635, B1 => n273, B2 => n641, C1
                           => n103, C2 => n644, ZN => n272);
   U484 : AOI222_X1 port map( A1 => A(30), A2 => n11, B1 => A(28), B2 => n30, 
                           C1 => A(29), C2 => n20, ZN => n273);
   U485 : NOR2_X1 port map( A1 => n490, A2 => B(18), ZN => n251);
   U486 : OAI22_X1 port map( A1 => B(2), A2 => n374, B1 => n639, B2 => n375, ZN
                           => n227);
   U487 : AOI21_X1 port map( B1 => n20, B2 => A(31), A => n533, ZN => n412);
   U488 : AOI21_X1 port map( B1 => n11, B2 => A(31), A => n580, ZN => n395);
   U489 : AOI21_X1 port map( B1 => B(1), B2 => A(31), A => n533, ZN => n417);
   U490 : AOI21_X1 port map( B1 => n8, B2 => A(31), A => n580, ZN => n400);
   U491 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n267);
   U492 : AOI211_X1 port map( C1 => n276, C2 => n330, A => n279, B => n331, ZN 
                           => n329);
   U493 : OAI21_X1 port map( B1 => n334, B2 => n281, A => n282, ZN => n330);
   U494 : NOR3_X1 port map( A1 => n332, A2 => B(3), A3 => n333, ZN => n331);
   U495 : AOI21_X1 port map( B1 => n283, B2 => n335, A => n285, ZN => n334);
   U496 : OAI221_X1 port map( B1 => n587, B2 => n436, C1 => n48, C2 => n32, A 
                           => n588, ZN => RES(0));
   U497 : AOI21_X1 port map( B1 => n242, B2 => n589, A => n244, ZN => n588);
   U498 : OAI21_X1 port map( B1 => n593, B2 => n249, A => n250, ZN => n589);
   U499 : AOI21_X1 port map( B1 => n251, B2 => n595, A => n253, ZN => n593);
   U500 : AND2_X1 port map( A1 => n491, A2 => n632, ZN => n276);
   U501 : NAND2_X1 port map( A1 => A(31), A2 => n490, ZN => n486);
   U502 : NOR2_X1 port map( A1 => B(2), A2 => B(3), ZN => n356);
   U503 : INV_X1 port map( A => A(10), ZN => n65);
   U504 : NAND2_X1 port map( A1 => n454, A2 => A(31), ZN => n401);
   U505 : OAI21_X1 port map( B1 => n489, B2 => n612, A => n162, ZN => n487);
   U506 : INV_X1 port map( A => B(3), ZN => n646);
   U507 : INV_X1 port map( A => A(11), ZN => n73);
   U508 : INV_X1 port map( A => A(15), ZN => n85);
   U509 : INV_X1 port map( A => A(16), ZN => n87);
   U510 : INV_X1 port map( A => A(9), ZN => n623);
   U511 : OAI21_X1 port map( B1 => n502, B2 => n152, A => n153, ZN => n501);
   U512 : AOI211_X1 port map( C1 => B(4), C2 => A(31), A => n503, B => n504, ZN
                           => n502);
   U513 : OAI22_X1 port map( A1 => n196, A2 => n505, B1 => n100, B2 => n157, ZN
                           => n504);
   U514 : OAI221_X1 port map( B1 => n126, B2 => n161, C1 => n115, C2 => n158, A
                           => n162, ZN => n503);
   U515 : NAND2_X1 port map( A1 => A(0), A2 => n7, ZN => n375);
   U516 : NOR2_X1 port map( A1 => n269, A2 => n38, ZN => n228);
   U517 : INV_X1 port map( A => A(30), ZN => n135);
   U518 : INV_X1 port map( A => A(12), ZN => n76);
   U519 : INV_X1 port map( A => A(13), ZN => n79);
   U520 : INV_X1 port map( A => A(14), ZN => n82);
   U521 : INV_X1 port map( A => A(19), ZN => n99);
   U522 : INV_X1 port map( A => A(20), ZN => n104);
   U523 : INV_X1 port map( A => A(21), ZN => n107);
   U524 : INV_X1 port map( A => A(22), ZN => n110);
   U525 : INV_X1 port map( A => A(23), ZN => n113);
   U526 : INV_X1 port map( A => A(24), ZN => n116);
   U527 : OR4_X1 port map( A1 => B(13), A2 => B(14), A3 => B(12), A4 => n596, 
                           ZN => n490);
   U528 : OR3_X1 port map( A1 => B(15), A2 => B(17), A3 => B(16), ZN => n596);
   U529 : INV_X1 port map( A => B(2), ZN => n639);
   U530 : INV_X1 port map( A => A(8), ZN => n622);
   U531 : INV_X1 port map( A => A(3), ZN => n614);
   U532 : AND3_X1 port map( A1 => n579, A2 => n591, A3 => n597, ZN => n445);
   U533 : NOR3_X1 port map( A1 => n152, A2 => n146, A3 => n629, ZN => n597);
   U534 : INV_X1 port map( A => n148, ZN => n629);
   U535 : AND2_X1 port map( A1 => n491, A2 => n648, ZN => n242);
   U536 : INV_X1 port map( A => A(17), ZN => n91);
   U537 : INV_X1 port map( A => A(7), ZN => n621);
   U538 : INV_X1 port map( A => A(18), ZN => n95);
   U539 : INV_X1 port map( A => A(25), ZN => n119);
   U540 : INV_X1 port map( A => A(29), ZN => n130);
   U541 : INV_X1 port map( A => B(25), ZN => n632);
   U542 : INV_X1 port map( A => A(4), ZN => n616);
   U543 : INV_X1 port map( A => A(27), ZN => n125);
   U544 : INV_X1 port map( A => A(26), ZN => n122);
   U545 : INV_X1 port map( A => A(6), ZN => n620);
   U546 : INV_X1 port map( A => A(5), ZN => n618);
   U547 : INV_X1 port map( A => A(28), ZN => n127);
   U548 : NAND2_X1 port map( A1 => n34, A2 => n648, ZN => n137);
   U549 : INV_X1 port map( A => A(2), ZN => n132);
   U550 : INV_X1 port map( A => n579, ZN => n647);
   U551 : OR2_X1 port map( A1 => n624, A2 => B(1), ZN => n1);
   U552 : INV_X1 port map( A => n436, ZN => n626);
   U553 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n263);
   U554 : NAND2_X1 port map( A1 => B(1), A2 => n624, ZN => n264);
   U555 : INV_X1 port map( A => A(1), ZN => n102);
   U556 : INV_X1 port map( A => B(11), ZN => n628);
   U557 : INV_X1 port map( A => A(0), ZN => n48);
   U558 : INV_X1 port map( A => B(18), ZN => n630);
   U559 : INV_X1 port map( A => B(0), ZN => n624);
   U560 : INV_X1 port map( A => B(4), ZN => n43);
   U561 : NOR3_X1 port map( A1 => B(9), A2 => B(8), A3 => B(10), ZN => n489);
   U562 : NOR3_X1 port map( A1 => B(7), A2 => B(6), A3 => B(5), ZN => n579);
   U563 : NOR3_X1 port map( A1 => B(28), A2 => B(27), A3 => B(26), ZN => n592);
   U564 : NAND3_X1 port map( A1 => n445, A2 => n34, A3 => LEFT_RIGHT, ZN => 
                           n269);
   U565 : NOR2_X1 port map( A1 => n481, A2 => LEFT_RIGHT, ZN => n244);
   U566 : AOI221_X1 port map( B1 => n140, B2 => n229, C1 => n142, C2 => n230, A
                           => n144, ZN => n225);
   U567 : OAI21_X1 port map( B1 => n231, B2 => n146, A => n147, ZN => n230);
   U568 : OAI221_X1 port map( B1 => n617, B2 => n641, C1 => n238, C2 => n40, A 
                           => n239, ZN => n229);
   U569 : AOI21_X1 port map( B1 => n148, B2 => n232, A => n150, ZN => n231);
   U570 : AOI221_X1 port map( B1 => n140, B2 => n498, C1 => n142, C2 => n499, A
                           => n144, ZN => n495);
   U571 : OAI21_X1 port map( B1 => n500, B2 => n146, A => n147, ZN => n499);
   U572 : OAI221_X1 port map( B1 => n100, B2 => n637, C1 => n196, C2 => n641, A
                           => n507, ZN => n498);
   U573 : AOI21_X1 port map( B1 => n148, B2 => n501, A => n150, ZN => n500);
   U574 : AOI221_X1 port map( B1 => n140, B2 => n69, C1 => n142, C2 => n215, A 
                           => n144, ZN => n213);
   U575 : INV_X1 port map( A => n222, ZN => n69);
   U576 : OAI21_X1 port map( B1 => n216, B2 => n146, A => n147, ZN => n215);
   U577 : AOI221_X1 port map( B1 => n219, B2 => n199, C1 => n223, C2 => n38, A 
                           => n224, ZN => n222);
   U578 : AOI221_X1 port map( B1 => n140, B2 => n66, C1 => n142, C2 => n203, A 
                           => n144, ZN => n201);
   U579 : INV_X1 port map( A => n210, ZN => n66);
   U580 : OAI21_X1 port map( B1 => n204, B2 => n146, A => n147, ZN => n203);
   U581 : AOI221_X1 port map( B1 => n207, B2 => n199, C1 => n211, C2 => n38, A 
                           => n212, ZN => n210);
   U582 : AOI221_X1 port map( B1 => n140, B2 => n60, C1 => n142, C2 => n189, A 
                           => n144, ZN => n187);
   U583 : INV_X1 port map( A => n198, ZN => n60);
   U584 : OAI21_X1 port map( B1 => n190, B2 => n146, A => n147, ZN => n189);
   U585 : AOI221_X1 port map( B1 => n193, B2 => n199, C1 => n114, C2 => n38, A 
                           => n200, ZN => n198);
   U586 : AOI221_X1 port map( B1 => n140, B2 => n173, C1 => n142, C2 => n174, A
                           => n144, ZN => n171);
   U587 : OAI21_X1 port map( B1 => n175, B2 => n146, A => n147, ZN => n174);
   U588 : OAI221_X1 port map( B1 => n64, B2 => n641, C1 => n182, C2 => n40, A 
                           => n183, ZN => n173);
   U589 : AOI21_X1 port map( B1 => n148, B2 => n176, A => n150, ZN => n175);
   U590 : AOI221_X1 port map( B1 => n140, B2 => n141, C1 => n142, C2 => n143, A
                           => n144, ZN => n136);
   U591 : OAI21_X1 port map( B1 => n145, B2 => n146, A => n147, ZN => n143);
   U592 : OAI221_X1 port map( B1 => n70, B2 => n641, C1 => n163, C2 => n41, A 
                           => n164, ZN => n141);
   U593 : AOI21_X1 port map( B1 => n148, B2 => n149, A => n150, ZN => n145);
   U594 : AOI221_X1 port map( B1 => n140, B2 => n572, C1 => n142, C2 => n573, A
                           => n144, ZN => n569);
   U595 : OAI21_X1 port map( B1 => n574, B2 => n146, A => n147, ZN => n573);
   U596 : OAI221_X1 port map( B1 => n67, B2 => n641, C1 => n344, C2 => n41, A 
                           => n581, ZN => n572);
   U597 : AOI21_X1 port map( B1 => n148, B2 => n575, A => n150, ZN => n574);
   U598 : AOI221_X1 port map( B1 => n140, B2 => n555, C1 => n142, C2 => n556, A
                           => n144, ZN => n551);
   U599 : OAI21_X1 port map( B1 => n557, B2 => n146, A => n147, ZN => n556);
   U600 : OAI221_X1 port map( B1 => n196, B2 => n637, C1 => n74, C2 => n641, A 
                           => n562, ZN => n555);
   U601 : AOI21_X1 port map( B1 => n148, B2 => n558, A => n150, ZN => n557);
   U602 : AOI221_X1 port map( B1 => n140, B2 => n543, C1 => n142, C2 => n544, A
                           => n144, ZN => n539);
   U603 : OAI21_X1 port map( B1 => n545, B2 => n146, A => n147, ZN => n544);
   U604 : OAI221_X1 port map( B1 => n89, B2 => n637, C1 => n77, C2 => n641, A 
                           => n550, ZN => n543);
   U605 : AOI21_X1 port map( B1 => n148, B2 => n546, A => n150, ZN => n545);
   U606 : AOI221_X1 port map( B1 => n140, B2 => n526, C1 => n142, C2 => n527, A
                           => n144, ZN => n521);
   U607 : OAI21_X1 port map( B1 => n528, B2 => n146, A => n147, ZN => n527);
   U608 : OAI221_X1 port map( B1 => n92, B2 => n637, C1 => n80, C2 => n641, A 
                           => n534, ZN => n526);
   U609 : AOI21_X1 port map( B1 => n148, B2 => n529, A => n150, ZN => n528);
   U610 : AOI221_X1 port map( B1 => n140, B2 => n511, C1 => n142, C2 => n512, A
                           => n144, ZN => n508);
   U611 : OAI21_X1 port map( B1 => n513, B2 => n146, A => n147, ZN => n512);
   U612 : OAI221_X1 port map( B1 => n96, B2 => n637, C1 => n83, C2 => n641, A 
                           => n520, ZN => n511);
   U613 : AOI21_X1 port map( B1 => n148, B2 => n514, A => n150, ZN => n513);
   U614 : AOI21_X1 port map( B1 => n633, B2 => n590, A => n144, ZN => n481);
   U615 : INV_X1 port map( A => n592, ZN => n633);
   U616 : NOR2_X1 port map( A1 => B(29), A2 => B(30), ZN => n591);
   U617 : INV_X1 port map( A => n590, ZN => n266);
   U618 : AND2_X1 port map( A1 => n140, A2 => n199, ZN => n278);
   U619 : NAND2_X1 port map( A1 => n140, A2 => n39, ZN => n332);
   U620 : NAND2_X1 port map( A1 => n140, A2 => n648, ZN => n436);
   U621 : INV_X1 port map( A => LEFT_RIGHT, ZN => n648);
   U622 : AND2_X1 port map( A1 => n142, A2 => n592, ZN => n491);
   U623 : NOR2_X2 port map( A1 => n634, A2 => LOGIC_ARITH, ZN => n142);
   U624 : INV_X1 port map( A => n591, ZN => n634);
   U625 : AND2_X1 port map( A1 => LOGIC_ARITH, A2 => n445, ZN => n140);
   U626 : NOR2_X1 port map( A1 => n612, A2 => LOGIC_ARITH, ZN => n590);
   U627 : OAI222_X1 port map( A1 => n268, A2 => n269, B1 => LEFT_RIGHT, B2 => 
                           n266, C1 => n612, C2 => n33, ZN => RES(31));
   U628 : OAI222_X1 port map( A1 => n187, A2 => n35, B1 => n188, B2 => n625, C1
                           => n621, C2 => n32, ZN => RES(7));
   U629 : OAI222_X1 port map( A1 => n171, A2 => n35, B1 => n54, B2 => n625, C1 
                           => n622, C2 => n32, ZN => RES(8));
   U630 : OAI222_X1 port map( A1 => n136, A2 => n35, B1 => n58, B2 => n625, C1 
                           => n623, C2 => n32, ZN => RES(9));
   U631 : OAI222_X1 port map( A1 => n539, A2 => n35, B1 => n327, B2 => n625, C1
                           => n76, C2 => n34, ZN => RES(12));
   U632 : OAI222_X1 port map( A1 => n521, A2 => n35, B1 => n56, B2 => n625, C1 
                           => n79, C2 => n34, ZN => RES(13));
   U633 : OAI222_X1 port map( A1 => n508, A2 => n35, B1 => n50, B2 => n625, C1 
                           => n82, C2 => n34, ZN => RES(14));
   U634 : OAI222_X1 port map( A1 => n468, A2 => n269, B1 => n469, B2 => n36, C1
                           => n91, C2 => n33, ZN => RES(17));
   U635 : OAI222_X1 port map( A1 => n495, A2 => n35, B1 => n46, B2 => n625, C1 
                           => n85, C2 => n34, ZN => RES(15));
   U636 : OAI222_X1 port map( A1 => n458, A2 => n269, B1 => n459, B2 => n37, C1
                           => n95, C2 => n33, ZN => RES(18));
   U640 : OAI222_X1 port map( A1 => n477, A2 => n269, B1 => n478, B2 => n37, C1
                           => n87, C2 => n34, ZN => RES(16));
   U643 : OAI222_X1 port map( A1 => n446, A2 => n269, B1 => n447, B2 => n36, C1
                           => n99, C2 => n33, ZN => RES(19));
   U644 : OAI222_X1 port map( A1 => n422, A2 => n269, B1 => n423, B2 => n36, C1
                           => n104, C2 => n33, ZN => RES(20));
   U645 : OAI222_X1 port map( A1 => n409, A2 => n269, B1 => n410, B2 => n36, C1
                           => n107, C2 => n33, ZN => RES(21));
   U646 : OAI222_X1 port map( A1 => n392, A2 => n269, B1 => n393, B2 => n36, C1
                           => n110, C2 => n33, ZN => RES(22));
   U647 : OAI222_X1 port map( A1 => n378, A2 => n269, B1 => n379, B2 => n36, C1
                           => n113, C2 => n33, ZN => RES(23));
   U648 : OAI222_X1 port map( A1 => n365, A2 => n269, B1 => n366, B2 => n36, C1
                           => n116, C2 => n33, ZN => RES(24));
   U649 : OAI222_X1 port map( A1 => n352, A2 => n269, B1 => n353, B2 => n36, C1
                           => n119, C2 => n33, ZN => RES(25));
   U650 : OAI222_X1 port map( A1 => n201, A2 => n35, B1 => n202, B2 => n625, C1
                           => n620, C2 => n32, ZN => RES(6));
   U651 : OAI222_X1 port map( A1 => n569, A2 => n35, B1 => n52, B2 => n625, C1 
                           => n65, C2 => n34, ZN => RES(10));
   U652 : OAI222_X1 port map( A1 => n551, A2 => n35, B1 => n44, B2 => n625, C1 
                           => n73, C2 => n34, ZN => RES(11));
   U653 : OAI222_X1 port map( A1 => n341, A2 => n269, B1 => n342, B2 => n36, C1
                           => n122, C2 => n33, ZN => RES(26));
   U654 : OAI222_X1 port map( A1 => n328, A2 => n269, B1 => n329, B2 => n36, C1
                           => n125, C2 => n33, ZN => RES(27));
   U655 : OAI222_X1 port map( A1 => n213, A2 => n35, B1 => n214, B2 => n625, C1
                           => n618, C2 => n32, ZN => RES(5));
   U656 : OAI222_X1 port map( A1 => n317, A2 => n269, B1 => n318, B2 => n36, C1
                           => n127, C2 => n33, ZN => RES(28));
   U657 : OAI222_X1 port map( A1 => n307, A2 => n269, B1 => n308, B2 => n36, C1
                           => n130, C2 => n32, ZN => RES(29));
   U658 : OAI222_X1 port map( A1 => n274, A2 => n269, B1 => n275, B2 => n37, C1
                           => n135, C2 => n32, ZN => RES(30));
   U659 : OAI221_X1 port map( B1 => n293, B2 => n240, C1 => n132, C2 => n32, A 
                           => n294, ZN => RES(2));
   U660 : OAI221_X1 port map( B1 => n362, B2 => n240, C1 => n102, C2 => n32, A 
                           => n431, ZN => RES(1));
   U661 : OAI221_X1 port map( B1 => n45, B2 => n240, C1 => n614, C2 => n32, A 
                           => n241, ZN => RES(3));
   U662 : OAI221_X1 port map( B1 => n225, B2 => n35, C1 => n616, C2 => n32, A 
                           => n226, ZN => RES(4));
   U663 : NOR4_X4 port map( A1 => B(16), A2 => B(17), A3 => B(15), A4 => n598, 
                           ZN => n148);
   U664 : INV_X1 port map( A => n8, ZN => n6);
   U665 : INV_X1 port map( A => n8, ZN => n7);
   U666 : INV_X1 port map( A => n1, ZN => n9);
   U667 : INV_X1 port map( A => n1, ZN => n10);
   U668 : INV_X1 port map( A => n1, ZN => n11);
   U669 : CLKBUF_X1 port map( A => n264, Z => n12);
   U670 : CLKBUF_X1 port map( A => n264, Z => n13);
   U671 : INV_X1 port map( A => n20, ZN => n17);
   U672 : INV_X1 port map( A => n12, ZN => n18);
   U673 : INV_X1 port map( A => n12, ZN => n19);
   U674 : INV_X1 port map( A => n12, ZN => n20);
   U675 : INV_X1 port map( A => n13, ZN => n21);
   U676 : CLKBUF_X1 port map( A => n263, Z => n22);
   U677 : CLKBUF_X1 port map( A => n263, Z => n23);
   U678 : INV_X1 port map( A => n22, ZN => n28);
   U679 : INV_X1 port map( A => n23, ZN => n29);
   U680 : INV_X1 port map( A => n23, ZN => n30);
   U681 : INV_X1 port map( A => n263, ZN => n31);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity comparator_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  OPSel : in std_logic_vector
         (0 to 2);  RES : out std_logic_vector (31 downto 0));

end comparator_NBIT32;

architecture SYN_bhv of comparator_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component comparator_NBIT32_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   signal X_Logic0_port, N26, N27, N28, N29, N30, N31, n10, n15, n16, n17, n18,
      n19, n20, RES_0_port, n2, n3, n4 : std_logic;

begin
   RES <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, RES_0_port 
      );
   
   X_Logic0_port <= '0';
   n10 <= '0';
   r57 : comparator_NBIT32_DW01_cmp6_0 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), TC => n10, LT => N30, GT => N28,
                           EQ => N26, LE => N31, GE => N29, NE => N27);
   U3 : INV_X1 port map( A => n15, ZN => RES_0_port);
   U4 : AOI21_X1 port map( B1 => n16, B2 => n4, A => n17, ZN => n15);
   U5 : NOR3_X1 port map( A1 => n4, A2 => OPSel(1), A3 => n18, ZN => n17);
   U6 : OAI22_X1 port map( A1 => n19, A2 => n3, B1 => OPSel(1), B2 => n20, ZN 
                           => n16);
   U7 : INV_X1 port map( A => OPSel(1), ZN => n3);
   U8 : AOI22_X1 port map( A1 => N28, A2 => n2, B1 => N29, B2 => OPSel(2), ZN 
                           => n19);
   U9 : INV_X1 port map( A => OPSel(2), ZN => n2);
   U10 : AOI22_X1 port map( A1 => N30, A2 => n2, B1 => OPSel(2), B2 => N31, ZN 
                           => n18);
   U11 : AOI22_X1 port map( A1 => N26, A2 => n2, B1 => N27, B2 => OPSel(2), ZN 
                           => n20);
   U12 : INV_X1 port map( A => OPSel(0), ZN => n4);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_NBIT32 is

   port( OP1, OP2 : in std_logic_vector (31 downto 0);  ALU_OPC : in 
         std_logic_vector (0 to 3);  ALU_RES : out std_logic_vector (31 downto 
         0));

end ALU_NBIT32;

architecture SYN_struct of ALU_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux21_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux41_NBIT32_1
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component P4Adder_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component shifter_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  LOGIC_ARITH, LEFT_RIGHT 
            : in std_logic;  RES : out std_logic_vector (31 downto 0));
   end component;
   
   component comparator_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  OPSel : in 
            std_logic_vector (0 to 2);  RES : out std_logic_vector (31 downto 
            0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, select_type_sig_1_port, select_type_sig_0_port, 
      select_zero_sig, A_SHF_31_port, A_SHF_30_port, A_SHF_29_port, 
      A_SHF_28_port, A_SHF_27_port, A_SHF_26_port, A_SHF_25_port, A_SHF_24_port
      , A_SHF_23_port, A_SHF_22_port, A_SHF_21_port, A_SHF_20_port, 
      A_SHF_19_port, A_SHF_18_port, A_SHF_17_port, A_SHF_16_port, A_SHF_15_port
      , A_SHF_14_port, A_SHF_13_port, A_SHF_12_port, A_SHF_11_port, 
      A_SHF_10_port, A_SHF_9_port, A_SHF_8_port, A_SHF_7_port, A_SHF_6_port, 
      A_SHF_5_port, A_SHF_4_port, A_SHF_3_port, A_SHF_2_port, A_SHF_1_port, 
      A_SHF_0_port, B_SHF_31_port, B_SHF_30_port, B_SHF_29_port, B_SHF_28_port,
      B_SHF_27_port, B_SHF_26_port, B_SHF_25_port, B_SHF_24_port, B_SHF_23_port
      , B_SHF_22_port, B_SHF_21_port, B_SHF_20_port, B_SHF_19_port, 
      B_SHF_18_port, B_SHF_17_port, B_SHF_16_port, B_SHF_15_port, B_SHF_14_port
      , B_SHF_13_port, B_SHF_12_port, B_SHF_11_port, B_SHF_10_port, 
      B_SHF_9_port, B_SHF_8_port, B_SHF_7_port, B_SHF_6_port, B_SHF_5_port, 
      B_SHF_4_port, B_SHF_3_port, B_SHF_2_port, B_SHF_1_port, B_SHF_0_port, 
      A_ADD_31_port, A_ADD_30_port, A_ADD_29_port, A_ADD_28_port, A_ADD_27_port
      , A_ADD_26_port, A_ADD_25_port, A_ADD_24_port, A_ADD_23_port, 
      A_ADD_22_port, A_ADD_21_port, A_ADD_20_port, A_ADD_19_port, A_ADD_18_port
      , A_ADD_17_port, A_ADD_16_port, A_ADD_15_port, A_ADD_14_port, 
      A_ADD_13_port, A_ADD_12_port, A_ADD_11_port, A_ADD_10_port, A_ADD_9_port,
      A_ADD_8_port, A_ADD_7_port, A_ADD_6_port, A_ADD_5_port, A_ADD_4_port, 
      A_ADD_3_port, A_ADD_2_port, A_ADD_1_port, A_ADD_0_port, B_ADD_31_port, 
      B_ADD_30_port, B_ADD_29_port, B_ADD_28_port, B_ADD_27_port, B_ADD_26_port
      , B_ADD_25_port, B_ADD_24_port, B_ADD_23_port, B_ADD_22_port, 
      B_ADD_21_port, B_ADD_20_port, B_ADD_19_port, B_ADD_18_port, B_ADD_17_port
      , B_ADD_16_port, B_ADD_15_port, B_ADD_14_port, B_ADD_13_port, 
      B_ADD_12_port, B_ADD_11_port, B_ADD_10_port, B_ADD_9_port, B_ADD_8_port, 
      B_ADD_7_port, B_ADD_6_port, B_ADD_5_port, B_ADD_4_port, B_ADD_3_port, 
      B_ADD_2_port, B_ADD_1_port, B_ADD_0_port, LOGIC_ARITH, OPSel_0_port, 
      LOGIC_RES_31_port, LOGIC_RES_30_port, LOGIC_RES_29_port, 
      LOGIC_RES_28_port, LOGIC_RES_27_port, LOGIC_RES_26_port, 
      LOGIC_RES_25_port, LOGIC_RES_24_port, LOGIC_RES_23_port, 
      LOGIC_RES_22_port, LOGIC_RES_21_port, LOGIC_RES_20_port, 
      LOGIC_RES_19_port, LOGIC_RES_18_port, LOGIC_RES_17_port, 
      LOGIC_RES_16_port, LOGIC_RES_15_port, LOGIC_RES_14_port, 
      LOGIC_RES_13_port, LOGIC_RES_12_port, LOGIC_RES_11_port, 
      LOGIC_RES_10_port, LOGIC_RES_9_port, LOGIC_RES_8_port, LOGIC_RES_7_port, 
      LOGIC_RES_6_port, LOGIC_RES_5_port, LOGIC_RES_4_port, LOGIC_RES_3_port, 
      LOGIC_RES_2_port, LOGIC_RES_1_port, LOGIC_RES_0_port, COMP_RES_31_port, 
      COMP_RES_30_port, COMP_RES_29_port, COMP_RES_28_port, COMP_RES_27_port, 
      COMP_RES_26_port, COMP_RES_25_port, COMP_RES_24_port, COMP_RES_23_port, 
      COMP_RES_22_port, COMP_RES_21_port, COMP_RES_20_port, COMP_RES_19_port, 
      COMP_RES_18_port, COMP_RES_17_port, COMP_RES_16_port, COMP_RES_15_port, 
      COMP_RES_14_port, COMP_RES_13_port, COMP_RES_12_port, COMP_RES_11_port, 
      COMP_RES_10_port, COMP_RES_9_port, COMP_RES_8_port, COMP_RES_7_port, 
      COMP_RES_6_port, COMP_RES_5_port, COMP_RES_4_port, COMP_RES_3_port, 
      COMP_RES_2_port, COMP_RES_1_port, COMP_RES_0_port, SHIFT_RES_31_port, 
      SHIFT_RES_30_port, SHIFT_RES_29_port, SHIFT_RES_28_port, 
      SHIFT_RES_27_port, SHIFT_RES_26_port, SHIFT_RES_25_port, 
      SHIFT_RES_24_port, SHIFT_RES_23_port, SHIFT_RES_22_port, 
      SHIFT_RES_21_port, SHIFT_RES_20_port, SHIFT_RES_19_port, 
      SHIFT_RES_18_port, SHIFT_RES_17_port, SHIFT_RES_16_port, 
      SHIFT_RES_15_port, SHIFT_RES_14_port, SHIFT_RES_13_port, 
      SHIFT_RES_12_port, SHIFT_RES_11_port, SHIFT_RES_10_port, SHIFT_RES_9_port
      , SHIFT_RES_8_port, SHIFT_RES_7_port, SHIFT_RES_6_port, SHIFT_RES_5_port,
      SHIFT_RES_4_port, SHIFT_RES_3_port, SHIFT_RES_2_port, SHIFT_RES_1_port, 
      SHIFT_RES_0_port, ADD_SUB_RES_31_port, ADD_SUB_RES_30_port, 
      ADD_SUB_RES_29_port, ADD_SUB_RES_28_port, ADD_SUB_RES_27_port, 
      ADD_SUB_RES_26_port, ADD_SUB_RES_25_port, ADD_SUB_RES_24_port, 
      ADD_SUB_RES_23_port, ADD_SUB_RES_22_port, ADD_SUB_RES_21_port, 
      ADD_SUB_RES_20_port, ADD_SUB_RES_19_port, ADD_SUB_RES_18_port, 
      ADD_SUB_RES_17_port, ADD_SUB_RES_16_port, ADD_SUB_RES_15_port, 
      ADD_SUB_RES_14_port, ADD_SUB_RES_13_port, ADD_SUB_RES_12_port, 
      ADD_SUB_RES_11_port, ADD_SUB_RES_10_port, ADD_SUB_RES_9_port, 
      ADD_SUB_RES_8_port, ADD_SUB_RES_7_port, ADD_SUB_RES_6_port, 
      ADD_SUB_RES_5_port, ADD_SUB_RES_4_port, ADD_SUB_RES_3_port, 
      ADD_SUB_RES_2_port, ADD_SUB_RES_1_port, ADD_SUB_RES_0_port, 
      sig_intraMux_31_port, sig_intraMux_30_port, sig_intraMux_29_port, 
      sig_intraMux_28_port, sig_intraMux_27_port, sig_intraMux_26_port, 
      sig_intraMux_25_port, sig_intraMux_24_port, sig_intraMux_23_port, 
      sig_intraMux_22_port, sig_intraMux_21_port, sig_intraMux_20_port, 
      sig_intraMux_19_port, sig_intraMux_18_port, sig_intraMux_17_port, 
      sig_intraMux_16_port, sig_intraMux_15_port, sig_intraMux_14_port, 
      sig_intraMux_13_port, sig_intraMux_12_port, sig_intraMux_11_port, 
      sig_intraMux_10_port, sig_intraMux_9_port, sig_intraMux_8_port, 
      sig_intraMux_7_port, sig_intraMux_6_port, sig_intraMux_5_port, 
      sig_intraMux_4_port, sig_intraMux_3_port, sig_intraMux_2_port, 
      sig_intraMux_1_port, sig_intraMux_0_port, n78, n79, n80, n81, n82, n83, 
      n84, n85, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99
      , n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n1, n2,
      n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n77, n86, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n_1122, n_1123, n_1124, n_1125, 
      n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, 
      n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, 
      n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, 
      n_1153 : std_logic;

begin
   
   X_Logic0_port <= '0';
   U177 : NOR2_X2 port map( A1 => n13, A2 => n55, ZN => A_SHF_31_port);
   U317 : NAND3_X1 port map( A1 => n185, A2 => n184, A3 => n186, ZN => n79);
   U318 : NAND3_X1 port map( A1 => n84, A2 => n83, A3 => n87, ZN => 
                           OPSel_0_port);
   U319 : NAND3_X1 port map( A1 => ALU_OPC(0), A2 => n186, A3 => n88, ZN => n87
                           );
   U320 : NAND3_X1 port map( A1 => ALU_OPC(0), A2 => n186, A3 => n89, ZN => n83
                           );
   U321 : NAND3_X1 port map( A1 => ALU_OPC(0), A2 => ALU_OPC(3), A3 => n89, ZN 
                           => n84);
   U322 : NAND3_X1 port map( A1 => ALU_OPC(1), A2 => ALU_OPC(2), A3 => n155, ZN
                           => n157);
   U323 : NAND3_X1 port map( A1 => ALU_OPC(1), A2 => ALU_OPC(2), A3 => n154, ZN
                           => n85);
   U324 : NAND3_X1 port map( A1 => n185, A2 => n184, A3 => n155, ZN => n156);
   Comp : comparator_NBIT32 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, OPSel(0) => n183, OPSel(1) => n182, 
                           OPSel(2) => OPSel_0_port, RES(31) => n_1122, RES(30)
                           => n_1123, RES(29) => n_1124, RES(28) => n_1125, 
                           RES(27) => n_1126, RES(26) => n_1127, RES(25) => 
                           n_1128, RES(24) => n_1129, RES(23) => n_1130, 
                           RES(22) => n_1131, RES(21) => n_1132, RES(20) => 
                           n_1133, RES(19) => n_1134, RES(18) => n_1135, 
                           RES(17) => n_1136, RES(16) => n_1137, RES(15) => 
                           n_1138, RES(14) => n_1139, RES(13) => n_1140, 
                           RES(12) => n_1141, RES(11) => n_1142, RES(10) => 
                           n_1143, RES(9) => n_1144, RES(8) => n_1145, RES(7) 
                           => n_1146, RES(6) => n_1147, RES(5) => n_1148, 
                           RES(4) => n_1149, RES(3) => n_1150, RES(2) => n_1151
                           , RES(1) => n_1152, RES(0) => COMP_RES_0_port);
   Shift : shifter_NBIT32 port map( A(31) => A_SHF_31_port, A(30) => 
                           A_SHF_30_port, A(29) => A_SHF_29_port, A(28) => 
                           A_SHF_28_port, A(27) => A_SHF_27_port, A(26) => 
                           A_SHF_26_port, A(25) => A_SHF_25_port, A(24) => 
                           A_SHF_24_port, A(23) => A_SHF_23_port, A(22) => 
                           A_SHF_22_port, A(21) => A_SHF_21_port, A(20) => 
                           A_SHF_20_port, A(19) => A_SHF_19_port, A(18) => 
                           A_SHF_18_port, A(17) => A_SHF_17_port, A(16) => 
                           A_SHF_16_port, A(15) => A_SHF_15_port, A(14) => 
                           A_SHF_14_port, A(13) => A_SHF_13_port, A(12) => 
                           A_SHF_12_port, A(11) => A_SHF_11_port, A(10) => 
                           A_SHF_10_port, A(9) => A_SHF_9_port, A(8) => 
                           A_SHF_8_port, A(7) => A_SHF_7_port, A(6) => 
                           A_SHF_6_port, A(5) => A_SHF_5_port, A(4) => 
                           A_SHF_4_port, A(3) => A_SHF_3_port, A(2) => 
                           A_SHF_2_port, A(1) => A_SHF_1_port, A(0) => 
                           A_SHF_0_port, B(31) => B_SHF_31_port, B(30) => 
                           B_SHF_30_port, B(29) => B_SHF_29_port, B(28) => 
                           B_SHF_28_port, B(27) => B_SHF_27_port, B(26) => 
                           B_SHF_26_port, B(25) => B_SHF_25_port, B(24) => 
                           B_SHF_24_port, B(23) => B_SHF_23_port, B(22) => 
                           B_SHF_22_port, B(21) => B_SHF_21_port, B(20) => 
                           B_SHF_20_port, B(19) => B_SHF_19_port, B(18) => 
                           B_SHF_18_port, B(17) => B_SHF_17_port, B(16) => 
                           B_SHF_16_port, B(15) => B_SHF_15_port, B(14) => 
                           B_SHF_14_port, B(13) => B_SHF_13_port, B(12) => 
                           B_SHF_12_port, B(11) => B_SHF_11_port, B(10) => 
                           B_SHF_10_port, B(9) => B_SHF_9_port, B(8) => 
                           B_SHF_8_port, B(7) => B_SHF_7_port, B(6) => 
                           B_SHF_6_port, B(5) => B_SHF_5_port, B(4) => 
                           B_SHF_4_port, B(3) => B_SHF_3_port, B(2) => 
                           B_SHF_2_port, B(1) => B_SHF_1_port, B(0) => 
                           B_SHF_0_port, LOGIC_ARITH => LOGIC_ARITH, LEFT_RIGHT
                           => n180, RES(31) => SHIFT_RES_31_port, RES(30) => 
                           SHIFT_RES_30_port, RES(29) => SHIFT_RES_29_port, 
                           RES(28) => SHIFT_RES_28_port, RES(27) => 
                           SHIFT_RES_27_port, RES(26) => SHIFT_RES_26_port, 
                           RES(25) => SHIFT_RES_25_port, RES(24) => 
                           SHIFT_RES_24_port, RES(23) => SHIFT_RES_23_port, 
                           RES(22) => SHIFT_RES_22_port, RES(21) => 
                           SHIFT_RES_21_port, RES(20) => SHIFT_RES_20_port, 
                           RES(19) => SHIFT_RES_19_port, RES(18) => 
                           SHIFT_RES_18_port, RES(17) => SHIFT_RES_17_port, 
                           RES(16) => SHIFT_RES_16_port, RES(15) => 
                           SHIFT_RES_15_port, RES(14) => SHIFT_RES_14_port, 
                           RES(13) => SHIFT_RES_13_port, RES(12) => 
                           SHIFT_RES_12_port, RES(11) => SHIFT_RES_11_port, 
                           RES(10) => SHIFT_RES_10_port, RES(9) => 
                           SHIFT_RES_9_port, RES(8) => SHIFT_RES_8_port, RES(7)
                           => SHIFT_RES_7_port, RES(6) => SHIFT_RES_6_port, 
                           RES(5) => SHIFT_RES_5_port, RES(4) => 
                           SHIFT_RES_4_port, RES(3) => SHIFT_RES_3_port, RES(2)
                           => SHIFT_RES_2_port, RES(1) => SHIFT_RES_1_port, 
                           RES(0) => SHIFT_RES_0_port);
   Add_Sub_unit : P4Adder_NBIT32 port map( A(31) => A_ADD_31_port, A(30) => 
                           A_ADD_30_port, A(29) => A_ADD_29_port, A(28) => 
                           A_ADD_28_port, A(27) => A_ADD_27_port, A(26) => 
                           A_ADD_26_port, A(25) => A_ADD_25_port, A(24) => 
                           A_ADD_24_port, A(23) => A_ADD_23_port, A(22) => 
                           A_ADD_22_port, A(21) => A_ADD_21_port, A(20) => 
                           A_ADD_20_port, A(19) => A_ADD_19_port, A(18) => 
                           A_ADD_18_port, A(17) => A_ADD_17_port, A(16) => 
                           A_ADD_16_port, A(15) => A_ADD_15_port, A(14) => 
                           A_ADD_14_port, A(13) => A_ADD_13_port, A(12) => 
                           A_ADD_12_port, A(11) => A_ADD_11_port, A(10) => 
                           A_ADD_10_port, A(9) => A_ADD_9_port, A(8) => 
                           A_ADD_8_port, A(7) => A_ADD_7_port, A(6) => 
                           A_ADD_6_port, A(5) => A_ADD_5_port, A(4) => 
                           A_ADD_4_port, A(3) => A_ADD_3_port, A(2) => 
                           A_ADD_2_port, A(1) => A_ADD_1_port, A(0) => 
                           A_ADD_0_port, B(31) => B_ADD_31_port, B(30) => 
                           B_ADD_30_port, B(29) => B_ADD_29_port, B(28) => 
                           B_ADD_28_port, B(27) => B_ADD_27_port, B(26) => 
                           B_ADD_26_port, B(25) => B_ADD_25_port, B(24) => 
                           B_ADD_24_port, B(23) => B_ADD_23_port, B(22) => 
                           B_ADD_22_port, B(21) => B_ADD_21_port, B(20) => 
                           B_ADD_20_port, B(19) => B_ADD_19_port, B(18) => 
                           B_ADD_18_port, B(17) => B_ADD_17_port, B(16) => 
                           B_ADD_16_port, B(15) => B_ADD_15_port, B(14) => 
                           B_ADD_14_port, B(13) => B_ADD_13_port, B(12) => 
                           B_ADD_12_port, B(11) => B_ADD_11_port, B(10) => 
                           B_ADD_10_port, B(9) => B_ADD_9_port, B(8) => 
                           B_ADD_8_port, B(7) => B_ADD_7_port, B(6) => 
                           B_ADD_6_port, B(5) => B_ADD_5_port, B(4) => 
                           B_ADD_4_port, B(3) => B_ADD_3_port, B(2) => 
                           B_ADD_2_port, B(1) => B_ADD_1_port, B(0) => 
                           B_ADD_0_port, Cin => n1, S(31) => 
                           ADD_SUB_RES_31_port, S(30) => ADD_SUB_RES_30_port, 
                           S(29) => ADD_SUB_RES_29_port, S(28) => 
                           ADD_SUB_RES_28_port, S(27) => ADD_SUB_RES_27_port, 
                           S(26) => ADD_SUB_RES_26_port, S(25) => 
                           ADD_SUB_RES_25_port, S(24) => ADD_SUB_RES_24_port, 
                           S(23) => ADD_SUB_RES_23_port, S(22) => 
                           ADD_SUB_RES_22_port, S(21) => ADD_SUB_RES_21_port, 
                           S(20) => ADD_SUB_RES_20_port, S(19) => 
                           ADD_SUB_RES_19_port, S(18) => ADD_SUB_RES_18_port, 
                           S(17) => ADD_SUB_RES_17_port, S(16) => 
                           ADD_SUB_RES_16_port, S(15) => ADD_SUB_RES_15_port, 
                           S(14) => ADD_SUB_RES_14_port, S(13) => 
                           ADD_SUB_RES_13_port, S(12) => ADD_SUB_RES_12_port, 
                           S(11) => ADD_SUB_RES_11_port, S(10) => 
                           ADD_SUB_RES_10_port, S(9) => ADD_SUB_RES_9_port, 
                           S(8) => ADD_SUB_RES_8_port, S(7) => 
                           ADD_SUB_RES_7_port, S(6) => ADD_SUB_RES_6_port, S(5)
                           => ADD_SUB_RES_5_port, S(4) => ADD_SUB_RES_4_port, 
                           S(3) => ADD_SUB_RES_3_port, S(2) => 
                           ADD_SUB_RES_2_port, S(1) => ADD_SUB_RES_1_port, S(0)
                           => ADD_SUB_RES_0_port, Cout => n_1153);
   Res_mux : mux41_NBIT32_1 port map( A(31) => ADD_SUB_RES_31_port, A(30) => 
                           ADD_SUB_RES_30_port, A(29) => ADD_SUB_RES_29_port, 
                           A(28) => ADD_SUB_RES_28_port, A(27) => 
                           ADD_SUB_RES_27_port, A(26) => ADD_SUB_RES_26_port, 
                           A(25) => ADD_SUB_RES_25_port, A(24) => 
                           ADD_SUB_RES_24_port, A(23) => ADD_SUB_RES_23_port, 
                           A(22) => ADD_SUB_RES_22_port, A(21) => 
                           ADD_SUB_RES_21_port, A(20) => ADD_SUB_RES_20_port, 
                           A(19) => ADD_SUB_RES_19_port, A(18) => 
                           ADD_SUB_RES_18_port, A(17) => ADD_SUB_RES_17_port, 
                           A(16) => ADD_SUB_RES_16_port, A(15) => 
                           ADD_SUB_RES_15_port, A(14) => ADD_SUB_RES_14_port, 
                           A(13) => ADD_SUB_RES_13_port, A(12) => 
                           ADD_SUB_RES_12_port, A(11) => ADD_SUB_RES_11_port, 
                           A(10) => ADD_SUB_RES_10_port, A(9) => 
                           ADD_SUB_RES_9_port, A(8) => ADD_SUB_RES_8_port, A(7)
                           => ADD_SUB_RES_7_port, A(6) => ADD_SUB_RES_6_port, 
                           A(5) => ADD_SUB_RES_5_port, A(4) => 
                           ADD_SUB_RES_4_port, A(3) => ADD_SUB_RES_3_port, A(2)
                           => ADD_SUB_RES_2_port, A(1) => ADD_SUB_RES_1_port, 
                           A(0) => ADD_SUB_RES_0_port, B(31) => 
                           LOGIC_RES_31_port, B(30) => LOGIC_RES_30_port, B(29)
                           => LOGIC_RES_29_port, B(28) => LOGIC_RES_28_port, 
                           B(27) => LOGIC_RES_27_port, B(26) => 
                           LOGIC_RES_26_port, B(25) => LOGIC_RES_25_port, B(24)
                           => LOGIC_RES_24_port, B(23) => LOGIC_RES_23_port, 
                           B(22) => LOGIC_RES_22_port, B(21) => 
                           LOGIC_RES_21_port, B(20) => LOGIC_RES_20_port, B(19)
                           => LOGIC_RES_19_port, B(18) => LOGIC_RES_18_port, 
                           B(17) => LOGIC_RES_17_port, B(16) => 
                           LOGIC_RES_16_port, B(15) => LOGIC_RES_15_port, B(14)
                           => LOGIC_RES_14_port, B(13) => LOGIC_RES_13_port, 
                           B(12) => LOGIC_RES_12_port, B(11) => 
                           LOGIC_RES_11_port, B(10) => LOGIC_RES_10_port, B(9) 
                           => LOGIC_RES_9_port, B(8) => LOGIC_RES_8_port, B(7) 
                           => LOGIC_RES_7_port, B(6) => LOGIC_RES_6_port, B(5) 
                           => LOGIC_RES_5_port, B(4) => LOGIC_RES_4_port, B(3) 
                           => LOGIC_RES_3_port, B(2) => LOGIC_RES_2_port, B(1) 
                           => LOGIC_RES_1_port, B(0) => LOGIC_RES_0_port, C(31)
                           => SHIFT_RES_31_port, C(30) => SHIFT_RES_30_port, 
                           C(29) => SHIFT_RES_29_port, C(28) => 
                           SHIFT_RES_28_port, C(27) => SHIFT_RES_27_port, C(26)
                           => SHIFT_RES_26_port, C(25) => SHIFT_RES_25_port, 
                           C(24) => SHIFT_RES_24_port, C(23) => 
                           SHIFT_RES_23_port, C(22) => SHIFT_RES_22_port, C(21)
                           => SHIFT_RES_21_port, C(20) => SHIFT_RES_20_port, 
                           C(19) => SHIFT_RES_19_port, C(18) => 
                           SHIFT_RES_18_port, C(17) => SHIFT_RES_17_port, C(16)
                           => SHIFT_RES_16_port, C(15) => SHIFT_RES_15_port, 
                           C(14) => SHIFT_RES_14_port, C(13) => 
                           SHIFT_RES_13_port, C(12) => SHIFT_RES_12_port, C(11)
                           => SHIFT_RES_11_port, C(10) => SHIFT_RES_10_port, 
                           C(9) => SHIFT_RES_9_port, C(8) => SHIFT_RES_8_port, 
                           C(7) => SHIFT_RES_7_port, C(6) => SHIFT_RES_6_port, 
                           C(5) => SHIFT_RES_5_port, C(4) => SHIFT_RES_4_port, 
                           C(3) => SHIFT_RES_3_port, C(2) => SHIFT_RES_2_port, 
                           C(1) => SHIFT_RES_1_port, C(0) => SHIFT_RES_0_port, 
                           D(31) => COMP_RES_31_port, D(30) => COMP_RES_30_port
                           , D(29) => COMP_RES_29_port, D(28) => 
                           COMP_RES_28_port, D(27) => COMP_RES_27_port, D(26) 
                           => COMP_RES_26_port, D(25) => COMP_RES_25_port, 
                           D(24) => COMP_RES_24_port, D(23) => COMP_RES_23_port
                           , D(22) => COMP_RES_22_port, D(21) => 
                           COMP_RES_21_port, D(20) => COMP_RES_20_port, D(19) 
                           => COMP_RES_19_port, D(18) => COMP_RES_18_port, 
                           D(17) => COMP_RES_17_port, D(16) => COMP_RES_16_port
                           , D(15) => COMP_RES_15_port, D(14) => 
                           COMP_RES_14_port, D(13) => COMP_RES_13_port, D(12) 
                           => COMP_RES_12_port, D(11) => COMP_RES_11_port, 
                           D(10) => COMP_RES_10_port, D(9) => COMP_RES_9_port, 
                           D(8) => COMP_RES_8_port, D(7) => COMP_RES_7_port, 
                           D(6) => COMP_RES_6_port, D(5) => COMP_RES_5_port, 
                           D(4) => COMP_RES_4_port, D(3) => COMP_RES_3_port, 
                           D(2) => COMP_RES_2_port, D(1) => COMP_RES_1_port, 
                           D(0) => COMP_RES_0_port, S(1) => 
                           select_type_sig_1_port, S(0) => 
                           select_type_sig_0_port, Z(31) => 
                           sig_intraMux_31_port, Z(30) => sig_intraMux_30_port,
                           Z(29) => sig_intraMux_29_port, Z(28) => 
                           sig_intraMux_28_port, Z(27) => sig_intraMux_27_port,
                           Z(26) => sig_intraMux_26_port, Z(25) => 
                           sig_intraMux_25_port, Z(24) => sig_intraMux_24_port,
                           Z(23) => sig_intraMux_23_port, Z(22) => 
                           sig_intraMux_22_port, Z(21) => sig_intraMux_21_port,
                           Z(20) => sig_intraMux_20_port, Z(19) => 
                           sig_intraMux_19_port, Z(18) => sig_intraMux_18_port,
                           Z(17) => sig_intraMux_17_port, Z(16) => 
                           sig_intraMux_16_port, Z(15) => sig_intraMux_15_port,
                           Z(14) => sig_intraMux_14_port, Z(13) => 
                           sig_intraMux_13_port, Z(12) => sig_intraMux_12_port,
                           Z(11) => sig_intraMux_11_port, Z(10) => 
                           sig_intraMux_10_port, Z(9) => sig_intraMux_9_port, 
                           Z(8) => sig_intraMux_8_port, Z(7) => 
                           sig_intraMux_7_port, Z(6) => sig_intraMux_6_port, 
                           Z(5) => sig_intraMux_5_port, Z(4) => 
                           sig_intraMux_4_port, Z(3) => sig_intraMux_3_port, 
                           Z(2) => sig_intraMux_2_port, Z(1) => 
                           sig_intraMux_1_port, Z(0) => sig_intraMux_0_port);
   Zeros_mux : mux21_NBIT32_1 port map( A(31) => sig_intraMux_31_port, A(30) =>
                           sig_intraMux_30_port, A(29) => sig_intraMux_29_port,
                           A(28) => sig_intraMux_28_port, A(27) => 
                           sig_intraMux_27_port, A(26) => sig_intraMux_26_port,
                           A(25) => sig_intraMux_25_port, A(24) => 
                           sig_intraMux_24_port, A(23) => sig_intraMux_23_port,
                           A(22) => sig_intraMux_22_port, A(21) => 
                           sig_intraMux_21_port, A(20) => sig_intraMux_20_port,
                           A(19) => sig_intraMux_19_port, A(18) => 
                           sig_intraMux_18_port, A(17) => sig_intraMux_17_port,
                           A(16) => sig_intraMux_16_port, A(15) => 
                           sig_intraMux_15_port, A(14) => sig_intraMux_14_port,
                           A(13) => sig_intraMux_13_port, A(12) => 
                           sig_intraMux_12_port, A(11) => sig_intraMux_11_port,
                           A(10) => sig_intraMux_10_port, A(9) => 
                           sig_intraMux_9_port, A(8) => sig_intraMux_8_port, 
                           A(7) => sig_intraMux_7_port, A(6) => 
                           sig_intraMux_6_port, A(5) => sig_intraMux_5_port, 
                           A(4) => sig_intraMux_4_port, A(3) => 
                           sig_intraMux_3_port, A(2) => sig_intraMux_2_port, 
                           A(1) => sig_intraMux_1_port, A(0) => 
                           sig_intraMux_0_port, B(31) => X_Logic0_port, B(30) 
                           => X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, S => select_zero_sig, Z(31) => 
                           ALU_RES(31), Z(30) => ALU_RES(30), Z(29) => 
                           ALU_RES(29), Z(28) => ALU_RES(28), Z(27) => 
                           ALU_RES(27), Z(26) => ALU_RES(26), Z(25) => 
                           ALU_RES(25), Z(24) => ALU_RES(24), Z(23) => 
                           ALU_RES(23), Z(22) => ALU_RES(22), Z(21) => 
                           ALU_RES(21), Z(20) => ALU_RES(20), Z(19) => 
                           ALU_RES(19), Z(18) => ALU_RES(18), Z(17) => 
                           ALU_RES(17), Z(16) => ALU_RES(16), Z(15) => 
                           ALU_RES(15), Z(14) => ALU_RES(14), Z(13) => 
                           ALU_RES(13), Z(12) => ALU_RES(12), Z(11) => 
                           ALU_RES(11), Z(10) => ALU_RES(10), Z(9) => 
                           ALU_RES(9), Z(8) => ALU_RES(8), Z(7) => ALU_RES(7), 
                           Z(6) => ALU_RES(6), Z(5) => ALU_RES(5), Z(4) => 
                           ALU_RES(4), Z(3) => ALU_RES(3), Z(2) => ALU_RES(2), 
                           Z(1) => ALU_RES(1), Z(0) => ALU_RES(0));
   U2 : NOR2_X1 port map( A1 => n13, A2 => n58, ZN => A_SHF_5_port);
   U3 : NOR2_X1 port map( A1 => n13, A2 => n59, ZN => A_SHF_6_port);
   U4 : BUF_X1 port map( A => n158, Z => n23);
   U5 : BUF_X1 port map( A => n158, Z => n24);
   U6 : BUF_X1 port map( A => n158, Z => n25);
   U7 : BUF_X1 port map( A => n177, Z => n5);
   U8 : BUF_X1 port map( A => n177, Z => n6);
   U9 : BUF_X1 port map( A => n177, Z => n7);
   U10 : BUF_X1 port map( A => n177, Z => n9);
   U11 : BUF_X1 port map( A => n177, Z => n8);
   U12 : BUF_X1 port map( A => n179, Z => n17);
   U13 : BUF_X1 port map( A => n179, Z => n18);
   U14 : BUF_X1 port map( A => n179, Z => n21);
   U15 : BUF_X1 port map( A => n179, Z => n20);
   U16 : BUF_X1 port map( A => n179, Z => n19);
   U17 : BUF_X1 port map( A => n176, Z => n2);
   U18 : BUF_X1 port map( A => n176, Z => n3);
   U19 : BUF_X1 port map( A => n176, Z => n4);
   U20 : AND2_X1 port map( A1 => n28, A2 => n29, ZN => n158);
   U21 : NOR2_X1 port map( A1 => n15, A2 => n168, ZN => B_SHF_3_port);
   U22 : NOR2_X1 port map( A1 => n12, A2 => n50, ZN => A_SHF_27_port);
   U23 : NOR2_X1 port map( A1 => n12, A2 => n49, ZN => A_SHF_26_port);
   U24 : NOR2_X1 port map( A1 => n13, A2 => n64, ZN => B_SHF_10_port);
   U25 : NOR2_X1 port map( A1 => n16, A2 => n174, ZN => B_SHF_9_port);
   U26 : NOR2_X1 port map( A1 => n16, A2 => n173, ZN => B_SHF_8_port);
   U27 : NOR2_X1 port map( A1 => n11, A2 => n39, ZN => A_SHF_17_port);
   U28 : NOR2_X1 port map( A1 => n13, A2 => n60, ZN => A_SHF_7_port);
   U29 : NOR2_X1 port map( A1 => n15, A2 => n165, ZN => B_SHF_2_port);
   U30 : NOR2_X1 port map( A1 => n11, A2 => n40, ZN => A_SHF_18_port);
   U31 : NOR2_X1 port map( A1 => n12, A2 => n48, ZN => A_SHF_25_port);
   U32 : NOR2_X1 port map( A1 => n13, A2 => n57, ZN => A_SHF_4_port);
   U33 : NOR2_X1 port map( A1 => n12, A2 => n51, ZN => A_SHF_28_port);
   U34 : NOR2_X1 port map( A1 => n15, A2 => n170, ZN => B_SHF_5_port);
   U35 : NOR2_X1 port map( A1 => n16, A2 => n172, ZN => B_SHF_7_port);
   U36 : NOR2_X1 port map( A1 => n16, A2 => n171, ZN => B_SHF_6_port);
   U37 : NOR2_X1 port map( A1 => n23, A2 => n31, ZN => A_ADD_0_port);
   U38 : NOR2_X1 port map( A1 => n13, A2 => n61, ZN => A_SHF_8_port);
   U39 : NOR2_X1 port map( A1 => n12, A2 => n53, ZN => A_SHF_2_port);
   U40 : NOR2_X1 port map( A1 => n25, A2 => n57, ZN => A_ADD_4_port);
   U41 : NOR2_X1 port map( A1 => n25, A2 => n58, ZN => A_ADD_5_port);
   U42 : NOR2_X1 port map( A1 => n25, A2 => n59, ZN => A_ADD_6_port);
   U43 : NOR2_X1 port map( A1 => n25, A2 => n61, ZN => A_ADD_8_port);
   U44 : NOR2_X1 port map( A1 => n25, A2 => n62, ZN => A_ADD_9_port);
   U45 : NOR2_X1 port map( A1 => n25, A2 => n56, ZN => A_ADD_3_port);
   U46 : NOR2_X1 port map( A1 => n25, A2 => n60, ZN => A_ADD_7_port);
   U47 : NOR2_X1 port map( A1 => n25, A2 => n55, ZN => A_ADD_31_port);
   U48 : NOR2_X1 port map( A1 => n23, A2 => n42, ZN => A_ADD_1_port);
   U49 : NOR2_X1 port map( A1 => n24, A2 => n53, ZN => A_ADD_2_port);
   U50 : NOR2_X1 port map( A1 => n23, A2 => n32, ZN => A_ADD_10_port);
   U51 : NOR2_X1 port map( A1 => n23, A2 => n34, ZN => A_ADD_12_port);
   U52 : NOR2_X1 port map( A1 => n23, A2 => n35, ZN => A_ADD_13_port);
   U53 : NOR2_X1 port map( A1 => n23, A2 => n36, ZN => A_ADD_14_port);
   U54 : NOR2_X1 port map( A1 => n23, A2 => n38, ZN => A_ADD_16_port);
   U55 : NOR2_X1 port map( A1 => n23, A2 => n39, ZN => A_ADD_17_port);
   U56 : NOR2_X1 port map( A1 => n23, A2 => n40, ZN => A_ADD_18_port);
   U57 : NOR2_X1 port map( A1 => n24, A2 => n43, ZN => A_ADD_20_port);
   U58 : NOR2_X1 port map( A1 => n24, A2 => n44, ZN => A_ADD_21_port);
   U59 : NOR2_X1 port map( A1 => n24, A2 => n45, ZN => A_ADD_22_port);
   U60 : NOR2_X1 port map( A1 => n24, A2 => n47, ZN => A_ADD_24_port);
   U61 : NOR2_X1 port map( A1 => n24, A2 => n48, ZN => A_ADD_25_port);
   U62 : NOR2_X1 port map( A1 => n24, A2 => n49, ZN => A_ADD_26_port);
   U63 : NOR2_X1 port map( A1 => n24, A2 => n51, ZN => A_ADD_28_port);
   U64 : NOR2_X1 port map( A1 => n24, A2 => n52, ZN => A_ADD_29_port);
   U65 : NOR2_X1 port map( A1 => n24, A2 => n54, ZN => A_ADD_30_port);
   U66 : NOR2_X1 port map( A1 => n23, A2 => n33, ZN => A_ADD_11_port);
   U67 : NOR2_X1 port map( A1 => n23, A2 => n37, ZN => A_ADD_15_port);
   U68 : NOR2_X1 port map( A1 => n23, A2 => n41, ZN => A_ADD_19_port);
   U69 : NOR2_X1 port map( A1 => n24, A2 => n46, ZN => A_ADD_23_port);
   U70 : NOR2_X1 port map( A1 => n24, A2 => n50, ZN => A_ADD_27_port);
   U71 : NOR2_X1 port map( A1 => n14, A2 => n74, ZN => B_SHF_1_port);
   U72 : NOR2_X1 port map( A1 => n12, A2 => n43, ZN => A_SHF_20_port);
   U73 : NOR2_X1 port map( A1 => n11, A2 => n34, ZN => A_SHF_12_port);
   U74 : NOR2_X1 port map( A1 => n12, A2 => n44, ZN => A_SHF_21_port);
   U75 : NOR2_X1 port map( A1 => n11, A2 => n35, ZN => A_SHF_13_port);
   U76 : NOR2_X1 port map( A1 => n11, A2 => n41, ZN => A_SHF_19_port);
   U77 : NOR2_X1 port map( A1 => n12, A2 => n45, ZN => A_SHF_22_port);
   U78 : NOR2_X1 port map( A1 => n11, A2 => n36, ZN => A_SHF_14_port);
   U79 : NOR2_X1 port map( A1 => n12, A2 => n46, ZN => A_SHF_23_port);
   U80 : NOR2_X1 port map( A1 => n12, A2 => n47, ZN => A_SHF_24_port);
   U81 : NOR2_X1 port map( A1 => n15, A2 => n163, ZN => B_SHF_28_port);
   U82 : NOR2_X1 port map( A1 => n15, A2 => n162, ZN => B_SHF_27_port);
   U83 : NOR2_X1 port map( A1 => n15, A2 => n161, ZN => B_SHF_26_port);
   U84 : NOR2_X1 port map( A1 => n11, A2 => n42, ZN => A_SHF_1_port);
   U85 : NOR2_X1 port map( A1 => n13, A2 => n65, ZN => B_SHF_11_port);
   U86 : NOR2_X1 port map( A1 => n13, A2 => n62, ZN => A_SHF_9_port);
   U87 : NOR2_X1 port map( A1 => n11, A2 => n31, ZN => A_SHF_0_port);
   U88 : NOR2_X1 port map( A1 => n11, A2 => n33, ZN => A_SHF_11_port);
   U89 : NOR2_X1 port map( A1 => n11, A2 => n37, ZN => A_SHF_15_port);
   U90 : NOR2_X1 port map( A1 => n12, A2 => n52, ZN => A_SHF_29_port);
   U91 : NOR2_X1 port map( A1 => n11, A2 => n38, ZN => A_SHF_16_port);
   U92 : NOR2_X1 port map( A1 => n13, A2 => n56, ZN => A_SHF_3_port);
   U93 : NOR2_X1 port map( A1 => n14, A2 => n72, ZN => B_SHF_18_port);
   U94 : BUF_X1 port map( A => n178, Z => n13);
   U95 : BUF_X1 port map( A => n178, Z => n14);
   U96 : BUF_X1 port map( A => n178, Z => n11);
   U97 : BUF_X1 port map( A => n178, Z => n12);
   U98 : BUF_X1 port map( A => n178, Z => n15);
   U99 : NOR2_X1 port map( A1 => n15, A2 => n164, ZN => B_SHF_29_port);
   U100 : NOR2_X1 port map( A1 => n15, A2 => n166, ZN => B_SHF_30_port);
   U101 : NOR2_X1 port map( A1 => n15, A2 => n160, ZN => B_SHF_25_port);
   U102 : NOR2_X1 port map( A1 => n13, A2 => n63, ZN => B_SHF_0_port);
   U103 : NOR2_X1 port map( A1 => n14, A2 => n70, ZN => B_SHF_16_port);
   U104 : NOR2_X1 port map( A1 => n11, A2 => n32, ZN => A_SHF_10_port);
   U105 : NOR2_X1 port map( A1 => n14, A2 => n71, ZN => B_SHF_17_port);
   U106 : NOR2_X1 port map( A1 => n14, A2 => n69, ZN => B_SHF_15_port);
   U107 : BUF_X1 port map( A => n156, Z => n27);
   U108 : BUF_X1 port map( A => n156, Z => n26);
   U109 : NOR2_X1 port map( A1 => n15, A2 => n159, ZN => B_SHF_24_port);
   U110 : NOR2_X1 port map( A1 => n14, A2 => n86, ZN => B_SHF_23_port);
   U111 : NOR2_X1 port map( A1 => n14, A2 => n77, ZN => B_SHF_22_port);
   U112 : NOR2_X1 port map( A1 => n15, A2 => n169, ZN => B_SHF_4_port);
   U113 : NAND4_X1 port map( A1 => n80, A2 => n81, A3 => n82, A4 => n181, ZN =>
                           select_type_sig_0_port);
   U114 : NOR2_X1 port map( A1 => n12, A2 => n54, ZN => A_SHF_30_port);
   U115 : INV_X1 port map( A => n81, ZN => n179);
   U116 : NOR2_X1 port map( A1 => n14, A2 => n73, ZN => B_SHF_19_port);
   U117 : NOR2_X1 port map( A1 => n14, A2 => n67, ZN => B_SHF_13_port);
   U118 : NOR2_X1 port map( A1 => n14, A2 => n76, ZN => B_SHF_21_port);
   U119 : NOR2_X1 port map( A1 => n14, A2 => n68, ZN => B_SHF_14_port);
   U120 : NOR2_X1 port map( A1 => n14, A2 => n75, ZN => B_SHF_20_port);
   U121 : NOR2_X1 port map( A1 => n13, A2 => n66, ZN => B_SHF_12_port);
   U122 : NAND2_X1 port map( A1 => n16, A2 => n181, ZN => 
                           select_type_sig_1_port);
   U123 : BUF_X1 port map( A => n156, Z => n28);
   U124 : INV_X1 port map( A => n80, ZN => n177);
   U125 : INV_X1 port map( A => n82, ZN => n176);
   U126 : NOR2_X1 port map( A1 => n15, A2 => n167, ZN => B_SHF_31_port);
   U127 : OAI22_X1 port map( A1 => n63, A2 => n28, B1 => OP2(0), B2 => n29, ZN 
                           => B_ADD_0_port);
   U128 : OAI22_X1 port map( A1 => n74, A2 => n27, B1 => OP2(1), B2 => n30, ZN 
                           => B_ADD_1_port);
   U129 : OAI22_X1 port map( A1 => n165, A2 => n26, B1 => OP2(2), B2 => n29, ZN
                           => B_ADD_2_port);
   U130 : OAI22_X1 port map( A1 => n169, A2 => n26, B1 => OP2(4), B2 => n29, ZN
                           => B_ADD_4_port);
   U131 : OAI22_X1 port map( A1 => n170, A2 => n26, B1 => OP2(5), B2 => n29, ZN
                           => B_ADD_5_port);
   U132 : OAI22_X1 port map( A1 => n171, A2 => n26, B1 => OP2(6), B2 => n29, ZN
                           => B_ADD_6_port);
   U133 : OAI22_X1 port map( A1 => n173, A2 => n26, B1 => OP2(8), B2 => n29, ZN
                           => B_ADD_8_port);
   U134 : OAI22_X1 port map( A1 => n174, A2 => n26, B1 => OP2(9), B2 => n29, ZN
                           => B_ADD_9_port);
   U135 : OAI22_X1 port map( A1 => n71, A2 => n27, B1 => OP2(17), B2 => n30, ZN
                           => B_ADD_17_port);
   U136 : OAI22_X1 port map( A1 => n72, A2 => n27, B1 => OP2(18), B2 => n30, ZN
                           => B_ADD_18_port);
   U137 : OAI22_X1 port map( A1 => n75, A2 => n27, B1 => OP2(20), B2 => n30, ZN
                           => B_ADD_20_port);
   U138 : OAI22_X1 port map( A1 => n76, A2 => n27, B1 => OP2(21), B2 => n30, ZN
                           => B_ADD_21_port);
   U139 : OAI22_X1 port map( A1 => n77, A2 => n27, B1 => OP2(22), B2 => n30, ZN
                           => B_ADD_22_port);
   U140 : OAI22_X1 port map( A1 => n159, A2 => n27, B1 => OP2(24), B2 => n30, 
                           ZN => B_ADD_24_port);
   U141 : OAI22_X1 port map( A1 => n160, A2 => n27, B1 => OP2(25), B2 => n30, 
                           ZN => B_ADD_25_port);
   U142 : OAI22_X1 port map( A1 => n161, A2 => n27, B1 => OP2(26), B2 => n30, 
                           ZN => B_ADD_26_port);
   U143 : OAI22_X1 port map( A1 => n163, A2 => n26, B1 => OP2(28), B2 => n29, 
                           ZN => B_ADD_28_port);
   U144 : OAI22_X1 port map( A1 => n164, A2 => n26, B1 => OP2(29), B2 => n29, 
                           ZN => B_ADD_29_port);
   U145 : OAI22_X1 port map( A1 => n166, A2 => n26, B1 => OP2(30), B2 => n29, 
                           ZN => B_ADD_30_port);
   U146 : OAI22_X1 port map( A1 => n168, A2 => n26, B1 => OP2(3), B2 => n29, ZN
                           => B_ADD_3_port);
   U147 : OAI22_X1 port map( A1 => n172, A2 => n26, B1 => OP2(7), B2 => n29, ZN
                           => B_ADD_7_port);
   U148 : OAI22_X1 port map( A1 => n73, A2 => n27, B1 => OP2(19), B2 => n30, ZN
                           => B_ADD_19_port);
   U149 : OAI22_X1 port map( A1 => n86, A2 => n27, B1 => OP2(23), B2 => n30, ZN
                           => B_ADD_23_port);
   U150 : OAI22_X1 port map( A1 => n162, A2 => n27, B1 => OP2(27), B2 => n30, 
                           ZN => B_ADD_27_port);
   U151 : OAI22_X1 port map( A1 => n167, A2 => n26, B1 => OP2(31), B2 => n29, 
                           ZN => B_ADD_31_port);
   U152 : OAI22_X1 port map( A1 => n64, A2 => n28, B1 => OP2(10), B2 => n30, ZN
                           => B_ADD_10_port);
   U153 : OAI22_X1 port map( A1 => n66, A2 => n28, B1 => OP2(12), B2 => n29, ZN
                           => B_ADD_12_port);
   U154 : OAI22_X1 port map( A1 => n67, A2 => n28, B1 => OP2(13), B2 => n30, ZN
                           => B_ADD_13_port);
   U155 : OAI22_X1 port map( A1 => n68, A2 => n28, B1 => OP2(14), B2 => n29, ZN
                           => B_ADD_14_port);
   U156 : OAI22_X1 port map( A1 => n70, A2 => n28, B1 => OP2(16), B2 => n30, ZN
                           => B_ADD_16_port);
   U157 : OAI22_X1 port map( A1 => n65, A2 => n28, B1 => OP2(11), B2 => n29, ZN
                           => B_ADD_11_port);
   U158 : OAI22_X1 port map( A1 => n69, A2 => n28, B1 => OP2(15), B2 => n30, ZN
                           => B_ADD_15_port);
   U159 : OAI22_X1 port map( A1 => n152, A2 => n63, B1 => n153, B2 => n31, ZN 
                           => LOGIC_RES_0_port);
   U160 : AOI21_X1 port map( B1 => n7, B2 => n63, A => n19, ZN => n153);
   U161 : AOI221_X1 port map( B1 => OP1(0), B2 => n4, C1 => n5, C2 => n31, A =>
                           n17, ZN => n152);
   U162 : OAI22_X1 port map( A1 => n130, A2 => n74, B1 => n131, B2 => n42, ZN 
                           => LOGIC_RES_1_port);
   U163 : AOI21_X1 port map( B1 => n9, B2 => n74, A => n21, ZN => n131);
   U164 : AOI221_X1 port map( B1 => OP1(1), B2 => n3, C1 => n6, C2 => n42, A =>
                           n18, ZN => n130);
   U165 : OAI22_X1 port map( A1 => n108, A2 => n165, B1 => n109, B2 => n53, ZN 
                           => LOGIC_RES_2_port);
   U166 : AOI21_X1 port map( B1 => n8, B2 => n165, A => n20, ZN => n109);
   U167 : AOI221_X1 port map( B1 => OP1(2), B2 => n2, C1 => n7, C2 => n53, A =>
                           n19, ZN => n108);
   U168 : OAI22_X1 port map( A1 => n102, A2 => n168, B1 => n103, B2 => n56, ZN 
                           => LOGIC_RES_3_port);
   U169 : AOI21_X1 port map( B1 => n8, B2 => n168, A => n20, ZN => n103);
   U170 : AOI221_X1 port map( B1 => OP1(3), B2 => n2, C1 => n6, C2 => n56, A =>
                           n18, ZN => n102);
   U171 : OAI22_X1 port map( A1 => n100, A2 => n169, B1 => n101, B2 => n57, ZN 
                           => LOGIC_RES_4_port);
   U172 : AOI21_X1 port map( B1 => n8, B2 => n169, A => n20, ZN => n101);
   U173 : AOI221_X1 port map( B1 => OP1(4), B2 => n2, C1 => n6, C2 => n57, A =>
                           n18, ZN => n100);
   U174 : OAI22_X1 port map( A1 => n98, A2 => n170, B1 => n99, B2 => n58, ZN =>
                           LOGIC_RES_5_port);
   U175 : AOI21_X1 port map( B1 => n7, B2 => n170, A => n19, ZN => n99);
   U176 : AOI221_X1 port map( B1 => OP1(5), B2 => n2, C1 => n6, C2 => n58, A =>
                           n18, ZN => n98);
   U178 : OAI22_X1 port map( A1 => n96, A2 => n171, B1 => n97, B2 => n59, ZN =>
                           LOGIC_RES_6_port);
   U179 : AOI21_X1 port map( B1 => n7, B2 => n171, A => n19, ZN => n97);
   U180 : AOI221_X1 port map( B1 => OP1(6), B2 => n2, C1 => n5, C2 => n59, A =>
                           n17, ZN => n96);
   U181 : OAI22_X1 port map( A1 => n94, A2 => n172, B1 => n95, B2 => n60, ZN =>
                           LOGIC_RES_7_port);
   U182 : AOI21_X1 port map( B1 => n8, B2 => n172, A => n20, ZN => n95);
   U183 : AOI221_X1 port map( B1 => OP1(7), B2 => n2, C1 => n5, C2 => n60, A =>
                           n17, ZN => n94);
   U184 : OAI22_X1 port map( A1 => n92, A2 => n173, B1 => n93, B2 => n61, ZN =>
                           LOGIC_RES_8_port);
   U185 : AOI21_X1 port map( B1 => n7, B2 => n173, A => n19, ZN => n93);
   U186 : AOI221_X1 port map( B1 => OP1(8), B2 => n2, C1 => n5, C2 => n61, A =>
                           n17, ZN => n92);
   U187 : OAI22_X1 port map( A1 => n90, A2 => n174, B1 => n91, B2 => n62, ZN =>
                           LOGIC_RES_9_port);
   U188 : AOI21_X1 port map( B1 => n8, B2 => n174, A => n20, ZN => n91);
   U189 : AOI221_X1 port map( B1 => n2, B2 => OP1(9), C1 => n5, C2 => n62, A =>
                           n17, ZN => n90);
   U190 : OAI22_X1 port map( A1 => n150, A2 => n64, B1 => n151, B2 => n32, ZN 
                           => LOGIC_RES_10_port);
   U191 : AOI21_X1 port map( B1 => n10, B2 => n64, A => n22, ZN => n151);
   U192 : AOI221_X1 port map( B1 => OP1(10), B2 => n4, C1 => n5, C2 => n32, A 
                           => n17, ZN => n150);
   U193 : OAI22_X1 port map( A1 => n148, A2 => n65, B1 => n149, B2 => n33, ZN 
                           => LOGIC_RES_11_port);
   U194 : AOI21_X1 port map( B1 => n10, B2 => n65, A => n22, ZN => n149);
   U195 : AOI221_X1 port map( B1 => OP1(11), B2 => n4, C1 => n5, C2 => n33, A 
                           => n17, ZN => n148);
   U196 : OAI22_X1 port map( A1 => n146, A2 => n66, B1 => n147, B2 => n34, ZN 
                           => LOGIC_RES_12_port);
   U197 : AOI21_X1 port map( B1 => n10, B2 => n66, A => n21, ZN => n147);
   U198 : AOI221_X1 port map( B1 => OP1(12), B2 => n4, C1 => n5, C2 => n34, A 
                           => n17, ZN => n146);
   U199 : OAI22_X1 port map( A1 => n144, A2 => n67, B1 => n145, B2 => n35, ZN 
                           => LOGIC_RES_13_port);
   U200 : AOI21_X1 port map( B1 => n10, B2 => n67, A => n21, ZN => n145);
   U201 : AOI221_X1 port map( B1 => OP1(13), B2 => n4, C1 => n5, C2 => n35, A 
                           => n17, ZN => n144);
   U202 : OAI22_X1 port map( A1 => n142, A2 => n68, B1 => n143, B2 => n36, ZN 
                           => LOGIC_RES_14_port);
   U203 : AOI21_X1 port map( B1 => n9, B2 => n68, A => n21, ZN => n143);
   U204 : AOI221_X1 port map( B1 => OP1(14), B2 => n4, C1 => n5, C2 => n36, A 
                           => n17, ZN => n142);
   U205 : OAI22_X1 port map( A1 => n140, A2 => n69, B1 => n141, B2 => n37, ZN 
                           => LOGIC_RES_15_port);
   U206 : AOI21_X1 port map( B1 => n9, B2 => n69, A => n21, ZN => n141);
   U207 : AOI221_X1 port map( B1 => OP1(15), B2 => n4, C1 => n5, C2 => n37, A 
                           => n17, ZN => n140);
   U208 : OAI22_X1 port map( A1 => n138, A2 => n70, B1 => n139, B2 => n38, ZN 
                           => LOGIC_RES_16_port);
   U209 : AOI21_X1 port map( B1 => n9, B2 => n70, A => n21, ZN => n139);
   U210 : AOI221_X1 port map( B1 => OP1(16), B2 => n4, C1 => n5, C2 => n38, A 
                           => n17, ZN => n138);
   U211 : OAI22_X1 port map( A1 => n136, A2 => n71, B1 => n137, B2 => n39, ZN 
                           => LOGIC_RES_17_port);
   U212 : AOI21_X1 port map( B1 => n9, B2 => n71, A => n21, ZN => n137);
   U213 : AOI221_X1 port map( B1 => OP1(17), B2 => n3, C1 => n6, C2 => n39, A 
                           => n18, ZN => n136);
   U214 : OAI22_X1 port map( A1 => n134, A2 => n72, B1 => n135, B2 => n40, ZN 
                           => LOGIC_RES_18_port);
   U215 : AOI21_X1 port map( B1 => n9, B2 => n72, A => n21, ZN => n135);
   U216 : AOI221_X1 port map( B1 => OP1(18), B2 => n3, C1 => n6, C2 => n40, A 
                           => n18, ZN => n134);
   U217 : OAI22_X1 port map( A1 => n132, A2 => n73, B1 => n133, B2 => n41, ZN 
                           => LOGIC_RES_19_port);
   U218 : AOI21_X1 port map( B1 => n9, B2 => n73, A => n21, ZN => n133);
   U219 : AOI221_X1 port map( B1 => OP1(19), B2 => n3, C1 => n6, C2 => n41, A 
                           => n18, ZN => n132);
   U220 : OAI22_X1 port map( A1 => n128, A2 => n75, B1 => n129, B2 => n43, ZN 
                           => LOGIC_RES_20_port);
   U221 : AOI21_X1 port map( B1 => n9, B2 => n75, A => n21, ZN => n129);
   U222 : AOI221_X1 port map( B1 => OP1(20), B2 => n3, C1 => n6, C2 => n43, A 
                           => n18, ZN => n128);
   U223 : OAI22_X1 port map( A1 => n126, A2 => n76, B1 => n127, B2 => n44, ZN 
                           => LOGIC_RES_21_port);
   U224 : AOI21_X1 port map( B1 => n9, B2 => n76, A => n21, ZN => n127);
   U225 : AOI221_X1 port map( B1 => OP1(21), B2 => n3, C1 => n6, C2 => n44, A 
                           => n18, ZN => n126);
   U226 : OAI22_X1 port map( A1 => n124, A2 => n77, B1 => n125, B2 => n45, ZN 
                           => LOGIC_RES_22_port);
   U227 : AOI21_X1 port map( B1 => n9, B2 => n77, A => n21, ZN => n125);
   U228 : AOI221_X1 port map( B1 => OP1(22), B2 => n3, C1 => n6, C2 => n45, A 
                           => n18, ZN => n124);
   U229 : OAI22_X1 port map( A1 => n122, A2 => n86, B1 => n123, B2 => n46, ZN 
                           => LOGIC_RES_23_port);
   U230 : AOI21_X1 port map( B1 => n9, B2 => n86, A => n21, ZN => n123);
   U231 : AOI221_X1 port map( B1 => OP1(23), B2 => n3, C1 => n6, C2 => n46, A 
                           => n18, ZN => n122);
   U232 : OAI22_X1 port map( A1 => n120, A2 => n159, B1 => n121, B2 => n47, ZN 
                           => LOGIC_RES_24_port);
   U233 : AOI21_X1 port map( B1 => n9, B2 => n159, A => n20, ZN => n121);
   U234 : AOI221_X1 port map( B1 => OP1(24), B2 => n3, C1 => n7, C2 => n47, A 
                           => n19, ZN => n120);
   U235 : OAI22_X1 port map( A1 => n118, A2 => n160, B1 => n119, B2 => n48, ZN 
                           => LOGIC_RES_25_port);
   U236 : AOI21_X1 port map( B1 => n8, B2 => n160, A => n20, ZN => n119);
   U237 : AOI221_X1 port map( B1 => OP1(25), B2 => n3, C1 => n7, C2 => n48, A 
                           => n19, ZN => n118);
   U238 : OAI22_X1 port map( A1 => n116, A2 => n161, B1 => n117, B2 => n49, ZN 
                           => LOGIC_RES_26_port);
   U239 : AOI21_X1 port map( B1 => n8, B2 => n161, A => n20, ZN => n117);
   U240 : AOI221_X1 port map( B1 => OP1(26), B2 => n3, C1 => n6, C2 => n49, A 
                           => n18, ZN => n116);
   U241 : OAI22_X1 port map( A1 => n114, A2 => n162, B1 => n115, B2 => n50, ZN 
                           => LOGIC_RES_27_port);
   U242 : AOI21_X1 port map( B1 => n8, B2 => n162, A => n20, ZN => n115);
   U243 : AOI221_X1 port map( B1 => OP1(27), B2 => n3, C1 => n7, C2 => n50, A 
                           => n19, ZN => n114);
   U244 : OAI22_X1 port map( A1 => n112, A2 => n163, B1 => n113, B2 => n51, ZN 
                           => LOGIC_RES_28_port);
   U245 : AOI21_X1 port map( B1 => n8, B2 => n163, A => n20, ZN => n113);
   U246 : AOI221_X1 port map( B1 => OP1(28), B2 => n2, C1 => n7, C2 => n51, A 
                           => n19, ZN => n112);
   U247 : OAI22_X1 port map( A1 => n110, A2 => n164, B1 => n111, B2 => n52, ZN 
                           => LOGIC_RES_29_port);
   U248 : AOI21_X1 port map( B1 => n8, B2 => n164, A => n20, ZN => n111);
   U249 : AOI221_X1 port map( B1 => OP1(29), B2 => n2, C1 => n7, C2 => n52, A 
                           => n19, ZN => n110);
   U250 : OAI22_X1 port map( A1 => n106, A2 => n166, B1 => n107, B2 => n54, ZN 
                           => LOGIC_RES_30_port);
   U251 : AOI21_X1 port map( B1 => n8, B2 => n166, A => n20, ZN => n107);
   U252 : AOI221_X1 port map( B1 => OP1(30), B2 => n2, C1 => n7, C2 => n54, A 
                           => n19, ZN => n106);
   U253 : OAI22_X1 port map( A1 => n104, A2 => n167, B1 => n105, B2 => n55, ZN 
                           => LOGIC_RES_31_port);
   U254 : AOI21_X1 port map( B1 => n8, B2 => n167, A => n20, ZN => n105);
   U255 : AOI221_X1 port map( B1 => OP1(31), B2 => n2, C1 => n7, C2 => n55, A 
                           => n19, ZN => n104);
   U256 : INV_X1 port map( A => n85, ZN => n180);
   U257 : INV_X1 port map( A => OPSel_0_port, ZN => n181);
   U258 : INV_X1 port map( A => OP1(10), ZN => n32);
   U259 : INV_X1 port map( A => OP1(16), ZN => n38);
   U260 : INV_X1 port map( A => OP1(20), ZN => n43);
   U261 : INV_X1 port map( A => OP1(4), ZN => n57);
   U262 : INV_X1 port map( A => OP1(12), ZN => n34);
   U263 : INV_X1 port map( A => OP1(21), ZN => n44);
   U264 : INV_X1 port map( A => OP1(13), ZN => n35);
   U265 : INV_X1 port map( A => OP1(22), ZN => n45);
   U266 : INV_X1 port map( A => OP1(14), ZN => n36);
   U267 : INV_X1 port map( A => OP1(0), ZN => n31);
   U268 : INV_X1 port map( A => OP1(1), ZN => n42);
   U269 : INV_X1 port map( A => OP1(2), ZN => n53);
   U270 : INV_X1 port map( A => OP1(17), ZN => n39);
   U271 : INV_X1 port map( A => OP1(18), ZN => n40);
   U272 : INV_X1 port map( A => OP1(5), ZN => n58);
   U273 : INV_X1 port map( A => OP1(6), ZN => n59);
   U274 : INV_X1 port map( A => OP1(24), ZN => n47);
   U275 : INV_X1 port map( A => OP1(25), ZN => n48);
   U276 : INV_X1 port map( A => OP1(28), ZN => n51);
   U277 : INV_X1 port map( A => OP1(29), ZN => n52);
   U278 : INV_X1 port map( A => OP1(30), ZN => n54);
   U279 : INV_X1 port map( A => OP1(8), ZN => n61);
   U280 : INV_X1 port map( A => OP1(9), ZN => n62);
   U281 : INV_X1 port map( A => OP1(26), ZN => n49);
   U282 : INV_X1 port map( A => OP1(3), ZN => n56);
   U283 : INV_X1 port map( A => OP1(7), ZN => n60);
   U284 : INV_X1 port map( A => OP1(11), ZN => n33);
   U285 : INV_X1 port map( A => OP1(15), ZN => n37);
   U286 : INV_X1 port map( A => OP1(19), ZN => n41);
   U287 : INV_X1 port map( A => OP1(23), ZN => n46);
   U288 : INV_X1 port map( A => OP1(27), ZN => n50);
   U289 : INV_X1 port map( A => OP1(31), ZN => n55);
   U290 : INV_X1 port map( A => OP2(1), ZN => n74);
   U291 : INV_X1 port map( A => OP2(0), ZN => n63);
   U292 : INV_X1 port map( A => OP2(2), ZN => n165);
   U293 : INV_X1 port map( A => OP2(6), ZN => n171);
   U294 : INV_X1 port map( A => OP2(5), ZN => n170);
   U295 : INV_X1 port map( A => OP2(4), ZN => n169);
   U296 : INV_X1 port map( A => OP2(13), ZN => n67);
   U297 : INV_X1 port map( A => OP2(14), ZN => n68);
   U298 : INV_X1 port map( A => OP2(12), ZN => n66);
   U299 : INV_X1 port map( A => OP2(16), ZN => n70);
   U300 : INV_X1 port map( A => OP2(17), ZN => n71);
   U301 : INV_X1 port map( A => OP2(8), ZN => n173);
   U302 : INV_X1 port map( A => OP2(9), ZN => n174);
   U303 : INV_X1 port map( A => OP2(10), ZN => n64);
   U304 : INV_X1 port map( A => OP2(18), ZN => n72);
   U305 : INV_X1 port map( A => OP2(21), ZN => n76);
   U306 : INV_X1 port map( A => OP2(20), ZN => n75);
   U307 : INV_X1 port map( A => OP2(30), ZN => n166);
   U308 : INV_X1 port map( A => OP2(29), ZN => n164);
   U309 : INV_X1 port map( A => OP2(24), ZN => n159);
   U310 : INV_X1 port map( A => OP2(22), ZN => n77);
   U311 : INV_X1 port map( A => OP2(25), ZN => n160);
   U312 : INV_X1 port map( A => OP2(26), ZN => n161);
   U313 : INV_X1 port map( A => OP2(28), ZN => n163);
   U314 : INV_X1 port map( A => OP2(3), ZN => n168);
   U315 : INV_X1 port map( A => OP2(7), ZN => n172);
   U316 : INV_X1 port map( A => OP2(11), ZN => n65);
   U325 : INV_X1 port map( A => OP2(15), ZN => n69);
   U326 : INV_X1 port map( A => OP2(19), ZN => n73);
   U327 : INV_X1 port map( A => OP2(23), ZN => n86);
   U328 : INV_X1 port map( A => OP2(27), ZN => n162);
   U329 : INV_X1 port map( A => OP2(31), ZN => n167);
   U330 : AND2_X1 port map( A1 => n154, A2 => n89, ZN => n1);
   U331 : INV_X1 port map( A => n83, ZN => n182);
   U332 : INV_X1 port map( A => LOGIC_ARITH, ZN => n178);
   U333 : NAND2_X1 port map( A1 => n155, A2 => n89, ZN => n82);
   U334 : NAND2_X1 port map( A1 => n155, A2 => n88, ZN => n80);
   U335 : NAND2_X1 port map( A1 => n154, A2 => n88, ZN => n81);
   U336 : INV_X1 port map( A => n84, ZN => n183);
   U337 : NOR2_X1 port map( A1 => n185, A2 => ALU_OPC(1), ZN => n89);
   U338 : NOR2_X1 port map( A1 => n186, A2 => ALU_OPC(0), ZN => n155);
   U339 : NOR2_X1 port map( A1 => n184, A2 => ALU_OPC(2), ZN => n88);
   U340 : NOR2_X1 port map( A1 => ALU_OPC(0), A2 => ALU_OPC(3), ZN => n154);
   U341 : NAND2_X1 port map( A1 => n85, A2 => n157, ZN => LOGIC_ARITH);
   U342 : OAI21_X1 port map( B1 => n78, B2 => n175, A => n79, ZN => 
                           select_zero_sig);
   U343 : INV_X1 port map( A => ALU_OPC(0), ZN => n175);
   U344 : AOI22_X1 port map( A1 => ALU_OPC(3), A2 => n185, B1 => ALU_OPC(1), B2
                           => ALU_OPC(2), ZN => n78);
   U345 : INV_X1 port map( A => ALU_OPC(2), ZN => n185);
   U346 : INV_X1 port map( A => ALU_OPC(3), ZN => n186);
   U347 : INV_X1 port map( A => ALU_OPC(1), ZN => n184);
   U348 : CLKBUF_X1 port map( A => n177, Z => n10);
   U349 : CLKBUF_X1 port map( A => n178, Z => n16);
   U350 : CLKBUF_X1 port map( A => n179, Z => n22);
   U351 : INV_X1 port map( A => n1, ZN => n29);
   U352 : INV_X1 port map( A => n1, ZN => n30);
   COMP_RES_1_port <= '0';
   COMP_RES_2_port <= '0';
   COMP_RES_3_port <= '0';
   COMP_RES_4_port <= '0';
   COMP_RES_5_port <= '0';
   COMP_RES_6_port <= '0';
   COMP_RES_7_port <= '0';
   COMP_RES_8_port <= '0';
   COMP_RES_9_port <= '0';
   COMP_RES_10_port <= '0';
   COMP_RES_11_port <= '0';
   COMP_RES_12_port <= '0';
   COMP_RES_13_port <= '0';
   COMP_RES_14_port <= '0';
   COMP_RES_15_port <= '0';
   COMP_RES_16_port <= '0';
   COMP_RES_17_port <= '0';
   COMP_RES_18_port <= '0';
   COMP_RES_19_port <= '0';
   COMP_RES_20_port <= '0';
   COMP_RES_21_port <= '0';
   COMP_RES_22_port <= '0';
   COMP_RES_23_port <= '0';
   COMP_RES_24_port <= '0';
   COMP_RES_25_port <= '0';
   COMP_RES_26_port <= '0';
   COMP_RES_27_port <= '0';
   COMP_RES_28_port <= '0';
   COMP_RES_29_port <= '0';
   COMP_RES_30_port <= '0';
   COMP_RES_31_port <= '0';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_0 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_0;

architecture SYN_bhv of mux41_NBIT32_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n1, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n6, Z => n72);
   U2 : BUF_X1 port map( A => n6, Z => n73);
   U3 : BUF_X1 port map( A => n4, Z => n78);
   U4 : BUF_X1 port map( A => n4, Z => n79);
   U5 : BUF_X1 port map( A => n7, Z => n1);
   U6 : BUF_X1 port map( A => n7, Z => n70);
   U7 : BUF_X1 port map( A => n5, Z => n75);
   U8 : BUF_X1 port map( A => n5, Z => n76);
   U9 : BUF_X1 port map( A => n6, Z => n74);
   U10 : BUF_X1 port map( A => n4, Z => n80);
   U11 : BUF_X1 port map( A => n7, Z => n71);
   U12 : BUF_X1 port map( A => n5, Z => n77);
   U13 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n6);
   U14 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n7);
   U15 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n4);
   U16 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n5);
   U17 : INV_X1 port map( A => S(0), ZN => n81);
   U18 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => Z(0));
   U19 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n69);
   U20 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n68);
   U21 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => Z(20));
   U22 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN 
                           => n45);
   U23 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN 
                           => n44);
   U24 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => Z(17));
   U25 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n53);
   U26 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n52);
   U27 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => Z(13));
   U28 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN 
                           => n61);
   U29 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n60);
   U30 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => Z(6));
   U31 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n13);
   U32 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n12);
   U33 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => Z(31));
   U34 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN 
                           => n21);
   U35 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN 
                           => n20);
   U36 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => Z(28));
   U37 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n29);
   U38 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n28);
   U39 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => Z(24));
   U40 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN 
                           => n37);
   U41 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN 
                           => n36);
   U42 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => Z(21));
   U43 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n43);
   U44 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n42);
   U45 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => Z(18));
   U46 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n51);
   U47 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n50);
   U48 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => Z(14));
   U49 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN 
                           => n59);
   U50 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n58);
   U51 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => Z(10));
   U52 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN 
                           => n67);
   U53 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n66);
   U54 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => Z(7));
   U55 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n11);
   U56 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n10);
   U57 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => Z(3));
   U58 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN =>
                           n19);
   U59 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN =>
                           n18);
   U60 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => Z(29));
   U61 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n27);
   U62 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n26);
   U63 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => Z(25));
   U64 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n35);
   U65 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n34);
   U66 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => Z(22));
   U67 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n41);
   U68 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n40);
   U69 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => Z(19));
   U70 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN 
                           => n49);
   U71 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n48);
   U72 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => Z(15));
   U73 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN 
                           => n57);
   U74 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n56);
   U75 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => Z(11));
   U76 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN 
                           => n65);
   U77 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n64);
   U78 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => Z(8));
   U79 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n9);
   U80 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n8);
   U81 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => Z(4));
   U82 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN =>
                           n17);
   U83 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN =>
                           n16);
   U84 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => Z(2));
   U85 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN =>
                           n25);
   U86 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN =>
                           n24);
   U87 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => Z(26));
   U88 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n33);
   U89 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n32);
   U90 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => Z(23));
   U91 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN 
                           => n39);
   U92 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN 
                           => n38);
   U93 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => Z(1));
   U94 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN =>
                           n47);
   U95 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN => 
                           n46);
   U96 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => Z(16));
   U97 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n55);
   U98 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n54);
   U99 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => Z(12));
   U100 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN
                           => n63);
   U101 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n62);
   U102 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Z(9));
   U103 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN 
                           => n3);
   U104 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN 
                           => n2);
   U105 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => Z(5));
   U106 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN 
                           => n15);
   U107 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN 
                           => n14);
   U108 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => Z(30));
   U109 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN
                           => n23);
   U110 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN
                           => n22);
   U111 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => Z(27));
   U112 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN
                           => n31);
   U113 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN
                           => n30);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FWD_Unit is

   port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB : in 
         std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;  
         FWDA, FWDB : out std_logic_vector (1 downto 0));

end FWD_Unit;

architecture SYN_bhv of FWD_Unit is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42 : std_logic;

begin
   
   U3 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => FWDB(1));
   U4 : AOI21_X1 port map( B1 => n3, B2 => n4, A => n5, ZN => n1);
   U5 : INV_X1 port map( A => n6, ZN => n3);
   U6 : NOR2_X1 port map( A1 => n2, A2 => n7, ZN => FWDB(0));
   U7 : MUX2_X1 port map( A => n6, B => n8, S => n5, Z => n7);
   U8 : AND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => n5);
   U9 : NOR2_X1 port map( A1 => n13, A2 => n14, ZN => n12);
   U10 : XOR2_X1 port map( A => ADD_WR_MEM(4), B => ADD_RS2(4), Z => n14);
   U11 : XOR2_X1 port map( A => ADD_WR_MEM(3), B => ADD_RS2(3), Z => n13);
   U12 : XNOR2_X1 port map( A => ADD_RS2(1), B => ADD_WR_MEM(1), ZN => n11);
   U13 : XNOR2_X1 port map( A => ADD_RS2(2), B => ADD_WR_MEM(2), ZN => n10);
   U14 : XNOR2_X1 port map( A => ADD_RS2(0), B => ADD_WR_MEM(0), ZN => n9);
   U15 : NAND4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           n6);
   U16 : NOR2_X1 port map( A1 => n19, A2 => n20, ZN => n18);
   U17 : XOR2_X1 port map( A => ADD_WR_WB(3), B => ADD_RS2(3), Z => n20);
   U18 : XOR2_X1 port map( A => ADD_WR_WB(2), B => ADD_RS2(2), Z => n19);
   U19 : XNOR2_X1 port map( A => ADD_RS2(4), B => ADD_WR_WB(4), ZN => n17);
   U20 : XNOR2_X1 port map( A => ADD_RS2(1), B => ADD_WR_WB(1), ZN => n16);
   U21 : XNOR2_X1 port map( A => ADD_RS2(0), B => ADD_WR_WB(0), ZN => n15);
   U22 : NOR2_X1 port map( A1 => n21, A2 => n2, ZN => FWDA(1));
   U23 : AOI21_X1 port map( B1 => n22, B2 => n4, A => n23, ZN => n21);
   U24 : OAI21_X1 port map( B1 => n24, B2 => n25, A => RF_WE_WB, ZN => n4);
   U25 : OR2_X1 port map( A1 => ADD_WR_WB(0), A2 => ADD_WR_WB(1), ZN => n25);
   U26 : OR3_X1 port map( A1 => ADD_WR_WB(3), A2 => ADD_WR_WB(4), A3 => 
                           ADD_WR_WB(2), ZN => n24);
   U27 : INV_X1 port map( A => n26, ZN => n22);
   U28 : NOR2_X1 port map( A1 => n2, A2 => n27, ZN => FWDA(0));
   U29 : MUX2_X1 port map( A => n26, B => n8, S => n23, Z => n27);
   U30 : AND4_X1 port map( A1 => n28, A2 => n29, A3 => n30, A4 => n31, ZN => 
                           n23);
   U31 : NOR2_X1 port map( A1 => n32, A2 => n33, ZN => n31);
   U32 : XOR2_X1 port map( A => ADD_WR_MEM(4), B => ADD_RS1(4), Z => n33);
   U33 : XOR2_X1 port map( A => ADD_WR_MEM(3), B => ADD_RS1(3), Z => n32);
   U34 : XNOR2_X1 port map( A => ADD_RS1(1), B => ADD_WR_MEM(1), ZN => n30);
   U35 : XNOR2_X1 port map( A => ADD_RS1(2), B => ADD_WR_MEM(2), ZN => n29);
   U36 : XNOR2_X1 port map( A => ADD_RS1(0), B => ADD_WR_MEM(0), ZN => n28);
   U37 : INV_X1 port map( A => n34, ZN => n8);
   U38 : OAI21_X1 port map( B1 => n35, B2 => n36, A => RF_WE_MEM, ZN => n34);
   U39 : OR2_X1 port map( A1 => ADD_WR_MEM(0), A2 => ADD_WR_MEM(1), ZN => n36);
   U40 : OR3_X1 port map( A1 => ADD_WR_MEM(3), A2 => ADD_WR_MEM(4), A3 => 
                           ADD_WR_MEM(2), ZN => n35);
   U41 : NAND4_X1 port map( A1 => n37, A2 => n38, A3 => n39, A4 => n40, ZN => 
                           n26);
   U42 : NOR2_X1 port map( A1 => n41, A2 => n42, ZN => n40);
   U43 : XOR2_X1 port map( A => ADD_WR_WB(3), B => ADD_RS1(3), Z => n42);
   U44 : XOR2_X1 port map( A => ADD_WR_WB(2), B => ADD_RS1(2), Z => n41);
   U45 : XNOR2_X1 port map( A => ADD_RS1(4), B => ADD_WR_WB(4), ZN => n39);
   U46 : XNOR2_X1 port map( A => ADD_RS1(1), B => ADD_WR_WB(1), ZN => n38);
   U47 : XNOR2_X1 port map( A => ADD_RS1(0), B => ADD_WR_WB(0), ZN => n37);
   U48 : INV_X1 port map( A => RST, ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N2 is

   port( DIN : in std_logic_vector (1 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (1 downto 0));

end regn_N2;

architecture SYN_bhv of regn_N2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   DOUT_reg_1_inst : DFFR_X1 port map( D => n6, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n4);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n5, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n3);
   U2 : OAI21_X1 port map( B1 => n3, B2 => EN, A => n1, ZN => n5);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n1);
   U4 : OAI21_X1 port map( B1 => n4, B2 => EN, A => n2, ZN => n6);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Branch_Cond_Unit_NBIT32 is

   port( RST : in std_logic;  A : in std_logic_vector (31 downto 0);  ALU_OPC :
         in std_logic_vector (0 to 3);  JUMP_TYPE : in std_logic_vector (1 
         downto 0);  PC_SEL : out std_logic_vector (1 downto 0);  ZERO : out 
         std_logic);

end Branch_Cond_Unit_NBIT32;

architecture SYN_bhv of Branch_Cond_Unit_NBIT32 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n1, n2 : std_logic;

begin
   
   U3 : NOR4_X1 port map( A1 => A(23), A2 => A(22), A3 => A(21), A4 => A(20), 
                           ZN => n15);
   U4 : NOR4_X1 port map( A1 => A(9), A2 => A(8), A3 => A(7), A4 => A(6), ZN =>
                           n19);
   U5 : NAND4_X1 port map( A1 => n12, A2 => n13, A3 => n14, A4 => n15, ZN => 
                           n11);
   U6 : NOR4_X1 port map( A1 => A(12), A2 => A(11), A3 => A(10), A4 => A(0), ZN
                           => n12);
   U7 : NOR4_X1 port map( A1 => A(16), A2 => A(15), A3 => A(14), A4 => A(13), 
                           ZN => n13);
   U8 : NOR4_X1 port map( A1 => A(1), A2 => A(19), A3 => A(18), A4 => A(17), ZN
                           => n14);
   U9 : NAND4_X1 port map( A1 => n16, A2 => n17, A3 => n18, A4 => n19, ZN => 
                           n10);
   U10 : NOR4_X1 port map( A1 => A(27), A2 => A(26), A3 => A(25), A4 => A(24), 
                           ZN => n16);
   U11 : NOR4_X1 port map( A1 => A(30), A2 => A(2), A3 => A(29), A4 => A(28), 
                           ZN => n17);
   U12 : NOR4_X1 port map( A1 => A(5), A2 => A(4), A3 => A(3), A4 => A(31), ZN 
                           => n18);
   U13 : NOR4_X1 port map( A1 => ALU_OPC(3), A2 => n1, A3 => ALU_OPC(1), A4 => 
                           ALU_OPC(2), ZN => n7);
   U14 : OAI211_X1 port map( C1 => n5, C2 => n6, A => JUMP_TYPE(0), B => RST, 
                           ZN => n4);
   U15 : AND2_X1 port map( A1 => n7, A2 => n8, ZN => n6);
   U16 : NOR4_X1 port map( A1 => n8, A2 => n9, A3 => n7, A4 => n1, ZN => n5);
   U17 : NOR2_X1 port map( A1 => n10, A2 => n11, ZN => n8);
   U18 : NAND2_X1 port map( A1 => JUMP_TYPE(1), A2 => RST, ZN => n3);
   U19 : INV_X1 port map( A => ALU_OPC(0), ZN => n1);
   U20 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => ZERO);
   U21 : OAI22_X1 port map( A1 => JUMP_TYPE(0), A2 => n3, B1 => JUMP_TYPE(1), 
                           B2 => n4, ZN => PC_SEL(0));
   U22 : NOR2_X1 port map( A1 => n2, A2 => n3, ZN => PC_SEL(1));
   U23 : INV_X1 port map( A => JUMP_TYPE(0), ZN => n2);
   U24 : OR2_X1 port map( A1 => ALU_OPC(2), A2 => ALU_OPC(1), ZN => n9);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity register_file_NBIT_ADD5_NBIT_DATA32 is

   port( CLK, RST, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RS1, 
         ADD_RS2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_NBIT_ADD5_NBIT_DATA32;

architecture SYN_bhv of register_file_NBIT_ADD5_NBIT_DATA32 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
      n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, 
      n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, 
      n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, 
      n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, 
      n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, 
      n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, 
      n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, 
      n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, 
      n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, 
      n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, 
      n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, 
      n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, 
      n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, 
      n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, 
      n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, 
      n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, 
      n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, 
      n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, 
      n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, 
      n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, 
      n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, 
      n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, 
      n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
      n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, 
      n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, 
      n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, 
      n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, 
      n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, 
      n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, 
      n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, 
      n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, 
      n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, 
      n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, 
      n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, 
      n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, 
      n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, 
      n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, 
      n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, 
      n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, 
      n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, 
      n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, 
      n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, 
      n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, 
      n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, 
      n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, 
      n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, 
      n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, 
      n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, 
      n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, 
      n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, 
      n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
      n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, 
      n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, 
      n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, 
      n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, 
      n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, 
      n3553, n3554, n3555, n3556, n3557, n3558, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
      n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
      n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
      n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
      n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
      n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
      n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
      n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
      n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, 
      n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, 
      n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, 
      n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, 
      n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, 
      n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, 
      n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, 
      n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, 
      n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, 
      n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, 
      n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, 
      n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, 
      n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, 
      n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
      n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, 
      n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, 
      n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, 
      n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, 
      n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, 
      n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, 
      n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, 
      n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, 
      n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, 
      n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, 
      n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, 
      n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, 
      n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, 
      n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, 
      n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, 
      n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, 
      n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, 
      n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, 
      n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, 
      n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, 
      n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, 
      n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, 
      n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, 
      n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, 
      n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, 
      n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, 
      n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, 
      n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, 
      n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, 
      n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, 
      n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, 
      n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, 
      n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, 
      n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, 
      n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, 
      n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, 
      n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, 
      n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, 
      n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, 
      n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, 
      n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, 
      n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
      n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
      n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, 
      n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, 
      n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, 
      n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, 
      n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, 
      n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, 
      n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, 
      n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, 
      n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, 
      n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, 
      n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, 
      n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, 
      n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, 
      n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, 
      n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, 
      n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, 
      n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, 
      n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, 
      n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, 
      n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, 
      n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
      n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, 
      n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, 
      n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, 
      n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, 
      n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, 
      n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, 
      n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, 
      n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, 
      n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, 
      n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, 
      n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, 
      n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, 
      n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, 
      n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, 
      n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, 
      n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, 
      n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, 
      n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, 
      n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, 
      n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, 
      n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, 
      n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, 
      n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, 
      n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, 
      n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, 
      n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, 
      n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, 
      n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, 
      n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, 
      n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, 
      n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, 
      n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, 
      n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, 
      n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, 
      n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, 
      n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, 
      n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, 
      n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, 
      n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, 
      n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, 
      n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, 
      n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, 
      n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, 
      n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, 
      n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, 
      n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, 
      n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, 
      n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, 
      n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, 
      n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, 
      n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, 
      n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, 
      n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, 
      n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, 
      n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, 
      n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, 
      n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, 
      n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, 
      n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, 
      n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, 
      n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, 
      n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, 
      n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, 
      n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, 
      n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, 
      n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, 
      n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, 
      n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, 
      n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, 
      n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, 
      n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, 
      n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, 
      n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, 
      n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
      n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
      n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
      n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, 
      n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
      n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
      n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, 
      n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, 
      n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, 
      n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, 
      n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
      n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, 
      n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, 
      n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, 
      n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
      n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, 
      n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, 
      n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, 
      n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, 
      n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, 
      n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, 
      n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, 
      n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, 
      n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, 
      n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, 
      n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, 
      n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, 
      n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, 
      n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, 
      n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, 
      n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, 
      n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, 
      n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, 
      n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, 
      n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, 
      n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, 
      n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, 
      n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, 
      n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, 
      n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, 
      n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, 
      n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, 
      n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, 
      n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, 
      n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, 
      n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, 
      n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, 
      n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, 
      n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, 
      n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, 
      n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, 
      n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, 
      n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, 
      n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, 
      n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, 
      n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, 
      n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, 
      n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, 
      n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, 
      n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, 
      n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, 
      n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, 
      n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, 
      n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, 
      n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, 
      n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, 
      n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, 
      n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, 
      n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, 
      n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, 
      n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, 
      n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, 
      n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, 
      n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, 
      n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, 
      n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, 
      n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, 
      n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, 
      n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, 
      n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, 
      n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, 
      n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, 
      n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, 
      n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, 
      n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, 
      n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, 
      n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, 
      n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, 
      n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, 
      n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, 
      n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, 
      n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, 
      n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, 
      n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, 
      n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, 
      n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, 
      n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, 
      n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, 
      n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, 
      n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, 
      n2978, n2979, n2980, n2981, n2982, n3559, n3560, n3561, n3562, n3563, 
      n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, 
      n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, 
      n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, 
      n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, 
      n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, 
      n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, 
      n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, 
      n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, 
      n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, 
      n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, 
      n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, 
      n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, 
      n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, 
      n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, 
      n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, 
      n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, 
      n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, 
      n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, 
      n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, 
      n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, 
      n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, 
      n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, 
      n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, 
      n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, 
      n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, 
      n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, 
      n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, 
      n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, 
      n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, 
      n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, 
      n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, 
      n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, 
      n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, 
      n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, 
      n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, 
      n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, 
      n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, 
      n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, 
      n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, 
      n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, 
      n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, 
      n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, 
      n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, 
      n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, 
      n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, 
      n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, 
      n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, 
      n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, 
      n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, 
      n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, 
      n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, 
      n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, 
      n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, 
      n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, 
      n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, 
      n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, 
      n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, 
      n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, 
      n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, 
      n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, 
      n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, 
      n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, 
      n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, 
      n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, 
      n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, 
      n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, 
      n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, 
      n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, 
      n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, 
      n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, 
      n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, 
      n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, 
      n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, 
      n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, 
      n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, 
      n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, 
      n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, 
      n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, 
      n4344, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, 
      n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, 
      n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, 
      n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, 
      n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, 
      n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, 
      n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, 
      n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, 
      n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, 
      n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, 
      n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, 
      n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, 
      n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, 
      n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, 
      n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, 
      n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, 
      n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, 
      n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, 
      n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, 
      n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, 
      n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, 
      n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, 
      n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, 
      n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, 
      n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, 
      n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, 
      n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, 
      n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, 
      n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, 
      n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, 
      n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, 
      n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, 
      n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, 
      n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, 
      n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, 
      n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, 
      n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, 
      n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, 
      n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, 
      n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, 
      n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, 
      n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, 
      n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, 
      n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, 
      n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, 
      n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, 
      n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, 
      n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, 
      n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, 
      n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, 
      n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, 
      n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, 
      n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, 
      n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, 
      n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, 
      n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, 
      n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, 
      n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, 
      n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, 
      n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, 
      n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, 
      n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, 
      n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, 
      n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, 
      n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, 
      n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, 
      n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, 
      n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, 
      n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, 
      n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, 
      n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, 
      n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, 
      n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, 
      n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, 
      n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, 
      n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, 
      n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, 
      n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, 
      n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, 
      n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, 
      n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, 
      n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, 
      n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, 
      n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, 
      n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, 
      n_1918, n_1919, n_1920, n_1921 : std_logic;

begin
   
   REGISTERS_reg_1_31_inst : DFFR_X1 port map( D => n4024, CK => CLK, RN => 
                           n378, Q => n603, QN => n_1154);
   REGISTERS_reg_1_30_inst : DFFR_X1 port map( D => n4023, CK => CLK, RN => 
                           n337, Q => n602, QN => n_1155);
   REGISTERS_reg_1_29_inst : DFFR_X1 port map( D => n4022, CK => CLK, RN => 
                           n368, Q => n601, QN => n_1156);
   REGISTERS_reg_1_28_inst : DFFR_X1 port map( D => n4021, CK => CLK, RN => 
                           n367, Q => n600, QN => n_1157);
   REGISTERS_reg_1_27_inst : DFFR_X1 port map( D => n4020, CK => CLK, RN => 
                           n367, Q => n599, QN => n_1158);
   REGISTERS_reg_1_26_inst : DFFR_X1 port map( D => n4019, CK => CLK, RN => 
                           n367, Q => n598, QN => n_1159);
   REGISTERS_reg_1_25_inst : DFFR_X1 port map( D => n4018, CK => CLK, RN => 
                           n367, Q => n597, QN => n_1160);
   REGISTERS_reg_1_24_inst : DFFR_X1 port map( D => n4017, CK => CLK, RN => 
                           n367, Q => n596, QN => n_1161);
   REGISTERS_reg_1_23_inst : DFFR_X1 port map( D => n4016, CK => CLK, RN => 
                           n367, Q => n595, QN => n_1162);
   REGISTERS_reg_1_22_inst : DFFR_X1 port map( D => n4015, CK => CLK, RN => 
                           n367, Q => n594, QN => n_1163);
   REGISTERS_reg_1_21_inst : DFFR_X1 port map( D => n4014, CK => CLK, RN => 
                           n367, Q => n593, QN => n_1164);
   REGISTERS_reg_1_20_inst : DFFR_X1 port map( D => n4013, CK => CLK, RN => 
                           n367, Q => n592, QN => n_1165);
   REGISTERS_reg_1_19_inst : DFFR_X1 port map( D => n4012, CK => CLK, RN => 
                           n367, Q => n591, QN => n_1166);
   REGISTERS_reg_1_18_inst : DFFR_X1 port map( D => n4011, CK => CLK, RN => 
                           n367, Q => n590, QN => n_1167);
   REGISTERS_reg_1_17_inst : DFFR_X1 port map( D => n4010, CK => CLK, RN => 
                           n367, Q => n589, QN => n_1168);
   REGISTERS_reg_1_16_inst : DFFR_X1 port map( D => n4009, CK => CLK, RN => 
                           n366, Q => n588, QN => n_1169);
   REGISTERS_reg_1_15_inst : DFFR_X1 port map( D => n4008, CK => CLK, RN => 
                           n366, Q => n587, QN => n_1170);
   REGISTERS_reg_1_14_inst : DFFR_X1 port map( D => n4007, CK => CLK, RN => 
                           n366, Q => n586, QN => n_1171);
   REGISTERS_reg_1_13_inst : DFFR_X1 port map( D => n4006, CK => CLK, RN => 
                           n366, Q => n585, QN => n_1172);
   REGISTERS_reg_1_12_inst : DFFR_X1 port map( D => n4005, CK => CLK, RN => 
                           n366, Q => n584, QN => n_1173);
   REGISTERS_reg_1_11_inst : DFFR_X1 port map( D => n4004, CK => CLK, RN => 
                           n366, Q => n583, QN => n_1174);
   REGISTERS_reg_1_10_inst : DFFR_X1 port map( D => n4003, CK => CLK, RN => 
                           n366, Q => n582, QN => n_1175);
   REGISTERS_reg_1_9_inst : DFFR_X1 port map( D => n4002, CK => CLK, RN => n366
                           , Q => n581, QN => n_1176);
   REGISTERS_reg_1_8_inst : DFFR_X1 port map( D => n4001, CK => CLK, RN => n366
                           , Q => n580, QN => n_1177);
   REGISTERS_reg_1_7_inst : DFFR_X1 port map( D => n4000, CK => CLK, RN => n366
                           , Q => n579, QN => n_1178);
   REGISTERS_reg_1_6_inst : DFFR_X1 port map( D => n3999, CK => CLK, RN => n366
                           , Q => n578, QN => n_1179);
   REGISTERS_reg_1_5_inst : DFFR_X1 port map( D => n3998, CK => CLK, RN => n366
                           , Q => n577, QN => n_1180);
   REGISTERS_reg_1_4_inst : DFFR_X1 port map( D => n3997, CK => CLK, RN => n365
                           , Q => n576, QN => n_1181);
   REGISTERS_reg_1_3_inst : DFFR_X1 port map( D => n3996, CK => CLK, RN => n365
                           , Q => n575, QN => n_1182);
   REGISTERS_reg_1_2_inst : DFFR_X1 port map( D => n3995, CK => CLK, RN => n365
                           , Q => n574, QN => n_1183);
   REGISTERS_reg_1_1_inst : DFFR_X1 port map( D => n3994, CK => CLK, RN => n365
                           , Q => n573, QN => n_1184);
   REGISTERS_reg_1_0_inst : DFFR_X1 port map( D => n3993, CK => CLK, RN => n365
                           , Q => n571, QN => n_1185);
   REGISTERS_reg_4_31_inst : DFFR_X1 port map( D => n4056, CK => CLK, RN => 
                           n360, Q => n637, QN => n_1186);
   REGISTERS_reg_4_30_inst : DFFR_X1 port map( D => n4055, CK => CLK, RN => 
                           n360, Q => n636, QN => n_1187);
   REGISTERS_reg_4_29_inst : DFFR_X1 port map( D => n4054, CK => CLK, RN => 
                           n359, Q => n635, QN => n_1188);
   REGISTERS_reg_4_28_inst : DFFR_X1 port map( D => n4053, CK => CLK, RN => 
                           n359, Q => n634, QN => n_1189);
   REGISTERS_reg_4_27_inst : DFFR_X1 port map( D => n4052, CK => CLK, RN => 
                           n359, Q => n633, QN => n_1190);
   REGISTERS_reg_4_26_inst : DFFR_X1 port map( D => n4051, CK => CLK, RN => 
                           n359, Q => n632, QN => n_1191);
   REGISTERS_reg_4_25_inst : DFFR_X1 port map( D => n4050, CK => CLK, RN => 
                           n359, Q => n631, QN => n_1192);
   REGISTERS_reg_4_24_inst : DFFR_X1 port map( D => n4049, CK => CLK, RN => 
                           n359, Q => n630, QN => n_1193);
   REGISTERS_reg_4_23_inst : DFFR_X1 port map( D => n4048, CK => CLK, RN => 
                           n359, Q => n629, QN => n_1194);
   REGISTERS_reg_4_22_inst : DFFR_X1 port map( D => n4047, CK => CLK, RN => 
                           n359, Q => n628, QN => n_1195);
   REGISTERS_reg_4_21_inst : DFFR_X1 port map( D => n4046, CK => CLK, RN => 
                           n359, Q => n627, QN => n_1196);
   REGISTERS_reg_4_20_inst : DFFR_X1 port map( D => n4045, CK => CLK, RN => 
                           n359, Q => n626, QN => n_1197);
   REGISTERS_reg_4_19_inst : DFFR_X1 port map( D => n4044, CK => CLK, RN => 
                           n359, Q => n625, QN => n_1198);
   REGISTERS_reg_4_18_inst : DFFR_X1 port map( D => n4043, CK => CLK, RN => 
                           n359, Q => n624, QN => n_1199);
   REGISTERS_reg_4_17_inst : DFFR_X1 port map( D => n4042, CK => CLK, RN => 
                           n358, Q => n623, QN => n_1200);
   REGISTERS_reg_4_16_inst : DFFR_X1 port map( D => n4041, CK => CLK, RN => 
                           n358, Q => n622, QN => n_1201);
   REGISTERS_reg_4_15_inst : DFFR_X1 port map( D => n4040, CK => CLK, RN => 
                           n358, Q => n621, QN => n_1202);
   REGISTERS_reg_4_14_inst : DFFR_X1 port map( D => n4039, CK => CLK, RN => 
                           n358, Q => n620, QN => n_1203);
   REGISTERS_reg_4_13_inst : DFFR_X1 port map( D => n4038, CK => CLK, RN => 
                           n358, Q => n619, QN => n_1204);
   REGISTERS_reg_4_12_inst : DFFR_X1 port map( D => n4037, CK => CLK, RN => 
                           n358, Q => n618, QN => n_1205);
   REGISTERS_reg_4_11_inst : DFFR_X1 port map( D => n4036, CK => CLK, RN => 
                           n358, Q => n617, QN => n_1206);
   REGISTERS_reg_4_10_inst : DFFR_X1 port map( D => n4035, CK => CLK, RN => 
                           n358, Q => n616, QN => n_1207);
   REGISTERS_reg_4_9_inst : DFFR_X1 port map( D => n4034, CK => CLK, RN => n358
                           , Q => n615, QN => n_1208);
   REGISTERS_reg_4_8_inst : DFFR_X1 port map( D => n4033, CK => CLK, RN => n358
                           , Q => n614, QN => n_1209);
   REGISTERS_reg_4_7_inst : DFFR_X1 port map( D => n4032, CK => CLK, RN => n358
                           , Q => n613, QN => n_1210);
   REGISTERS_reg_4_6_inst : DFFR_X1 port map( D => n4031, CK => CLK, RN => n358
                           , Q => n612, QN => n_1211);
   REGISTERS_reg_4_5_inst : DFFR_X1 port map( D => n4030, CK => CLK, RN => n357
                           , Q => n611, QN => n_1212);
   REGISTERS_reg_4_4_inst : DFFR_X1 port map( D => n4029, CK => CLK, RN => n357
                           , Q => n610, QN => n_1213);
   REGISTERS_reg_4_3_inst : DFFR_X1 port map( D => n4028, CK => CLK, RN => n357
                           , Q => n609, QN => n_1214);
   REGISTERS_reg_4_2_inst : DFFR_X1 port map( D => n4027, CK => CLK, RN => n362
                           , Q => n608, QN => n_1215);
   REGISTERS_reg_4_1_inst : DFFR_X1 port map( D => n4026, CK => CLK, RN => n378
                           , Q => n607, QN => n_1216);
   REGISTERS_reg_4_0_inst : DFFR_X1 port map( D => n4025, CK => CLK, RN => n378
                           , Q => n605, QN => n_1217);
   REGISTERS_reg_5_31_inst : DFFR_X1 port map( D => n4088, CK => CLK, RN => 
                           n378, Q => n670, QN => n_1218);
   REGISTERS_reg_5_30_inst : DFFR_X1 port map( D => n4087, CK => CLK, RN => 
                           n378, Q => n669, QN => n_1219);
   REGISTERS_reg_5_29_inst : DFFR_X1 port map( D => n4086, CK => CLK, RN => 
                           n377, Q => n668, QN => n_1220);
   REGISTERS_reg_5_28_inst : DFFR_X1 port map( D => n4085, CK => CLK, RN => 
                           n377, Q => n667, QN => n_1221);
   REGISTERS_reg_5_27_inst : DFFR_X1 port map( D => n4084, CK => CLK, RN => 
                           n377, Q => n666, QN => n_1222);
   REGISTERS_reg_5_26_inst : DFFR_X1 port map( D => n4083, CK => CLK, RN => 
                           n377, Q => n665, QN => n_1223);
   REGISTERS_reg_5_25_inst : DFFR_X1 port map( D => n4082, CK => CLK, RN => 
                           n377, Q => n664, QN => n_1224);
   REGISTERS_reg_5_24_inst : DFFR_X1 port map( D => n4081, CK => CLK, RN => 
                           n377, Q => n663, QN => n_1225);
   REGISTERS_reg_5_23_inst : DFFR_X1 port map( D => n4080, CK => CLK, RN => 
                           n377, Q => n662, QN => n_1226);
   REGISTERS_reg_5_22_inst : DFFR_X1 port map( D => n4079, CK => CLK, RN => 
                           n377, Q => n661, QN => n_1227);
   REGISTERS_reg_5_21_inst : DFFR_X1 port map( D => n4078, CK => CLK, RN => 
                           n377, Q => n660, QN => n_1228);
   REGISTERS_reg_5_20_inst : DFFR_X1 port map( D => n4077, CK => CLK, RN => 
                           n377, Q => n659, QN => n_1229);
   REGISTERS_reg_5_19_inst : DFFR_X1 port map( D => n4076, CK => CLK, RN => 
                           n377, Q => n658, QN => n_1230);
   REGISTERS_reg_5_18_inst : DFFR_X1 port map( D => n4075, CK => CLK, RN => 
                           n377, Q => n657, QN => n_1231);
   REGISTERS_reg_5_17_inst : DFFR_X1 port map( D => n4074, CK => CLK, RN => 
                           n376, Q => n656, QN => n_1232);
   REGISTERS_reg_5_16_inst : DFFR_X1 port map( D => n4073, CK => CLK, RN => 
                           n376, Q => n655, QN => n_1233);
   REGISTERS_reg_5_15_inst : DFFR_X1 port map( D => n4072, CK => CLK, RN => 
                           n376, Q => n654, QN => n_1234);
   REGISTERS_reg_5_14_inst : DFFR_X1 port map( D => n4071, CK => CLK, RN => 
                           n376, Q => n653, QN => n_1235);
   REGISTERS_reg_5_13_inst : DFFR_X1 port map( D => n4070, CK => CLK, RN => 
                           n376, Q => n652, QN => n_1236);
   REGISTERS_reg_5_12_inst : DFFR_X1 port map( D => n4069, CK => CLK, RN => 
                           n376, Q => n651, QN => n_1237);
   REGISTERS_reg_5_11_inst : DFFR_X1 port map( D => n4068, CK => CLK, RN => 
                           n376, Q => n650, QN => n_1238);
   REGISTERS_reg_5_10_inst : DFFR_X1 port map( D => n4067, CK => CLK, RN => 
                           n376, Q => n649, QN => n_1239);
   REGISTERS_reg_5_9_inst : DFFR_X1 port map( D => n4066, CK => CLK, RN => n376
                           , Q => n648, QN => n_1240);
   REGISTERS_reg_5_8_inst : DFFR_X1 port map( D => n4065, CK => CLK, RN => n376
                           , Q => n647, QN => n_1241);
   REGISTERS_reg_5_7_inst : DFFR_X1 port map( D => n4064, CK => CLK, RN => n376
                           , Q => n646, QN => n_1242);
   REGISTERS_reg_5_6_inst : DFFR_X1 port map( D => n4063, CK => CLK, RN => n376
                           , Q => n645, QN => n_1243);
   REGISTERS_reg_5_5_inst : DFFR_X1 port map( D => n4062, CK => CLK, RN => n375
                           , Q => n644, QN => n_1244);
   REGISTERS_reg_5_4_inst : DFFR_X1 port map( D => n4061, CK => CLK, RN => n375
                           , Q => n643, QN => n_1245);
   REGISTERS_reg_5_3_inst : DFFR_X1 port map( D => n4060, CK => CLK, RN => n375
                           , Q => n642, QN => n_1246);
   REGISTERS_reg_5_2_inst : DFFR_X1 port map( D => n4059, CK => CLK, RN => n375
                           , Q => n641, QN => n_1247);
   REGISTERS_reg_5_1_inst : DFFR_X1 port map( D => n4058, CK => CLK, RN => n375
                           , Q => n640, QN => n_1248);
   REGISTERS_reg_5_0_inst : DFFR_X1 port map( D => n4057, CK => CLK, RN => n375
                           , Q => n638, QN => n_1249);
   REGISTERS_reg_8_31_inst : DFFR_X1 port map( D => n3896, CK => CLK, RN => 
                           n370, Q => n_1250, QN => n2494);
   REGISTERS_reg_8_30_inst : DFFR_X1 port map( D => n3895, CK => CLK, RN => 
                           n369, Q => n_1251, QN => n2515);
   REGISTERS_reg_8_29_inst : DFFR_X1 port map( D => n3894, CK => CLK, RN => 
                           n369, Q => n_1252, QN => n2536);
   REGISTERS_reg_8_28_inst : DFFR_X1 port map( D => n3893, CK => CLK, RN => 
                           n369, Q => n_1253, QN => n2557);
   REGISTERS_reg_8_27_inst : DFFR_X1 port map( D => n3892, CK => CLK, RN => 
                           n369, Q => n_1254, QN => n2578);
   REGISTERS_reg_8_26_inst : DFFR_X1 port map( D => n3891, CK => CLK, RN => 
                           n369, Q => n_1255, QN => n2599);
   REGISTERS_reg_8_25_inst : DFFR_X1 port map( D => n3890, CK => CLK, RN => 
                           n369, Q => n_1256, QN => n2620);
   REGISTERS_reg_8_24_inst : DFFR_X1 port map( D => n3889, CK => CLK, RN => 
                           n369, Q => n_1257, QN => n2641);
   REGISTERS_reg_8_23_inst : DFFR_X1 port map( D => n3888, CK => CLK, RN => 
                           n369, Q => n_1258, QN => n2662);
   REGISTERS_reg_8_22_inst : DFFR_X1 port map( D => n3887, CK => CLK, RN => 
                           n369, Q => n_1259, QN => n2683);
   REGISTERS_reg_8_21_inst : DFFR_X1 port map( D => n3886, CK => CLK, RN => 
                           n369, Q => n_1260, QN => n2704);
   REGISTERS_reg_8_20_inst : DFFR_X1 port map( D => n3885, CK => CLK, RN => 
                           n369, Q => n_1261, QN => n2725);
   REGISTERS_reg_8_19_inst : DFFR_X1 port map( D => n3884, CK => CLK, RN => 
                           n369, Q => n_1262, QN => n2746);
   REGISTERS_reg_8_18_inst : DFFR_X1 port map( D => n3883, CK => CLK, RN => 
                           n368, Q => n_1263, QN => n2767);
   REGISTERS_reg_8_17_inst : DFFR_X1 port map( D => n3882, CK => CLK, RN => 
                           n368, Q => n_1264, QN => n2788);
   REGISTERS_reg_8_16_inst : DFFR_X1 port map( D => n3881, CK => CLK, RN => 
                           n368, Q => n_1265, QN => n2809);
   REGISTERS_reg_8_15_inst : DFFR_X1 port map( D => n3880, CK => CLK, RN => 
                           n368, Q => n_1266, QN => n2830);
   REGISTERS_reg_8_14_inst : DFFR_X1 port map( D => n3879, CK => CLK, RN => 
                           n368, Q => n_1267, QN => n2851);
   REGISTERS_reg_8_13_inst : DFFR_X1 port map( D => n3878, CK => CLK, RN => 
                           n368, Q => n_1268, QN => n2872);
   REGISTERS_reg_8_12_inst : DFFR_X1 port map( D => n3877, CK => CLK, RN => 
                           n368, Q => n_1269, QN => n2893);
   REGISTERS_reg_8_11_inst : DFFR_X1 port map( D => n3876, CK => CLK, RN => 
                           n368, Q => n_1270, QN => n2914);
   REGISTERS_reg_8_10_inst : DFFR_X1 port map( D => n3875, CK => CLK, RN => 
                           n368, Q => n_1271, QN => n2935);
   REGISTERS_reg_8_9_inst : DFFR_X1 port map( D => n3874, CK => CLK, RN => n368
                           , Q => n_1272, QN => n2956);
   REGISTERS_reg_8_8_inst : DFFR_X1 port map( D => n3873, CK => CLK, RN => n368
                           , Q => n_1273, QN => n2977);
   REGISTERS_reg_8_7_inst : DFFR_X1 port map( D => n3872, CK => CLK, RN => n373
                           , Q => n_1274, QN => n3574);
   REGISTERS_reg_8_6_inst : DFFR_X1 port map( D => n3871, CK => CLK, RN => n347
                           , Q => n_1275, QN => n3595);
   REGISTERS_reg_8_5_inst : DFFR_X1 port map( D => n3870, CK => CLK, RN => n347
                           , Q => n_1276, QN => n3616);
   REGISTERS_reg_8_4_inst : DFFR_X1 port map( D => n3869, CK => CLK, RN => n347
                           , Q => n_1277, QN => n3637);
   REGISTERS_reg_8_3_inst : DFFR_X1 port map( D => n3868, CK => CLK, RN => n347
                           , Q => n_1278, QN => n3658);
   REGISTERS_reg_8_2_inst : DFFR_X1 port map( D => n3867, CK => CLK, RN => n347
                           , Q => n_1279, QN => n3679);
   REGISTERS_reg_8_1_inst : DFFR_X1 port map( D => n3866, CK => CLK, RN => n346
                           , Q => n_1280, QN => n3700);
   REGISTERS_reg_8_0_inst : DFFR_X1 port map( D => n3865, CK => CLK, RN => n346
                           , Q => n_1281, QN => n3721);
   REGISTERS_reg_9_31_inst : DFFR_X1 port map( D => n3928, CK => CLK, RN => 
                           n346, Q => n_1282, QN => n2495);
   REGISTERS_reg_9_30_inst : DFFR_X1 port map( D => n3927, CK => CLK, RN => 
                           n346, Q => n_1283, QN => n2516);
   REGISTERS_reg_9_29_inst : DFFR_X1 port map( D => n3926, CK => CLK, RN => 
                           n346, Q => n_1284, QN => n2537);
   REGISTERS_reg_9_28_inst : DFFR_X1 port map( D => n3925, CK => CLK, RN => 
                           n346, Q => n_1285, QN => n2558);
   REGISTERS_reg_9_27_inst : DFFR_X1 port map( D => n3924, CK => CLK, RN => 
                           n346, Q => n_1286, QN => n2579);
   REGISTERS_reg_9_26_inst : DFFR_X1 port map( D => n3923, CK => CLK, RN => 
                           n346, Q => n_1287, QN => n2600);
   REGISTERS_reg_9_25_inst : DFFR_X1 port map( D => n3922, CK => CLK, RN => 
                           n346, Q => n_1288, QN => n2621);
   REGISTERS_reg_9_24_inst : DFFR_X1 port map( D => n3921, CK => CLK, RN => 
                           n346, Q => n_1289, QN => n2642);
   REGISTERS_reg_9_23_inst : DFFR_X1 port map( D => n3920, CK => CLK, RN => 
                           n346, Q => n_1290, QN => n2663);
   REGISTERS_reg_9_22_inst : DFFR_X1 port map( D => n3919, CK => CLK, RN => 
                           n346, Q => n_1291, QN => n2684);
   REGISTERS_reg_9_21_inst : DFFR_X1 port map( D => n3918, CK => CLK, RN => 
                           n345, Q => n_1292, QN => n2705);
   REGISTERS_reg_9_20_inst : DFFR_X1 port map( D => n3917, CK => CLK, RN => 
                           n345, Q => n_1293, QN => n2726);
   REGISTERS_reg_9_19_inst : DFFR_X1 port map( D => n3916, CK => CLK, RN => 
                           n345, Q => n_1294, QN => n2747);
   REGISTERS_reg_9_18_inst : DFFR_X1 port map( D => n3915, CK => CLK, RN => 
                           n345, Q => n_1295, QN => n2768);
   REGISTERS_reg_9_17_inst : DFFR_X1 port map( D => n3914, CK => CLK, RN => 
                           n345, Q => n_1296, QN => n2789);
   REGISTERS_reg_9_16_inst : DFFR_X1 port map( D => n3913, CK => CLK, RN => 
                           n345, Q => n_1297, QN => n2810);
   REGISTERS_reg_9_15_inst : DFFR_X1 port map( D => n3912, CK => CLK, RN => 
                           n345, Q => n_1298, QN => n2831);
   REGISTERS_reg_9_14_inst : DFFR_X1 port map( D => n3911, CK => CLK, RN => 
                           n345, Q => n_1299, QN => n2852);
   REGISTERS_reg_9_13_inst : DFFR_X1 port map( D => n3910, CK => CLK, RN => 
                           n345, Q => n_1300, QN => n2873);
   REGISTERS_reg_9_12_inst : DFFR_X1 port map( D => n3909, CK => CLK, RN => 
                           n345, Q => n_1301, QN => n2894);
   REGISTERS_reg_9_11_inst : DFFR_X1 port map( D => n3908, CK => CLK, RN => 
                           n345, Q => n_1302, QN => n2915);
   REGISTERS_reg_9_10_inst : DFFR_X1 port map( D => n3907, CK => CLK, RN => 
                           n345, Q => n_1303, QN => n2936);
   REGISTERS_reg_9_9_inst : DFFR_X1 port map( D => n3906, CK => CLK, RN => n344
                           , Q => n_1304, QN => n2957);
   REGISTERS_reg_9_8_inst : DFFR_X1 port map( D => n3905, CK => CLK, RN => n344
                           , Q => n_1305, QN => n2978);
   REGISTERS_reg_9_7_inst : DFFR_X1 port map( D => n3904, CK => CLK, RN => n344
                           , Q => n_1306, QN => n3575);
   REGISTERS_reg_9_6_inst : DFFR_X1 port map( D => n3903, CK => CLK, RN => n344
                           , Q => n_1307, QN => n3596);
   REGISTERS_reg_9_5_inst : DFFR_X1 port map( D => n3902, CK => CLK, RN => n344
                           , Q => n_1308, QN => n3617);
   REGISTERS_reg_9_4_inst : DFFR_X1 port map( D => n3901, CK => CLK, RN => n344
                           , Q => n_1309, QN => n3638);
   REGISTERS_reg_9_3_inst : DFFR_X1 port map( D => n3900, CK => CLK, RN => n344
                           , Q => n_1310, QN => n3659);
   REGISTERS_reg_9_2_inst : DFFR_X1 port map( D => n3899, CK => CLK, RN => n344
                           , Q => n_1311, QN => n3680);
   REGISTERS_reg_9_1_inst : DFFR_X1 port map( D => n3898, CK => CLK, RN => n344
                           , Q => n_1312, QN => n3701);
   REGISTERS_reg_9_0_inst : DFFR_X1 port map( D => n3897, CK => CLK, RN => n344
                           , Q => n_1313, QN => n3722);
   REGISTERS_reg_10_31_inst : DFFR_X1 port map( D => n3430, CK => CLK, RN => 
                           n344, Q => n2497, QN => n_1314);
   REGISTERS_reg_10_30_inst : DFFR_X1 port map( D => n3429, CK => CLK, RN => 
                           n344, Q => n2518, QN => n_1315);
   REGISTERS_reg_10_29_inst : DFFR_X1 port map( D => n3428, CK => CLK, RN => 
                           n343, Q => n2539, QN => n_1316);
   REGISTERS_reg_10_28_inst : DFFR_X1 port map( D => n3427, CK => CLK, RN => 
                           n343, Q => n2560, QN => n_1317);
   REGISTERS_reg_10_27_inst : DFFR_X1 port map( D => n3426, CK => CLK, RN => 
                           n343, Q => n2581, QN => n_1318);
   REGISTERS_reg_10_26_inst : DFFR_X1 port map( D => n3425, CK => CLK, RN => 
                           n343, Q => n2602, QN => n_1319);
   REGISTERS_reg_10_25_inst : DFFR_X1 port map( D => n3424, CK => CLK, RN => 
                           n343, Q => n2623, QN => n_1320);
   REGISTERS_reg_10_24_inst : DFFR_X1 port map( D => n3423, CK => CLK, RN => 
                           n343, Q => n2644, QN => n_1321);
   REGISTERS_reg_10_23_inst : DFFR_X1 port map( D => n3422, CK => CLK, RN => 
                           n343, Q => n2665, QN => n_1322);
   REGISTERS_reg_10_22_inst : DFFR_X1 port map( D => n3421, CK => CLK, RN => 
                           n343, Q => n2686, QN => n_1323);
   REGISTERS_reg_10_21_inst : DFFR_X1 port map( D => n3420, CK => CLK, RN => 
                           n343, Q => n2707, QN => n_1324);
   REGISTERS_reg_10_20_inst : DFFR_X1 port map( D => n3419, CK => CLK, RN => 
                           n343, Q => n2728, QN => n_1325);
   REGISTERS_reg_10_19_inst : DFFR_X1 port map( D => n3418, CK => CLK, RN => 
                           n343, Q => n2749, QN => n_1326);
   REGISTERS_reg_10_18_inst : DFFR_X1 port map( D => n3417, CK => CLK, RN => 
                           n343, Q => n2770, QN => n_1327);
   REGISTERS_reg_10_17_inst : DFFR_X1 port map( D => n3416, CK => CLK, RN => 
                           n342, Q => n2791, QN => n_1328);
   REGISTERS_reg_10_16_inst : DFFR_X1 port map( D => n3415, CK => CLK, RN => 
                           n342, Q => n2812, QN => n_1329);
   REGISTERS_reg_10_15_inst : DFFR_X1 port map( D => n3414, CK => CLK, RN => 
                           n342, Q => n2833, QN => n_1330);
   REGISTERS_reg_10_14_inst : DFFR_X1 port map( D => n3413, CK => CLK, RN => 
                           n342, Q => n2854, QN => n_1331);
   REGISTERS_reg_10_13_inst : DFFR_X1 port map( D => n3412, CK => CLK, RN => 
                           n342, Q => n2875, QN => n_1332);
   REGISTERS_reg_10_12_inst : DFFR_X1 port map( D => n3411, CK => CLK, RN => 
                           n342, Q => n2896, QN => n_1333);
   REGISTERS_reg_10_11_inst : DFFR_X1 port map( D => n3410, CK => CLK, RN => 
                           n342, Q => n2917, QN => n_1334);
   REGISTERS_reg_10_10_inst : DFFR_X1 port map( D => n3409, CK => CLK, RN => 
                           n342, Q => n2938, QN => n_1335);
   REGISTERS_reg_10_9_inst : DFFR_X1 port map( D => n3408, CK => CLK, RN => 
                           n342, Q => n2959, QN => n_1336);
   REGISTERS_reg_10_8_inst : DFFR_X1 port map( D => n3407, CK => CLK, RN => 
                           n342, Q => n2980, QN => n_1337);
   REGISTERS_reg_10_7_inst : DFFR_X1 port map( D => n3406, CK => CLK, RN => 
                           n342, Q => n3577, QN => n_1338);
   REGISTERS_reg_10_6_inst : DFFR_X1 port map( D => n3405, CK => CLK, RN => 
                           n341, Q => n3598, QN => n_1339);
   REGISTERS_reg_10_5_inst : DFFR_X1 port map( D => n3404, CK => CLK, RN => 
                           n341, Q => n3619, QN => n_1340);
   REGISTERS_reg_10_4_inst : DFFR_X1 port map( D => n3403, CK => CLK, RN => 
                           n341, Q => n3640, QN => n_1341);
   REGISTERS_reg_10_3_inst : DFFR_X1 port map( D => n3402, CK => CLK, RN => 
                           n341, Q => n3661, QN => n_1342);
   REGISTERS_reg_10_2_inst : DFFR_X1 port map( D => n3401, CK => CLK, RN => 
                           n341, Q => n3682, QN => n_1343);
   REGISTERS_reg_10_1_inst : DFFR_X1 port map( D => n3400, CK => CLK, RN => 
                           n341, Q => n3703, QN => n_1344);
   REGISTERS_reg_10_0_inst : DFFR_X1 port map( D => n3399, CK => CLK, RN => 
                           n341, Q => n3724, QN => n_1345);
   REGISTERS_reg_11_31_inst : DFFR_X1 port map( D => n3398, CK => CLK, RN => 
                           n341, Q => n2496, QN => n_1346);
   REGISTERS_reg_11_30_inst : DFFR_X1 port map( D => n3397, CK => CLK, RN => 
                           n341, Q => n2517, QN => n_1347);
   REGISTERS_reg_11_29_inst : DFFR_X1 port map( D => n3396, CK => CLK, RN => 
                           n341, Q => n2538, QN => n_1348);
   REGISTERS_reg_11_28_inst : DFFR_X1 port map( D => n3395, CK => CLK, RN => 
                           n341, Q => n2559, QN => n_1349);
   REGISTERS_reg_11_27_inst : DFFR_X1 port map( D => n3394, CK => CLK, RN => 
                           n341, Q => n2580, QN => n_1350);
   REGISTERS_reg_11_26_inst : DFFR_X1 port map( D => n3393, CK => CLK, RN => 
                           n340, Q => n2601, QN => n_1351);
   REGISTERS_reg_11_25_inst : DFFR_X1 port map( D => n3392, CK => CLK, RN => 
                           n340, Q => n2622, QN => n_1352);
   REGISTERS_reg_11_24_inst : DFFR_X1 port map( D => n3391, CK => CLK, RN => 
                           n340, Q => n2643, QN => n_1353);
   REGISTERS_reg_11_23_inst : DFFR_X1 port map( D => n3390, CK => CLK, RN => 
                           n340, Q => n2664, QN => n_1354);
   REGISTERS_reg_11_22_inst : DFFR_X1 port map( D => n3389, CK => CLK, RN => 
                           n340, Q => n2685, QN => n_1355);
   REGISTERS_reg_11_21_inst : DFFR_X1 port map( D => n3388, CK => CLK, RN => 
                           n340, Q => n2706, QN => n_1356);
   REGISTERS_reg_11_20_inst : DFFR_X1 port map( D => n3387, CK => CLK, RN => 
                           n340, Q => n2727, QN => n_1357);
   REGISTERS_reg_11_19_inst : DFFR_X1 port map( D => n3386, CK => CLK, RN => 
                           n340, Q => n2748, QN => n_1358);
   REGISTERS_reg_11_18_inst : DFFR_X1 port map( D => n3385, CK => CLK, RN => 
                           n340, Q => n2769, QN => n_1359);
   REGISTERS_reg_11_17_inst : DFFR_X1 port map( D => n3384, CK => CLK, RN => 
                           n340, Q => n2790, QN => n_1360);
   REGISTERS_reg_11_16_inst : DFFR_X1 port map( D => n3383, CK => CLK, RN => 
                           n340, Q => n2811, QN => n_1361);
   REGISTERS_reg_11_15_inst : DFFR_X1 port map( D => n3382, CK => CLK, RN => 
                           n340, Q => n2832, QN => n_1362);
   REGISTERS_reg_11_14_inst : DFFR_X1 port map( D => n3381, CK => CLK, RN => 
                           n339, Q => n2853, QN => n_1363);
   REGISTERS_reg_11_13_inst : DFFR_X1 port map( D => n3380, CK => CLK, RN => 
                           n339, Q => n2874, QN => n_1364);
   REGISTERS_reg_11_12_inst : DFFR_X1 port map( D => n3379, CK => CLK, RN => 
                           n339, Q => n2895, QN => n_1365);
   REGISTERS_reg_11_11_inst : DFFR_X1 port map( D => n3378, CK => CLK, RN => 
                           n339, Q => n2916, QN => n_1366);
   REGISTERS_reg_11_10_inst : DFFR_X1 port map( D => n3377, CK => CLK, RN => 
                           n339, Q => n2937, QN => n_1367);
   REGISTERS_reg_11_9_inst : DFFR_X1 port map( D => n3376, CK => CLK, RN => 
                           n339, Q => n2958, QN => n_1368);
   REGISTERS_reg_11_8_inst : DFFR_X1 port map( D => n3375, CK => CLK, RN => 
                           n339, Q => n2979, QN => n_1369);
   REGISTERS_reg_11_7_inst : DFFR_X1 port map( D => n3374, CK => CLK, RN => 
                           n339, Q => n3576, QN => n_1370);
   REGISTERS_reg_11_6_inst : DFFR_X1 port map( D => n3373, CK => CLK, RN => 
                           n339, Q => n3597, QN => n_1371);
   REGISTERS_reg_11_5_inst : DFFR_X1 port map( D => n3372, CK => CLK, RN => 
                           n339, Q => n3618, QN => n_1372);
   REGISTERS_reg_11_4_inst : DFFR_X1 port map( D => n3371, CK => CLK, RN => 
                           n339, Q => n3639, QN => n_1373);
   REGISTERS_reg_11_3_inst : DFFR_X1 port map( D => n3370, CK => CLK, RN => 
                           n339, Q => n3660, QN => n_1374);
   REGISTERS_reg_11_2_inst : DFFR_X1 port map( D => n3369, CK => CLK, RN => 
                           n338, Q => n3681, QN => n_1375);
   REGISTERS_reg_11_1_inst : DFFR_X1 port map( D => n3368, CK => CLK, RN => 
                           n338, Q => n3702, QN => n_1376);
   REGISTERS_reg_11_0_inst : DFFR_X1 port map( D => n3367, CK => CLK, RN => 
                           n338, Q => n3723, QN => n_1377);
   REGISTERS_reg_12_31_inst : DFFR_X1 port map( D => n3960, CK => CLK, RN => 
                           n338, Q => n_1378, QN => n2490);
   REGISTERS_reg_12_30_inst : DFFR_X1 port map( D => n3959, CK => CLK, RN => 
                           n338, Q => n_1379, QN => n2511);
   REGISTERS_reg_12_29_inst : DFFR_X1 port map( D => n3958, CK => CLK, RN => 
                           n338, Q => n_1380, QN => n2532);
   REGISTERS_reg_12_28_inst : DFFR_X1 port map( D => n3957, CK => CLK, RN => 
                           n338, Q => n_1381, QN => n2553);
   REGISTERS_reg_12_27_inst : DFFR_X1 port map( D => n3956, CK => CLK, RN => 
                           n338, Q => n_1382, QN => n2574);
   REGISTERS_reg_12_26_inst : DFFR_X1 port map( D => n3955, CK => CLK, RN => 
                           n338, Q => n_1383, QN => n2595);
   REGISTERS_reg_12_25_inst : DFFR_X1 port map( D => n3954, CK => CLK, RN => 
                           n338, Q => n_1384, QN => n2616);
   REGISTERS_reg_12_24_inst : DFFR_X1 port map( D => n3953, CK => CLK, RN => 
                           n338, Q => n_1385, QN => n2637);
   REGISTERS_reg_12_23_inst : DFFR_X1 port map( D => n3952, CK => CLK, RN => 
                           n338, Q => n_1386, QN => n2658);
   REGISTERS_reg_12_22_inst : DFFR_X1 port map( D => n3951, CK => CLK, RN => 
                           n337, Q => n_1387, QN => n2679);
   REGISTERS_reg_12_21_inst : DFFR_X1 port map( D => n3950, CK => CLK, RN => 
                           n337, Q => n_1388, QN => n2700);
   REGISTERS_reg_12_20_inst : DFFR_X1 port map( D => n3949, CK => CLK, RN => 
                           n337, Q => n_1389, QN => n2721);
   REGISTERS_reg_12_19_inst : DFFR_X1 port map( D => n3948, CK => CLK, RN => 
                           n337, Q => n_1390, QN => n2742);
   REGISTERS_reg_12_18_inst : DFFR_X1 port map( D => n3947, CK => CLK, RN => 
                           n337, Q => n_1391, QN => n2763);
   REGISTERS_reg_12_17_inst : DFFR_X1 port map( D => n3946, CK => CLK, RN => 
                           n337, Q => n_1392, QN => n2784);
   REGISTERS_reg_12_16_inst : DFFR_X1 port map( D => n3945, CK => CLK, RN => 
                           n337, Q => n_1393, QN => n2805);
   REGISTERS_reg_12_15_inst : DFFR_X1 port map( D => n3944, CK => CLK, RN => 
                           n337, Q => n_1394, QN => n2826);
   REGISTERS_reg_12_14_inst : DFFR_X1 port map( D => n3943, CK => CLK, RN => 
                           n337, Q => n_1395, QN => n2847);
   REGISTERS_reg_12_13_inst : DFFR_X1 port map( D => n3942, CK => CLK, RN => 
                           n337, Q => n_1396, QN => n2868);
   REGISTERS_reg_12_12_inst : DFFR_X1 port map( D => n3941, CK => CLK, RN => 
                           n337, Q => n_1397, QN => n2889);
   REGISTERS_reg_12_11_inst : DFFR_X1 port map( D => n3940, CK => CLK, RN => 
                           n342, Q => n_1398, QN => n2910);
   REGISTERS_reg_12_10_inst : DFFR_X1 port map( D => n3939, CK => CLK, RN => 
                           n357, Q => n_1399, QN => n2931);
   REGISTERS_reg_12_9_inst : DFFR_X1 port map( D => n3938, CK => CLK, RN => 
                           n357, Q => n_1400, QN => n2952);
   REGISTERS_reg_12_8_inst : DFFR_X1 port map( D => n3937, CK => CLK, RN => 
                           n357, Q => n_1401, QN => n2973);
   REGISTERS_reg_12_7_inst : DFFR_X1 port map( D => n3936, CK => CLK, RN => 
                           n357, Q => n_1402, QN => n3570);
   REGISTERS_reg_12_6_inst : DFFR_X1 port map( D => n3935, CK => CLK, RN => 
                           n357, Q => n_1403, QN => n3591);
   REGISTERS_reg_12_5_inst : DFFR_X1 port map( D => n3934, CK => CLK, RN => 
                           n357, Q => n_1404, QN => n3612);
   REGISTERS_reg_12_4_inst : DFFR_X1 port map( D => n3933, CK => CLK, RN => 
                           n357, Q => n_1405, QN => n3633);
   REGISTERS_reg_12_3_inst : DFFR_X1 port map( D => n3932, CK => CLK, RN => 
                           n357, Q => n_1406, QN => n3654);
   REGISTERS_reg_12_2_inst : DFFR_X1 port map( D => n3931, CK => CLK, RN => 
                           n356, Q => n_1407, QN => n3675);
   REGISTERS_reg_12_1_inst : DFFR_X1 port map( D => n3930, CK => CLK, RN => 
                           n356, Q => n_1408, QN => n3696);
   REGISTERS_reg_12_0_inst : DFFR_X1 port map( D => n3929, CK => CLK, RN => 
                           n356, Q => n_1409, QN => n3717);
   REGISTERS_reg_13_31_inst : DFFR_X1 port map( D => n3992, CK => CLK, RN => 
                           n356, Q => n_1410, QN => n2491);
   REGISTERS_reg_13_30_inst : DFFR_X1 port map( D => n3991, CK => CLK, RN => 
                           n356, Q => n_1411, QN => n2512);
   REGISTERS_reg_13_29_inst : DFFR_X1 port map( D => n3990, CK => CLK, RN => 
                           n356, Q => n_1412, QN => n2533);
   REGISTERS_reg_13_28_inst : DFFR_X1 port map( D => n3989, CK => CLK, RN => 
                           n356, Q => n_1413, QN => n2554);
   REGISTERS_reg_13_27_inst : DFFR_X1 port map( D => n3988, CK => CLK, RN => 
                           n356, Q => n_1414, QN => n2575);
   REGISTERS_reg_13_26_inst : DFFR_X1 port map( D => n3987, CK => CLK, RN => 
                           n356, Q => n_1415, QN => n2596);
   REGISTERS_reg_13_25_inst : DFFR_X1 port map( D => n3986, CK => CLK, RN => 
                           n356, Q => n_1416, QN => n2617);
   REGISTERS_reg_13_24_inst : DFFR_X1 port map( D => n3985, CK => CLK, RN => 
                           n356, Q => n_1417, QN => n2638);
   REGISTERS_reg_13_23_inst : DFFR_X1 port map( D => n3984, CK => CLK, RN => 
                           n356, Q => n_1418, QN => n2659);
   REGISTERS_reg_13_22_inst : DFFR_X1 port map( D => n3983, CK => CLK, RN => 
                           n355, Q => n_1419, QN => n2680);
   REGISTERS_reg_13_21_inst : DFFR_X1 port map( D => n3982, CK => CLK, RN => 
                           n355, Q => n_1420, QN => n2701);
   REGISTERS_reg_13_20_inst : DFFR_X1 port map( D => n3981, CK => CLK, RN => 
                           n355, Q => n_1421, QN => n2722);
   REGISTERS_reg_13_19_inst : DFFR_X1 port map( D => n3980, CK => CLK, RN => 
                           n355, Q => n_1422, QN => n2743);
   REGISTERS_reg_13_18_inst : DFFR_X1 port map( D => n3979, CK => CLK, RN => 
                           n355, Q => n_1423, QN => n2764);
   REGISTERS_reg_13_17_inst : DFFR_X1 port map( D => n3978, CK => CLK, RN => 
                           n355, Q => n_1424, QN => n2785);
   REGISTERS_reg_13_16_inst : DFFR_X1 port map( D => n3977, CK => CLK, RN => 
                           n355, Q => n_1425, QN => n2806);
   REGISTERS_reg_13_15_inst : DFFR_X1 port map( D => n3976, CK => CLK, RN => 
                           n355, Q => n_1426, QN => n2827);
   REGISTERS_reg_13_14_inst : DFFR_X1 port map( D => n3975, CK => CLK, RN => 
                           n355, Q => n_1427, QN => n2848);
   REGISTERS_reg_13_13_inst : DFFR_X1 port map( D => n3974, CK => CLK, RN => 
                           n355, Q => n_1428, QN => n2869);
   REGISTERS_reg_13_12_inst : DFFR_X1 port map( D => n3973, CK => CLK, RN => 
                           n355, Q => n_1429, QN => n2890);
   REGISTERS_reg_13_11_inst : DFFR_X1 port map( D => n3972, CK => CLK, RN => 
                           n355, Q => n_1430, QN => n2911);
   REGISTERS_reg_13_10_inst : DFFR_X1 port map( D => n3971, CK => CLK, RN => 
                           n354, Q => n_1431, QN => n2932);
   REGISTERS_reg_13_9_inst : DFFR_X1 port map( D => n3970, CK => CLK, RN => 
                           n354, Q => n_1432, QN => n2953);
   REGISTERS_reg_13_8_inst : DFFR_X1 port map( D => n3969, CK => CLK, RN => 
                           n354, Q => n_1433, QN => n2974);
   REGISTERS_reg_13_7_inst : DFFR_X1 port map( D => n3968, CK => CLK, RN => 
                           n354, Q => n_1434, QN => n3571);
   REGISTERS_reg_13_6_inst : DFFR_X1 port map( D => n3967, CK => CLK, RN => 
                           n354, Q => n_1435, QN => n3592);
   REGISTERS_reg_13_5_inst : DFFR_X1 port map( D => n3966, CK => CLK, RN => 
                           n354, Q => n_1436, QN => n3613);
   REGISTERS_reg_13_4_inst : DFFR_X1 port map( D => n3965, CK => CLK, RN => 
                           n354, Q => n_1437, QN => n3634);
   REGISTERS_reg_13_3_inst : DFFR_X1 port map( D => n3964, CK => CLK, RN => 
                           n354, Q => n_1438, QN => n3655);
   REGISTERS_reg_13_2_inst : DFFR_X1 port map( D => n3963, CK => CLK, RN => 
                           n354, Q => n_1439, QN => n3676);
   REGISTERS_reg_13_1_inst : DFFR_X1 port map( D => n3962, CK => CLK, RN => 
                           n354, Q => n_1440, QN => n3697);
   REGISTERS_reg_13_0_inst : DFFR_X1 port map( D => n3961, CK => CLK, RN => 
                           n354, Q => n_1441, QN => n3718);
   REGISTERS_reg_14_31_inst : DFFR_X1 port map( D => n3366, CK => CLK, RN => 
                           n354, Q => n2493, QN => n_1442);
   REGISTERS_reg_14_30_inst : DFFR_X1 port map( D => n3365, CK => CLK, RN => 
                           n353, Q => n2514, QN => n_1443);
   REGISTERS_reg_14_29_inst : DFFR_X1 port map( D => n3364, CK => CLK, RN => 
                           n353, Q => n2535, QN => n_1444);
   REGISTERS_reg_14_28_inst : DFFR_X1 port map( D => n3363, CK => CLK, RN => 
                           n353, Q => n2556, QN => n_1445);
   REGISTERS_reg_14_27_inst : DFFR_X1 port map( D => n3362, CK => CLK, RN => 
                           n353, Q => n2577, QN => n_1446);
   REGISTERS_reg_14_26_inst : DFFR_X1 port map( D => n3361, CK => CLK, RN => 
                           n353, Q => n2598, QN => n_1447);
   REGISTERS_reg_14_25_inst : DFFR_X1 port map( D => n3360, CK => CLK, RN => 
                           n353, Q => n2619, QN => n_1448);
   REGISTERS_reg_14_24_inst : DFFR_X1 port map( D => n3359, CK => CLK, RN => 
                           n353, Q => n2640, QN => n_1449);
   REGISTERS_reg_14_23_inst : DFFR_X1 port map( D => n3358, CK => CLK, RN => 
                           n353, Q => n2661, QN => n_1450);
   REGISTERS_reg_14_22_inst : DFFR_X1 port map( D => n3357, CK => CLK, RN => 
                           n353, Q => n2682, QN => n_1451);
   REGISTERS_reg_14_21_inst : DFFR_X1 port map( D => n3356, CK => CLK, RN => 
                           n353, Q => n2703, QN => n_1452);
   REGISTERS_reg_14_20_inst : DFFR_X1 port map( D => n3355, CK => CLK, RN => 
                           n353, Q => n2724, QN => n_1453);
   REGISTERS_reg_14_19_inst : DFFR_X1 port map( D => n3354, CK => CLK, RN => 
                           n353, Q => n2745, QN => n_1454);
   REGISTERS_reg_14_18_inst : DFFR_X1 port map( D => n3353, CK => CLK, RN => 
                           n352, Q => n2766, QN => n_1455);
   REGISTERS_reg_14_17_inst : DFFR_X1 port map( D => n3352, CK => CLK, RN => 
                           n352, Q => n2787, QN => n_1456);
   REGISTERS_reg_14_16_inst : DFFR_X1 port map( D => n3351, CK => CLK, RN => 
                           n352, Q => n2808, QN => n_1457);
   REGISTERS_reg_14_15_inst : DFFR_X1 port map( D => n3350, CK => CLK, RN => 
                           n352, Q => n2829, QN => n_1458);
   REGISTERS_reg_14_14_inst : DFFR_X1 port map( D => n3349, CK => CLK, RN => 
                           n352, Q => n2850, QN => n_1459);
   REGISTERS_reg_14_13_inst : DFFR_X1 port map( D => n3348, CK => CLK, RN => 
                           n352, Q => n2871, QN => n_1460);
   REGISTERS_reg_14_12_inst : DFFR_X1 port map( D => n3347, CK => CLK, RN => 
                           n352, Q => n2892, QN => n_1461);
   REGISTERS_reg_14_11_inst : DFFR_X1 port map( D => n3346, CK => CLK, RN => 
                           n352, Q => n2913, QN => n_1462);
   REGISTERS_reg_14_10_inst : DFFR_X1 port map( D => n3345, CK => CLK, RN => 
                           n352, Q => n2934, QN => n_1463);
   REGISTERS_reg_14_9_inst : DFFR_X1 port map( D => n3344, CK => CLK, RN => 
                           n352, Q => n2955, QN => n_1464);
   REGISTERS_reg_14_8_inst : DFFR_X1 port map( D => n3343, CK => CLK, RN => 
                           n352, Q => n2976, QN => n_1465);
   REGISTERS_reg_14_7_inst : DFFR_X1 port map( D => n3342, CK => CLK, RN => 
                           n351, Q => n3573, QN => n_1466);
   REGISTERS_reg_14_6_inst : DFFR_X1 port map( D => n3341, CK => CLK, RN => 
                           n351, Q => n3594, QN => n_1467);
   REGISTERS_reg_14_5_inst : DFFR_X1 port map( D => n3340, CK => CLK, RN => 
                           n351, Q => n3615, QN => n_1468);
   REGISTERS_reg_14_4_inst : DFFR_X1 port map( D => n3339, CK => CLK, RN => 
                           n351, Q => n3636, QN => n_1469);
   REGISTERS_reg_14_3_inst : DFFR_X1 port map( D => n3338, CK => CLK, RN => 
                           n351, Q => n3657, QN => n_1470);
   REGISTERS_reg_14_2_inst : DFFR_X1 port map( D => n3337, CK => CLK, RN => 
                           n351, Q => n3678, QN => n_1471);
   REGISTERS_reg_14_1_inst : DFFR_X1 port map( D => n3336, CK => CLK, RN => 
                           n351, Q => n3699, QN => n_1472);
   REGISTERS_reg_14_0_inst : DFFR_X1 port map( D => n3335, CK => CLK, RN => 
                           n351, Q => n3720, QN => n_1473);
   REGISTERS_reg_15_31_inst : DFFR_X1 port map( D => n3334, CK => CLK, RN => 
                           n351, Q => n2492, QN => n_1474);
   REGISTERS_reg_15_30_inst : DFFR_X1 port map( D => n3333, CK => CLK, RN => 
                           n351, Q => n2513, QN => n_1475);
   REGISTERS_reg_15_29_inst : DFFR_X1 port map( D => n3332, CK => CLK, RN => 
                           n351, Q => n2534, QN => n_1476);
   REGISTERS_reg_15_28_inst : DFFR_X1 port map( D => n3331, CK => CLK, RN => 
                           n351, Q => n2555, QN => n_1477);
   REGISTERS_reg_15_27_inst : DFFR_X1 port map( D => n3330, CK => CLK, RN => 
                           n350, Q => n2576, QN => n_1478);
   REGISTERS_reg_15_26_inst : DFFR_X1 port map( D => n3329, CK => CLK, RN => 
                           n350, Q => n2597, QN => n_1479);
   REGISTERS_reg_15_25_inst : DFFR_X1 port map( D => n3328, CK => CLK, RN => 
                           n350, Q => n2618, QN => n_1480);
   REGISTERS_reg_15_24_inst : DFFR_X1 port map( D => n3327, CK => CLK, RN => 
                           n350, Q => n2639, QN => n_1481);
   REGISTERS_reg_15_23_inst : DFFR_X1 port map( D => n3326, CK => CLK, RN => 
                           n350, Q => n2660, QN => n_1482);
   REGISTERS_reg_15_22_inst : DFFR_X1 port map( D => n3325, CK => CLK, RN => 
                           n350, Q => n2681, QN => n_1483);
   REGISTERS_reg_15_21_inst : DFFR_X1 port map( D => n3324, CK => CLK, RN => 
                           n350, Q => n2702, QN => n_1484);
   REGISTERS_reg_15_20_inst : DFFR_X1 port map( D => n3323, CK => CLK, RN => 
                           n350, Q => n2723, QN => n_1485);
   REGISTERS_reg_15_19_inst : DFFR_X1 port map( D => n3322, CK => CLK, RN => 
                           n350, Q => n2744, QN => n_1486);
   REGISTERS_reg_15_18_inst : DFFR_X1 port map( D => n3321, CK => CLK, RN => 
                           n350, Q => n2765, QN => n_1487);
   REGISTERS_reg_15_17_inst : DFFR_X1 port map( D => n3320, CK => CLK, RN => 
                           n350, Q => n2786, QN => n_1488);
   REGISTERS_reg_15_16_inst : DFFR_X1 port map( D => n3319, CK => CLK, RN => 
                           n350, Q => n2807, QN => n_1489);
   REGISTERS_reg_15_15_inst : DFFR_X1 port map( D => n3318, CK => CLK, RN => 
                           n349, Q => n2828, QN => n_1490);
   REGISTERS_reg_15_14_inst : DFFR_X1 port map( D => n3317, CK => CLK, RN => 
                           n349, Q => n2849, QN => n_1491);
   REGISTERS_reg_15_13_inst : DFFR_X1 port map( D => n3316, CK => CLK, RN => 
                           n349, Q => n2870, QN => n_1492);
   REGISTERS_reg_15_12_inst : DFFR_X1 port map( D => n3315, CK => CLK, RN => 
                           n349, Q => n2891, QN => n_1493);
   REGISTERS_reg_15_11_inst : DFFR_X1 port map( D => n3314, CK => CLK, RN => 
                           n349, Q => n2912, QN => n_1494);
   REGISTERS_reg_15_10_inst : DFFR_X1 port map( D => n3313, CK => CLK, RN => 
                           n349, Q => n2933, QN => n_1495);
   REGISTERS_reg_15_9_inst : DFFR_X1 port map( D => n3312, CK => CLK, RN => 
                           n349, Q => n2954, QN => n_1496);
   REGISTERS_reg_15_8_inst : DFFR_X1 port map( D => n3311, CK => CLK, RN => 
                           n349, Q => n2975, QN => n_1497);
   REGISTERS_reg_15_7_inst : DFFR_X1 port map( D => n3310, CK => CLK, RN => 
                           n349, Q => n3572, QN => n_1498);
   REGISTERS_reg_15_6_inst : DFFR_X1 port map( D => n3309, CK => CLK, RN => 
                           n349, Q => n3593, QN => n_1499);
   REGISTERS_reg_15_5_inst : DFFR_X1 port map( D => n3308, CK => CLK, RN => 
                           n349, Q => n3614, QN => n_1500);
   REGISTERS_reg_15_4_inst : DFFR_X1 port map( D => n3307, CK => CLK, RN => 
                           n349, Q => n3635, QN => n_1501);
   REGISTERS_reg_15_3_inst : DFFR_X1 port map( D => n3306, CK => CLK, RN => 
                           n348, Q => n3656, QN => n_1502);
   REGISTERS_reg_15_2_inst : DFFR_X1 port map( D => n3305, CK => CLK, RN => 
                           n348, Q => n3677, QN => n_1503);
   REGISTERS_reg_15_1_inst : DFFR_X1 port map( D => n3304, CK => CLK, RN => 
                           n348, Q => n3698, QN => n_1504);
   REGISTERS_reg_15_0_inst : DFFR_X1 port map( D => n3303, CK => CLK, RN => 
                           n348, Q => n3719, QN => n_1505);
   REGISTERS_reg_16_31_inst : DFFR_X1 port map( D => n4248, CK => CLK, RN => 
                           n348, Q => n840, QN => n_1506);
   REGISTERS_reg_16_30_inst : DFFR_X1 port map( D => n4247, CK => CLK, RN => 
                           n348, Q => n839, QN => n_1507);
   REGISTERS_reg_16_29_inst : DFFR_X1 port map( D => n4246, CK => CLK, RN => 
                           n348, Q => n838, QN => n_1508);
   REGISTERS_reg_16_28_inst : DFFR_X1 port map( D => n4245, CK => CLK, RN => 
                           n348, Q => n837, QN => n_1509);
   REGISTERS_reg_16_27_inst : DFFR_X1 port map( D => n4244, CK => CLK, RN => 
                           n348, Q => n836, QN => n_1510);
   REGISTERS_reg_16_26_inst : DFFR_X1 port map( D => n4243, CK => CLK, RN => 
                           n348, Q => n835, QN => n_1511);
   REGISTERS_reg_16_25_inst : DFFR_X1 port map( D => n4242, CK => CLK, RN => 
                           n348, Q => n834, QN => n_1512);
   REGISTERS_reg_16_24_inst : DFFR_X1 port map( D => n4241, CK => CLK, RN => 
                           n348, Q => n833, QN => n_1513);
   REGISTERS_reg_16_23_inst : DFFR_X1 port map( D => n4240, CK => CLK, RN => 
                           n347, Q => n832, QN => n_1514);
   REGISTERS_reg_16_22_inst : DFFR_X1 port map( D => n4239, CK => CLK, RN => 
                           n347, Q => n831, QN => n_1515);
   REGISTERS_reg_16_21_inst : DFFR_X1 port map( D => n4238, CK => CLK, RN => 
                           n347, Q => n830, QN => n_1516);
   REGISTERS_reg_16_20_inst : DFFR_X1 port map( D => n4237, CK => CLK, RN => 
                           n347, Q => n829, QN => n_1517);
   REGISTERS_reg_16_19_inst : DFFR_X1 port map( D => n4236, CK => CLK, RN => 
                           n347, Q => n828, QN => n_1518);
   REGISTERS_reg_16_18_inst : DFFR_X1 port map( D => n4235, CK => CLK, RN => 
                           n347, Q => n827, QN => n_1519);
   REGISTERS_reg_16_17_inst : DFFR_X1 port map( D => n4234, CK => CLK, RN => 
                           n347, Q => n826, QN => n_1520);
   REGISTERS_reg_16_16_inst : DFFR_X1 port map( D => n4233, CK => CLK, RN => 
                           n352, Q => n825, QN => n_1521);
   REGISTERS_reg_16_15_inst : DFFR_X1 port map( D => n4232, CK => CLK, RN => 
                           n357, Q => n824, QN => n_1522);
   REGISTERS_reg_16_14_inst : DFFR_X1 port map( D => n4231, CK => CLK, RN => 
                           n409, Q => n823, QN => n_1523);
   REGISTERS_reg_16_13_inst : DFFR_X1 port map( D => n4230, CK => CLK, RN => 
                           n409, Q => n822, QN => n_1524);
   REGISTERS_reg_16_12_inst : DFFR_X1 port map( D => n4229, CK => CLK, RN => 
                           n409, Q => n821, QN => n_1525);
   REGISTERS_reg_16_11_inst : DFFR_X1 port map( D => n4228, CK => CLK, RN => 
                           n409, Q => n820, QN => n_1526);
   REGISTERS_reg_16_10_inst : DFFR_X1 port map( D => n4227, CK => CLK, RN => 
                           n409, Q => n819, QN => n_1527);
   REGISTERS_reg_16_9_inst : DFFR_X1 port map( D => n4226, CK => CLK, RN => 
                           n408, Q => n818, QN => n_1528);
   REGISTERS_reg_16_8_inst : DFFR_X1 port map( D => n4225, CK => CLK, RN => 
                           n408, Q => n817, QN => n_1529);
   REGISTERS_reg_16_7_inst : DFFR_X1 port map( D => n4224, CK => CLK, RN => 
                           n408, Q => n816, QN => n_1530);
   REGISTERS_reg_16_6_inst : DFFR_X1 port map( D => n4223, CK => CLK, RN => 
                           n408, Q => n815, QN => n_1531);
   REGISTERS_reg_16_5_inst : DFFR_X1 port map( D => n4222, CK => CLK, RN => 
                           n408, Q => n814, QN => n_1532);
   REGISTERS_reg_16_4_inst : DFFR_X1 port map( D => n4221, CK => CLK, RN => 
                           n408, Q => n813, QN => n_1533);
   REGISTERS_reg_16_3_inst : DFFR_X1 port map( D => n4220, CK => CLK, RN => 
                           n408, Q => n812, QN => n_1534);
   REGISTERS_reg_16_2_inst : DFFR_X1 port map( D => n4219, CK => CLK, RN => 
                           n408, Q => n811, QN => n_1535);
   REGISTERS_reg_16_1_inst : DFFR_X1 port map( D => n4218, CK => CLK, RN => 
                           n408, Q => n810, QN => n_1536);
   REGISTERS_reg_16_0_inst : DFFR_X1 port map( D => n4217, CK => CLK, RN => 
                           n408, Q => n808, QN => n_1537);
   REGISTERS_reg_17_31_inst : DFFR_X1 port map( D => n4280, CK => CLK, RN => 
                           n408, Q => n_1538, QN => n2507);
   REGISTERS_reg_17_30_inst : DFFR_X1 port map( D => n4279, CK => CLK, RN => 
                           n408, Q => n_1539, QN => n2528);
   REGISTERS_reg_17_29_inst : DFFR_X1 port map( D => n4278, CK => CLK, RN => 
                           n407, Q => n_1540, QN => n2549);
   REGISTERS_reg_17_28_inst : DFFR_X1 port map( D => n4277, CK => CLK, RN => 
                           n407, Q => n_1541, QN => n2570);
   REGISTERS_reg_17_27_inst : DFFR_X1 port map( D => n4276, CK => CLK, RN => 
                           n407, Q => n_1542, QN => n2591);
   REGISTERS_reg_17_26_inst : DFFR_X1 port map( D => n4275, CK => CLK, RN => 
                           n407, Q => n_1543, QN => n2612);
   REGISTERS_reg_17_25_inst : DFFR_X1 port map( D => n4274, CK => CLK, RN => 
                           n407, Q => n_1544, QN => n2633);
   REGISTERS_reg_17_24_inst : DFFR_X1 port map( D => n4273, CK => CLK, RN => 
                           n407, Q => n_1545, QN => n2654);
   REGISTERS_reg_17_23_inst : DFFR_X1 port map( D => n4272, CK => CLK, RN => 
                           n407, Q => n_1546, QN => n2675);
   REGISTERS_reg_17_22_inst : DFFR_X1 port map( D => n4271, CK => CLK, RN => 
                           n407, Q => n_1547, QN => n2696);
   REGISTERS_reg_17_21_inst : DFFR_X1 port map( D => n4270, CK => CLK, RN => 
                           n407, Q => n_1548, QN => n2717);
   REGISTERS_reg_17_20_inst : DFFR_X1 port map( D => n4269, CK => CLK, RN => 
                           n407, Q => n_1549, QN => n2738);
   REGISTERS_reg_17_19_inst : DFFR_X1 port map( D => n4268, CK => CLK, RN => 
                           n407, Q => n_1550, QN => n2759);
   REGISTERS_reg_17_18_inst : DFFR_X1 port map( D => n4267, CK => CLK, RN => 
                           n407, Q => n_1551, QN => n2780);
   REGISTERS_reg_17_17_inst : DFFR_X1 port map( D => n4266, CK => CLK, RN => 
                           n406, Q => n_1552, QN => n2801);
   REGISTERS_reg_17_16_inst : DFFR_X1 port map( D => n4265, CK => CLK, RN => 
                           n406, Q => n_1553, QN => n2822);
   REGISTERS_reg_17_15_inst : DFFR_X1 port map( D => n4264, CK => CLK, RN => 
                           n406, Q => n_1554, QN => n2843);
   REGISTERS_reg_17_14_inst : DFFR_X1 port map( D => n4263, CK => CLK, RN => 
                           n406, Q => n_1555, QN => n2864);
   REGISTERS_reg_17_13_inst : DFFR_X1 port map( D => n4262, CK => CLK, RN => 
                           n406, Q => n_1556, QN => n2885);
   REGISTERS_reg_17_12_inst : DFFR_X1 port map( D => n4261, CK => CLK, RN => 
                           n406, Q => n_1557, QN => n2906);
   REGISTERS_reg_17_11_inst : DFFR_X1 port map( D => n4260, CK => CLK, RN => 
                           n406, Q => n_1558, QN => n2927);
   REGISTERS_reg_17_10_inst : DFFR_X1 port map( D => n4259, CK => CLK, RN => 
                           n406, Q => n_1559, QN => n2948);
   REGISTERS_reg_17_9_inst : DFFR_X1 port map( D => n4258, CK => CLK, RN => 
                           n406, Q => n_1560, QN => n2969);
   REGISTERS_reg_17_8_inst : DFFR_X1 port map( D => n4257, CK => CLK, RN => 
                           n406, Q => n_1561, QN => n3566);
   REGISTERS_reg_17_7_inst : DFFR_X1 port map( D => n4256, CK => CLK, RN => 
                           n406, Q => n_1562, QN => n3587);
   REGISTERS_reg_17_6_inst : DFFR_X1 port map( D => n4255, CK => CLK, RN => 
                           n406, Q => n_1563, QN => n3608);
   REGISTERS_reg_17_5_inst : DFFR_X1 port map( D => n4254, CK => CLK, RN => 
                           n405, Q => n_1564, QN => n3629);
   REGISTERS_reg_17_4_inst : DFFR_X1 port map( D => n4253, CK => CLK, RN => 
                           n405, Q => n_1565, QN => n3650);
   REGISTERS_reg_17_3_inst : DFFR_X1 port map( D => n4252, CK => CLK, RN => 
                           n405, Q => n_1566, QN => n3671);
   REGISTERS_reg_17_2_inst : DFFR_X1 port map( D => n4251, CK => CLK, RN => 
                           n405, Q => n_1567, QN => n3692);
   REGISTERS_reg_17_1_inst : DFFR_X1 port map( D => n4250, CK => CLK, RN => 
                           n405, Q => n_1568, QN => n3713);
   REGISTERS_reg_17_0_inst : DFFR_X1 port map( D => n4249, CK => CLK, RN => 
                           n405, Q => n_1569, QN => n3734);
   REGISTERS_reg_18_31_inst : DFFR_X1 port map( D => n3302, CK => CLK, RN => 
                           n405, Q => n2509, QN => n_1570);
   REGISTERS_reg_18_30_inst : DFFR_X1 port map( D => n3301, CK => CLK, RN => 
                           n405, Q => n2530, QN => n_1571);
   REGISTERS_reg_18_29_inst : DFFR_X1 port map( D => n3300, CK => CLK, RN => 
                           n405, Q => n2551, QN => n_1572);
   REGISTERS_reg_18_28_inst : DFFR_X1 port map( D => n3299, CK => CLK, RN => 
                           n405, Q => n2572, QN => n_1573);
   REGISTERS_reg_18_27_inst : DFFR_X1 port map( D => n3298, CK => CLK, RN => 
                           n405, Q => n2593, QN => n_1574);
   REGISTERS_reg_18_26_inst : DFFR_X1 port map( D => n3297, CK => CLK, RN => 
                           n405, Q => n2614, QN => n_1575);
   REGISTERS_reg_18_25_inst : DFFR_X1 port map( D => n3296, CK => CLK, RN => 
                           n404, Q => n2635, QN => n_1576);
   REGISTERS_reg_18_24_inst : DFFR_X1 port map( D => n3295, CK => CLK, RN => 
                           n404, Q => n2656, QN => n_1577);
   REGISTERS_reg_18_23_inst : DFFR_X1 port map( D => n3294, CK => CLK, RN => 
                           n404, Q => n2677, QN => n_1578);
   REGISTERS_reg_18_22_inst : DFFR_X1 port map( D => n3293, CK => CLK, RN => 
                           n404, Q => n2698, QN => n_1579);
   REGISTERS_reg_18_21_inst : DFFR_X1 port map( D => n3292, CK => CLK, RN => 
                           n404, Q => n2719, QN => n_1580);
   REGISTERS_reg_18_20_inst : DFFR_X1 port map( D => n3291, CK => CLK, RN => 
                           n404, Q => n2740, QN => n_1581);
   REGISTERS_reg_18_19_inst : DFFR_X1 port map( D => n3290, CK => CLK, RN => 
                           n404, Q => n2761, QN => n_1582);
   REGISTERS_reg_18_18_inst : DFFR_X1 port map( D => n3289, CK => CLK, RN => 
                           n404, Q => n2782, QN => n_1583);
   REGISTERS_reg_18_17_inst : DFFR_X1 port map( D => n3288, CK => CLK, RN => 
                           n404, Q => n2803, QN => n_1584);
   REGISTERS_reg_18_16_inst : DFFR_X1 port map( D => n3287, CK => CLK, RN => 
                           n404, Q => n2824, QN => n_1585);
   REGISTERS_reg_18_15_inst : DFFR_X1 port map( D => n3286, CK => CLK, RN => 
                           n404, Q => n2845, QN => n_1586);
   REGISTERS_reg_18_14_inst : DFFR_X1 port map( D => n3285, CK => CLK, RN => 
                           n403, Q => n2866, QN => n_1587);
   REGISTERS_reg_18_13_inst : DFFR_X1 port map( D => n3284, CK => CLK, RN => 
                           n403, Q => n2887, QN => n_1588);
   REGISTERS_reg_18_12_inst : DFFR_X1 port map( D => n3283, CK => CLK, RN => 
                           n403, Q => n2908, QN => n_1589);
   REGISTERS_reg_18_11_inst : DFFR_X1 port map( D => n3282, CK => CLK, RN => 
                           n403, Q => n2929, QN => n_1590);
   REGISTERS_reg_18_10_inst : DFFR_X1 port map( D => n3281, CK => CLK, RN => 
                           n403, Q => n2950, QN => n_1591);
   REGISTERS_reg_18_9_inst : DFFR_X1 port map( D => n3280, CK => CLK, RN => 
                           n403, Q => n2971, QN => n_1592);
   REGISTERS_reg_18_8_inst : DFFR_X1 port map( D => n3279, CK => CLK, RN => 
                           n403, Q => n3568, QN => n_1593);
   REGISTERS_reg_18_7_inst : DFFR_X1 port map( D => n3278, CK => CLK, RN => 
                           n403, Q => n3589, QN => n_1594);
   REGISTERS_reg_18_6_inst : DFFR_X1 port map( D => n3277, CK => CLK, RN => 
                           n403, Q => n3610, QN => n_1595);
   REGISTERS_reg_18_5_inst : DFFR_X1 port map( D => n3276, CK => CLK, RN => 
                           n403, Q => n3631, QN => n_1596);
   REGISTERS_reg_18_4_inst : DFFR_X1 port map( D => n3275, CK => CLK, RN => 
                           n403, Q => n3652, QN => n_1597);
   REGISTERS_reg_18_3_inst : DFFR_X1 port map( D => n3274, CK => CLK, RN => 
                           n403, Q => n3673, QN => n_1598);
   REGISTERS_reg_18_2_inst : DFFR_X1 port map( D => n3273, CK => CLK, RN => 
                           n402, Q => n3694, QN => n_1599);
   REGISTERS_reg_18_1_inst : DFFR_X1 port map( D => n3272, CK => CLK, RN => 
                           n402, Q => n3715, QN => n_1600);
   REGISTERS_reg_18_0_inst : DFFR_X1 port map( D => n3271, CK => CLK, RN => 
                           n402, Q => n3736, QN => n_1601);
   REGISTERS_reg_19_31_inst : DFFR_X1 port map( D => n3270, CK => CLK, RN => 
                           n402, Q => n2508, QN => n_1602);
   REGISTERS_reg_19_30_inst : DFFR_X1 port map( D => n3269, CK => CLK, RN => 
                           n402, Q => n2529, QN => n_1603);
   REGISTERS_reg_19_29_inst : DFFR_X1 port map( D => n3268, CK => CLK, RN => 
                           n402, Q => n2550, QN => n_1604);
   REGISTERS_reg_19_28_inst : DFFR_X1 port map( D => n3267, CK => CLK, RN => 
                           n402, Q => n2571, QN => n_1605);
   REGISTERS_reg_19_27_inst : DFFR_X1 port map( D => n3266, CK => CLK, RN => 
                           n402, Q => n2592, QN => n_1606);
   REGISTERS_reg_19_26_inst : DFFR_X1 port map( D => n3265, CK => CLK, RN => 
                           n402, Q => n2613, QN => n_1607);
   REGISTERS_reg_19_25_inst : DFFR_X1 port map( D => n3264, CK => CLK, RN => 
                           n402, Q => n2634, QN => n_1608);
   REGISTERS_reg_19_24_inst : DFFR_X1 port map( D => n3263, CK => CLK, RN => 
                           n402, Q => n2655, QN => n_1609);
   REGISTERS_reg_19_23_inst : DFFR_X1 port map( D => n3262, CK => CLK, RN => 
                           n402, Q => n2676, QN => n_1610);
   REGISTERS_reg_19_22_inst : DFFR_X1 port map( D => n3261, CK => CLK, RN => 
                           n401, Q => n2697, QN => n_1611);
   REGISTERS_reg_19_21_inst : DFFR_X1 port map( D => n3260, CK => CLK, RN => 
                           n401, Q => n2718, QN => n_1612);
   REGISTERS_reg_19_20_inst : DFFR_X1 port map( D => n3259, CK => CLK, RN => 
                           n401, Q => n2739, QN => n_1613);
   REGISTERS_reg_19_19_inst : DFFR_X1 port map( D => n3258, CK => CLK, RN => 
                           n401, Q => n2760, QN => n_1614);
   REGISTERS_reg_19_18_inst : DFFR_X1 port map( D => n3257, CK => CLK, RN => 
                           n401, Q => n2781, QN => n_1615);
   REGISTERS_reg_19_17_inst : DFFR_X1 port map( D => n3256, CK => CLK, RN => 
                           n401, Q => n2802, QN => n_1616);
   REGISTERS_reg_19_16_inst : DFFR_X1 port map( D => n3255, CK => CLK, RN => 
                           n401, Q => n2823, QN => n_1617);
   REGISTERS_reg_19_15_inst : DFFR_X1 port map( D => n3254, CK => CLK, RN => 
                           n401, Q => n2844, QN => n_1618);
   REGISTERS_reg_19_14_inst : DFFR_X1 port map( D => n3253, CK => CLK, RN => 
                           n401, Q => n2865, QN => n_1619);
   REGISTERS_reg_19_13_inst : DFFR_X1 port map( D => n3252, CK => CLK, RN => 
                           n401, Q => n2886, QN => n_1620);
   REGISTERS_reg_19_12_inst : DFFR_X1 port map( D => n3251, CK => CLK, RN => 
                           n401, Q => n2907, QN => n_1621);
   REGISTERS_reg_19_11_inst : DFFR_X1 port map( D => n3250, CK => CLK, RN => 
                           n401, Q => n2928, QN => n_1622);
   REGISTERS_reg_19_10_inst : DFFR_X1 port map( D => n3249, CK => CLK, RN => 
                           n400, Q => n2949, QN => n_1623);
   REGISTERS_reg_19_9_inst : DFFR_X1 port map( D => n3248, CK => CLK, RN => 
                           n400, Q => n2970, QN => n_1624);
   REGISTERS_reg_19_8_inst : DFFR_X1 port map( D => n3247, CK => CLK, RN => 
                           n400, Q => n3567, QN => n_1625);
   REGISTERS_reg_19_7_inst : DFFR_X1 port map( D => n3246, CK => CLK, RN => 
                           n400, Q => n3588, QN => n_1626);
   REGISTERS_reg_19_6_inst : DFFR_X1 port map( D => n3245, CK => CLK, RN => 
                           n400, Q => n3609, QN => n_1627);
   REGISTERS_reg_19_5_inst : DFFR_X1 port map( D => n3244, CK => CLK, RN => 
                           n400, Q => n3630, QN => n_1628);
   REGISTERS_reg_19_4_inst : DFFR_X1 port map( D => n3243, CK => CLK, RN => 
                           n400, Q => n3651, QN => n_1629);
   REGISTERS_reg_19_3_inst : DFFR_X1 port map( D => n3242, CK => CLK, RN => 
                           n400, Q => n3672, QN => n_1630);
   REGISTERS_reg_19_2_inst : DFFR_X1 port map( D => n3241, CK => CLK, RN => 
                           n400, Q => n3693, QN => n_1631);
   REGISTERS_reg_19_1_inst : DFFR_X1 port map( D => n3240, CK => CLK, RN => 
                           n400, Q => n3714, QN => n_1632);
   REGISTERS_reg_19_0_inst : DFFR_X1 port map( D => n3239, CK => CLK, RN => 
                           n400, Q => n3735, QN => n_1633);
   REGISTERS_reg_20_31_inst : DFFR_X1 port map( D => n4312, CK => CLK, RN => 
                           n400, Q => n_1634, QN => n2504);
   REGISTERS_reg_20_30_inst : DFFR_X1 port map( D => n4311, CK => CLK, RN => 
                           n399, Q => n_1635, QN => n2525);
   REGISTERS_reg_20_29_inst : DFFR_X1 port map( D => n4310, CK => CLK, RN => 
                           n399, Q => n_1636, QN => n2546);
   REGISTERS_reg_20_28_inst : DFFR_X1 port map( D => n4309, CK => CLK, RN => 
                           n399, Q => n_1637, QN => n2567);
   REGISTERS_reg_20_27_inst : DFFR_X1 port map( D => n4308, CK => CLK, RN => 
                           n399, Q => n_1638, QN => n2588);
   REGISTERS_reg_20_26_inst : DFFR_X1 port map( D => n4307, CK => CLK, RN => 
                           n399, Q => n_1639, QN => n2609);
   REGISTERS_reg_20_25_inst : DFFR_X1 port map( D => n4306, CK => CLK, RN => 
                           n399, Q => n_1640, QN => n2630);
   REGISTERS_reg_20_24_inst : DFFR_X1 port map( D => n4305, CK => CLK, RN => 
                           n399, Q => n_1641, QN => n2651);
   REGISTERS_reg_20_23_inst : DFFR_X1 port map( D => n4304, CK => CLK, RN => 
                           n399, Q => n_1642, QN => n2672);
   REGISTERS_reg_20_22_inst : DFFR_X1 port map( D => n4303, CK => CLK, RN => 
                           n399, Q => n_1643, QN => n2693);
   REGISTERS_reg_20_21_inst : DFFR_X1 port map( D => n4302, CK => CLK, RN => 
                           n399, Q => n_1644, QN => n2714);
   REGISTERS_reg_20_20_inst : DFFR_X1 port map( D => n4301, CK => CLK, RN => 
                           n399, Q => n_1645, QN => n2735);
   REGISTERS_reg_20_19_inst : DFFR_X1 port map( D => n4300, CK => CLK, RN => 
                           n404, Q => n_1646, QN => n2756);
   REGISTERS_reg_20_18_inst : DFFR_X1 port map( D => n4299, CK => CLK, RN => 
                           n419, Q => n_1647, QN => n2777);
   REGISTERS_reg_20_17_inst : DFFR_X1 port map( D => n4298, CK => CLK, RN => 
                           n419, Q => n_1648, QN => n2798);
   REGISTERS_reg_20_16_inst : DFFR_X1 port map( D => n4297, CK => CLK, RN => 
                           n419, Q => n_1649, QN => n2819);
   REGISTERS_reg_20_15_inst : DFFR_X1 port map( D => n4296, CK => CLK, RN => 
                           n419, Q => n_1650, QN => n2840);
   REGISTERS_reg_20_14_inst : DFFR_X1 port map( D => n4295, CK => CLK, RN => 
                           n419, Q => n_1651, QN => n2861);
   REGISTERS_reg_20_13_inst : DFFR_X1 port map( D => n4294, CK => CLK, RN => 
                           n419, Q => n_1652, QN => n2882);
   REGISTERS_reg_20_12_inst : DFFR_X1 port map( D => n4293, CK => CLK, RN => 
                           n419, Q => n_1653, QN => n2903);
   REGISTERS_reg_20_11_inst : DFFR_X1 port map( D => n4292, CK => CLK, RN => 
                           n419, Q => n_1654, QN => n2924);
   REGISTERS_reg_20_10_inst : DFFR_X1 port map( D => n4291, CK => CLK, RN => 
                           n418, Q => n_1655, QN => n2945);
   REGISTERS_reg_20_9_inst : DFFR_X1 port map( D => n4290, CK => CLK, RN => 
                           n418, Q => n_1656, QN => n2966);
   REGISTERS_reg_20_8_inst : DFFR_X1 port map( D => n4289, CK => CLK, RN => 
                           n418, Q => n_1657, QN => n3563);
   REGISTERS_reg_20_7_inst : DFFR_X1 port map( D => n4288, CK => CLK, RN => 
                           n418, Q => n_1658, QN => n3584);
   REGISTERS_reg_20_6_inst : DFFR_X1 port map( D => n4287, CK => CLK, RN => 
                           n418, Q => n_1659, QN => n3605);
   REGISTERS_reg_20_5_inst : DFFR_X1 port map( D => n4286, CK => CLK, RN => 
                           n418, Q => n_1660, QN => n3626);
   REGISTERS_reg_20_4_inst : DFFR_X1 port map( D => n4285, CK => CLK, RN => 
                           n418, Q => n_1661, QN => n3647);
   REGISTERS_reg_20_3_inst : DFFR_X1 port map( D => n4284, CK => CLK, RN => 
                           n418, Q => n_1662, QN => n3668);
   REGISTERS_reg_20_2_inst : DFFR_X1 port map( D => n4283, CK => CLK, RN => 
                           n418, Q => n_1663, QN => n3689);
   REGISTERS_reg_20_1_inst : DFFR_X1 port map( D => n4282, CK => CLK, RN => 
                           n418, Q => n_1664, QN => n3710);
   REGISTERS_reg_20_0_inst : DFFR_X1 port map( D => n4281, CK => CLK, RN => 
                           n418, Q => n_1665, QN => n3731);
   REGISTERS_reg_21_31_inst : DFFR_X1 port map( D => n4344, CK => CLK, RN => 
                           n418, Q => n940, QN => n_1666);
   REGISTERS_reg_21_30_inst : DFFR_X1 port map( D => n4343, CK => CLK, RN => 
                           n417, Q => n939, QN => n_1667);
   REGISTERS_reg_21_29_inst : DFFR_X1 port map( D => n4342, CK => CLK, RN => 
                           n417, Q => n938, QN => n_1668);
   REGISTERS_reg_21_28_inst : DFFR_X1 port map( D => n4341, CK => CLK, RN => 
                           n417, Q => n937, QN => n_1669);
   REGISTERS_reg_21_27_inst : DFFR_X1 port map( D => n4340, CK => CLK, RN => 
                           n417, Q => n936, QN => n_1670);
   REGISTERS_reg_21_26_inst : DFFR_X1 port map( D => n4339, CK => CLK, RN => 
                           n417, Q => n935, QN => n_1671);
   REGISTERS_reg_21_25_inst : DFFR_X1 port map( D => n4338, CK => CLK, RN => 
                           n417, Q => n934, QN => n_1672);
   REGISTERS_reg_21_24_inst : DFFR_X1 port map( D => n4337, CK => CLK, RN => 
                           n417, Q => n933, QN => n_1673);
   REGISTERS_reg_21_23_inst : DFFR_X1 port map( D => n4336, CK => CLK, RN => 
                           n417, Q => n932, QN => n_1674);
   REGISTERS_reg_21_22_inst : DFFR_X1 port map( D => n4335, CK => CLK, RN => 
                           n417, Q => n931, QN => n_1675);
   REGISTERS_reg_21_21_inst : DFFR_X1 port map( D => n4334, CK => CLK, RN => 
                           n417, Q => n930, QN => n_1676);
   REGISTERS_reg_21_20_inst : DFFR_X1 port map( D => n4333, CK => CLK, RN => 
                           n417, Q => n929, QN => n_1677);
   REGISTERS_reg_21_19_inst : DFFR_X1 port map( D => n4332, CK => CLK, RN => 
                           n417, Q => n928, QN => n_1678);
   REGISTERS_reg_21_18_inst : DFFR_X1 port map( D => n4331, CK => CLK, RN => 
                           n416, Q => n927, QN => n_1679);
   REGISTERS_reg_21_17_inst : DFFR_X1 port map( D => n4330, CK => CLK, RN => 
                           n416, Q => n926, QN => n_1680);
   REGISTERS_reg_21_16_inst : DFFR_X1 port map( D => n4329, CK => CLK, RN => 
                           n416, Q => n925, QN => n_1681);
   REGISTERS_reg_21_15_inst : DFFR_X1 port map( D => n4328, CK => CLK, RN => 
                           n416, Q => n924, QN => n_1682);
   REGISTERS_reg_21_14_inst : DFFR_X1 port map( D => n4327, CK => CLK, RN => 
                           n416, Q => n923, QN => n_1683);
   REGISTERS_reg_21_13_inst : DFFR_X1 port map( D => n4326, CK => CLK, RN => 
                           n416, Q => n922, QN => n_1684);
   REGISTERS_reg_21_12_inst : DFFR_X1 port map( D => n4325, CK => CLK, RN => 
                           n416, Q => n921, QN => n_1685);
   REGISTERS_reg_21_11_inst : DFFR_X1 port map( D => n4324, CK => CLK, RN => 
                           n416, Q => n920, QN => n_1686);
   REGISTERS_reg_21_10_inst : DFFR_X1 port map( D => n4323, CK => CLK, RN => 
                           n416, Q => n919, QN => n_1687);
   REGISTERS_reg_21_9_inst : DFFR_X1 port map( D => n4322, CK => CLK, RN => 
                           n416, Q => n918, QN => n_1688);
   REGISTERS_reg_21_8_inst : DFFR_X1 port map( D => n4321, CK => CLK, RN => 
                           n416, Q => n917, QN => n_1689);
   REGISTERS_reg_21_7_inst : DFFR_X1 port map( D => n4320, CK => CLK, RN => 
                           n416, Q => n916, QN => n_1690);
   REGISTERS_reg_21_6_inst : DFFR_X1 port map( D => n4319, CK => CLK, RN => 
                           n415, Q => n915, QN => n_1691);
   REGISTERS_reg_21_5_inst : DFFR_X1 port map( D => n4318, CK => CLK, RN => 
                           n415, Q => n914, QN => n_1692);
   REGISTERS_reg_21_4_inst : DFFR_X1 port map( D => n4317, CK => CLK, RN => 
                           n415, Q => n913, QN => n_1693);
   REGISTERS_reg_21_3_inst : DFFR_X1 port map( D => n4316, CK => CLK, RN => 
                           n415, Q => n912, QN => n_1694);
   REGISTERS_reg_21_2_inst : DFFR_X1 port map( D => n4315, CK => CLK, RN => 
                           n415, Q => n911, QN => n_1695);
   REGISTERS_reg_21_1_inst : DFFR_X1 port map( D => n4314, CK => CLK, RN => 
                           n415, Q => n910, QN => n_1696);
   REGISTERS_reg_21_0_inst : DFFR_X1 port map( D => n4313, CK => CLK, RN => 
                           n415, Q => n908, QN => n_1697);
   REGISTERS_reg_24_31_inst : DFFR_X1 port map( D => n3174, CK => CLK, RN => 
                           n409, Q => n2503, QN => n_1698);
   REGISTERS_reg_24_30_inst : DFFR_X1 port map( D => n3173, CK => CLK, RN => 
                           n409, Q => n2524, QN => n_1699);
   REGISTERS_reg_24_29_inst : DFFR_X1 port map( D => n3172, CK => CLK, RN => 
                           n409, Q => n2545, QN => n_1700);
   REGISTERS_reg_24_28_inst : DFFR_X1 port map( D => n3171, CK => CLK, RN => 
                           n409, Q => n2566, QN => n_1701);
   REGISTERS_reg_24_27_inst : DFFR_X1 port map( D => n3170, CK => CLK, RN => 
                           n409, Q => n2587, QN => n_1702);
   REGISTERS_reg_24_26_inst : DFFR_X1 port map( D => n3169, CK => CLK, RN => 
                           n409, Q => n2608, QN => n_1703);
   REGISTERS_reg_24_25_inst : DFFR_X1 port map( D => n3168, CK => CLK, RN => 
                           n409, Q => n2629, QN => n_1704);
   REGISTERS_reg_24_24_inst : DFFR_X1 port map( D => n3167, CK => CLK, RN => 
                           n414, Q => n2650, QN => n_1705);
   REGISTERS_reg_24_23_inst : DFFR_X1 port map( D => n3166, CK => CLK, RN => 
                           n388, Q => n2671, QN => n_1706);
   REGISTERS_reg_24_22_inst : DFFR_X1 port map( D => n3165, CK => CLK, RN => 
                           n388, Q => n2692, QN => n_1707);
   REGISTERS_reg_24_21_inst : DFFR_X1 port map( D => n3164, CK => CLK, RN => 
                           n388, Q => n2713, QN => n_1708);
   REGISTERS_reg_24_20_inst : DFFR_X1 port map( D => n3163, CK => CLK, RN => 
                           n388, Q => n2734, QN => n_1709);
   REGISTERS_reg_24_19_inst : DFFR_X1 port map( D => n3162, CK => CLK, RN => 
                           n388, Q => n2755, QN => n_1710);
   REGISTERS_reg_24_18_inst : DFFR_X1 port map( D => n3161, CK => CLK, RN => 
                           n388, Q => n2776, QN => n_1711);
   REGISTERS_reg_24_17_inst : DFFR_X1 port map( D => n3160, CK => CLK, RN => 
                           n388, Q => n2797, QN => n_1712);
   REGISTERS_reg_24_16_inst : DFFR_X1 port map( D => n3159, CK => CLK, RN => 
                           n388, Q => n2818, QN => n_1713);
   REGISTERS_reg_24_15_inst : DFFR_X1 port map( D => n3158, CK => CLK, RN => 
                           n388, Q => n2839, QN => n_1714);
   REGISTERS_reg_24_14_inst : DFFR_X1 port map( D => n3157, CK => CLK, RN => 
                           n387, Q => n2860, QN => n_1715);
   REGISTERS_reg_24_13_inst : DFFR_X1 port map( D => n3156, CK => CLK, RN => 
                           n387, Q => n2881, QN => n_1716);
   REGISTERS_reg_24_12_inst : DFFR_X1 port map( D => n3155, CK => CLK, RN => 
                           n387, Q => n2902, QN => n_1717);
   REGISTERS_reg_24_11_inst : DFFR_X1 port map( D => n3154, CK => CLK, RN => 
                           n387, Q => n2923, QN => n_1718);
   REGISTERS_reg_24_10_inst : DFFR_X1 port map( D => n3153, CK => CLK, RN => 
                           n387, Q => n2944, QN => n_1719);
   REGISTERS_reg_24_9_inst : DFFR_X1 port map( D => n3152, CK => CLK, RN => 
                           n387, Q => n2965, QN => n_1720);
   REGISTERS_reg_24_8_inst : DFFR_X1 port map( D => n3151, CK => CLK, RN => 
                           n387, Q => n3562, QN => n_1721);
   REGISTERS_reg_24_7_inst : DFFR_X1 port map( D => n3150, CK => CLK, RN => 
                           n387, Q => n3583, QN => n_1722);
   REGISTERS_reg_24_6_inst : DFFR_X1 port map( D => n3149, CK => CLK, RN => 
                           n387, Q => n3604, QN => n_1723);
   REGISTERS_reg_24_5_inst : DFFR_X1 port map( D => n3148, CK => CLK, RN => 
                           n387, Q => n3625, QN => n_1724);
   REGISTERS_reg_24_4_inst : DFFR_X1 port map( D => n3147, CK => CLK, RN => 
                           n387, Q => n3646, QN => n_1725);
   REGISTERS_reg_24_3_inst : DFFR_X1 port map( D => n3146, CK => CLK, RN => 
                           n387, Q => n3667, QN => n_1726);
   REGISTERS_reg_24_2_inst : DFFR_X1 port map( D => n3145, CK => CLK, RN => 
                           n386, Q => n3688, QN => n_1727);
   REGISTERS_reg_24_1_inst : DFFR_X1 port map( D => n3144, CK => CLK, RN => 
                           n386, Q => n3709, QN => n_1728);
   REGISTERS_reg_24_0_inst : DFFR_X1 port map( D => n3143, CK => CLK, RN => 
                           n386, Q => n3730, QN => n_1729);
   REGISTERS_reg_25_3_inst : DFFR_X1 port map( D => n3114, CK => CLK, RN => 
                           n384, Q => n3666, QN => n_1730);
   REGISTERS_reg_25_2_inst : DFFR_X1 port map( D => n3113, CK => CLK, RN => 
                           n384, Q => n3687, QN => n_1731);
   REGISTERS_reg_25_1_inst : DFFR_X1 port map( D => n3112, CK => CLK, RN => 
                           n384, Q => n3708, QN => n_1732);
   REGISTERS_reg_25_0_inst : DFFR_X1 port map( D => n3111, CK => CLK, RN => 
                           n384, Q => n3729, QN => n_1733);
   REGISTERS_reg_26_31_inst : DFFR_X1 port map( D => n4089, CK => CLK, RN => 
                           n384, Q => n671, QN => n_1734);
   REGISTERS_reg_26_30_inst : DFFR_X1 port map( D => n4120, CK => CLK, RN => 
                           n383, Q => n703, QN => n_1735);
   REGISTERS_reg_26_29_inst : DFFR_X1 port map( D => n4119, CK => CLK, RN => 
                           n383, Q => n702, QN => n_1736);
   REGISTERS_reg_26_28_inst : DFFR_X1 port map( D => n4118, CK => CLK, RN => 
                           n383, Q => n701, QN => n_1737);
   REGISTERS_reg_26_27_inst : DFFR_X1 port map( D => n4117, CK => CLK, RN => 
                           n383, Q => n700, QN => n_1738);
   REGISTERS_reg_26_26_inst : DFFR_X1 port map( D => n4116, CK => CLK, RN => 
                           n383, Q => n699, QN => n_1739);
   REGISTERS_reg_26_25_inst : DFFR_X1 port map( D => n4115, CK => CLK, RN => 
                           n383, Q => n698, QN => n_1740);
   REGISTERS_reg_26_24_inst : DFFR_X1 port map( D => n4114, CK => CLK, RN => 
                           n383, Q => n697, QN => n_1741);
   REGISTERS_reg_26_23_inst : DFFR_X1 port map( D => n4113, CK => CLK, RN => 
                           n383, Q => n696, QN => n_1742);
   REGISTERS_reg_26_22_inst : DFFR_X1 port map( D => n4112, CK => CLK, RN => 
                           n383, Q => n695, QN => n_1743);
   REGISTERS_reg_26_21_inst : DFFR_X1 port map( D => n4111, CK => CLK, RN => 
                           n383, Q => n694, QN => n_1744);
   REGISTERS_reg_26_20_inst : DFFR_X1 port map( D => n4110, CK => CLK, RN => 
                           n383, Q => n693, QN => n_1745);
   REGISTERS_reg_26_19_inst : DFFR_X1 port map( D => n4109, CK => CLK, RN => 
                           n382, Q => n692, QN => n_1746);
   REGISTERS_reg_26_18_inst : DFFR_X1 port map( D => n4108, CK => CLK, RN => 
                           n382, Q => n691, QN => n_1747);
   REGISTERS_reg_26_17_inst : DFFR_X1 port map( D => n4107, CK => CLK, RN => 
                           n382, Q => n690, QN => n_1748);
   REGISTERS_reg_26_16_inst : DFFR_X1 port map( D => n4106, CK => CLK, RN => 
                           n382, Q => n689, QN => n_1749);
   REGISTERS_reg_26_15_inst : DFFR_X1 port map( D => n4105, CK => CLK, RN => 
                           n382, Q => n688, QN => n_1750);
   REGISTERS_reg_26_14_inst : DFFR_X1 port map( D => n4104, CK => CLK, RN => 
                           n382, Q => n687, QN => n_1751);
   REGISTERS_reg_26_13_inst : DFFR_X1 port map( D => n4103, CK => CLK, RN => 
                           n382, Q => n686, QN => n_1752);
   REGISTERS_reg_26_12_inst : DFFR_X1 port map( D => n4102, CK => CLK, RN => 
                           n382, Q => n685, QN => n_1753);
   REGISTERS_reg_26_11_inst : DFFR_X1 port map( D => n4101, CK => CLK, RN => 
                           n382, Q => n684, QN => n_1754);
   REGISTERS_reg_26_10_inst : DFFR_X1 port map( D => n4100, CK => CLK, RN => 
                           n382, Q => n683, QN => n_1755);
   REGISTERS_reg_26_9_inst : DFFR_X1 port map( D => n4099, CK => CLK, RN => 
                           n382, Q => n682, QN => n_1756);
   REGISTERS_reg_26_8_inst : DFFR_X1 port map( D => n4098, CK => CLK, RN => 
                           n382, Q => n681, QN => n_1757);
   REGISTERS_reg_26_7_inst : DFFR_X1 port map( D => n4097, CK => CLK, RN => 
                           n381, Q => n680, QN => n_1758);
   REGISTERS_reg_26_6_inst : DFFR_X1 port map( D => n4096, CK => CLK, RN => 
                           n381, Q => n679, QN => n_1759);
   REGISTERS_reg_26_5_inst : DFFR_X1 port map( D => n4095, CK => CLK, RN => 
                           n381, Q => n678, QN => n_1760);
   REGISTERS_reg_26_4_inst : DFFR_X1 port map( D => n4094, CK => CLK, RN => 
                           n381, Q => n677, QN => n_1761);
   REGISTERS_reg_26_3_inst : DFFR_X1 port map( D => n4093, CK => CLK, RN => 
                           n381, Q => n676, QN => n_1762);
   REGISTERS_reg_26_2_inst : DFFR_X1 port map( D => n4092, CK => CLK, RN => 
                           n381, Q => n675, QN => n_1763);
   REGISTERS_reg_26_1_inst : DFFR_X1 port map( D => n4091, CK => CLK, RN => 
                           n381, Q => n674, QN => n_1764);
   REGISTERS_reg_26_0_inst : DFFR_X1 port map( D => n4090, CK => CLK, RN => 
                           n381, Q => n673, QN => n_1765);
   REGISTERS_reg_27_31_inst : DFFR_X1 port map( D => n4152, CK => CLK, RN => 
                           n381, Q => n_1766, QN => n3864);
   REGISTERS_reg_27_30_inst : DFFR_X1 port map( D => n4151, CK => CLK, RN => 
                           n381, Q => n_1767, QN => n3863);
   REGISTERS_reg_27_29_inst : DFFR_X1 port map( D => n4150, CK => CLK, RN => 
                           n381, Q => n_1768, QN => n3862);
   REGISTERS_reg_27_28_inst : DFFR_X1 port map( D => n4149, CK => CLK, RN => 
                           n381, Q => n_1769, QN => n3861);
   REGISTERS_reg_27_27_inst : DFFR_X1 port map( D => n4148, CK => CLK, RN => 
                           n380, Q => n_1770, QN => n3860);
   REGISTERS_reg_27_26_inst : DFFR_X1 port map( D => n4147, CK => CLK, RN => 
                           n380, Q => n_1771, QN => n3859);
   REGISTERS_reg_27_25_inst : DFFR_X1 port map( D => n4146, CK => CLK, RN => 
                           n380, Q => n_1772, QN => n3858);
   REGISTERS_reg_27_24_inst : DFFR_X1 port map( D => n4145, CK => CLK, RN => 
                           n380, Q => n_1773, QN => n3857);
   REGISTERS_reg_27_23_inst : DFFR_X1 port map( D => n4144, CK => CLK, RN => 
                           n380, Q => n_1774, QN => n3856);
   REGISTERS_reg_27_22_inst : DFFR_X1 port map( D => n4143, CK => CLK, RN => 
                           n380, Q => n_1775, QN => n3855);
   REGISTERS_reg_27_21_inst : DFFR_X1 port map( D => n4142, CK => CLK, RN => 
                           n380, Q => n_1776, QN => n3854);
   REGISTERS_reg_27_20_inst : DFFR_X1 port map( D => n4141, CK => CLK, RN => 
                           n380, Q => n_1777, QN => n3853);
   REGISTERS_reg_27_19_inst : DFFR_X1 port map( D => n4140, CK => CLK, RN => 
                           n380, Q => n_1778, QN => n3852);
   REGISTERS_reg_27_18_inst : DFFR_X1 port map( D => n4139, CK => CLK, RN => 
                           n380, Q => n_1779, QN => n3851);
   REGISTERS_reg_27_17_inst : DFFR_X1 port map( D => n4138, CK => CLK, RN => 
                           n380, Q => n_1780, QN => n3850);
   REGISTERS_reg_27_16_inst : DFFR_X1 port map( D => n4137, CK => CLK, RN => 
                           n380, Q => n_1781, QN => n3849);
   REGISTERS_reg_27_15_inst : DFFR_X1 port map( D => n4136, CK => CLK, RN => 
                           n379, Q => n_1782, QN => n3848);
   REGISTERS_reg_27_14_inst : DFFR_X1 port map( D => n4135, CK => CLK, RN => 
                           n379, Q => n_1783, QN => n3847);
   REGISTERS_reg_27_13_inst : DFFR_X1 port map( D => n4134, CK => CLK, RN => 
                           n379, Q => n_1784, QN => n3846);
   REGISTERS_reg_27_12_inst : DFFR_X1 port map( D => n4133, CK => CLK, RN => 
                           n379, Q => n_1785, QN => n3845);
   REGISTERS_reg_27_11_inst : DFFR_X1 port map( D => n4132, CK => CLK, RN => 
                           n379, Q => n_1786, QN => n3844);
   REGISTERS_reg_27_10_inst : DFFR_X1 port map( D => n4131, CK => CLK, RN => 
                           n379, Q => n_1787, QN => n3843);
   REGISTERS_reg_27_9_inst : DFFR_X1 port map( D => n4130, CK => CLK, RN => 
                           n379, Q => n_1788, QN => n3842);
   REGISTERS_reg_27_8_inst : DFFR_X1 port map( D => n4129, CK => CLK, RN => 
                           n379, Q => n_1789, QN => n3841);
   REGISTERS_reg_27_7_inst : DFFR_X1 port map( D => n4128, CK => CLK, RN => 
                           n379, Q => n_1790, QN => n3840);
   REGISTERS_reg_27_6_inst : DFFR_X1 port map( D => n4127, CK => CLK, RN => 
                           n379, Q => n_1791, QN => n3839);
   REGISTERS_reg_27_5_inst : DFFR_X1 port map( D => n4126, CK => CLK, RN => 
                           n379, Q => n_1792, QN => n3838);
   REGISTERS_reg_27_4_inst : DFFR_X1 port map( D => n4125, CK => CLK, RN => 
                           n379, Q => n_1793, QN => n3837);
   REGISTERS_reg_27_3_inst : DFFR_X1 port map( D => n4124, CK => CLK, RN => 
                           n378, Q => n_1794, QN => n3836);
   REGISTERS_reg_27_2_inst : DFFR_X1 port map( D => n4123, CK => CLK, RN => 
                           n378, Q => n_1795, QN => n3835);
   REGISTERS_reg_27_1_inst : DFFR_X1 port map( D => n4122, CK => CLK, RN => 
                           n378, Q => n_1796, QN => n3834);
   REGISTERS_reg_27_0_inst : DFFR_X1 port map( D => n4121, CK => CLK, RN => 
                           n378, Q => n_1797, QN => n3833);
   REGISTERS_reg_29_31_inst : DFFR_X1 port map( D => n3078, CK => CLK, RN => 
                           n396, Q => n3800, QN => n_1798);
   REGISTERS_reg_29_30_inst : DFFR_X1 port map( D => n3077, CK => CLK, RN => 
                           n396, Q => n3799, QN => n_1799);
   REGISTERS_reg_29_29_inst : DFFR_X1 port map( D => n3076, CK => CLK, RN => 
                           n396, Q => n3798, QN => n_1800);
   REGISTERS_reg_29_28_inst : DFFR_X1 port map( D => n3075, CK => CLK, RN => 
                           n396, Q => n3797, QN => n_1801);
   REGISTERS_reg_29_27_inst : DFFR_X1 port map( D => n3074, CK => CLK, RN => 
                           n396, Q => n3796, QN => n_1802);
   REGISTERS_reg_29_26_inst : DFFR_X1 port map( D => n3073, CK => CLK, RN => 
                           n396, Q => n3795, QN => n_1803);
   REGISTERS_reg_29_25_inst : DFFR_X1 port map( D => n3072, CK => CLK, RN => 
                           n396, Q => n3794, QN => n_1804);
   REGISTERS_reg_29_24_inst : DFFR_X1 port map( D => n3071, CK => CLK, RN => 
                           n396, Q => n3793, QN => n_1805);
   REGISTERS_reg_29_23_inst : DFFR_X1 port map( D => n3070, CK => CLK, RN => 
                           n396, Q => n3792, QN => n_1806);
   REGISTERS_reg_29_22_inst : DFFR_X1 port map( D => n3069, CK => CLK, RN => 
                           n395, Q => n3791, QN => n_1807);
   REGISTERS_reg_29_21_inst : DFFR_X1 port map( D => n3068, CK => CLK, RN => 
                           n395, Q => n3790, QN => n_1808);
   REGISTERS_reg_29_20_inst : DFFR_X1 port map( D => n3067, CK => CLK, RN => 
                           n395, Q => n3789, QN => n_1809);
   REGISTERS_reg_29_19_inst : DFFR_X1 port map( D => n3066, CK => CLK, RN => 
                           n395, Q => n3788, QN => n_1810);
   REGISTERS_reg_29_18_inst : DFFR_X1 port map( D => n3065, CK => CLK, RN => 
                           n395, Q => n3787, QN => n_1811);
   REGISTERS_reg_29_17_inst : DFFR_X1 port map( D => n3064, CK => CLK, RN => 
                           n395, Q => n3786, QN => n_1812);
   REGISTERS_reg_29_16_inst : DFFR_X1 port map( D => n3063, CK => CLK, RN => 
                           n395, Q => n3785, QN => n_1813);
   REGISTERS_reg_29_15_inst : DFFR_X1 port map( D => n3062, CK => CLK, RN => 
                           n395, Q => n3784, QN => n_1814);
   REGISTERS_reg_29_14_inst : DFFR_X1 port map( D => n3061, CK => CLK, RN => 
                           n395, Q => n3783, QN => n_1815);
   REGISTERS_reg_29_13_inst : DFFR_X1 port map( D => n3060, CK => CLK, RN => 
                           n395, Q => n3782, QN => n_1816);
   REGISTERS_reg_29_12_inst : DFFR_X1 port map( D => n3059, CK => CLK, RN => 
                           n395, Q => n3781, QN => n_1817);
   REGISTERS_reg_29_11_inst : DFFR_X1 port map( D => n3058, CK => CLK, RN => 
                           n395, Q => n3780, QN => n_1818);
   REGISTERS_reg_29_10_inst : DFFR_X1 port map( D => n3057, CK => CLK, RN => 
                           n394, Q => n3779, QN => n_1819);
   REGISTERS_reg_29_9_inst : DFFR_X1 port map( D => n3056, CK => CLK, RN => 
                           n394, Q => n3778, QN => n_1820);
   REGISTERS_reg_29_8_inst : DFFR_X1 port map( D => n3055, CK => CLK, RN => 
                           n394, Q => n3777, QN => n_1821);
   REGISTERS_reg_29_7_inst : DFFR_X1 port map( D => n3054, CK => CLK, RN => 
                           n394, Q => n3776, QN => n_1822);
   REGISTERS_reg_29_6_inst : DFFR_X1 port map( D => n3053, CK => CLK, RN => 
                           n394, Q => n3775, QN => n_1823);
   REGISTERS_reg_29_5_inst : DFFR_X1 port map( D => n3052, CK => CLK, RN => 
                           n394, Q => n3774, QN => n_1824);
   REGISTERS_reg_29_4_inst : DFFR_X1 port map( D => n3051, CK => CLK, RN => 
                           n394, Q => n3773, QN => n_1825);
   REGISTERS_reg_29_3_inst : DFFR_X1 port map( D => n3050, CK => CLK, RN => 
                           n394, Q => n3772, QN => n_1826);
   REGISTERS_reg_29_2_inst : DFFR_X1 port map( D => n3049, CK => CLK, RN => 
                           n394, Q => n3771, QN => n_1827);
   REGISTERS_reg_29_1_inst : DFFR_X1 port map( D => n3048, CK => CLK, RN => 
                           n394, Q => n3770, QN => n_1828);
   REGISTERS_reg_29_0_inst : DFFR_X1 port map( D => n3047, CK => CLK, RN => 
                           n394, Q => n3769, QN => n_1829);
   REGISTERS_reg_30_31_inst : DFFR_X1 port map( D => n4184, CK => CLK, RN => 
                           n394, Q => n_1830, QN => n3768);
   REGISTERS_reg_30_30_inst : DFFR_X1 port map( D => n4183, CK => CLK, RN => 
                           n393, Q => n_1831, QN => n3767);
   REGISTERS_reg_30_29_inst : DFFR_X1 port map( D => n4182, CK => CLK, RN => 
                           n393, Q => n_1832, QN => n3766);
   REGISTERS_reg_30_28_inst : DFFR_X1 port map( D => n4181, CK => CLK, RN => 
                           n393, Q => n_1833, QN => n3765);
   REGISTERS_reg_30_27_inst : DFFR_X1 port map( D => n4180, CK => CLK, RN => 
                           n393, Q => n_1834, QN => n3764);
   REGISTERS_reg_30_26_inst : DFFR_X1 port map( D => n4179, CK => CLK, RN => 
                           n393, Q => n_1835, QN => n3763);
   REGISTERS_reg_30_25_inst : DFFR_X1 port map( D => n4178, CK => CLK, RN => 
                           n393, Q => n_1836, QN => n3762);
   REGISTERS_reg_30_24_inst : DFFR_X1 port map( D => n4177, CK => CLK, RN => 
                           n393, Q => n_1837, QN => n3761);
   REGISTERS_reg_30_23_inst : DFFR_X1 port map( D => n4176, CK => CLK, RN => 
                           n393, Q => n_1838, QN => n3760);
   REGISTERS_reg_30_22_inst : DFFR_X1 port map( D => n4175, CK => CLK, RN => 
                           n393, Q => n_1839, QN => n3759);
   REGISTERS_reg_30_21_inst : DFFR_X1 port map( D => n4174, CK => CLK, RN => 
                           n393, Q => n_1840, QN => n3758);
   REGISTERS_reg_30_20_inst : DFFR_X1 port map( D => n4173, CK => CLK, RN => 
                           n393, Q => n_1841, QN => n3757);
   REGISTERS_reg_30_19_inst : DFFR_X1 port map( D => n4172, CK => CLK, RN => 
                           n392, Q => n_1842, QN => n3756);
   REGISTERS_reg_30_18_inst : DFFR_X1 port map( D => n4171, CK => CLK, RN => 
                           n392, Q => n_1843, QN => n3755);
   REGISTERS_reg_30_17_inst : DFFR_X1 port map( D => n4170, CK => CLK, RN => 
                           n392, Q => n_1844, QN => n3754);
   REGISTERS_reg_30_16_inst : DFFR_X1 port map( D => n4169, CK => CLK, RN => 
                           n392, Q => n_1845, QN => n3753);
   REGISTERS_reg_30_15_inst : DFFR_X1 port map( D => n4168, CK => CLK, RN => 
                           n392, Q => n_1846, QN => n3752);
   REGISTERS_reg_30_14_inst : DFFR_X1 port map( D => n4167, CK => CLK, RN => 
                           n392, Q => n_1847, QN => n3751);
   REGISTERS_reg_30_13_inst : DFFR_X1 port map( D => n4166, CK => CLK, RN => 
                           n392, Q => n_1848, QN => n3750);
   REGISTERS_reg_30_12_inst : DFFR_X1 port map( D => n4165, CK => CLK, RN => 
                           n392, Q => n_1849, QN => n3749);
   REGISTERS_reg_30_11_inst : DFFR_X1 port map( D => n4164, CK => CLK, RN => 
                           n392, Q => n_1850, QN => n3748);
   REGISTERS_reg_30_10_inst : DFFR_X1 port map( D => n4163, CK => CLK, RN => 
                           n392, Q => n_1851, QN => n3747);
   REGISTERS_reg_30_9_inst : DFFR_X1 port map( D => n4162, CK => CLK, RN => 
                           n392, Q => n_1852, QN => n3746);
   REGISTERS_reg_30_8_inst : DFFR_X1 port map( D => n4161, CK => CLK, RN => 
                           n392, Q => n_1853, QN => n3745);
   REGISTERS_reg_30_7_inst : DFFR_X1 port map( D => n4160, CK => CLK, RN => 
                           n391, Q => n_1854, QN => n3744);
   REGISTERS_reg_30_6_inst : DFFR_X1 port map( D => n4159, CK => CLK, RN => 
                           n391, Q => n_1855, QN => n3743);
   REGISTERS_reg_30_5_inst : DFFR_X1 port map( D => n4158, CK => CLK, RN => 
                           n391, Q => n_1856, QN => n3742);
   REGISTERS_reg_30_4_inst : DFFR_X1 port map( D => n4157, CK => CLK, RN => 
                           n391, Q => n_1857, QN => n3741);
   REGISTERS_reg_30_3_inst : DFFR_X1 port map( D => n4156, CK => CLK, RN => 
                           n391, Q => n_1858, QN => n3740);
   REGISTERS_reg_30_2_inst : DFFR_X1 port map( D => n4155, CK => CLK, RN => 
                           n391, Q => n_1859, QN => n3739);
   REGISTERS_reg_30_1_inst : DFFR_X1 port map( D => n4154, CK => CLK, RN => 
                           n391, Q => n_1860, QN => n3738);
   REGISTERS_reg_30_0_inst : DFFR_X1 port map( D => n4153, CK => CLK, RN => 
                           n391, Q => n_1861, QN => n3737);
   REGISTERS_reg_31_31_inst : DFFR_X1 port map( D => n4216, CK => CLK, RN => 
                           n391, Q => n806, QN => n_1862);
   OUT2_reg_31_inst : DFF_X1 port map( D => n3015, CK => CLK, Q => OUT2(31), QN
                           => n2489);
   REGISTERS_reg_31_30_inst : DFFR_X1 port map( D => n4215, CK => CLK, RN => 
                           n391, Q => n805, QN => n_1863);
   OUT2_reg_30_inst : DFF_X1 port map( D => n3016, CK => CLK, Q => OUT2(30), QN
                           => n2510);
   REGISTERS_reg_31_29_inst : DFFR_X1 port map( D => n4214, CK => CLK, RN => 
                           n391, Q => n804, QN => n_1864);
   OUT2_reg_29_inst : DFF_X1 port map( D => n3017, CK => CLK, Q => OUT2(29), QN
                           => n2531);
   REGISTERS_reg_31_28_inst : DFFR_X1 port map( D => n4213, CK => CLK, RN => 
                           n391, Q => n803, QN => n_1865);
   OUT2_reg_28_inst : DFF_X1 port map( D => n3018, CK => CLK, Q => OUT2(28), QN
                           => n2552);
   REGISTERS_reg_31_27_inst : DFFR_X1 port map( D => n4212, CK => CLK, RN => 
                           n390, Q => n802, QN => n_1866);
   OUT2_reg_27_inst : DFF_X1 port map( D => n3019, CK => CLK, Q => OUT2(27), QN
                           => n2573);
   REGISTERS_reg_31_26_inst : DFFR_X1 port map( D => n4211, CK => CLK, RN => 
                           n390, Q => n801, QN => n_1867);
   OUT2_reg_26_inst : DFF_X1 port map( D => n3020, CK => CLK, Q => OUT2(26), QN
                           => n2594);
   REGISTERS_reg_31_25_inst : DFFR_X1 port map( D => n4210, CK => CLK, RN => 
                           n390, Q => n800, QN => n_1868);
   OUT2_reg_25_inst : DFF_X1 port map( D => n3021, CK => CLK, Q => OUT2(25), QN
                           => n2615);
   REGISTERS_reg_31_24_inst : DFFR_X1 port map( D => n4209, CK => CLK, RN => 
                           n390, Q => n799, QN => n_1869);
   OUT2_reg_24_inst : DFF_X1 port map( D => n3022, CK => CLK, Q => OUT2(24), QN
                           => n2636);
   REGISTERS_reg_31_23_inst : DFFR_X1 port map( D => n4208, CK => CLK, RN => 
                           n390, Q => n798, QN => n_1870);
   OUT2_reg_23_inst : DFF_X1 port map( D => n3023, CK => CLK, Q => OUT2(23), QN
                           => n2657);
   REGISTERS_reg_31_22_inst : DFFR_X1 port map( D => n4207, CK => CLK, RN => 
                           n390, Q => n797, QN => n_1871);
   OUT2_reg_22_inst : DFF_X1 port map( D => n3024, CK => CLK, Q => OUT2(22), QN
                           => n2678);
   REGISTERS_reg_31_21_inst : DFFR_X1 port map( D => n4206, CK => CLK, RN => 
                           n390, Q => n796, QN => n_1872);
   OUT2_reg_21_inst : DFF_X1 port map( D => n3025, CK => CLK, Q => OUT2(21), QN
                           => n2699);
   REGISTERS_reg_31_20_inst : DFFR_X1 port map( D => n4205, CK => CLK, RN => 
                           n390, Q => n795, QN => n_1873);
   OUT2_reg_20_inst : DFF_X1 port map( D => n3026, CK => CLK, Q => OUT2(20), QN
                           => n2720);
   REGISTERS_reg_31_19_inst : DFFR_X1 port map( D => n4204, CK => CLK, RN => 
                           n390, Q => n794, QN => n_1874);
   OUT2_reg_19_inst : DFF_X1 port map( D => n3027, CK => CLK, Q => OUT2(19), QN
                           => n2741);
   REGISTERS_reg_31_18_inst : DFFR_X1 port map( D => n4203, CK => CLK, RN => 
                           n390, Q => n793, QN => n_1875);
   OUT2_reg_18_inst : DFF_X1 port map( D => n3028, CK => CLK, Q => OUT2(18), QN
                           => n2762);
   REGISTERS_reg_31_17_inst : DFFR_X1 port map( D => n4202, CK => CLK, RN => 
                           n390, Q => n792, QN => n_1876);
   OUT2_reg_17_inst : DFF_X1 port map( D => n3029, CK => CLK, Q => OUT2(17), QN
                           => n2783);
   REGISTERS_reg_31_16_inst : DFFR_X1 port map( D => n4201, CK => CLK, RN => 
                           n390, Q => n791, QN => n_1877);
   OUT2_reg_16_inst : DFF_X1 port map( D => n3030, CK => CLK, Q => OUT2(16), QN
                           => n2804);
   REGISTERS_reg_31_15_inst : DFFR_X1 port map( D => n4200, CK => CLK, RN => 
                           n389, Q => n790, QN => n_1878);
   OUT2_reg_15_inst : DFF_X1 port map( D => n3031, CK => CLK, Q => OUT2(15), QN
                           => n2825);
   REGISTERS_reg_31_14_inst : DFFR_X1 port map( D => n4199, CK => CLK, RN => 
                           n389, Q => n789, QN => n_1879);
   OUT2_reg_14_inst : DFF_X1 port map( D => n3032, CK => CLK, Q => OUT2(14), QN
                           => n2846);
   REGISTERS_reg_31_13_inst : DFFR_X1 port map( D => n4198, CK => CLK, RN => 
                           n389, Q => n788, QN => n_1880);
   OUT2_reg_13_inst : DFF_X1 port map( D => n3033, CK => CLK, Q => OUT2(13), QN
                           => n2867);
   REGISTERS_reg_31_12_inst : DFFR_X1 port map( D => n4197, CK => CLK, RN => 
                           n389, Q => n787, QN => n_1881);
   OUT2_reg_12_inst : DFF_X1 port map( D => n3034, CK => CLK, Q => OUT2(12), QN
                           => n2888);
   REGISTERS_reg_31_11_inst : DFFR_X1 port map( D => n4196, CK => CLK, RN => 
                           n389, Q => n786, QN => n_1882);
   OUT2_reg_11_inst : DFF_X1 port map( D => n3035, CK => CLK, Q => OUT2(11), QN
                           => n2909);
   REGISTERS_reg_31_10_inst : DFFR_X1 port map( D => n4195, CK => CLK, RN => 
                           n389, Q => n785, QN => n_1883);
   OUT2_reg_10_inst : DFF_X1 port map( D => n3036, CK => CLK, Q => OUT2(10), QN
                           => n2930);
   REGISTERS_reg_31_9_inst : DFFR_X1 port map( D => n4194, CK => CLK, RN => 
                           n389, Q => n784, QN => n_1884);
   OUT2_reg_9_inst : DFF_X1 port map( D => n3037, CK => CLK, Q => OUT2(9), QN 
                           => n2951);
   REGISTERS_reg_31_8_inst : DFFR_X1 port map( D => n4193, CK => CLK, RN => 
                           n389, Q => n783, QN => n_1885);
   OUT2_reg_8_inst : DFF_X1 port map( D => n3038, CK => CLK, Q => OUT2(8), QN 
                           => n2972);
   REGISTERS_reg_31_7_inst : DFFR_X1 port map( D => n4192, CK => CLK, RN => 
                           n389, Q => n782, QN => n_1886);
   OUT2_reg_7_inst : DFF_X1 port map( D => n3039, CK => CLK, Q => OUT2(7), QN 
                           => n3569);
   REGISTERS_reg_31_6_inst : DFFR_X1 port map( D => n4191, CK => CLK, RN => 
                           n389, Q => n781, QN => n_1887);
   OUT2_reg_6_inst : DFF_X1 port map( D => n3040, CK => CLK, Q => OUT2(6), QN 
                           => n3590);
   REGISTERS_reg_31_5_inst : DFFR_X1 port map( D => n4190, CK => CLK, RN => 
                           n389, Q => n780, QN => n_1888);
   OUT2_reg_5_inst : DFF_X1 port map( D => n3041, CK => CLK, Q => OUT2(5), QN 
                           => n3611);
   REGISTERS_reg_31_4_inst : DFFR_X1 port map( D => n4189, CK => CLK, RN => 
                           n389, Q => n779, QN => n_1889);
   OUT2_reg_4_inst : DFF_X1 port map( D => n3042, CK => CLK, Q => OUT2(4), QN 
                           => n3632);
   REGISTERS_reg_31_3_inst : DFFR_X1 port map( D => n4188, CK => CLK, RN => 
                           n388, Q => n778, QN => n_1890);
   OUT2_reg_3_inst : DFF_X1 port map( D => n3043, CK => CLK, Q => OUT2(3), QN 
                           => n3653);
   REGISTERS_reg_31_2_inst : DFFR_X1 port map( D => n4187, CK => CLK, RN => 
                           n388, Q => n777, QN => n_1891);
   OUT2_reg_2_inst : DFF_X1 port map( D => n3044, CK => CLK, Q => OUT2(2), QN 
                           => n3674);
   REGISTERS_reg_31_1_inst : DFFR_X1 port map( D => n4186, CK => CLK, RN => 
                           n388, Q => n776, QN => n_1892);
   OUT2_reg_1_inst : DFF_X1 port map( D => n3045, CK => CLK, Q => OUT2(1), QN 
                           => n3695);
   REGISTERS_reg_31_0_inst : DFFR_X1 port map( D => n4185, CK => CLK, RN => 
                           n393, Q => n774, QN => n_1893);
   OUT2_reg_0_inst : DFF_X1 port map( D => n3046, CK => CLK, Q => OUT2(0), QN 
                           => n3716);
   OUT1_reg_31_inst : DFF_X1 port map( D => n3014, CK => CLK, Q => OUT1(31), QN
                           => n2488);
   OUT1_reg_30_inst : DFF_X1 port map( D => n3013, CK => CLK, Q => OUT1(30), QN
                           => n2487);
   OUT1_reg_29_inst : DFF_X1 port map( D => n3012, CK => CLK, Q => OUT1(29), QN
                           => n2486);
   OUT1_reg_28_inst : DFF_X1 port map( D => n3011, CK => CLK, Q => OUT1(28), QN
                           => n2485);
   OUT1_reg_27_inst : DFF_X1 port map( D => n3010, CK => CLK, Q => OUT1(27), QN
                           => n2484);
   OUT1_reg_26_inst : DFF_X1 port map( D => n3009, CK => CLK, Q => OUT1(26), QN
                           => n2483);
   OUT1_reg_25_inst : DFF_X1 port map( D => n3008, CK => CLK, Q => OUT1(25), QN
                           => n2482);
   OUT1_reg_24_inst : DFF_X1 port map( D => n3007, CK => CLK, Q => OUT1(24), QN
                           => n2481);
   OUT1_reg_23_inst : DFF_X1 port map( D => n3006, CK => CLK, Q => OUT1(23), QN
                           => n2480);
   OUT1_reg_22_inst : DFF_X1 port map( D => n3005, CK => CLK, Q => OUT1(22), QN
                           => n2479);
   OUT1_reg_21_inst : DFF_X1 port map( D => n3004, CK => CLK, Q => OUT1(21), QN
                           => n2478);
   OUT1_reg_20_inst : DFF_X1 port map( D => n3003, CK => CLK, Q => OUT1(20), QN
                           => n2477);
   OUT1_reg_19_inst : DFF_X1 port map( D => n3002, CK => CLK, Q => OUT1(19), QN
                           => n2476);
   OUT1_reg_18_inst : DFF_X1 port map( D => n3001, CK => CLK, Q => OUT1(18), QN
                           => n2475);
   OUT1_reg_17_inst : DFF_X1 port map( D => n3000, CK => CLK, Q => OUT1(17), QN
                           => n2474);
   OUT1_reg_16_inst : DFF_X1 port map( D => n2999, CK => CLK, Q => OUT1(16), QN
                           => n2473);
   OUT1_reg_15_inst : DFF_X1 port map( D => n2998, CK => CLK, Q => OUT1(15), QN
                           => n2472);
   OUT1_reg_14_inst : DFF_X1 port map( D => n2997, CK => CLK, Q => OUT1(14), QN
                           => n2471);
   OUT1_reg_13_inst : DFF_X1 port map( D => n2996, CK => CLK, Q => OUT1(13), QN
                           => n2470);
   OUT1_reg_12_inst : DFF_X1 port map( D => n2995, CK => CLK, Q => OUT1(12), QN
                           => n2469);
   OUT1_reg_11_inst : DFF_X1 port map( D => n2994, CK => CLK, Q => OUT1(11), QN
                           => n2468);
   OUT1_reg_10_inst : DFF_X1 port map( D => n2993, CK => CLK, Q => OUT1(10), QN
                           => n2467);
   OUT1_reg_9_inst : DFF_X1 port map( D => n2992, CK => CLK, Q => OUT1(9), QN 
                           => n2466);
   OUT1_reg_8_inst : DFF_X1 port map( D => n2991, CK => CLK, Q => OUT1(8), QN 
                           => n2465);
   OUT1_reg_7_inst : DFF_X1 port map( D => n2990, CK => CLK, Q => OUT1(7), QN 
                           => n2464);
   OUT1_reg_6_inst : DFF_X1 port map( D => n2989, CK => CLK, Q => OUT1(6), QN 
                           => n2463);
   OUT1_reg_5_inst : DFF_X1 port map( D => n2988, CK => CLK, Q => OUT1(5), QN 
                           => n2462);
   OUT1_reg_4_inst : DFF_X1 port map( D => n2987, CK => CLK, Q => OUT1(4), QN 
                           => n2461);
   OUT1_reg_3_inst : DFF_X1 port map( D => n2986, CK => CLK, Q => OUT1(3), QN 
                           => n2460);
   OUT1_reg_2_inst : DFF_X1 port map( D => n2985, CK => CLK, Q => OUT1(2), QN 
                           => n2459);
   OUT1_reg_1_inst : DFF_X1 port map( D => n2984, CK => CLK, Q => OUT1(1), QN 
                           => n2458);
   OUT1_reg_0_inst : DFF_X1 port map( D => n2983, CK => CLK, Q => OUT1(0), QN 
                           => n2457);
   REGISTERS_reg_28_31_inst : DFFR_X1 port map( D => n3110, CK => CLK, RN => 
                           n378, Q => n3832, QN => n1785);
   REGISTERS_reg_28_30_inst : DFFR_X1 port map( D => n3109, CK => CLK, RN => 
                           n378, Q => n3831, QN => n1753);
   REGISTERS_reg_28_29_inst : DFFR_X1 port map( D => n3108, CK => CLK, RN => 
                           n378, Q => n3830, QN => n1728);
   REGISTERS_reg_28_28_inst : DFFR_X1 port map( D => n3107, CK => CLK, RN => 
                           n383, Q => n3829, QN => n1703);
   REGISTERS_reg_28_27_inst : DFFR_X1 port map( D => n3106, CK => CLK, RN => 
                           n398, Q => n3828, QN => n1678);
   REGISTERS_reg_28_26_inst : DFFR_X1 port map( D => n3105, CK => CLK, RN => 
                           n399, Q => n3827, QN => n1653);
   REGISTERS_reg_28_25_inst : DFFR_X1 port map( D => n3104, CK => CLK, RN => 
                           n398, Q => n3826, QN => n1628);
   REGISTERS_reg_28_24_inst : DFFR_X1 port map( D => n3103, CK => CLK, RN => 
                           n398, Q => n3825, QN => n1603);
   REGISTERS_reg_28_23_inst : DFFR_X1 port map( D => n3102, CK => CLK, RN => 
                           n398, Q => n3824, QN => n1578);
   REGISTERS_reg_28_22_inst : DFFR_X1 port map( D => n3101, CK => CLK, RN => 
                           n398, Q => n3823, QN => n1553);
   REGISTERS_reg_28_21_inst : DFFR_X1 port map( D => n3100, CK => CLK, RN => 
                           n398, Q => n3822, QN => n1528);
   REGISTERS_reg_28_20_inst : DFFR_X1 port map( D => n3099, CK => CLK, RN => 
                           n398, Q => n3821, QN => n1503);
   REGISTERS_reg_28_19_inst : DFFR_X1 port map( D => n3098, CK => CLK, RN => 
                           n398, Q => n3820, QN => n1478);
   REGISTERS_reg_28_18_inst : DFFR_X1 port map( D => n3097, CK => CLK, RN => 
                           n398, Q => n3819, QN => n1453);
   REGISTERS_reg_28_17_inst : DFFR_X1 port map( D => n3096, CK => CLK, RN => 
                           n398, Q => n3818, QN => n1428);
   REGISTERS_reg_28_16_inst : DFFR_X1 port map( D => n3095, CK => CLK, RN => 
                           n398, Q => n3817, QN => n1403);
   REGISTERS_reg_28_15_inst : DFFR_X1 port map( D => n3094, CK => CLK, RN => 
                           n398, Q => n3816, QN => n1378);
   REGISTERS_reg_28_14_inst : DFFR_X1 port map( D => n3093, CK => CLK, RN => 
                           n397, Q => n3815, QN => n1353);
   REGISTERS_reg_28_13_inst : DFFR_X1 port map( D => n3092, CK => CLK, RN => 
                           n397, Q => n3814, QN => n1328);
   REGISTERS_reg_28_12_inst : DFFR_X1 port map( D => n3091, CK => CLK, RN => 
                           n397, Q => n3813, QN => n1303);
   REGISTERS_reg_28_11_inst : DFFR_X1 port map( D => n3090, CK => CLK, RN => 
                           n397, Q => n3812, QN => n1278);
   REGISTERS_reg_28_10_inst : DFFR_X1 port map( D => n3089, CK => CLK, RN => 
                           n397, Q => n3811, QN => n1253);
   REGISTERS_reg_28_9_inst : DFFR_X1 port map( D => n3088, CK => CLK, RN => 
                           n397, Q => n3810, QN => n1228);
   REGISTERS_reg_28_8_inst : DFFR_X1 port map( D => n3087, CK => CLK, RN => 
                           n397, Q => n3809, QN => n1203);
   REGISTERS_reg_28_7_inst : DFFR_X1 port map( D => n3086, CK => CLK, RN => 
                           n397, Q => n3808, QN => n1178);
   REGISTERS_reg_28_6_inst : DFFR_X1 port map( D => n3085, CK => CLK, RN => 
                           n397, Q => n3807, QN => n1153);
   REGISTERS_reg_28_5_inst : DFFR_X1 port map( D => n3084, CK => CLK, RN => 
                           n397, Q => n3806, QN => n1128);
   REGISTERS_reg_28_4_inst : DFFR_X1 port map( D => n3083, CK => CLK, RN => 
                           n397, Q => n3805, QN => n1103);
   REGISTERS_reg_28_3_inst : DFFR_X1 port map( D => n3082, CK => CLK, RN => 
                           n397, Q => n3804, QN => n1078);
   REGISTERS_reg_28_2_inst : DFFR_X1 port map( D => n3081, CK => CLK, RN => 
                           n396, Q => n3803, QN => n1053);
   REGISTERS_reg_28_1_inst : DFFR_X1 port map( D => n3080, CK => CLK, RN => 
                           n396, Q => n3802, QN => n1028);
   REGISTERS_reg_28_0_inst : DFFR_X1 port map( D => n3079, CK => CLK, RN => 
                           n396, Q => n3801, QN => n976);
   REGISTERS_reg_23_31_inst : DFFR_X1 port map( D => n3206, CK => CLK, RN => 
                           n412, Q => n2505, QN => n1777);
   REGISTERS_reg_23_30_inst : DFFR_X1 port map( D => n3205, CK => CLK, RN => 
                           n412, Q => n2526, QN => n1751);
   REGISTERS_reg_23_29_inst : DFFR_X1 port map( D => n3204, CK => CLK, RN => 
                           n412, Q => n2547, QN => n1726);
   REGISTERS_reg_23_28_inst : DFFR_X1 port map( D => n3203, CK => CLK, RN => 
                           n412, Q => n2568, QN => n1701);
   REGISTERS_reg_23_27_inst : DFFR_X1 port map( D => n3202, CK => CLK, RN => 
                           n412, Q => n2589, QN => n1676);
   REGISTERS_reg_23_26_inst : DFFR_X1 port map( D => n3201, CK => CLK, RN => 
                           n412, Q => n2610, QN => n1651);
   REGISTERS_reg_23_25_inst : DFFR_X1 port map( D => n3200, CK => CLK, RN => 
                           n412, Q => n2631, QN => n1626);
   REGISTERS_reg_23_24_inst : DFFR_X1 port map( D => n3199, CK => CLK, RN => 
                           n412, Q => n2652, QN => n1601);
   REGISTERS_reg_23_23_inst : DFFR_X1 port map( D => n3198, CK => CLK, RN => 
                           n411, Q => n2673, QN => n1576);
   REGISTERS_reg_23_22_inst : DFFR_X1 port map( D => n3197, CK => CLK, RN => 
                           n411, Q => n2694, QN => n1551);
   REGISTERS_reg_23_21_inst : DFFR_X1 port map( D => n3196, CK => CLK, RN => 
                           n411, Q => n2715, QN => n1526);
   REGISTERS_reg_23_20_inst : DFFR_X1 port map( D => n3195, CK => CLK, RN => 
                           n411, Q => n2736, QN => n1501);
   REGISTERS_reg_23_19_inst : DFFR_X1 port map( D => n3194, CK => CLK, RN => 
                           n411, Q => n2757, QN => n1476);
   REGISTERS_reg_23_18_inst : DFFR_X1 port map( D => n3193, CK => CLK, RN => 
                           n411, Q => n2778, QN => n1451);
   REGISTERS_reg_23_17_inst : DFFR_X1 port map( D => n3192, CK => CLK, RN => 
                           n411, Q => n2799, QN => n1426);
   REGISTERS_reg_23_16_inst : DFFR_X1 port map( D => n3191, CK => CLK, RN => 
                           n411, Q => n2820, QN => n1401);
   REGISTERS_reg_23_15_inst : DFFR_X1 port map( D => n3190, CK => CLK, RN => 
                           n411, Q => n2841, QN => n1376);
   REGISTERS_reg_23_14_inst : DFFR_X1 port map( D => n3189, CK => CLK, RN => 
                           n411, Q => n2862, QN => n1351);
   REGISTERS_reg_23_13_inst : DFFR_X1 port map( D => n3188, CK => CLK, RN => 
                           n411, Q => n2883, QN => n1326);
   REGISTERS_reg_23_12_inst : DFFR_X1 port map( D => n3187, CK => CLK, RN => 
                           n411, Q => n2904, QN => n1301);
   REGISTERS_reg_23_11_inst : DFFR_X1 port map( D => n3186, CK => CLK, RN => 
                           n410, Q => n2925, QN => n1276);
   REGISTERS_reg_23_10_inst : DFFR_X1 port map( D => n3185, CK => CLK, RN => 
                           n410, Q => n2946, QN => n1251);
   REGISTERS_reg_23_9_inst : DFFR_X1 port map( D => n3184, CK => CLK, RN => 
                           n410, Q => n2967, QN => n1226);
   REGISTERS_reg_23_8_inst : DFFR_X1 port map( D => n3183, CK => CLK, RN => 
                           n410, Q => n3564, QN => n1201);
   REGISTERS_reg_23_7_inst : DFFR_X1 port map( D => n3182, CK => CLK, RN => 
                           n410, Q => n3585, QN => n1176);
   REGISTERS_reg_23_6_inst : DFFR_X1 port map( D => n3181, CK => CLK, RN => 
                           n410, Q => n3606, QN => n1151);
   REGISTERS_reg_23_5_inst : DFFR_X1 port map( D => n3180, CK => CLK, RN => 
                           n410, Q => n3627, QN => n1126);
   REGISTERS_reg_23_4_inst : DFFR_X1 port map( D => n3179, CK => CLK, RN => 
                           n410, Q => n3648, QN => n1101);
   REGISTERS_reg_23_3_inst : DFFR_X1 port map( D => n3178, CK => CLK, RN => 
                           n410, Q => n3669, QN => n1076);
   REGISTERS_reg_23_2_inst : DFFR_X1 port map( D => n3177, CK => CLK, RN => 
                           n410, Q => n3690, QN => n1051);
   REGISTERS_reg_23_1_inst : DFFR_X1 port map( D => n3176, CK => CLK, RN => 
                           n410, Q => n3711, QN => n1026);
   REGISTERS_reg_23_0_inst : DFFR_X1 port map( D => n3175, CK => CLK, RN => 
                           n410, Q => n3732, QN => n971);
   REGISTERS_reg_22_31_inst : DFFR_X1 port map( D => n3238, CK => CLK, RN => 
                           n415, Q => n2506, QN => n1793);
   REGISTERS_reg_22_30_inst : DFFR_X1 port map( D => n3237, CK => CLK, RN => 
                           n415, Q => n2527, QN => n1758);
   REGISTERS_reg_22_29_inst : DFFR_X1 port map( D => n3236, CK => CLK, RN => 
                           n415, Q => n2548, QN => n1733);
   REGISTERS_reg_22_28_inst : DFFR_X1 port map( D => n3235, CK => CLK, RN => 
                           n415, Q => n2569, QN => n1708);
   REGISTERS_reg_22_27_inst : DFFR_X1 port map( D => n3234, CK => CLK, RN => 
                           n415, Q => n2590, QN => n1683);
   REGISTERS_reg_22_26_inst : DFFR_X1 port map( D => n3233, CK => CLK, RN => 
                           n414, Q => n2611, QN => n1658);
   REGISTERS_reg_22_25_inst : DFFR_X1 port map( D => n3232, CK => CLK, RN => 
                           n414, Q => n2632, QN => n1633);
   REGISTERS_reg_22_24_inst : DFFR_X1 port map( D => n3231, CK => CLK, RN => 
                           n414, Q => n2653, QN => n1608);
   REGISTERS_reg_22_23_inst : DFFR_X1 port map( D => n3230, CK => CLK, RN => 
                           n414, Q => n2674, QN => n1583);
   REGISTERS_reg_22_22_inst : DFFR_X1 port map( D => n3229, CK => CLK, RN => 
                           n414, Q => n2695, QN => n1558);
   REGISTERS_reg_22_21_inst : DFFR_X1 port map( D => n3228, CK => CLK, RN => 
                           n414, Q => n2716, QN => n1533);
   REGISTERS_reg_22_20_inst : DFFR_X1 port map( D => n3227, CK => CLK, RN => 
                           n414, Q => n2737, QN => n1508);
   REGISTERS_reg_22_19_inst : DFFR_X1 port map( D => n3226, CK => CLK, RN => 
                           n414, Q => n2758, QN => n1483);
   REGISTERS_reg_22_18_inst : DFFR_X1 port map( D => n3225, CK => CLK, RN => 
                           n414, Q => n2779, QN => n1458);
   REGISTERS_reg_22_17_inst : DFFR_X1 port map( D => n3224, CK => CLK, RN => 
                           n414, Q => n2800, QN => n1433);
   REGISTERS_reg_22_16_inst : DFFR_X1 port map( D => n3223, CK => CLK, RN => 
                           n414, Q => n2821, QN => n1408);
   REGISTERS_reg_22_15_inst : DFFR_X1 port map( D => n3222, CK => CLK, RN => 
                           n413, Q => n2842, QN => n1383);
   REGISTERS_reg_22_14_inst : DFFR_X1 port map( D => n3221, CK => CLK, RN => 
                           n413, Q => n2863, QN => n1358);
   REGISTERS_reg_22_13_inst : DFFR_X1 port map( D => n3220, CK => CLK, RN => 
                           n413, Q => n2884, QN => n1333);
   REGISTERS_reg_22_12_inst : DFFR_X1 port map( D => n3219, CK => CLK, RN => 
                           n413, Q => n2905, QN => n1308);
   REGISTERS_reg_22_11_inst : DFFR_X1 port map( D => n3218, CK => CLK, RN => 
                           n413, Q => n2926, QN => n1283);
   REGISTERS_reg_22_10_inst : DFFR_X1 port map( D => n3217, CK => CLK, RN => 
                           n413, Q => n2947, QN => n1258);
   REGISTERS_reg_22_9_inst : DFFR_X1 port map( D => n3216, CK => CLK, RN => 
                           n413, Q => n2968, QN => n1233);
   REGISTERS_reg_22_8_inst : DFFR_X1 port map( D => n3215, CK => CLK, RN => 
                           n413, Q => n3565, QN => n1208);
   REGISTERS_reg_22_7_inst : DFFR_X1 port map( D => n3214, CK => CLK, RN => 
                           n413, Q => n3586, QN => n1183);
   REGISTERS_reg_22_6_inst : DFFR_X1 port map( D => n3213, CK => CLK, RN => 
                           n413, Q => n3607, QN => n1158);
   REGISTERS_reg_22_5_inst : DFFR_X1 port map( D => n3212, CK => CLK, RN => 
                           n413, Q => n3628, QN => n1133);
   REGISTERS_reg_22_4_inst : DFFR_X1 port map( D => n3211, CK => CLK, RN => 
                           n413, Q => n3649, QN => n1108);
   REGISTERS_reg_22_3_inst : DFFR_X1 port map( D => n3210, CK => CLK, RN => 
                           n412, Q => n3670, QN => n1083);
   REGISTERS_reg_22_2_inst : DFFR_X1 port map( D => n3209, CK => CLK, RN => 
                           n412, Q => n3691, QN => n1058);
   REGISTERS_reg_22_1_inst : DFFR_X1 port map( D => n3208, CK => CLK, RN => 
                           n412, Q => n3712, QN => n1033);
   REGISTERS_reg_22_0_inst : DFFR_X1 port map( D => n3207, CK => CLK, RN => 
                           n412, Q => n3733, QN => n989);
   REGISTERS_reg_7_31_inst : DFFR_X1 port map( D => n3462, CK => CLK, RN => 
                           n372, Q => n2498, QN => n1806);
   REGISTERS_reg_7_30_inst : DFFR_X1 port map( D => n3461, CK => CLK, RN => 
                           n372, Q => n2519, QN => n1767);
   REGISTERS_reg_7_29_inst : DFFR_X1 port map( D => n3460, CK => CLK, RN => 
                           n372, Q => n2540, QN => n1742);
   REGISTERS_reg_7_28_inst : DFFR_X1 port map( D => n3459, CK => CLK, RN => 
                           n372, Q => n2561, QN => n1717);
   REGISTERS_reg_7_27_inst : DFFR_X1 port map( D => n3458, CK => CLK, RN => 
                           n372, Q => n2582, QN => n1692);
   REGISTERS_reg_7_26_inst : DFFR_X1 port map( D => n3457, CK => CLK, RN => 
                           n372, Q => n2603, QN => n1667);
   REGISTERS_reg_7_25_inst : DFFR_X1 port map( D => n3456, CK => CLK, RN => 
                           n372, Q => n2624, QN => n1642);
   REGISTERS_reg_7_24_inst : DFFR_X1 port map( D => n3455, CK => CLK, RN => 
                           n372, Q => n2645, QN => n1617);
   REGISTERS_reg_7_23_inst : DFFR_X1 port map( D => n3454, CK => CLK, RN => 
                           n372, Q => n2666, QN => n1592);
   REGISTERS_reg_7_22_inst : DFFR_X1 port map( D => n3453, CK => CLK, RN => 
                           n371, Q => n2687, QN => n1567);
   REGISTERS_reg_7_21_inst : DFFR_X1 port map( D => n3452, CK => CLK, RN => 
                           n371, Q => n2708, QN => n1542);
   REGISTERS_reg_7_20_inst : DFFR_X1 port map( D => n3451, CK => CLK, RN => 
                           n371, Q => n2729, QN => n1517);
   REGISTERS_reg_7_19_inst : DFFR_X1 port map( D => n3450, CK => CLK, RN => 
                           n371, Q => n2750, QN => n1492);
   REGISTERS_reg_7_18_inst : DFFR_X1 port map( D => n3449, CK => CLK, RN => 
                           n371, Q => n2771, QN => n1467);
   REGISTERS_reg_7_17_inst : DFFR_X1 port map( D => n3448, CK => CLK, RN => 
                           n371, Q => n2792, QN => n1442);
   REGISTERS_reg_7_16_inst : DFFR_X1 port map( D => n3447, CK => CLK, RN => 
                           n371, Q => n2813, QN => n1417);
   REGISTERS_reg_7_15_inst : DFFR_X1 port map( D => n3446, CK => CLK, RN => 
                           n371, Q => n2834, QN => n1392);
   REGISTERS_reg_7_14_inst : DFFR_X1 port map( D => n3445, CK => CLK, RN => 
                           n371, Q => n2855, QN => n1367);
   REGISTERS_reg_7_13_inst : DFFR_X1 port map( D => n3444, CK => CLK, RN => 
                           n371, Q => n2876, QN => n1342);
   REGISTERS_reg_7_12_inst : DFFR_X1 port map( D => n3443, CK => CLK, RN => 
                           n371, Q => n2897, QN => n1317);
   REGISTERS_reg_7_11_inst : DFFR_X1 port map( D => n3442, CK => CLK, RN => 
                           n371, Q => n2918, QN => n1292);
   REGISTERS_reg_7_10_inst : DFFR_X1 port map( D => n3441, CK => CLK, RN => 
                           n370, Q => n2939, QN => n1267);
   REGISTERS_reg_7_9_inst : DFFR_X1 port map( D => n3440, CK => CLK, RN => n370
                           , Q => n2960, QN => n1242);
   REGISTERS_reg_7_8_inst : DFFR_X1 port map( D => n3439, CK => CLK, RN => n370
                           , Q => n2981, QN => n1217);
   REGISTERS_reg_7_7_inst : DFFR_X1 port map( D => n3438, CK => CLK, RN => n370
                           , Q => n3578, QN => n1192);
   REGISTERS_reg_7_6_inst : DFFR_X1 port map( D => n3437, CK => CLK, RN => n370
                           , Q => n3599, QN => n1167);
   REGISTERS_reg_7_5_inst : DFFR_X1 port map( D => n3436, CK => CLK, RN => n370
                           , Q => n3620, QN => n1142);
   REGISTERS_reg_7_4_inst : DFFR_X1 port map( D => n3435, CK => CLK, RN => n370
                           , Q => n3641, QN => n1117);
   REGISTERS_reg_7_3_inst : DFFR_X1 port map( D => n3434, CK => CLK, RN => n370
                           , Q => n3662, QN => n1092);
   REGISTERS_reg_7_2_inst : DFFR_X1 port map( D => n3433, CK => CLK, RN => n370
                           , Q => n3683, QN => n1067);
   REGISTERS_reg_7_1_inst : DFFR_X1 port map( D => n3432, CK => CLK, RN => n370
                           , Q => n3704, QN => n1042);
   REGISTERS_reg_7_0_inst : DFFR_X1 port map( D => n3431, CK => CLK, RN => n370
                           , Q => n3725, QN => n1012);
   REGISTERS_reg_6_31_inst : DFFR_X1 port map( D => n3494, CK => CLK, RN => 
                           n375, Q => n2499, QN => n1805);
   REGISTERS_reg_6_30_inst : DFFR_X1 port map( D => n3493, CK => CLK, RN => 
                           n375, Q => n2520, QN => n1766);
   REGISTERS_reg_6_29_inst : DFFR_X1 port map( D => n3492, CK => CLK, RN => 
                           n375, Q => n2541, QN => n1741);
   REGISTERS_reg_6_28_inst : DFFR_X1 port map( D => n3491, CK => CLK, RN => 
                           n375, Q => n2562, QN => n1716);
   REGISTERS_reg_6_27_inst : DFFR_X1 port map( D => n3490, CK => CLK, RN => 
                           n375, Q => n2583, QN => n1691);
   REGISTERS_reg_6_26_inst : DFFR_X1 port map( D => n3489, CK => CLK, RN => 
                           n375, Q => n2604, QN => n1666);
   REGISTERS_reg_6_25_inst : DFFR_X1 port map( D => n3488, CK => CLK, RN => 
                           n374, Q => n2625, QN => n1641);
   REGISTERS_reg_6_24_inst : DFFR_X1 port map( D => n3487, CK => CLK, RN => 
                           n374, Q => n2646, QN => n1616);
   REGISTERS_reg_6_23_inst : DFFR_X1 port map( D => n3486, CK => CLK, RN => 
                           n374, Q => n2667, QN => n1591);
   REGISTERS_reg_6_22_inst : DFFR_X1 port map( D => n3485, CK => CLK, RN => 
                           n374, Q => n2688, QN => n1566);
   REGISTERS_reg_6_21_inst : DFFR_X1 port map( D => n3484, CK => CLK, RN => 
                           n374, Q => n2709, QN => n1541);
   REGISTERS_reg_6_20_inst : DFFR_X1 port map( D => n3483, CK => CLK, RN => 
                           n374, Q => n2730, QN => n1516);
   REGISTERS_reg_6_19_inst : DFFR_X1 port map( D => n3482, CK => CLK, RN => 
                           n374, Q => n2751, QN => n1491);
   REGISTERS_reg_6_18_inst : DFFR_X1 port map( D => n3481, CK => CLK, RN => 
                           n374, Q => n2772, QN => n1466);
   REGISTERS_reg_6_17_inst : DFFR_X1 port map( D => n3480, CK => CLK, RN => 
                           n374, Q => n2793, QN => n1441);
   REGISTERS_reg_6_16_inst : DFFR_X1 port map( D => n3479, CK => CLK, RN => 
                           n374, Q => n2814, QN => n1416);
   REGISTERS_reg_6_15_inst : DFFR_X1 port map( D => n3478, CK => CLK, RN => 
                           n374, Q => n2835, QN => n1391);
   REGISTERS_reg_6_14_inst : DFFR_X1 port map( D => n3477, CK => CLK, RN => 
                           n374, Q => n2856, QN => n1366);
   REGISTERS_reg_6_13_inst : DFFR_X1 port map( D => n3476, CK => CLK, RN => 
                           n373, Q => n2877, QN => n1341);
   REGISTERS_reg_6_12_inst : DFFR_X1 port map( D => n3475, CK => CLK, RN => 
                           n373, Q => n2898, QN => n1316);
   REGISTERS_reg_6_11_inst : DFFR_X1 port map( D => n3474, CK => CLK, RN => 
                           n373, Q => n2919, QN => n1291);
   REGISTERS_reg_6_10_inst : DFFR_X1 port map( D => n3473, CK => CLK, RN => 
                           n373, Q => n2940, QN => n1266);
   REGISTERS_reg_6_9_inst : DFFR_X1 port map( D => n3472, CK => CLK, RN => n373
                           , Q => n2961, QN => n1241);
   REGISTERS_reg_6_8_inst : DFFR_X1 port map( D => n3471, CK => CLK, RN => n373
                           , Q => n2982, QN => n1216);
   REGISTERS_reg_6_7_inst : DFFR_X1 port map( D => n3470, CK => CLK, RN => n373
                           , Q => n3579, QN => n1191);
   REGISTERS_reg_6_6_inst : DFFR_X1 port map( D => n3469, CK => CLK, RN => n373
                           , Q => n3600, QN => n1166);
   REGISTERS_reg_6_5_inst : DFFR_X1 port map( D => n3468, CK => CLK, RN => n373
                           , Q => n3621, QN => n1141);
   REGISTERS_reg_6_4_inst : DFFR_X1 port map( D => n3467, CK => CLK, RN => n373
                           , Q => n3642, QN => n1116);
   REGISTERS_reg_6_3_inst : DFFR_X1 port map( D => n3466, CK => CLK, RN => n373
                           , Q => n3663, QN => n1091);
   REGISTERS_reg_6_2_inst : DFFR_X1 port map( D => n3465, CK => CLK, RN => n372
                           , Q => n3684, QN => n1066);
   REGISTERS_reg_6_1_inst : DFFR_X1 port map( D => n3464, CK => CLK, RN => n372
                           , Q => n3705, QN => n1041);
   REGISTERS_reg_6_0_inst : DFFR_X1 port map( D => n3463, CK => CLK, RN => n372
                           , Q => n3726, QN => n1010);
   REGISTERS_reg_3_31_inst : DFFR_X1 port map( D => n3526, CK => CLK, RN => 
                           n362, Q => n2500, QN => n1813);
   REGISTERS_reg_3_30_inst : DFFR_X1 port map( D => n3525, CK => CLK, RN => 
                           n362, Q => n2521, QN => n1770);
   REGISTERS_reg_3_29_inst : DFFR_X1 port map( D => n3524, CK => CLK, RN => 
                           n362, Q => n2542, QN => n1745);
   REGISTERS_reg_3_28_inst : DFFR_X1 port map( D => n3523, CK => CLK, RN => 
                           n362, Q => n2563, QN => n1720);
   REGISTERS_reg_3_27_inst : DFFR_X1 port map( D => n3522, CK => CLK, RN => 
                           n362, Q => n2584, QN => n1695);
   REGISTERS_reg_3_26_inst : DFFR_X1 port map( D => n3521, CK => CLK, RN => 
                           n362, Q => n2605, QN => n1670);
   REGISTERS_reg_3_25_inst : DFFR_X1 port map( D => n3520, CK => CLK, RN => 
                           n362, Q => n2626, QN => n1645);
   REGISTERS_reg_3_24_inst : DFFR_X1 port map( D => n3519, CK => CLK, RN => 
                           n362, Q => n2647, QN => n1620);
   REGISTERS_reg_3_23_inst : DFFR_X1 port map( D => n3518, CK => CLK, RN => 
                           n362, Q => n2668, QN => n1595);
   REGISTERS_reg_3_22_inst : DFFR_X1 port map( D => n3517, CK => CLK, RN => 
                           n362, Q => n2689, QN => n1570);
   REGISTERS_reg_3_21_inst : DFFR_X1 port map( D => n3516, CK => CLK, RN => 
                           n361, Q => n2710, QN => n1545);
   REGISTERS_reg_3_20_inst : DFFR_X1 port map( D => n3515, CK => CLK, RN => 
                           n361, Q => n2731, QN => n1520);
   REGISTERS_reg_3_19_inst : DFFR_X1 port map( D => n3514, CK => CLK, RN => 
                           n361, Q => n2752, QN => n1495);
   REGISTERS_reg_3_18_inst : DFFR_X1 port map( D => n3513, CK => CLK, RN => 
                           n361, Q => n2773, QN => n1470);
   REGISTERS_reg_3_17_inst : DFFR_X1 port map( D => n3512, CK => CLK, RN => 
                           n361, Q => n2794, QN => n1445);
   REGISTERS_reg_3_16_inst : DFFR_X1 port map( D => n3511, CK => CLK, RN => 
                           n361, Q => n2815, QN => n1420);
   REGISTERS_reg_3_15_inst : DFFR_X1 port map( D => n3510, CK => CLK, RN => 
                           n361, Q => n2836, QN => n1395);
   REGISTERS_reg_3_14_inst : DFFR_X1 port map( D => n3509, CK => CLK, RN => 
                           n361, Q => n2857, QN => n1370);
   REGISTERS_reg_3_13_inst : DFFR_X1 port map( D => n3508, CK => CLK, RN => 
                           n361, Q => n2878, QN => n1345);
   REGISTERS_reg_3_12_inst : DFFR_X1 port map( D => n3507, CK => CLK, RN => 
                           n361, Q => n2899, QN => n1320);
   REGISTERS_reg_3_11_inst : DFFR_X1 port map( D => n3506, CK => CLK, RN => 
                           n361, Q => n2920, QN => n1295);
   REGISTERS_reg_3_10_inst : DFFR_X1 port map( D => n3505, CK => CLK, RN => 
                           n361, Q => n2941, QN => n1270);
   REGISTERS_reg_3_9_inst : DFFR_X1 port map( D => n3504, CK => CLK, RN => n360
                           , Q => n2962, QN => n1245);
   REGISTERS_reg_3_8_inst : DFFR_X1 port map( D => n3503, CK => CLK, RN => n360
                           , Q => n3559, QN => n1220);
   REGISTERS_reg_3_7_inst : DFFR_X1 port map( D => n3502, CK => CLK, RN => n360
                           , Q => n3580, QN => n1195);
   REGISTERS_reg_3_6_inst : DFFR_X1 port map( D => n3501, CK => CLK, RN => n360
                           , Q => n3601, QN => n1170);
   REGISTERS_reg_3_5_inst : DFFR_X1 port map( D => n3500, CK => CLK, RN => n360
                           , Q => n3622, QN => n1145);
   REGISTERS_reg_3_4_inst : DFFR_X1 port map( D => n3499, CK => CLK, RN => n360
                           , Q => n3643, QN => n1120);
   REGISTERS_reg_3_3_inst : DFFR_X1 port map( D => n3498, CK => CLK, RN => n360
                           , Q => n3664, QN => n1095);
   REGISTERS_reg_3_2_inst : DFFR_X1 port map( D => n3497, CK => CLK, RN => n360
                           , Q => n3685, QN => n1070);
   REGISTERS_reg_3_1_inst : DFFR_X1 port map( D => n3496, CK => CLK, RN => n360
                           , Q => n3706, QN => n1045);
   REGISTERS_reg_3_0_inst : DFFR_X1 port map( D => n3495, CK => CLK, RN => n360
                           , Q => n3727, QN => n1019);
   REGISTERS_reg_2_31_inst : DFFR_X1 port map( D => n3558, CK => CLK, RN => 
                           n365, Q => n2501, QN => n1812);
   REGISTERS_reg_2_30_inst : DFFR_X1 port map( D => n3557, CK => CLK, RN => 
                           n365, Q => n2522, QN => n1769);
   REGISTERS_reg_2_29_inst : DFFR_X1 port map( D => n3556, CK => CLK, RN => 
                           n365, Q => n2543, QN => n1744);
   REGISTERS_reg_2_28_inst : DFFR_X1 port map( D => n3555, CK => CLK, RN => 
                           n365, Q => n2564, QN => n1719);
   REGISTERS_reg_2_27_inst : DFFR_X1 port map( D => n3554, CK => CLK, RN => 
                           n365, Q => n2585, QN => n1694);
   REGISTERS_reg_2_26_inst : DFFR_X1 port map( D => n3553, CK => CLK, RN => 
                           n365, Q => n2606, QN => n1669);
   REGISTERS_reg_2_25_inst : DFFR_X1 port map( D => n3552, CK => CLK, RN => 
                           n365, Q => n2627, QN => n1644);
   REGISTERS_reg_2_24_inst : DFFR_X1 port map( D => n3551, CK => CLK, RN => 
                           n364, Q => n2648, QN => n1619);
   REGISTERS_reg_2_23_inst : DFFR_X1 port map( D => n3550, CK => CLK, RN => 
                           n364, Q => n2669, QN => n1594);
   REGISTERS_reg_2_22_inst : DFFR_X1 port map( D => n3549, CK => CLK, RN => 
                           n364, Q => n2690, QN => n1569);
   REGISTERS_reg_2_21_inst : DFFR_X1 port map( D => n3548, CK => CLK, RN => 
                           n364, Q => n2711, QN => n1544);
   REGISTERS_reg_2_20_inst : DFFR_X1 port map( D => n3547, CK => CLK, RN => 
                           n364, Q => n2732, QN => n1519);
   REGISTERS_reg_2_19_inst : DFFR_X1 port map( D => n3546, CK => CLK, RN => 
                           n364, Q => n2753, QN => n1494);
   REGISTERS_reg_2_18_inst : DFFR_X1 port map( D => n3545, CK => CLK, RN => 
                           n364, Q => n2774, QN => n1469);
   REGISTERS_reg_2_17_inst : DFFR_X1 port map( D => n3544, CK => CLK, RN => 
                           n364, Q => n2795, QN => n1444);
   REGISTERS_reg_2_16_inst : DFFR_X1 port map( D => n3543, CK => CLK, RN => 
                           n364, Q => n2816, QN => n1419);
   REGISTERS_reg_2_15_inst : DFFR_X1 port map( D => n3542, CK => CLK, RN => 
                           n364, Q => n2837, QN => n1394);
   REGISTERS_reg_2_14_inst : DFFR_X1 port map( D => n3541, CK => CLK, RN => 
                           n364, Q => n2858, QN => n1369);
   REGISTERS_reg_2_13_inst : DFFR_X1 port map( D => n3540, CK => CLK, RN => 
                           n364, Q => n2879, QN => n1344);
   REGISTERS_reg_2_12_inst : DFFR_X1 port map( D => n3539, CK => CLK, RN => 
                           n363, Q => n2900, QN => n1319);
   REGISTERS_reg_2_11_inst : DFFR_X1 port map( D => n3538, CK => CLK, RN => 
                           n363, Q => n2921, QN => n1294);
   REGISTERS_reg_2_10_inst : DFFR_X1 port map( D => n3537, CK => CLK, RN => 
                           n363, Q => n2942, QN => n1269);
   REGISTERS_reg_2_9_inst : DFFR_X1 port map( D => n3536, CK => CLK, RN => n363
                           , Q => n2963, QN => n1244);
   REGISTERS_reg_2_8_inst : DFFR_X1 port map( D => n3535, CK => CLK, RN => n363
                           , Q => n3560, QN => n1219);
   REGISTERS_reg_2_7_inst : DFFR_X1 port map( D => n3534, CK => CLK, RN => n363
                           , Q => n3581, QN => n1194);
   REGISTERS_reg_2_6_inst : DFFR_X1 port map( D => n3533, CK => CLK, RN => n363
                           , Q => n3602, QN => n1169);
   REGISTERS_reg_2_5_inst : DFFR_X1 port map( D => n3532, CK => CLK, RN => n363
                           , Q => n3623, QN => n1144);
   REGISTERS_reg_2_4_inst : DFFR_X1 port map( D => n3531, CK => CLK, RN => n363
                           , Q => n3644, QN => n1119);
   REGISTERS_reg_2_3_inst : DFFR_X1 port map( D => n3530, CK => CLK, RN => n363
                           , Q => n3665, QN => n1094);
   REGISTERS_reg_2_2_inst : DFFR_X1 port map( D => n3529, CK => CLK, RN => n363
                           , Q => n3686, QN => n1069);
   REGISTERS_reg_2_1_inst : DFFR_X1 port map( D => n3528, CK => CLK, RN => n363
                           , Q => n3707, QN => n1044);
   REGISTERS_reg_2_0_inst : DFFR_X1 port map( D => n3527, CK => CLK, RN => n362
                           , Q => n3728, QN => n1017);
   REGISTERS_reg_25_31_inst : DFFR_X1 port map( D => n3142, CK => CLK, RN => 
                           n386, Q => n2502, QN => n_1894);
   REGISTERS_reg_25_30_inst : DFFR_X1 port map( D => n3141, CK => CLK, RN => 
                           n386, Q => n2523, QN => n_1895);
   REGISTERS_reg_25_29_inst : DFFR_X1 port map( D => n3140, CK => CLK, RN => 
                           n386, Q => n2544, QN => n_1896);
   REGISTERS_reg_25_28_inst : DFFR_X1 port map( D => n3139, CK => CLK, RN => 
                           n386, Q => n2565, QN => n_1897);
   REGISTERS_reg_25_27_inst : DFFR_X1 port map( D => n3138, CK => CLK, RN => 
                           n386, Q => n2586, QN => n_1898);
   REGISTERS_reg_25_26_inst : DFFR_X1 port map( D => n3137, CK => CLK, RN => 
                           n386, Q => n2607, QN => n_1899);
   REGISTERS_reg_25_25_inst : DFFR_X1 port map( D => n3136, CK => CLK, RN => 
                           n386, Q => n2628, QN => n_1900);
   REGISTERS_reg_25_24_inst : DFFR_X1 port map( D => n3135, CK => CLK, RN => 
                           n386, Q => n2649, QN => n_1901);
   REGISTERS_reg_25_23_inst : DFFR_X1 port map( D => n3134, CK => CLK, RN => 
                           n386, Q => n2670, QN => n_1902);
   REGISTERS_reg_25_22_inst : DFFR_X1 port map( D => n3133, CK => CLK, RN => 
                           n385, Q => n2691, QN => n_1903);
   REGISTERS_reg_25_21_inst : DFFR_X1 port map( D => n3132, CK => CLK, RN => 
                           n385, Q => n2712, QN => n_1904);
   REGISTERS_reg_25_20_inst : DFFR_X1 port map( D => n3131, CK => CLK, RN => 
                           n385, Q => n2733, QN => n_1905);
   REGISTERS_reg_25_19_inst : DFFR_X1 port map( D => n3130, CK => CLK, RN => 
                           n385, Q => n2754, QN => n_1906);
   REGISTERS_reg_25_18_inst : DFFR_X1 port map( D => n3129, CK => CLK, RN => 
                           n385, Q => n2775, QN => n_1907);
   REGISTERS_reg_25_17_inst : DFFR_X1 port map( D => n3128, CK => CLK, RN => 
                           n385, Q => n2796, QN => n_1908);
   REGISTERS_reg_25_16_inst : DFFR_X1 port map( D => n3127, CK => CLK, RN => 
                           n385, Q => n2817, QN => n_1909);
   REGISTERS_reg_25_15_inst : DFFR_X1 port map( D => n3126, CK => CLK, RN => 
                           n385, Q => n2838, QN => n_1910);
   REGISTERS_reg_25_14_inst : DFFR_X1 port map( D => n3125, CK => CLK, RN => 
                           n385, Q => n2859, QN => n_1911);
   REGISTERS_reg_25_13_inst : DFFR_X1 port map( D => n3124, CK => CLK, RN => 
                           n385, Q => n2880, QN => n_1912);
   REGISTERS_reg_25_12_inst : DFFR_X1 port map( D => n3123, CK => CLK, RN => 
                           n385, Q => n2901, QN => n_1913);
   REGISTERS_reg_25_11_inst : DFFR_X1 port map( D => n3122, CK => CLK, RN => 
                           n385, Q => n2922, QN => n_1914);
   REGISTERS_reg_25_10_inst : DFFR_X1 port map( D => n3121, CK => CLK, RN => 
                           n384, Q => n2943, QN => n_1915);
   REGISTERS_reg_25_9_inst : DFFR_X1 port map( D => n3120, CK => CLK, RN => 
                           n384, Q => n2964, QN => n_1916);
   REGISTERS_reg_25_8_inst : DFFR_X1 port map( D => n3119, CK => CLK, RN => 
                           n384, Q => n3561, QN => n_1917);
   REGISTERS_reg_25_7_inst : DFFR_X1 port map( D => n3118, CK => CLK, RN => 
                           n384, Q => n3582, QN => n_1918);
   REGISTERS_reg_25_6_inst : DFFR_X1 port map( D => n3117, CK => CLK, RN => 
                           n384, Q => n3603, QN => n_1919);
   REGISTERS_reg_25_5_inst : DFFR_X1 port map( D => n3116, CK => CLK, RN => 
                           n384, Q => n3624, QN => n_1920);
   REGISTERS_reg_25_4_inst : DFFR_X1 port map( D => n3115, CK => CLK, RN => 
                           n384, Q => n3645, QN => n_1921);
   U2 : BUF_X1 port map( A => n420, Z => n419);
   U3 : BUF_X1 port map( A => n980, Z => n122);
   U4 : BUF_X1 port map( A => n980, Z => n121);
   U5 : BUF_X1 port map( A => n980, Z => n123);
   U6 : BUF_X1 port map( A => n1838, Z => n223);
   U7 : BUF_X1 port map( A => n1833, Z => n211);
   U8 : BUF_X1 port map( A => n1848, Z => n244);
   U9 : BUF_X1 port map( A => n1838, Z => n224);
   U10 : BUF_X1 port map( A => n1833, Z => n212);
   U11 : BUF_X1 port map( A => n1848, Z => n245);
   U12 : BUF_X1 port map( A => n974, Z => n110);
   U13 : BUF_X1 port map( A => n991, Z => n143);
   U14 : BUF_X1 port map( A => n974, Z => n109);
   U15 : BUF_X1 port map( A => n991, Z => n142);
   U16 : BUF_X1 port map( A => n1003, Z => n164);
   U17 : BUF_X1 port map( A => n1003, Z => n163);
   U18 : BUF_X1 port map( A => n1844, Z => n235);
   U19 : BUF_X1 port map( A => n1870, Z => n289);
   U20 : BUF_X1 port map( A => n1844, Z => n236);
   U21 : BUF_X1 port map( A => n1870, Z => n290);
   U22 : BUF_X1 port map( A => n986, Z => n134);
   U23 : BUF_X1 port map( A => n998, Z => n152);
   U24 : BUF_X1 port map( A => n1008, Z => n176);
   U25 : BUF_X1 port map( A => n1015, Z => n188);
   U26 : BUF_X1 port map( A => n986, Z => n133);
   U27 : BUF_X1 port map( A => n998, Z => n151);
   U28 : BUF_X1 port map( A => n1008, Z => n175);
   U29 : BUF_X1 port map( A => n1015, Z => n187);
   U30 : BUF_X1 port map( A => n1020, Z => n194);
   U31 : BUF_X1 port map( A => n1020, Z => n193);
   U32 : BUF_X1 port map( A => n1001, Z => n158);
   U33 : BUF_X1 port map( A => n1006, Z => n170);
   U34 : BUF_X1 port map( A => n1001, Z => n157);
   U35 : BUF_X1 port map( A => n1006, Z => n169);
   U36 : BUF_X1 port map( A => n1847, Z => n241);
   U37 : BUF_X1 port map( A => n1847, Z => n242);
   U38 : BUF_X1 port map( A => n990, Z => n140);
   U39 : BUF_X1 port map( A => n1013, Z => n182);
   U40 : BUF_X1 port map( A => n990, Z => n139);
   U41 : BUF_X1 port map( A => n1013, Z => n181);
   U42 : BUF_X1 port map( A => n1830, Z => n205);
   U43 : BUF_X1 port map( A => n1830, Z => n206);
   U44 : BUF_X1 port map( A => n970, Z => n104);
   U45 : BUF_X1 port map( A => n970, Z => n103);
   U46 : BUF_X1 port map( A => n1835, Z => n217);
   U47 : BUF_X1 port map( A => n1835, Z => n218);
   U48 : BUF_X1 port map( A => n977, Z => n116);
   U49 : BUF_X1 port map( A => n977, Z => n115);
   U50 : BUF_X1 port map( A => n1018, Z => n191);
   U51 : BUF_X1 port map( A => n1018, Z => n190);
   U52 : BUF_X1 port map( A => n1846, Z => n238);
   U53 : BUF_X1 port map( A => n1846, Z => n239);
   U54 : BUF_X1 port map( A => n988, Z => n137);
   U55 : BUF_X1 port map( A => n988, Z => n136);
   U56 : BUF_X1 port map( A => n1000, Z => n155);
   U57 : BUF_X1 port map( A => n1005, Z => n167);
   U58 : BUF_X1 port map( A => n1000, Z => n154);
   U59 : BUF_X1 port map( A => n1005, Z => n166);
   U60 : BUF_X1 port map( A => n1011, Z => n179);
   U61 : BUF_X1 port map( A => n1011, Z => n178);
   U62 : BUF_X1 port map( A => n1836, Z => n220);
   U63 : BUF_X1 port map( A => n1831, Z => n208);
   U64 : BUF_X1 port map( A => n1836, Z => n221);
   U65 : BUF_X1 port map( A => n1831, Z => n209);
   U66 : BUF_X1 port map( A => n978, Z => n119);
   U67 : BUF_X1 port map( A => n972, Z => n107);
   U68 : BUF_X1 port map( A => n978, Z => n118);
   U69 : BUF_X1 port map( A => n972, Z => n106);
   U70 : BUF_X1 port map( A => n1839, Z => n226);
   U71 : BUF_X1 port map( A => n1834, Z => n214);
   U72 : BUF_X1 port map( A => n1849, Z => n247);
   U73 : BUF_X1 port map( A => n1839, Z => n227);
   U74 : BUF_X1 port map( A => n1834, Z => n215);
   U75 : BUF_X1 port map( A => n1849, Z => n248);
   U76 : BUF_X1 port map( A => n981, Z => n125);
   U77 : BUF_X1 port map( A => n975, Z => n113);
   U78 : BUF_X1 port map( A => n992, Z => n146);
   U79 : BUF_X1 port map( A => n981, Z => n124);
   U80 : BUF_X1 port map( A => n975, Z => n112);
   U81 : BUF_X1 port map( A => n992, Z => n145);
   U82 : BUF_X1 port map( A => n997, Z => n149);
   U83 : BUF_X1 port map( A => n997, Z => n148);
   U84 : BUF_X1 port map( A => n1002, Z => n161);
   U85 : BUF_X1 port map( A => n1002, Z => n160);
   U86 : BUF_X1 port map( A => n1843, Z => n232);
   U87 : BUF_X1 port map( A => n1843, Z => n233);
   U88 : BUF_X1 port map( A => n985, Z => n131);
   U89 : BUF_X1 port map( A => n1007, Z => n173);
   U90 : BUF_X1 port map( A => n1014, Z => n185);
   U91 : BUF_X1 port map( A => n985, Z => n130);
   U92 : BUF_X1 port map( A => n1007, Z => n172);
   U93 : BUF_X1 port map( A => n1014, Z => n184);
   U94 : BUF_X1 port map( A => n1840, Z => n229);
   U95 : BUF_X1 port map( A => n1840, Z => n230);
   U96 : BUF_X1 port map( A => n982, Z => n128);
   U97 : BUF_X1 port map( A => n982, Z => n127);
   U98 : BUF_X1 port map( A => n1838, Z => n225);
   U99 : BUF_X1 port map( A => n1833, Z => n213);
   U100 : BUF_X1 port map( A => n1848, Z => n246);
   U101 : BUF_X1 port map( A => n974, Z => n111);
   U102 : BUF_X1 port map( A => n991, Z => n144);
   U103 : BUF_X1 port map( A => n1003, Z => n165);
   U104 : BUF_X1 port map( A => n998, Z => n153);
   U105 : BUF_X1 port map( A => n1844, Z => n237);
   U106 : BUF_X1 port map( A => n1870, Z => n291);
   U107 : BUF_X1 port map( A => n986, Z => n135);
   U108 : BUF_X1 port map( A => n1008, Z => n177);
   U109 : BUF_X1 port map( A => n1015, Z => n189);
   U110 : BUF_X1 port map( A => n1020, Z => n195);
   U111 : BUF_X1 port map( A => n1001, Z => n159);
   U112 : BUF_X1 port map( A => n1006, Z => n171);
   U113 : BUF_X1 port map( A => n1847, Z => n243);
   U114 : BUF_X1 port map( A => n990, Z => n141);
   U115 : BUF_X1 port map( A => n1013, Z => n183);
   U116 : BUF_X1 port map( A => n1830, Z => n207);
   U117 : BUF_X1 port map( A => n970, Z => n105);
   U118 : BUF_X1 port map( A => n1835, Z => n219);
   U119 : BUF_X1 port map( A => n977, Z => n117);
   U120 : BUF_X1 port map( A => n1018, Z => n192);
   U121 : BUF_X1 port map( A => n1846, Z => n240);
   U122 : BUF_X1 port map( A => n988, Z => n138);
   U123 : BUF_X1 port map( A => n1000, Z => n156);
   U124 : BUF_X1 port map( A => n1005, Z => n168);
   U125 : BUF_X1 port map( A => n1011, Z => n180);
   U126 : BUF_X1 port map( A => n1836, Z => n222);
   U127 : BUF_X1 port map( A => n1831, Z => n210);
   U128 : BUF_X1 port map( A => n978, Z => n120);
   U129 : BUF_X1 port map( A => n972, Z => n108);
   U130 : BUF_X1 port map( A => n1839, Z => n228);
   U131 : BUF_X1 port map( A => n1834, Z => n216);
   U132 : BUF_X1 port map( A => n1849, Z => n249);
   U133 : BUF_X1 port map( A => n981, Z => n126);
   U134 : BUF_X1 port map( A => n975, Z => n114);
   U135 : BUF_X1 port map( A => n992, Z => n147);
   U136 : BUF_X1 port map( A => n997, Z => n150);
   U137 : BUF_X1 port map( A => n1002, Z => n162);
   U138 : BUF_X1 port map( A => n1843, Z => n234);
   U139 : BUF_X1 port map( A => n985, Z => n132);
   U140 : BUF_X1 port map( A => n1007, Z => n174);
   U141 : BUF_X1 port map( A => n1014, Z => n186);
   U142 : BUF_X1 port map( A => n1840, Z => n231);
   U143 : BUF_X1 port map( A => n982, Z => n129);
   U144 : BUF_X1 port map( A => n330, Z => n420);
   U145 : BUF_X1 port map( A => n331, Z => n424);
   U146 : BUF_X1 port map( A => n331, Z => n425);
   U147 : BUF_X1 port map( A => n331, Z => n423);
   U148 : BUF_X1 port map( A => n330, Z => n422);
   U149 : BUF_X1 port map( A => n330, Z => n421);
   U150 : BUF_X1 port map( A => n333, Z => n431);
   U151 : BUF_X1 port map( A => n332, Z => n427);
   U152 : BUF_X1 port map( A => n333, Z => n430);
   U153 : BUF_X1 port map( A => n333, Z => n429);
   U154 : BUF_X1 port map( A => n332, Z => n428);
   U155 : BUF_X1 port map( A => n332, Z => n426);
   U156 : BUF_X1 port map( A => n334, Z => n432);
   U157 : BUF_X1 port map( A => n334, Z => n433);
   U158 : BUF_X1 port map( A => n1860, Z => n265);
   U159 : BUF_X1 port map( A => n1860, Z => n266);
   U160 : BUF_X1 port map( A => n1855, Z => n253);
   U161 : BUF_X1 port map( A => n1865, Z => n277);
   U162 : BUF_X1 port map( A => n1855, Z => n254);
   U163 : BUF_X1 port map( A => n1865, Z => n278);
   U164 : BUF_X1 port map( A => n1873, Z => n295);
   U165 : BUF_X1 port map( A => n1873, Z => n296);
   U166 : BUF_X1 port map( A => n1858, Z => n259);
   U167 : BUF_X1 port map( A => n1863, Z => n271);
   U168 : BUF_X1 port map( A => n1858, Z => n260);
   U169 : BUF_X1 port map( A => n1863, Z => n272);
   U170 : BUF_X1 port map( A => n1868, Z => n283);
   U171 : BUF_X1 port map( A => n1868, Z => n284);
   U172 : BUF_X1 port map( A => n1872, Z => n292);
   U173 : BUF_X1 port map( A => n1872, Z => n293);
   U174 : BUF_X1 port map( A => n1857, Z => n256);
   U175 : BUF_X1 port map( A => n1862, Z => n268);
   U176 : BUF_X1 port map( A => n1857, Z => n257);
   U177 : BUF_X1 port map( A => n1862, Z => n269);
   U178 : BUF_X1 port map( A => n1867, Z => n280);
   U179 : BUF_X1 port map( A => n1867, Z => n281);
   U180 : BUF_X1 port map( A => n1854, Z => n250);
   U181 : BUF_X1 port map( A => n1854, Z => n251);
   U182 : BUF_X1 port map( A => n1859, Z => n262);
   U183 : BUF_X1 port map( A => n1859, Z => n263);
   U184 : BUF_X1 port map( A => n1864, Z => n274);
   U185 : BUF_X1 port map( A => n1869, Z => n286);
   U186 : BUF_X1 port map( A => n1864, Z => n275);
   U187 : BUF_X1 port map( A => n1869, Z => n287);
   U188 : BUF_X1 port map( A => n1860, Z => n267);
   U189 : BUF_X1 port map( A => n1855, Z => n255);
   U190 : BUF_X1 port map( A => n1865, Z => n279);
   U191 : BUF_X1 port map( A => n1873, Z => n297);
   U192 : BUF_X1 port map( A => n1858, Z => n261);
   U193 : BUF_X1 port map( A => n1863, Z => n273);
   U194 : BUF_X1 port map( A => n1868, Z => n285);
   U195 : BUF_X1 port map( A => n1872, Z => n294);
   U196 : BUF_X1 port map( A => n1857, Z => n258);
   U197 : BUF_X1 port map( A => n1862, Z => n270);
   U198 : BUF_X1 port map( A => n1867, Z => n282);
   U199 : BUF_X1 port map( A => n1854, Z => n252);
   U200 : BUF_X1 port map( A => n1859, Z => n264);
   U201 : BUF_X1 port map( A => n1864, Z => n276);
   U202 : BUF_X1 port map( A => n1869, Z => n288);
   U203 : BUF_X1 port map( A => n335, Z => n333);
   U204 : BUF_X1 port map( A => n335, Z => n332);
   U205 : BUF_X1 port map( A => n336, Z => n331);
   U206 : BUF_X1 port map( A => n336, Z => n330);
   U207 : BUF_X1 port map( A => n335, Z => n334);
   U208 : BUF_X1 port map( A => n741, Z => n29);
   U209 : BUF_X1 port map( A => n741, Z => n28);
   U210 : BUF_X1 port map( A => n707, Z => n26);
   U211 : BUF_X1 port map( A => n707, Z => n25);
   U212 : BUF_X1 port map( A => n876, Z => n41);
   U213 : BUF_X1 port map( A => n876, Z => n40);
   U214 : BUF_X1 port map( A => n843, Z => n38);
   U215 : BUF_X1 port map( A => n843, Z => n37);
   U216 : BUF_X1 port map( A => n538, Z => n11);
   U217 : BUF_X1 port map( A => n538, Z => n10);
   U218 : BUF_X1 port map( A => n504, Z => n8);
   U219 : BUF_X1 port map( A => n504, Z => n7);
   U220 : BUF_X1 port map( A => n470, Z => n5);
   U221 : BUF_X1 port map( A => n470, Z => n4);
   U222 : BUF_X1 port map( A => n435, Z => n2);
   U223 : BUF_X1 port map( A => n435, Z => n1);
   U224 : BUF_X1 port map( A => n775, Z => n32);
   U225 : BUF_X1 port map( A => n775, Z => n31);
   U226 : BUF_X1 port map( A => n961, Z => n91);
   U227 : BUF_X1 port map( A => n961, Z => n92);
   U228 : BUF_X1 port map( A => n960, Z => n88);
   U229 : BUF_X1 port map( A => n960, Z => n89);
   U230 : BUF_X1 port map( A => n672, Z => n23);
   U231 : BUF_X1 port map( A => n672, Z => n22);
   U232 : BUF_X1 port map( A => n959, Z => n85);
   U233 : BUF_X1 port map( A => n959, Z => n86);
   U234 : BUF_X1 port map( A => n958, Z => n82);
   U235 : BUF_X1 port map( A => n958, Z => n83);
   U236 : BUF_X1 port map( A => n957, Z => n79);
   U237 : BUF_X1 port map( A => n957, Z => n80);
   U238 : BUF_X1 port map( A => n956, Z => n76);
   U239 : BUF_X1 port map( A => n956, Z => n77);
   U240 : BUF_X1 port map( A => n909, Z => n44);
   U241 : BUF_X1 port map( A => n909, Z => n43);
   U242 : BUF_X1 port map( A => n955, Z => n73);
   U243 : BUF_X1 port map( A => n955, Z => n74);
   U244 : BUF_X1 port map( A => n952, Z => n70);
   U245 : BUF_X1 port map( A => n952, Z => n71);
   U246 : BUF_X1 port map( A => n809, Z => n35);
   U247 : BUF_X1 port map( A => n809, Z => n34);
   U248 : BUF_X1 port map( A => n951, Z => n67);
   U249 : BUF_X1 port map( A => n951, Z => n68);
   U250 : BUF_X1 port map( A => n950, Z => n64);
   U251 : BUF_X1 port map( A => n950, Z => n65);
   U252 : BUF_X1 port map( A => n949, Z => n61);
   U253 : BUF_X1 port map( A => n949, Z => n62);
   U254 : BUF_X1 port map( A => n948, Z => n58);
   U255 : BUF_X1 port map( A => n948, Z => n59);
   U256 : BUF_X1 port map( A => n944, Z => n55);
   U257 : BUF_X1 port map( A => n944, Z => n56);
   U258 : BUF_X1 port map( A => n943, Z => n52);
   U259 : BUF_X1 port map( A => n943, Z => n53);
   U260 : BUF_X1 port map( A => n639, Z => n20);
   U261 : BUF_X1 port map( A => n639, Z => n19);
   U262 : BUF_X1 port map( A => n606, Z => n17);
   U263 : BUF_X1 port map( A => n606, Z => n16);
   U264 : BUF_X1 port map( A => n942, Z => n49);
   U265 : BUF_X1 port map( A => n942, Z => n50);
   U266 : BUF_X1 port map( A => n941, Z => n46);
   U267 : BUF_X1 port map( A => n941, Z => n47);
   U268 : BUF_X1 port map( A => n572, Z => n14);
   U269 : BUF_X1 port map( A => n572, Z => n13);
   U270 : BUF_X1 port map( A => n1824, Z => n199);
   U271 : BUF_X1 port map( A => n1824, Z => n200);
   U272 : BUF_X1 port map( A => n964, Z => n98);
   U273 : BUF_X1 port map( A => n964, Z => n97);
   U274 : BUF_X1 port map( A => n1822, Z => n196);
   U275 : BUF_X1 port map( A => n1822, Z => n197);
   U276 : BUF_X1 port map( A => n962, Z => n95);
   U277 : BUF_X1 port map( A => n962, Z => n94);
   U278 : BUF_X1 port map( A => n876, Z => n42);
   U279 : BUF_X1 port map( A => n843, Z => n39);
   U280 : BUF_X1 port map( A => n538, Z => n12);
   U281 : BUF_X1 port map( A => n504, Z => n9);
   U282 : BUF_X1 port map( A => n470, Z => n6);
   U283 : BUF_X1 port map( A => n435, Z => n3);
   U284 : BUF_X1 port map( A => n961, Z => n93);
   U285 : BUF_X1 port map( A => n960, Z => n90);
   U286 : BUF_X1 port map( A => n959, Z => n87);
   U287 : BUF_X1 port map( A => n707, Z => n27);
   U288 : BUF_X1 port map( A => n775, Z => n33);
   U289 : BUF_X1 port map( A => n672, Z => n24);
   U290 : BUF_X1 port map( A => n958, Z => n84);
   U291 : BUF_X1 port map( A => n957, Z => n81);
   U292 : BUF_X1 port map( A => n956, Z => n78);
   U293 : BUF_X1 port map( A => n909, Z => n45);
   U294 : BUF_X1 port map( A => n955, Z => n75);
   U295 : BUF_X1 port map( A => n952, Z => n72);
   U296 : BUF_X1 port map( A => n809, Z => n36);
   U297 : BUF_X1 port map( A => n639, Z => n21);
   U298 : BUF_X1 port map( A => n606, Z => n18);
   U299 : BUF_X1 port map( A => n572, Z => n15);
   U300 : BUF_X1 port map( A => n741, Z => n30);
   U301 : BUF_X1 port map( A => n951, Z => n69);
   U302 : BUF_X1 port map( A => n950, Z => n66);
   U303 : BUF_X1 port map( A => n949, Z => n63);
   U304 : BUF_X1 port map( A => n948, Z => n60);
   U305 : BUF_X1 port map( A => n944, Z => n57);
   U306 : BUF_X1 port map( A => n943, Z => n54);
   U307 : BUF_X1 port map( A => n942, Z => n51);
   U308 : BUF_X1 port map( A => n941, Z => n48);
   U309 : BUF_X1 port map( A => n1824, Z => n201);
   U310 : BUF_X1 port map( A => n964, Z => n99);
   U311 : BUF_X1 port map( A => n1822, Z => n198);
   U312 : BUF_X1 port map( A => n962, Z => n96);
   U313 : BUF_X1 port map( A => RST, Z => n335);
   U314 : BUF_X1 port map( A => RST, Z => n336);
   U315 : BUF_X1 port map( A => n1825, Z => n202);
   U316 : BUF_X1 port map( A => n965, Z => n100);
   U317 : BUF_X1 port map( A => n1825, Z => n203);
   U318 : BUF_X1 port map( A => n965, Z => n101);
   U319 : BUF_X1 port map( A => n1825, Z => n204);
   U320 : BUF_X1 port map( A => n965, Z => n102);
   U321 : INV_X1 port map( A => DATAIN(0), ZN => n298);
   U322 : INV_X1 port map( A => DATAIN(1), ZN => n299);
   U323 : INV_X1 port map( A => DATAIN(2), ZN => n300);
   U324 : INV_X1 port map( A => DATAIN(3), ZN => n301);
   U325 : INV_X1 port map( A => DATAIN(4), ZN => n302);
   U326 : INV_X1 port map( A => DATAIN(5), ZN => n303);
   U327 : INV_X1 port map( A => DATAIN(6), ZN => n304);
   U328 : INV_X1 port map( A => DATAIN(7), ZN => n305);
   U329 : INV_X1 port map( A => DATAIN(8), ZN => n306);
   U330 : INV_X1 port map( A => DATAIN(10), ZN => n308);
   U331 : INV_X1 port map( A => DATAIN(11), ZN => n309);
   U332 : INV_X1 port map( A => DATAIN(12), ZN => n310);
   U333 : INV_X1 port map( A => DATAIN(13), ZN => n311);
   U334 : INV_X1 port map( A => DATAIN(14), ZN => n312);
   U335 : INV_X1 port map( A => DATAIN(15), ZN => n313);
   U336 : INV_X1 port map( A => DATAIN(16), ZN => n314);
   U337 : INV_X1 port map( A => DATAIN(17), ZN => n315);
   U338 : INV_X1 port map( A => DATAIN(18), ZN => n316);
   U339 : INV_X1 port map( A => DATAIN(19), ZN => n317);
   U340 : INV_X1 port map( A => DATAIN(20), ZN => n318);
   U341 : INV_X1 port map( A => DATAIN(21), ZN => n319);
   U342 : INV_X1 port map( A => DATAIN(22), ZN => n320);
   U343 : INV_X1 port map( A => DATAIN(23), ZN => n321);
   U344 : INV_X1 port map( A => DATAIN(24), ZN => n322);
   U345 : INV_X1 port map( A => DATAIN(25), ZN => n323);
   U346 : INV_X1 port map( A => DATAIN(26), ZN => n324);
   U347 : INV_X1 port map( A => DATAIN(27), ZN => n325);
   U348 : INV_X1 port map( A => DATAIN(28), ZN => n326);
   U349 : INV_X1 port map( A => DATAIN(29), ZN => n327);
   U350 : INV_X1 port map( A => DATAIN(30), ZN => n328);
   U351 : INV_X1 port map( A => DATAIN(31), ZN => n329);
   U352 : INV_X1 port map( A => DATAIN(9), ZN => n307);
   U353 : CLKBUF_X1 port map( A => n433, Z => n337);
   U354 : CLKBUF_X1 port map( A => n433, Z => n338);
   U355 : CLKBUF_X1 port map( A => n433, Z => n339);
   U356 : CLKBUF_X1 port map( A => n433, Z => n340);
   U357 : CLKBUF_X1 port map( A => n433, Z => n341);
   U358 : CLKBUF_X1 port map( A => n432, Z => n342);
   U359 : CLKBUF_X1 port map( A => n432, Z => n343);
   U360 : CLKBUF_X1 port map( A => n432, Z => n344);
   U361 : CLKBUF_X1 port map( A => n432, Z => n345);
   U362 : CLKBUF_X1 port map( A => n432, Z => n346);
   U363 : CLKBUF_X1 port map( A => n432, Z => n347);
   U364 : CLKBUF_X1 port map( A => n431, Z => n348);
   U365 : CLKBUF_X1 port map( A => n431, Z => n349);
   U366 : CLKBUF_X1 port map( A => n431, Z => n350);
   U367 : CLKBUF_X1 port map( A => n431, Z => n351);
   U368 : CLKBUF_X1 port map( A => n431, Z => n352);
   U369 : CLKBUF_X1 port map( A => n431, Z => n353);
   U370 : CLKBUF_X1 port map( A => n430, Z => n354);
   U371 : CLKBUF_X1 port map( A => n430, Z => n355);
   U372 : CLKBUF_X1 port map( A => n430, Z => n356);
   U373 : CLKBUF_X1 port map( A => n430, Z => n357);
   U374 : CLKBUF_X1 port map( A => n430, Z => n358);
   U375 : CLKBUF_X1 port map( A => n430, Z => n359);
   U376 : CLKBUF_X1 port map( A => n429, Z => n360);
   U377 : CLKBUF_X1 port map( A => n429, Z => n361);
   U378 : CLKBUF_X1 port map( A => n429, Z => n362);
   U379 : CLKBUF_X1 port map( A => n429, Z => n363);
   U380 : CLKBUF_X1 port map( A => n429, Z => n364);
   U381 : CLKBUF_X1 port map( A => n429, Z => n365);
   U382 : CLKBUF_X1 port map( A => n428, Z => n366);
   U383 : CLKBUF_X1 port map( A => n428, Z => n367);
   U384 : CLKBUF_X1 port map( A => n428, Z => n368);
   U385 : CLKBUF_X1 port map( A => n428, Z => n369);
   U386 : CLKBUF_X1 port map( A => n428, Z => n370);
   U387 : CLKBUF_X1 port map( A => n428, Z => n371);
   U388 : CLKBUF_X1 port map( A => n427, Z => n372);
   U389 : CLKBUF_X1 port map( A => n427, Z => n373);
   U390 : CLKBUF_X1 port map( A => n427, Z => n374);
   U391 : CLKBUF_X1 port map( A => n427, Z => n375);
   U392 : CLKBUF_X1 port map( A => n427, Z => n376);
   U393 : CLKBUF_X1 port map( A => n427, Z => n377);
   U394 : CLKBUF_X1 port map( A => n426, Z => n378);
   U395 : CLKBUF_X1 port map( A => n426, Z => n379);
   U396 : CLKBUF_X1 port map( A => n426, Z => n380);
   U397 : CLKBUF_X1 port map( A => n426, Z => n381);
   U398 : CLKBUF_X1 port map( A => n426, Z => n382);
   U399 : CLKBUF_X1 port map( A => n426, Z => n383);
   U400 : CLKBUF_X1 port map( A => n425, Z => n384);
   U401 : CLKBUF_X1 port map( A => n425, Z => n385);
   U402 : CLKBUF_X1 port map( A => n425, Z => n386);
   U403 : CLKBUF_X1 port map( A => n425, Z => n387);
   U404 : CLKBUF_X1 port map( A => n425, Z => n388);
   U405 : CLKBUF_X1 port map( A => n425, Z => n389);
   U406 : CLKBUF_X1 port map( A => n424, Z => n390);
   U407 : CLKBUF_X1 port map( A => n424, Z => n391);
   U408 : CLKBUF_X1 port map( A => n424, Z => n392);
   U409 : CLKBUF_X1 port map( A => n424, Z => n393);
   U410 : CLKBUF_X1 port map( A => n424, Z => n394);
   U411 : CLKBUF_X1 port map( A => n424, Z => n395);
   U412 : CLKBUF_X1 port map( A => n423, Z => n396);
   U413 : CLKBUF_X1 port map( A => n423, Z => n397);
   U414 : CLKBUF_X1 port map( A => n423, Z => n398);
   U415 : CLKBUF_X1 port map( A => n423, Z => n399);
   U416 : CLKBUF_X1 port map( A => n423, Z => n400);
   U417 : CLKBUF_X1 port map( A => n423, Z => n401);
   U418 : CLKBUF_X1 port map( A => n422, Z => n402);
   U419 : CLKBUF_X1 port map( A => n422, Z => n403);
   U420 : CLKBUF_X1 port map( A => n422, Z => n404);
   U421 : CLKBUF_X1 port map( A => n422, Z => n405);
   U422 : CLKBUF_X1 port map( A => n422, Z => n406);
   U423 : CLKBUF_X1 port map( A => n422, Z => n407);
   U424 : CLKBUF_X1 port map( A => n421, Z => n408);
   U425 : CLKBUF_X1 port map( A => n421, Z => n409);
   U426 : CLKBUF_X1 port map( A => n421, Z => n410);
   U427 : CLKBUF_X1 port map( A => n421, Z => n411);
   U428 : CLKBUF_X1 port map( A => n421, Z => n412);
   U429 : CLKBUF_X1 port map( A => n421, Z => n413);
   U430 : CLKBUF_X1 port map( A => n420, Z => n414);
   U431 : CLKBUF_X1 port map( A => n420, Z => n415);
   U432 : CLKBUF_X1 port map( A => n420, Z => n416);
   U433 : CLKBUF_X1 port map( A => n420, Z => n417);
   U434 : CLKBUF_X1 port map( A => n420, Z => n418);
   U435 : INV_X1 port map( A => n434, ZN => n3865);
   U436 : MUX2_X1 port map( A => n3721, B => n298, S => n3, Z => n434);
   U437 : INV_X1 port map( A => n436, ZN => n3866);
   U438 : MUX2_X1 port map( A => n3700, B => n299, S => n3, Z => n436);
   U439 : INV_X1 port map( A => n437, ZN => n3867);
   U440 : MUX2_X1 port map( A => n3679, B => n300, S => n3, Z => n437);
   U441 : INV_X1 port map( A => n438, ZN => n3868);
   U442 : MUX2_X1 port map( A => n3658, B => n301, S => n3, Z => n438);
   U443 : INV_X1 port map( A => n439, ZN => n3869);
   U444 : MUX2_X1 port map( A => n3637, B => n302, S => n3, Z => n439);
   U445 : INV_X1 port map( A => n440, ZN => n3870);
   U446 : MUX2_X1 port map( A => n3616, B => n303, S => n3, Z => n440);
   U447 : INV_X1 port map( A => n441, ZN => n3871);
   U448 : MUX2_X1 port map( A => n3595, B => n304, S => n3, Z => n441);
   U449 : INV_X1 port map( A => n442, ZN => n3872);
   U450 : MUX2_X1 port map( A => n3574, B => n305, S => n3, Z => n442);
   U451 : INV_X1 port map( A => n443, ZN => n3873);
   U452 : MUX2_X1 port map( A => n2977, B => n306, S => n2, Z => n443);
   U453 : INV_X1 port map( A => n444, ZN => n3874);
   U454 : MUX2_X1 port map( A => n2956, B => n307, S => n2, Z => n444);
   U455 : INV_X1 port map( A => n445, ZN => n3875);
   U456 : MUX2_X1 port map( A => n2935, B => n308, S => n2, Z => n445);
   U457 : INV_X1 port map( A => n446, ZN => n3876);
   U458 : MUX2_X1 port map( A => n2914, B => n309, S => n2, Z => n446);
   U459 : INV_X1 port map( A => n447, ZN => n3877);
   U460 : MUX2_X1 port map( A => n2893, B => n310, S => n2, Z => n447);
   U461 : INV_X1 port map( A => n448, ZN => n3878);
   U462 : MUX2_X1 port map( A => n2872, B => n311, S => n2, Z => n448);
   U463 : INV_X1 port map( A => n449, ZN => n3879);
   U464 : MUX2_X1 port map( A => n2851, B => n312, S => n2, Z => n449);
   U465 : INV_X1 port map( A => n450, ZN => n3880);
   U466 : MUX2_X1 port map( A => n2830, B => n313, S => n2, Z => n450);
   U467 : INV_X1 port map( A => n451, ZN => n3881);
   U468 : MUX2_X1 port map( A => n2809, B => n314, S => n2, Z => n451);
   U469 : INV_X1 port map( A => n452, ZN => n3882);
   U470 : MUX2_X1 port map( A => n2788, B => n315, S => n2, Z => n452);
   U471 : INV_X1 port map( A => n453, ZN => n3883);
   U472 : MUX2_X1 port map( A => n2767, B => n316, S => n2, Z => n453);
   U473 : INV_X1 port map( A => n454, ZN => n3884);
   U474 : MUX2_X1 port map( A => n2746, B => n317, S => n2, Z => n454);
   U475 : INV_X1 port map( A => n455, ZN => n3885);
   U476 : MUX2_X1 port map( A => n2725, B => n318, S => n1, Z => n455);
   U477 : INV_X1 port map( A => n456, ZN => n3886);
   U478 : MUX2_X1 port map( A => n2704, B => n319, S => n1, Z => n456);
   U479 : INV_X1 port map( A => n457, ZN => n3887);
   U480 : MUX2_X1 port map( A => n2683, B => n320, S => n1, Z => n457);
   U481 : INV_X1 port map( A => n458, ZN => n3888);
   U482 : MUX2_X1 port map( A => n2662, B => n321, S => n1, Z => n458);
   U483 : INV_X1 port map( A => n459, ZN => n3889);
   U484 : MUX2_X1 port map( A => n2641, B => n322, S => n1, Z => n459);
   U485 : INV_X1 port map( A => n460, ZN => n3890);
   U486 : MUX2_X1 port map( A => n2620, B => n323, S => n1, Z => n460);
   U487 : INV_X1 port map( A => n461, ZN => n3891);
   U488 : MUX2_X1 port map( A => n2599, B => n324, S => n1, Z => n461);
   U489 : INV_X1 port map( A => n462, ZN => n3892);
   U490 : MUX2_X1 port map( A => n2578, B => n325, S => n1, Z => n462);
   U491 : INV_X1 port map( A => n463, ZN => n3893);
   U492 : MUX2_X1 port map( A => n2557, B => n326, S => n1, Z => n463);
   U493 : INV_X1 port map( A => n464, ZN => n3894);
   U494 : MUX2_X1 port map( A => n2536, B => n327, S => n1, Z => n464);
   U495 : INV_X1 port map( A => n465, ZN => n3895);
   U496 : MUX2_X1 port map( A => n2515, B => n328, S => n1, Z => n465);
   U497 : INV_X1 port map( A => n466, ZN => n3896);
   U498 : MUX2_X1 port map( A => n2494, B => n329, S => n1, Z => n466);
   U499 : AND2_X1 port map( A1 => n467, A2 => n468, ZN => n435);
   U500 : INV_X1 port map( A => n469, ZN => n3897);
   U501 : MUX2_X1 port map( A => n3722, B => n298, S => n6, Z => n469);
   U502 : INV_X1 port map( A => n471, ZN => n3898);
   U503 : MUX2_X1 port map( A => n3701, B => n299, S => n6, Z => n471);
   U504 : INV_X1 port map( A => n472, ZN => n3899);
   U505 : MUX2_X1 port map( A => n3680, B => n300, S => n6, Z => n472);
   U506 : INV_X1 port map( A => n473, ZN => n3900);
   U507 : MUX2_X1 port map( A => n3659, B => n301, S => n6, Z => n473);
   U508 : INV_X1 port map( A => n474, ZN => n3901);
   U509 : MUX2_X1 port map( A => n3638, B => n302, S => n6, Z => n474);
   U510 : INV_X1 port map( A => n475, ZN => n3902);
   U511 : MUX2_X1 port map( A => n3617, B => n303, S => n6, Z => n475);
   U512 : INV_X1 port map( A => n476, ZN => n3903);
   U513 : MUX2_X1 port map( A => n3596, B => n304, S => n6, Z => n476);
   U514 : INV_X1 port map( A => n477, ZN => n3904);
   U515 : MUX2_X1 port map( A => n3575, B => n305, S => n6, Z => n477);
   U516 : INV_X1 port map( A => n478, ZN => n3905);
   U517 : MUX2_X1 port map( A => n2978, B => n306, S => n5, Z => n478);
   U518 : INV_X1 port map( A => n479, ZN => n3906);
   U519 : MUX2_X1 port map( A => n2957, B => n307, S => n5, Z => n479);
   U520 : INV_X1 port map( A => n480, ZN => n3907);
   U521 : MUX2_X1 port map( A => n2936, B => n308, S => n5, Z => n480);
   U522 : INV_X1 port map( A => n481, ZN => n3908);
   U523 : MUX2_X1 port map( A => n2915, B => n309, S => n5, Z => n481);
   U524 : INV_X1 port map( A => n482, ZN => n3909);
   U525 : MUX2_X1 port map( A => n2894, B => n310, S => n5, Z => n482);
   U526 : INV_X1 port map( A => n483, ZN => n3910);
   U527 : MUX2_X1 port map( A => n2873, B => n311, S => n5, Z => n483);
   U528 : INV_X1 port map( A => n484, ZN => n3911);
   U529 : MUX2_X1 port map( A => n2852, B => n312, S => n5, Z => n484);
   U530 : INV_X1 port map( A => n485, ZN => n3912);
   U531 : MUX2_X1 port map( A => n2831, B => n313, S => n5, Z => n485);
   U532 : INV_X1 port map( A => n486, ZN => n3913);
   U533 : MUX2_X1 port map( A => n2810, B => n314, S => n5, Z => n486);
   U534 : INV_X1 port map( A => n487, ZN => n3914);
   U535 : MUX2_X1 port map( A => n2789, B => n315, S => n5, Z => n487);
   U536 : INV_X1 port map( A => n488, ZN => n3915);
   U537 : MUX2_X1 port map( A => n2768, B => n316, S => n5, Z => n488);
   U538 : INV_X1 port map( A => n489, ZN => n3916);
   U539 : MUX2_X1 port map( A => n2747, B => n317, S => n5, Z => n489);
   U540 : INV_X1 port map( A => n490, ZN => n3917);
   U541 : MUX2_X1 port map( A => n2726, B => n318, S => n4, Z => n490);
   U542 : INV_X1 port map( A => n491, ZN => n3918);
   U543 : MUX2_X1 port map( A => n2705, B => n319, S => n4, Z => n491);
   U544 : INV_X1 port map( A => n492, ZN => n3919);
   U545 : MUX2_X1 port map( A => n2684, B => n320, S => n4, Z => n492);
   U546 : INV_X1 port map( A => n493, ZN => n3920);
   U547 : MUX2_X1 port map( A => n2663, B => n321, S => n4, Z => n493);
   U548 : INV_X1 port map( A => n494, ZN => n3921);
   U549 : MUX2_X1 port map( A => n2642, B => n322, S => n4, Z => n494);
   U550 : INV_X1 port map( A => n495, ZN => n3922);
   U551 : MUX2_X1 port map( A => n2621, B => n323, S => n4, Z => n495);
   U552 : INV_X1 port map( A => n496, ZN => n3923);
   U553 : MUX2_X1 port map( A => n2600, B => n324, S => n4, Z => n496);
   U554 : INV_X1 port map( A => n497, ZN => n3924);
   U555 : MUX2_X1 port map( A => n2579, B => n325, S => n4, Z => n497);
   U556 : INV_X1 port map( A => n498, ZN => n3925);
   U557 : MUX2_X1 port map( A => n2558, B => n326, S => n4, Z => n498);
   U558 : INV_X1 port map( A => n499, ZN => n3926);
   U559 : MUX2_X1 port map( A => n2537, B => n327, S => n4, Z => n499);
   U560 : INV_X1 port map( A => n500, ZN => n3927);
   U561 : MUX2_X1 port map( A => n2516, B => n328, S => n4, Z => n500);
   U562 : INV_X1 port map( A => n501, ZN => n3928);
   U563 : MUX2_X1 port map( A => n2495, B => n329, S => n4, Z => n501);
   U564 : AND2_X1 port map( A1 => n502, A2 => n467, ZN => n470);
   U565 : INV_X1 port map( A => n503, ZN => n3929);
   U566 : MUX2_X1 port map( A => n3717, B => n298, S => n9, Z => n503);
   U567 : INV_X1 port map( A => n505, ZN => n3930);
   U568 : MUX2_X1 port map( A => n3696, B => n299, S => n9, Z => n505);
   U569 : INV_X1 port map( A => n506, ZN => n3931);
   U570 : MUX2_X1 port map( A => n3675, B => n300, S => n9, Z => n506);
   U571 : INV_X1 port map( A => n507, ZN => n3932);
   U572 : MUX2_X1 port map( A => n3654, B => n301, S => n9, Z => n507);
   U573 : INV_X1 port map( A => n508, ZN => n3933);
   U574 : MUX2_X1 port map( A => n3633, B => n302, S => n9, Z => n508);
   U575 : INV_X1 port map( A => n509, ZN => n3934);
   U576 : MUX2_X1 port map( A => n3612, B => n303, S => n9, Z => n509);
   U577 : INV_X1 port map( A => n510, ZN => n3935);
   U578 : MUX2_X1 port map( A => n3591, B => n304, S => n9, Z => n510);
   U579 : INV_X1 port map( A => n511, ZN => n3936);
   U580 : MUX2_X1 port map( A => n3570, B => n305, S => n9, Z => n511);
   U581 : INV_X1 port map( A => n512, ZN => n3937);
   U582 : MUX2_X1 port map( A => n2973, B => n306, S => n8, Z => n512);
   U583 : INV_X1 port map( A => n513, ZN => n3938);
   U584 : MUX2_X1 port map( A => n2952, B => n307, S => n8, Z => n513);
   U585 : INV_X1 port map( A => n514, ZN => n3939);
   U586 : MUX2_X1 port map( A => n2931, B => n308, S => n8, Z => n514);
   U587 : INV_X1 port map( A => n515, ZN => n3940);
   U588 : MUX2_X1 port map( A => n2910, B => n309, S => n8, Z => n515);
   U589 : INV_X1 port map( A => n516, ZN => n3941);
   U590 : MUX2_X1 port map( A => n2889, B => n310, S => n8, Z => n516);
   U591 : INV_X1 port map( A => n517, ZN => n3942);
   U592 : MUX2_X1 port map( A => n2868, B => n311, S => n8, Z => n517);
   U593 : INV_X1 port map( A => n518, ZN => n3943);
   U594 : MUX2_X1 port map( A => n2847, B => n312, S => n8, Z => n518);
   U595 : INV_X1 port map( A => n519, ZN => n3944);
   U596 : MUX2_X1 port map( A => n2826, B => n313, S => n8, Z => n519);
   U597 : INV_X1 port map( A => n520, ZN => n3945);
   U598 : MUX2_X1 port map( A => n2805, B => n314, S => n8, Z => n520);
   U599 : INV_X1 port map( A => n521, ZN => n3946);
   U600 : MUX2_X1 port map( A => n2784, B => n315, S => n8, Z => n521);
   U601 : INV_X1 port map( A => n522, ZN => n3947);
   U602 : MUX2_X1 port map( A => n2763, B => n316, S => n8, Z => n522);
   U603 : INV_X1 port map( A => n523, ZN => n3948);
   U604 : MUX2_X1 port map( A => n2742, B => n317, S => n8, Z => n523);
   U605 : INV_X1 port map( A => n524, ZN => n3949);
   U606 : MUX2_X1 port map( A => n2721, B => n318, S => n7, Z => n524);
   U607 : INV_X1 port map( A => n525, ZN => n3950);
   U608 : MUX2_X1 port map( A => n2700, B => n319, S => n7, Z => n525);
   U609 : INV_X1 port map( A => n526, ZN => n3951);
   U610 : MUX2_X1 port map( A => n2679, B => n320, S => n7, Z => n526);
   U611 : INV_X1 port map( A => n527, ZN => n3952);
   U612 : MUX2_X1 port map( A => n2658, B => n321, S => n7, Z => n527);
   U613 : INV_X1 port map( A => n528, ZN => n3953);
   U614 : MUX2_X1 port map( A => n2637, B => n322, S => n7, Z => n528);
   U615 : INV_X1 port map( A => n529, ZN => n3954);
   U616 : MUX2_X1 port map( A => n2616, B => n323, S => n7, Z => n529);
   U617 : INV_X1 port map( A => n530, ZN => n3955);
   U618 : MUX2_X1 port map( A => n2595, B => n324, S => n7, Z => n530);
   U619 : INV_X1 port map( A => n531, ZN => n3956);
   U620 : MUX2_X1 port map( A => n2574, B => n325, S => n7, Z => n531);
   U621 : INV_X1 port map( A => n532, ZN => n3957);
   U622 : MUX2_X1 port map( A => n2553, B => n326, S => n7, Z => n532);
   U623 : INV_X1 port map( A => n533, ZN => n3958);
   U624 : MUX2_X1 port map( A => n2532, B => n327, S => n7, Z => n533);
   U625 : INV_X1 port map( A => n534, ZN => n3959);
   U626 : MUX2_X1 port map( A => n2511, B => n328, S => n7, Z => n534);
   U627 : INV_X1 port map( A => n535, ZN => n3960);
   U628 : MUX2_X1 port map( A => n2490, B => n329, S => n7, Z => n535);
   U629 : AND2_X1 port map( A1 => n536, A2 => n467, ZN => n504);
   U630 : INV_X1 port map( A => n537, ZN => n3961);
   U631 : MUX2_X1 port map( A => n3718, B => n298, S => n12, Z => n537);
   U632 : INV_X1 port map( A => n539, ZN => n3962);
   U633 : MUX2_X1 port map( A => n3697, B => n299, S => n12, Z => n539);
   U634 : INV_X1 port map( A => n540, ZN => n3963);
   U635 : MUX2_X1 port map( A => n3676, B => n300, S => n12, Z => n540);
   U636 : INV_X1 port map( A => n541, ZN => n3964);
   U637 : MUX2_X1 port map( A => n3655, B => n301, S => n12, Z => n541);
   U638 : INV_X1 port map( A => n542, ZN => n3965);
   U639 : MUX2_X1 port map( A => n3634, B => n302, S => n12, Z => n542);
   U640 : INV_X1 port map( A => n543, ZN => n3966);
   U641 : MUX2_X1 port map( A => n3613, B => n303, S => n12, Z => n543);
   U642 : INV_X1 port map( A => n544, ZN => n3967);
   U643 : MUX2_X1 port map( A => n3592, B => n304, S => n12, Z => n544);
   U644 : INV_X1 port map( A => n545, ZN => n3968);
   U645 : MUX2_X1 port map( A => n3571, B => n305, S => n12, Z => n545);
   U646 : INV_X1 port map( A => n546, ZN => n3969);
   U647 : MUX2_X1 port map( A => n2974, B => n306, S => n11, Z => n546);
   U648 : INV_X1 port map( A => n547, ZN => n3970);
   U649 : MUX2_X1 port map( A => n2953, B => n307, S => n11, Z => n547);
   U650 : INV_X1 port map( A => n548, ZN => n3971);
   U651 : MUX2_X1 port map( A => n2932, B => n308, S => n11, Z => n548);
   U652 : INV_X1 port map( A => n549, ZN => n3972);
   U653 : MUX2_X1 port map( A => n2911, B => n309, S => n11, Z => n549);
   U654 : INV_X1 port map( A => n550, ZN => n3973);
   U655 : MUX2_X1 port map( A => n2890, B => n310, S => n11, Z => n550);
   U656 : INV_X1 port map( A => n551, ZN => n3974);
   U657 : MUX2_X1 port map( A => n2869, B => n311, S => n11, Z => n551);
   U658 : INV_X1 port map( A => n552, ZN => n3975);
   U659 : MUX2_X1 port map( A => n2848, B => n312, S => n11, Z => n552);
   U660 : INV_X1 port map( A => n553, ZN => n3976);
   U661 : MUX2_X1 port map( A => n2827, B => n313, S => n11, Z => n553);
   U662 : INV_X1 port map( A => n554, ZN => n3977);
   U663 : MUX2_X1 port map( A => n2806, B => n314, S => n11, Z => n554);
   U664 : INV_X1 port map( A => n555, ZN => n3978);
   U665 : MUX2_X1 port map( A => n2785, B => n315, S => n11, Z => n555);
   U666 : INV_X1 port map( A => n556, ZN => n3979);
   U667 : MUX2_X1 port map( A => n2764, B => n316, S => n11, Z => n556);
   U668 : INV_X1 port map( A => n557, ZN => n3980);
   U669 : MUX2_X1 port map( A => n2743, B => n317, S => n11, Z => n557);
   U670 : INV_X1 port map( A => n558, ZN => n3981);
   U671 : MUX2_X1 port map( A => n2722, B => n318, S => n10, Z => n558);
   U672 : INV_X1 port map( A => n559, ZN => n3982);
   U673 : MUX2_X1 port map( A => n2701, B => n319, S => n10, Z => n559);
   U674 : INV_X1 port map( A => n560, ZN => n3983);
   U675 : MUX2_X1 port map( A => n2680, B => n320, S => n10, Z => n560);
   U676 : INV_X1 port map( A => n561, ZN => n3984);
   U677 : MUX2_X1 port map( A => n2659, B => n321, S => n10, Z => n561);
   U678 : INV_X1 port map( A => n562, ZN => n3985);
   U679 : MUX2_X1 port map( A => n2638, B => n322, S => n10, Z => n562);
   U680 : INV_X1 port map( A => n563, ZN => n3986);
   U681 : MUX2_X1 port map( A => n2617, B => n323, S => n10, Z => n563);
   U682 : INV_X1 port map( A => n564, ZN => n3987);
   U683 : MUX2_X1 port map( A => n2596, B => n324, S => n10, Z => n564);
   U684 : INV_X1 port map( A => n565, ZN => n3988);
   U685 : MUX2_X1 port map( A => n2575, B => n325, S => n10, Z => n565);
   U686 : INV_X1 port map( A => n566, ZN => n3989);
   U687 : MUX2_X1 port map( A => n2554, B => n326, S => n10, Z => n566);
   U688 : INV_X1 port map( A => n567, ZN => n3990);
   U689 : MUX2_X1 port map( A => n2533, B => n327, S => n10, Z => n567);
   U690 : INV_X1 port map( A => n568, ZN => n3991);
   U691 : MUX2_X1 port map( A => n2512, B => n328, S => n10, Z => n568);
   U692 : INV_X1 port map( A => n569, ZN => n3992);
   U693 : MUX2_X1 port map( A => n2491, B => n329, S => n10, Z => n569);
   U694 : AND2_X1 port map( A1 => n570, A2 => n467, ZN => n538);
   U695 : MUX2_X1 port map( A => n571, B => DATAIN(0), S => n15, Z => n3993);
   U696 : MUX2_X1 port map( A => n573, B => DATAIN(1), S => n15, Z => n3994);
   U697 : MUX2_X1 port map( A => n574, B => DATAIN(2), S => n15, Z => n3995);
   U698 : MUX2_X1 port map( A => n575, B => DATAIN(3), S => n15, Z => n3996);
   U699 : MUX2_X1 port map( A => n576, B => DATAIN(4), S => n15, Z => n3997);
   U700 : MUX2_X1 port map( A => n577, B => DATAIN(5), S => n15, Z => n3998);
   U701 : MUX2_X1 port map( A => n578, B => DATAIN(6), S => n15, Z => n3999);
   U702 : MUX2_X1 port map( A => n579, B => DATAIN(7), S => n15, Z => n4000);
   U703 : MUX2_X1 port map( A => n580, B => DATAIN(8), S => n14, Z => n4001);
   U704 : MUX2_X1 port map( A => n581, B => DATAIN(9), S => n14, Z => n4002);
   U705 : MUX2_X1 port map( A => n582, B => DATAIN(10), S => n14, Z => n4003);
   U706 : MUX2_X1 port map( A => n583, B => DATAIN(11), S => n14, Z => n4004);
   U707 : MUX2_X1 port map( A => n584, B => DATAIN(12), S => n14, Z => n4005);
   U708 : MUX2_X1 port map( A => n585, B => DATAIN(13), S => n14, Z => n4006);
   U709 : MUX2_X1 port map( A => n586, B => DATAIN(14), S => n14, Z => n4007);
   U710 : MUX2_X1 port map( A => n587, B => DATAIN(15), S => n14, Z => n4008);
   U711 : MUX2_X1 port map( A => n588, B => DATAIN(16), S => n14, Z => n4009);
   U712 : MUX2_X1 port map( A => n589, B => DATAIN(17), S => n14, Z => n4010);
   U713 : MUX2_X1 port map( A => n590, B => DATAIN(18), S => n14, Z => n4011);
   U714 : MUX2_X1 port map( A => n591, B => DATAIN(19), S => n14, Z => n4012);
   U715 : MUX2_X1 port map( A => n592, B => DATAIN(20), S => n13, Z => n4013);
   U716 : MUX2_X1 port map( A => n593, B => DATAIN(21), S => n13, Z => n4014);
   U717 : MUX2_X1 port map( A => n594, B => DATAIN(22), S => n13, Z => n4015);
   U718 : MUX2_X1 port map( A => n595, B => DATAIN(23), S => n13, Z => n4016);
   U719 : MUX2_X1 port map( A => n596, B => DATAIN(24), S => n13, Z => n4017);
   U720 : MUX2_X1 port map( A => n597, B => DATAIN(25), S => n13, Z => n4018);
   U721 : MUX2_X1 port map( A => n598, B => DATAIN(26), S => n13, Z => n4019);
   U722 : MUX2_X1 port map( A => n599, B => DATAIN(27), S => n13, Z => n4020);
   U723 : MUX2_X1 port map( A => n600, B => DATAIN(28), S => n13, Z => n4021);
   U724 : MUX2_X1 port map( A => n601, B => DATAIN(29), S => n13, Z => n4022);
   U725 : MUX2_X1 port map( A => n602, B => DATAIN(30), S => n13, Z => n4023);
   U726 : MUX2_X1 port map( A => n603, B => DATAIN(31), S => n13, Z => n4024);
   U727 : AND2_X1 port map( A1 => n604, A2 => n502, ZN => n572);
   U728 : MUX2_X1 port map( A => n605, B => DATAIN(0), S => n18, Z => n4025);
   U729 : MUX2_X1 port map( A => n607, B => DATAIN(1), S => n18, Z => n4026);
   U730 : MUX2_X1 port map( A => n608, B => DATAIN(2), S => n18, Z => n4027);
   U731 : MUX2_X1 port map( A => n609, B => DATAIN(3), S => n18, Z => n4028);
   U732 : MUX2_X1 port map( A => n610, B => DATAIN(4), S => n18, Z => n4029);
   U733 : MUX2_X1 port map( A => n611, B => DATAIN(5), S => n18, Z => n4030);
   U734 : MUX2_X1 port map( A => n612, B => DATAIN(6), S => n18, Z => n4031);
   U735 : MUX2_X1 port map( A => n613, B => DATAIN(7), S => n18, Z => n4032);
   U736 : MUX2_X1 port map( A => n614, B => DATAIN(8), S => n17, Z => n4033);
   U737 : MUX2_X1 port map( A => n615, B => DATAIN(9), S => n17, Z => n4034);
   U738 : MUX2_X1 port map( A => n616, B => DATAIN(10), S => n17, Z => n4035);
   U739 : MUX2_X1 port map( A => n617, B => DATAIN(11), S => n17, Z => n4036);
   U740 : MUX2_X1 port map( A => n618, B => DATAIN(12), S => n17, Z => n4037);
   U741 : MUX2_X1 port map( A => n619, B => DATAIN(13), S => n17, Z => n4038);
   U742 : MUX2_X1 port map( A => n620, B => DATAIN(14), S => n17, Z => n4039);
   U743 : MUX2_X1 port map( A => n621, B => DATAIN(15), S => n17, Z => n4040);
   U744 : MUX2_X1 port map( A => n622, B => DATAIN(16), S => n17, Z => n4041);
   U745 : MUX2_X1 port map( A => n623, B => DATAIN(17), S => n17, Z => n4042);
   U746 : MUX2_X1 port map( A => n624, B => DATAIN(18), S => n17, Z => n4043);
   U747 : MUX2_X1 port map( A => n625, B => DATAIN(19), S => n17, Z => n4044);
   U748 : MUX2_X1 port map( A => n626, B => DATAIN(20), S => n16, Z => n4045);
   U749 : MUX2_X1 port map( A => n627, B => DATAIN(21), S => n16, Z => n4046);
   U750 : MUX2_X1 port map( A => n628, B => DATAIN(22), S => n16, Z => n4047);
   U751 : MUX2_X1 port map( A => n629, B => DATAIN(23), S => n16, Z => n4048);
   U752 : MUX2_X1 port map( A => n630, B => DATAIN(24), S => n16, Z => n4049);
   U753 : MUX2_X1 port map( A => n631, B => DATAIN(25), S => n16, Z => n4050);
   U754 : MUX2_X1 port map( A => n632, B => DATAIN(26), S => n16, Z => n4051);
   U755 : MUX2_X1 port map( A => n633, B => DATAIN(27), S => n16, Z => n4052);
   U756 : MUX2_X1 port map( A => n634, B => DATAIN(28), S => n16, Z => n4053);
   U757 : MUX2_X1 port map( A => n635, B => DATAIN(29), S => n16, Z => n4054);
   U758 : MUX2_X1 port map( A => n636, B => DATAIN(30), S => n16, Z => n4055);
   U759 : MUX2_X1 port map( A => n637, B => DATAIN(31), S => n16, Z => n4056);
   U760 : AND2_X1 port map( A1 => n604, A2 => n536, ZN => n606);
   U761 : MUX2_X1 port map( A => n638, B => DATAIN(0), S => n21, Z => n4057);
   U762 : MUX2_X1 port map( A => n640, B => DATAIN(1), S => n21, Z => n4058);
   U763 : MUX2_X1 port map( A => n641, B => DATAIN(2), S => n21, Z => n4059);
   U764 : MUX2_X1 port map( A => n642, B => DATAIN(3), S => n21, Z => n4060);
   U765 : MUX2_X1 port map( A => n643, B => DATAIN(4), S => n21, Z => n4061);
   U766 : MUX2_X1 port map( A => n644, B => DATAIN(5), S => n21, Z => n4062);
   U767 : MUX2_X1 port map( A => n645, B => DATAIN(6), S => n21, Z => n4063);
   U768 : MUX2_X1 port map( A => n646, B => DATAIN(7), S => n21, Z => n4064);
   U769 : MUX2_X1 port map( A => n647, B => DATAIN(8), S => n20, Z => n4065);
   U770 : MUX2_X1 port map( A => n648, B => DATAIN(9), S => n20, Z => n4066);
   U771 : MUX2_X1 port map( A => n649, B => DATAIN(10), S => n20, Z => n4067);
   U772 : MUX2_X1 port map( A => n650, B => DATAIN(11), S => n20, Z => n4068);
   U773 : MUX2_X1 port map( A => n651, B => DATAIN(12), S => n20, Z => n4069);
   U774 : MUX2_X1 port map( A => n652, B => DATAIN(13), S => n20, Z => n4070);
   U775 : MUX2_X1 port map( A => n653, B => DATAIN(14), S => n20, Z => n4071);
   U776 : MUX2_X1 port map( A => n654, B => DATAIN(15), S => n20, Z => n4072);
   U777 : MUX2_X1 port map( A => n655, B => DATAIN(16), S => n20, Z => n4073);
   U778 : MUX2_X1 port map( A => n656, B => DATAIN(17), S => n20, Z => n4074);
   U779 : MUX2_X1 port map( A => n657, B => DATAIN(18), S => n20, Z => n4075);
   U780 : MUX2_X1 port map( A => n658, B => DATAIN(19), S => n20, Z => n4076);
   U781 : MUX2_X1 port map( A => n659, B => DATAIN(20), S => n19, Z => n4077);
   U782 : MUX2_X1 port map( A => n660, B => DATAIN(21), S => n19, Z => n4078);
   U783 : MUX2_X1 port map( A => n661, B => DATAIN(22), S => n19, Z => n4079);
   U784 : MUX2_X1 port map( A => n662, B => DATAIN(23), S => n19, Z => n4080);
   U785 : MUX2_X1 port map( A => n663, B => DATAIN(24), S => n19, Z => n4081);
   U786 : MUX2_X1 port map( A => n664, B => DATAIN(25), S => n19, Z => n4082);
   U787 : MUX2_X1 port map( A => n665, B => DATAIN(26), S => n19, Z => n4083);
   U788 : MUX2_X1 port map( A => n666, B => DATAIN(27), S => n19, Z => n4084);
   U789 : MUX2_X1 port map( A => n667, B => DATAIN(28), S => n19, Z => n4085);
   U790 : MUX2_X1 port map( A => n668, B => DATAIN(29), S => n19, Z => n4086);
   U791 : MUX2_X1 port map( A => n669, B => DATAIN(30), S => n19, Z => n4087);
   U792 : MUX2_X1 port map( A => n670, B => DATAIN(31), S => n19, Z => n4088);
   U793 : AND2_X1 port map( A1 => n604, A2 => n570, ZN => n639);
   U794 : MUX2_X1 port map( A => n671, B => DATAIN(31), S => n24, Z => n4089);
   U795 : MUX2_X1 port map( A => n673, B => DATAIN(0), S => n24, Z => n4090);
   U796 : MUX2_X1 port map( A => n674, B => DATAIN(1), S => n24, Z => n4091);
   U797 : MUX2_X1 port map( A => n675, B => DATAIN(2), S => n24, Z => n4092);
   U798 : MUX2_X1 port map( A => n676, B => DATAIN(3), S => n24, Z => n4093);
   U799 : MUX2_X1 port map( A => n677, B => DATAIN(4), S => n24, Z => n4094);
   U800 : MUX2_X1 port map( A => n678, B => DATAIN(5), S => n24, Z => n4095);
   U801 : MUX2_X1 port map( A => n679, B => DATAIN(6), S => n24, Z => n4096);
   U802 : MUX2_X1 port map( A => n680, B => DATAIN(7), S => n23, Z => n4097);
   U803 : MUX2_X1 port map( A => n681, B => DATAIN(8), S => n23, Z => n4098);
   U804 : MUX2_X1 port map( A => n682, B => DATAIN(9), S => n23, Z => n4099);
   U805 : MUX2_X1 port map( A => n683, B => DATAIN(10), S => n23, Z => n4100);
   U806 : MUX2_X1 port map( A => n684, B => DATAIN(11), S => n23, Z => n4101);
   U807 : MUX2_X1 port map( A => n685, B => DATAIN(12), S => n23, Z => n4102);
   U808 : MUX2_X1 port map( A => n686, B => DATAIN(13), S => n23, Z => n4103);
   U809 : MUX2_X1 port map( A => n687, B => DATAIN(14), S => n23, Z => n4104);
   U810 : MUX2_X1 port map( A => n688, B => DATAIN(15), S => n23, Z => n4105);
   U811 : MUX2_X1 port map( A => n689, B => DATAIN(16), S => n23, Z => n4106);
   U812 : MUX2_X1 port map( A => n690, B => DATAIN(17), S => n23, Z => n4107);
   U813 : MUX2_X1 port map( A => n691, B => DATAIN(18), S => n23, Z => n4108);
   U814 : MUX2_X1 port map( A => n692, B => DATAIN(19), S => n22, Z => n4109);
   U815 : MUX2_X1 port map( A => n693, B => DATAIN(20), S => n22, Z => n4110);
   U816 : MUX2_X1 port map( A => n694, B => DATAIN(21), S => n22, Z => n4111);
   U817 : MUX2_X1 port map( A => n695, B => DATAIN(22), S => n22, Z => n4112);
   U818 : MUX2_X1 port map( A => n696, B => DATAIN(23), S => n22, Z => n4113);
   U819 : MUX2_X1 port map( A => n697, B => DATAIN(24), S => n22, Z => n4114);
   U820 : MUX2_X1 port map( A => n698, B => DATAIN(25), S => n22, Z => n4115);
   U821 : MUX2_X1 port map( A => n699, B => DATAIN(26), S => n22, Z => n4116);
   U822 : MUX2_X1 port map( A => n700, B => DATAIN(27), S => n22, Z => n4117);
   U823 : MUX2_X1 port map( A => n701, B => DATAIN(28), S => n22, Z => n4118);
   U824 : MUX2_X1 port map( A => n702, B => DATAIN(29), S => n22, Z => n4119);
   U825 : MUX2_X1 port map( A => n703, B => DATAIN(30), S => n22, Z => n4120);
   U826 : AND2_X1 port map( A1 => n704, A2 => n705, ZN => n672);
   U827 : INV_X1 port map( A => n706, ZN => n4121);
   U828 : MUX2_X1 port map( A => n3833, B => n298, S => n27, Z => n706);
   U829 : INV_X1 port map( A => n708, ZN => n4122);
   U830 : MUX2_X1 port map( A => n3834, B => n299, S => n27, Z => n708);
   U831 : INV_X1 port map( A => n709, ZN => n4123);
   U832 : MUX2_X1 port map( A => n3835, B => n300, S => n27, Z => n709);
   U833 : INV_X1 port map( A => n710, ZN => n4124);
   U834 : MUX2_X1 port map( A => n3836, B => n301, S => n27, Z => n710);
   U835 : INV_X1 port map( A => n711, ZN => n4125);
   U836 : MUX2_X1 port map( A => n3837, B => n302, S => n27, Z => n711);
   U837 : INV_X1 port map( A => n712, ZN => n4126);
   U838 : MUX2_X1 port map( A => n3838, B => n303, S => n27, Z => n712);
   U839 : INV_X1 port map( A => n713, ZN => n4127);
   U840 : MUX2_X1 port map( A => n3839, B => n304, S => n27, Z => n713);
   U841 : INV_X1 port map( A => n714, ZN => n4128);
   U842 : MUX2_X1 port map( A => n3840, B => n305, S => n27, Z => n714);
   U843 : INV_X1 port map( A => n715, ZN => n4129);
   U844 : MUX2_X1 port map( A => n3841, B => n306, S => n26, Z => n715);
   U845 : INV_X1 port map( A => n716, ZN => n4130);
   U846 : MUX2_X1 port map( A => n3842, B => n307, S => n26, Z => n716);
   U847 : INV_X1 port map( A => n717, ZN => n4131);
   U848 : MUX2_X1 port map( A => n3843, B => n308, S => n26, Z => n717);
   U849 : INV_X1 port map( A => n718, ZN => n4132);
   U850 : MUX2_X1 port map( A => n3844, B => n309, S => n26, Z => n718);
   U851 : INV_X1 port map( A => n719, ZN => n4133);
   U852 : MUX2_X1 port map( A => n3845, B => n310, S => n26, Z => n719);
   U853 : INV_X1 port map( A => n720, ZN => n4134);
   U854 : MUX2_X1 port map( A => n3846, B => n311, S => n26, Z => n720);
   U855 : INV_X1 port map( A => n721, ZN => n4135);
   U856 : MUX2_X1 port map( A => n3847, B => n312, S => n26, Z => n721);
   U857 : INV_X1 port map( A => n722, ZN => n4136);
   U858 : MUX2_X1 port map( A => n3848, B => n313, S => n26, Z => n722);
   U859 : INV_X1 port map( A => n723, ZN => n4137);
   U860 : MUX2_X1 port map( A => n3849, B => n314, S => n26, Z => n723);
   U861 : INV_X1 port map( A => n724, ZN => n4138);
   U862 : MUX2_X1 port map( A => n3850, B => n315, S => n26, Z => n724);
   U863 : INV_X1 port map( A => n725, ZN => n4139);
   U864 : MUX2_X1 port map( A => n3851, B => n316, S => n26, Z => n725);
   U865 : INV_X1 port map( A => n726, ZN => n4140);
   U866 : MUX2_X1 port map( A => n3852, B => n317, S => n26, Z => n726);
   U867 : INV_X1 port map( A => n727, ZN => n4141);
   U868 : MUX2_X1 port map( A => n3853, B => n318, S => n25, Z => n727);
   U869 : INV_X1 port map( A => n728, ZN => n4142);
   U870 : MUX2_X1 port map( A => n3854, B => n319, S => n25, Z => n728);
   U871 : INV_X1 port map( A => n729, ZN => n4143);
   U872 : MUX2_X1 port map( A => n3855, B => n320, S => n25, Z => n729);
   U873 : INV_X1 port map( A => n730, ZN => n4144);
   U874 : MUX2_X1 port map( A => n3856, B => n321, S => n25, Z => n730);
   U875 : INV_X1 port map( A => n731, ZN => n4145);
   U876 : MUX2_X1 port map( A => n3857, B => n322, S => n25, Z => n731);
   U877 : INV_X1 port map( A => n732, ZN => n4146);
   U878 : MUX2_X1 port map( A => n3858, B => n323, S => n25, Z => n732);
   U879 : INV_X1 port map( A => n733, ZN => n4147);
   U880 : MUX2_X1 port map( A => n3859, B => n324, S => n25, Z => n733);
   U881 : INV_X1 port map( A => n734, ZN => n4148);
   U882 : MUX2_X1 port map( A => n3860, B => n325, S => n25, Z => n734);
   U883 : INV_X1 port map( A => n735, ZN => n4149);
   U884 : MUX2_X1 port map( A => n3861, B => n326, S => n25, Z => n735);
   U885 : INV_X1 port map( A => n736, ZN => n4150);
   U886 : MUX2_X1 port map( A => n3862, B => n327, S => n25, Z => n736);
   U887 : INV_X1 port map( A => n737, ZN => n4151);
   U888 : MUX2_X1 port map( A => n3863, B => n328, S => n25, Z => n737);
   U889 : INV_X1 port map( A => n738, ZN => n4152);
   U890 : MUX2_X1 port map( A => n3864, B => n329, S => n25, Z => n738);
   U891 : AND2_X1 port map( A1 => n739, A2 => n704, ZN => n707);
   U892 : INV_X1 port map( A => n740, ZN => n4153);
   U893 : MUX2_X1 port map( A => n3737, B => n298, S => n30, Z => n740);
   U894 : INV_X1 port map( A => n742, ZN => n4154);
   U895 : MUX2_X1 port map( A => n3738, B => n299, S => n30, Z => n742);
   U896 : INV_X1 port map( A => n743, ZN => n4155);
   U897 : MUX2_X1 port map( A => n3739, B => n300, S => n30, Z => n743);
   U898 : INV_X1 port map( A => n744, ZN => n4156);
   U899 : MUX2_X1 port map( A => n3740, B => n301, S => n30, Z => n744);
   U900 : INV_X1 port map( A => n745, ZN => n4157);
   U901 : MUX2_X1 port map( A => n3741, B => n302, S => n30, Z => n745);
   U902 : INV_X1 port map( A => n746, ZN => n4158);
   U903 : MUX2_X1 port map( A => n3742, B => n303, S => n30, Z => n746);
   U904 : INV_X1 port map( A => n747, ZN => n4159);
   U905 : MUX2_X1 port map( A => n3743, B => n304, S => n30, Z => n747);
   U906 : INV_X1 port map( A => n748, ZN => n4160);
   U907 : MUX2_X1 port map( A => n3744, B => n305, S => n30, Z => n748);
   U908 : INV_X1 port map( A => n749, ZN => n4161);
   U909 : MUX2_X1 port map( A => n3745, B => n306, S => n29, Z => n749);
   U910 : INV_X1 port map( A => n750, ZN => n4162);
   U911 : MUX2_X1 port map( A => n3746, B => n307, S => n29, Z => n750);
   U912 : INV_X1 port map( A => n751, ZN => n4163);
   U913 : MUX2_X1 port map( A => n3747, B => n308, S => n29, Z => n751);
   U914 : INV_X1 port map( A => n752, ZN => n4164);
   U915 : MUX2_X1 port map( A => n3748, B => n309, S => n29, Z => n752);
   U916 : INV_X1 port map( A => n753, ZN => n4165);
   U917 : MUX2_X1 port map( A => n3749, B => n310, S => n29, Z => n753);
   U918 : INV_X1 port map( A => n754, ZN => n4166);
   U919 : MUX2_X1 port map( A => n3750, B => n311, S => n29, Z => n754);
   U920 : INV_X1 port map( A => n755, ZN => n4167);
   U921 : MUX2_X1 port map( A => n3751, B => n312, S => n29, Z => n755);
   U922 : INV_X1 port map( A => n756, ZN => n4168);
   U923 : MUX2_X1 port map( A => n3752, B => n313, S => n29, Z => n756);
   U924 : INV_X1 port map( A => n757, ZN => n4169);
   U925 : MUX2_X1 port map( A => n3753, B => n314, S => n29, Z => n757);
   U926 : INV_X1 port map( A => n758, ZN => n4170);
   U927 : MUX2_X1 port map( A => n3754, B => n315, S => n29, Z => n758);
   U928 : INV_X1 port map( A => n759, ZN => n4171);
   U929 : MUX2_X1 port map( A => n3755, B => n316, S => n29, Z => n759);
   U930 : INV_X1 port map( A => n760, ZN => n4172);
   U931 : MUX2_X1 port map( A => n3756, B => n317, S => n29, Z => n760);
   U932 : INV_X1 port map( A => n761, ZN => n4173);
   U933 : MUX2_X1 port map( A => n3757, B => n318, S => n28, Z => n761);
   U934 : INV_X1 port map( A => n762, ZN => n4174);
   U935 : MUX2_X1 port map( A => n3758, B => n319, S => n28, Z => n762);
   U936 : INV_X1 port map( A => n763, ZN => n4175);
   U937 : MUX2_X1 port map( A => n3759, B => n320, S => n28, Z => n763);
   U938 : INV_X1 port map( A => n764, ZN => n4176);
   U939 : MUX2_X1 port map( A => n3760, B => n321, S => n28, Z => n764);
   U940 : INV_X1 port map( A => n765, ZN => n4177);
   U941 : MUX2_X1 port map( A => n3761, B => n322, S => n28, Z => n765);
   U942 : INV_X1 port map( A => n766, ZN => n4178);
   U943 : MUX2_X1 port map( A => n3762, B => n323, S => n28, Z => n766);
   U944 : INV_X1 port map( A => n767, ZN => n4179);
   U945 : MUX2_X1 port map( A => n3763, B => n324, S => n28, Z => n767);
   U946 : INV_X1 port map( A => n768, ZN => n4180);
   U947 : MUX2_X1 port map( A => n3764, B => n325, S => n28, Z => n768);
   U948 : INV_X1 port map( A => n769, ZN => n4181);
   U949 : MUX2_X1 port map( A => n3765, B => n326, S => n28, Z => n769);
   U950 : INV_X1 port map( A => n770, ZN => n4182);
   U951 : MUX2_X1 port map( A => n3766, B => n327, S => n28, Z => n770);
   U952 : INV_X1 port map( A => n771, ZN => n4183);
   U953 : MUX2_X1 port map( A => n3767, B => n328, S => n28, Z => n771);
   U954 : INV_X1 port map( A => n772, ZN => n4184);
   U955 : MUX2_X1 port map( A => n3768, B => n329, S => n28, Z => n772);
   U956 : AND2_X1 port map( A1 => n773, A2 => n704, ZN => n741);
   U957 : MUX2_X1 port map( A => n774, B => DATAIN(0), S => n33, Z => n4185);
   U958 : MUX2_X1 port map( A => n776, B => DATAIN(1), S => n33, Z => n4186);
   U959 : MUX2_X1 port map( A => n777, B => DATAIN(2), S => n33, Z => n4187);
   U960 : MUX2_X1 port map( A => n778, B => DATAIN(3), S => n33, Z => n4188);
   U961 : MUX2_X1 port map( A => n779, B => DATAIN(4), S => n33, Z => n4189);
   U962 : MUX2_X1 port map( A => n780, B => DATAIN(5), S => n33, Z => n4190);
   U963 : MUX2_X1 port map( A => n781, B => DATAIN(6), S => n33, Z => n4191);
   U964 : MUX2_X1 port map( A => n782, B => DATAIN(7), S => n33, Z => n4192);
   U965 : MUX2_X1 port map( A => n783, B => DATAIN(8), S => n32, Z => n4193);
   U966 : MUX2_X1 port map( A => n784, B => DATAIN(9), S => n32, Z => n4194);
   U967 : MUX2_X1 port map( A => n785, B => DATAIN(10), S => n32, Z => n4195);
   U968 : MUX2_X1 port map( A => n786, B => DATAIN(11), S => n32, Z => n4196);
   U969 : MUX2_X1 port map( A => n787, B => DATAIN(12), S => n32, Z => n4197);
   U970 : MUX2_X1 port map( A => n788, B => DATAIN(13), S => n32, Z => n4198);
   U971 : MUX2_X1 port map( A => n789, B => DATAIN(14), S => n32, Z => n4199);
   U972 : MUX2_X1 port map( A => n790, B => DATAIN(15), S => n32, Z => n4200);
   U973 : MUX2_X1 port map( A => n791, B => DATAIN(16), S => n32, Z => n4201);
   U974 : MUX2_X1 port map( A => n792, B => DATAIN(17), S => n32, Z => n4202);
   U975 : MUX2_X1 port map( A => n793, B => DATAIN(18), S => n32, Z => n4203);
   U976 : MUX2_X1 port map( A => n794, B => DATAIN(19), S => n32, Z => n4204);
   U977 : MUX2_X1 port map( A => n795, B => DATAIN(20), S => n31, Z => n4205);
   U978 : MUX2_X1 port map( A => n796, B => DATAIN(21), S => n31, Z => n4206);
   U979 : MUX2_X1 port map( A => n797, B => DATAIN(22), S => n31, Z => n4207);
   U980 : MUX2_X1 port map( A => n798, B => DATAIN(23), S => n31, Z => n4208);
   U981 : MUX2_X1 port map( A => n799, B => DATAIN(24), S => n31, Z => n4209);
   U982 : MUX2_X1 port map( A => n800, B => DATAIN(25), S => n31, Z => n4210);
   U983 : MUX2_X1 port map( A => n801, B => DATAIN(26), S => n31, Z => n4211);
   U984 : MUX2_X1 port map( A => n802, B => DATAIN(27), S => n31, Z => n4212);
   U985 : MUX2_X1 port map( A => n803, B => DATAIN(28), S => n31, Z => n4213);
   U986 : MUX2_X1 port map( A => n804, B => DATAIN(29), S => n31, Z => n4214);
   U987 : MUX2_X1 port map( A => n805, B => DATAIN(30), S => n31, Z => n4215);
   U988 : MUX2_X1 port map( A => n806, B => DATAIN(31), S => n31, Z => n4216);
   U989 : AND2_X1 port map( A1 => n807, A2 => n704, ZN => n775);
   U990 : MUX2_X1 port map( A => n808, B => DATAIN(0), S => n36, Z => n4217);
   U991 : MUX2_X1 port map( A => n810, B => DATAIN(1), S => n36, Z => n4218);
   U992 : MUX2_X1 port map( A => n811, B => DATAIN(2), S => n36, Z => n4219);
   U993 : MUX2_X1 port map( A => n812, B => DATAIN(3), S => n36, Z => n4220);
   U994 : MUX2_X1 port map( A => n813, B => DATAIN(4), S => n36, Z => n4221);
   U995 : MUX2_X1 port map( A => n814, B => DATAIN(5), S => n36, Z => n4222);
   U996 : MUX2_X1 port map( A => n815, B => DATAIN(6), S => n36, Z => n4223);
   U997 : MUX2_X1 port map( A => n816, B => DATAIN(7), S => n36, Z => n4224);
   U998 : MUX2_X1 port map( A => n817, B => DATAIN(8), S => n35, Z => n4225);
   U999 : MUX2_X1 port map( A => n818, B => DATAIN(9), S => n35, Z => n4226);
   U1000 : MUX2_X1 port map( A => n819, B => DATAIN(10), S => n35, Z => n4227);
   U1001 : MUX2_X1 port map( A => n820, B => DATAIN(11), S => n35, Z => n4228);
   U1002 : MUX2_X1 port map( A => n821, B => DATAIN(12), S => n35, Z => n4229);
   U1003 : MUX2_X1 port map( A => n822, B => DATAIN(13), S => n35, Z => n4230);
   U1004 : MUX2_X1 port map( A => n823, B => DATAIN(14), S => n35, Z => n4231);
   U1005 : MUX2_X1 port map( A => n824, B => DATAIN(15), S => n35, Z => n4232);
   U1006 : MUX2_X1 port map( A => n825, B => DATAIN(16), S => n35, Z => n4233);
   U1007 : MUX2_X1 port map( A => n826, B => DATAIN(17), S => n35, Z => n4234);
   U1008 : MUX2_X1 port map( A => n827, B => DATAIN(18), S => n35, Z => n4235);
   U1009 : MUX2_X1 port map( A => n828, B => DATAIN(19), S => n35, Z => n4236);
   U1010 : MUX2_X1 port map( A => n829, B => DATAIN(20), S => n34, Z => n4237);
   U1011 : MUX2_X1 port map( A => n830, B => DATAIN(21), S => n34, Z => n4238);
   U1012 : MUX2_X1 port map( A => n831, B => DATAIN(22), S => n34, Z => n4239);
   U1013 : MUX2_X1 port map( A => n832, B => DATAIN(23), S => n34, Z => n4240);
   U1014 : MUX2_X1 port map( A => n833, B => DATAIN(24), S => n34, Z => n4241);
   U1015 : MUX2_X1 port map( A => n834, B => DATAIN(25), S => n34, Z => n4242);
   U1016 : MUX2_X1 port map( A => n835, B => DATAIN(26), S => n34, Z => n4243);
   U1017 : MUX2_X1 port map( A => n836, B => DATAIN(27), S => n34, Z => n4244);
   U1018 : MUX2_X1 port map( A => n837, B => DATAIN(28), S => n34, Z => n4245);
   U1019 : MUX2_X1 port map( A => n838, B => DATAIN(29), S => n34, Z => n4246);
   U1020 : MUX2_X1 port map( A => n839, B => DATAIN(30), S => n34, Z => n4247);
   U1021 : MUX2_X1 port map( A => n840, B => DATAIN(31), S => n34, Z => n4248);
   U1022 : AND2_X1 port map( A1 => n841, A2 => n468, ZN => n809);
   U1023 : INV_X1 port map( A => n842, ZN => n4249);
   U1024 : MUX2_X1 port map( A => n3734, B => n298, S => n39, Z => n842);
   U1025 : INV_X1 port map( A => n844, ZN => n4250);
   U1026 : MUX2_X1 port map( A => n3713, B => n299, S => n39, Z => n844);
   U1027 : INV_X1 port map( A => n845, ZN => n4251);
   U1028 : MUX2_X1 port map( A => n3692, B => n300, S => n39, Z => n845);
   U1029 : INV_X1 port map( A => n846, ZN => n4252);
   U1030 : MUX2_X1 port map( A => n3671, B => n301, S => n39, Z => n846);
   U1031 : INV_X1 port map( A => n847, ZN => n4253);
   U1032 : MUX2_X1 port map( A => n3650, B => n302, S => n39, Z => n847);
   U1033 : INV_X1 port map( A => n848, ZN => n4254);
   U1034 : MUX2_X1 port map( A => n3629, B => n303, S => n39, Z => n848);
   U1035 : INV_X1 port map( A => n849, ZN => n4255);
   U1036 : MUX2_X1 port map( A => n3608, B => n304, S => n39, Z => n849);
   U1037 : INV_X1 port map( A => n850, ZN => n4256);
   U1038 : MUX2_X1 port map( A => n3587, B => n305, S => n39, Z => n850);
   U1039 : INV_X1 port map( A => n851, ZN => n4257);
   U1040 : MUX2_X1 port map( A => n3566, B => n306, S => n38, Z => n851);
   U1041 : INV_X1 port map( A => n852, ZN => n4258);
   U1042 : MUX2_X1 port map( A => n2969, B => n307, S => n38, Z => n852);
   U1043 : INV_X1 port map( A => n853, ZN => n4259);
   U1044 : MUX2_X1 port map( A => n2948, B => n308, S => n38, Z => n853);
   U1045 : INV_X1 port map( A => n854, ZN => n4260);
   U1046 : MUX2_X1 port map( A => n2927, B => n309, S => n38, Z => n854);
   U1047 : INV_X1 port map( A => n855, ZN => n4261);
   U1048 : MUX2_X1 port map( A => n2906, B => n310, S => n38, Z => n855);
   U1049 : INV_X1 port map( A => n856, ZN => n4262);
   U1050 : MUX2_X1 port map( A => n2885, B => n311, S => n38, Z => n856);
   U1051 : INV_X1 port map( A => n857, ZN => n4263);
   U1052 : MUX2_X1 port map( A => n2864, B => n312, S => n38, Z => n857);
   U1053 : INV_X1 port map( A => n858, ZN => n4264);
   U1054 : MUX2_X1 port map( A => n2843, B => n313, S => n38, Z => n858);
   U1055 : INV_X1 port map( A => n859, ZN => n4265);
   U1056 : MUX2_X1 port map( A => n2822, B => n314, S => n38, Z => n859);
   U1057 : INV_X1 port map( A => n860, ZN => n4266);
   U1058 : MUX2_X1 port map( A => n2801, B => n315, S => n38, Z => n860);
   U1059 : INV_X1 port map( A => n861, ZN => n4267);
   U1060 : MUX2_X1 port map( A => n2780, B => n316, S => n38, Z => n861);
   U1061 : INV_X1 port map( A => n862, ZN => n4268);
   U1062 : MUX2_X1 port map( A => n2759, B => n317, S => n38, Z => n862);
   U1063 : INV_X1 port map( A => n863, ZN => n4269);
   U1064 : MUX2_X1 port map( A => n2738, B => n318, S => n37, Z => n863);
   U1065 : INV_X1 port map( A => n864, ZN => n4270);
   U1066 : MUX2_X1 port map( A => n2717, B => n319, S => n37, Z => n864);
   U1067 : INV_X1 port map( A => n865, ZN => n4271);
   U1068 : MUX2_X1 port map( A => n2696, B => n320, S => n37, Z => n865);
   U1069 : INV_X1 port map( A => n866, ZN => n4272);
   U1070 : MUX2_X1 port map( A => n2675, B => n321, S => n37, Z => n866);
   U1071 : INV_X1 port map( A => n867, ZN => n4273);
   U1072 : MUX2_X1 port map( A => n2654, B => n322, S => n37, Z => n867);
   U1073 : INV_X1 port map( A => n868, ZN => n4274);
   U1074 : MUX2_X1 port map( A => n2633, B => n323, S => n37, Z => n868);
   U1075 : INV_X1 port map( A => n869, ZN => n4275);
   U1076 : MUX2_X1 port map( A => n2612, B => n324, S => n37, Z => n869);
   U1077 : INV_X1 port map( A => n870, ZN => n4276);
   U1078 : MUX2_X1 port map( A => n2591, B => n325, S => n37, Z => n870);
   U1079 : INV_X1 port map( A => n871, ZN => n4277);
   U1080 : MUX2_X1 port map( A => n2570, B => n326, S => n37, Z => n871);
   U1081 : INV_X1 port map( A => n872, ZN => n4278);
   U1082 : MUX2_X1 port map( A => n2549, B => n327, S => n37, Z => n872);
   U1083 : INV_X1 port map( A => n873, ZN => n4279);
   U1084 : MUX2_X1 port map( A => n2528, B => n328, S => n37, Z => n873);
   U1085 : INV_X1 port map( A => n874, ZN => n4280);
   U1086 : MUX2_X1 port map( A => n2507, B => n329, S => n37, Z => n874);
   U1087 : AND2_X1 port map( A1 => n841, A2 => n502, ZN => n843);
   U1088 : INV_X1 port map( A => n875, ZN => n4281);
   U1089 : MUX2_X1 port map( A => n3731, B => n298, S => n42, Z => n875);
   U1090 : INV_X1 port map( A => n877, ZN => n4282);
   U1091 : MUX2_X1 port map( A => n3710, B => n299, S => n42, Z => n877);
   U1092 : INV_X1 port map( A => n878, ZN => n4283);
   U1093 : MUX2_X1 port map( A => n3689, B => n300, S => n42, Z => n878);
   U1094 : INV_X1 port map( A => n879, ZN => n4284);
   U1095 : MUX2_X1 port map( A => n3668, B => n301, S => n42, Z => n879);
   U1096 : INV_X1 port map( A => n880, ZN => n4285);
   U1097 : MUX2_X1 port map( A => n3647, B => n302, S => n42, Z => n880);
   U1098 : INV_X1 port map( A => n881, ZN => n4286);
   U1099 : MUX2_X1 port map( A => n3626, B => n303, S => n42, Z => n881);
   U1100 : INV_X1 port map( A => n882, ZN => n4287);
   U1101 : MUX2_X1 port map( A => n3605, B => n304, S => n42, Z => n882);
   U1102 : INV_X1 port map( A => n883, ZN => n4288);
   U1103 : MUX2_X1 port map( A => n3584, B => n305, S => n42, Z => n883);
   U1104 : INV_X1 port map( A => n884, ZN => n4289);
   U1105 : MUX2_X1 port map( A => n3563, B => n306, S => n41, Z => n884);
   U1106 : INV_X1 port map( A => n885, ZN => n4290);
   U1107 : MUX2_X1 port map( A => n2966, B => n307, S => n41, Z => n885);
   U1108 : INV_X1 port map( A => n886, ZN => n4291);
   U1109 : MUX2_X1 port map( A => n2945, B => n308, S => n41, Z => n886);
   U1110 : INV_X1 port map( A => n887, ZN => n4292);
   U1111 : MUX2_X1 port map( A => n2924, B => n309, S => n41, Z => n887);
   U1112 : INV_X1 port map( A => n888, ZN => n4293);
   U1113 : MUX2_X1 port map( A => n2903, B => n310, S => n41, Z => n888);
   U1114 : INV_X1 port map( A => n889, ZN => n4294);
   U1115 : MUX2_X1 port map( A => n2882, B => n311, S => n41, Z => n889);
   U1116 : INV_X1 port map( A => n890, ZN => n4295);
   U1117 : MUX2_X1 port map( A => n2861, B => n312, S => n41, Z => n890);
   U1118 : INV_X1 port map( A => n891, ZN => n4296);
   U1119 : MUX2_X1 port map( A => n2840, B => n313, S => n41, Z => n891);
   U1120 : INV_X1 port map( A => n892, ZN => n4297);
   U1121 : MUX2_X1 port map( A => n2819, B => n314, S => n41, Z => n892);
   U1122 : INV_X1 port map( A => n893, ZN => n4298);
   U1123 : MUX2_X1 port map( A => n2798, B => n315, S => n41, Z => n893);
   U1124 : INV_X1 port map( A => n894, ZN => n4299);
   U1125 : MUX2_X1 port map( A => n2777, B => n316, S => n41, Z => n894);
   U1126 : INV_X1 port map( A => n895, ZN => n4300);
   U1127 : MUX2_X1 port map( A => n2756, B => n317, S => n41, Z => n895);
   U1128 : INV_X1 port map( A => n896, ZN => n4301);
   U1129 : MUX2_X1 port map( A => n2735, B => n318, S => n40, Z => n896);
   U1130 : INV_X1 port map( A => n897, ZN => n4302);
   U1131 : MUX2_X1 port map( A => n2714, B => n319, S => n40, Z => n897);
   U1132 : INV_X1 port map( A => n898, ZN => n4303);
   U1133 : MUX2_X1 port map( A => n2693, B => n320, S => n40, Z => n898);
   U1134 : INV_X1 port map( A => n899, ZN => n4304);
   U1135 : MUX2_X1 port map( A => n2672, B => n321, S => n40, Z => n899);
   U1136 : INV_X1 port map( A => n900, ZN => n4305);
   U1137 : MUX2_X1 port map( A => n2651, B => n322, S => n40, Z => n900);
   U1138 : INV_X1 port map( A => n901, ZN => n4306);
   U1139 : MUX2_X1 port map( A => n2630, B => n323, S => n40, Z => n901);
   U1140 : INV_X1 port map( A => n902, ZN => n4307);
   U1141 : MUX2_X1 port map( A => n2609, B => n324, S => n40, Z => n902);
   U1142 : INV_X1 port map( A => n903, ZN => n4308);
   U1143 : MUX2_X1 port map( A => n2588, B => n325, S => n40, Z => n903);
   U1144 : INV_X1 port map( A => n904, ZN => n4309);
   U1145 : MUX2_X1 port map( A => n2567, B => n326, S => n40, Z => n904);
   U1146 : INV_X1 port map( A => n905, ZN => n4310);
   U1147 : MUX2_X1 port map( A => n2546, B => n327, S => n40, Z => n905);
   U1148 : INV_X1 port map( A => n906, ZN => n4311);
   U1149 : MUX2_X1 port map( A => n2525, B => n328, S => n40, Z => n906);
   U1150 : INV_X1 port map( A => n907, ZN => n4312);
   U1151 : MUX2_X1 port map( A => n2504, B => n329, S => n40, Z => n907);
   U1152 : AND2_X1 port map( A1 => n841, A2 => n536, ZN => n876);
   U1153 : MUX2_X1 port map( A => n908, B => DATAIN(0), S => n45, Z => n4313);
   U1154 : MUX2_X1 port map( A => n910, B => DATAIN(1), S => n45, Z => n4314);
   U1155 : MUX2_X1 port map( A => n911, B => DATAIN(2), S => n45, Z => n4315);
   U1156 : MUX2_X1 port map( A => n912, B => DATAIN(3), S => n45, Z => n4316);
   U1157 : MUX2_X1 port map( A => n913, B => DATAIN(4), S => n45, Z => n4317);
   U1158 : MUX2_X1 port map( A => n914, B => DATAIN(5), S => n45, Z => n4318);
   U1159 : MUX2_X1 port map( A => n915, B => DATAIN(6), S => n45, Z => n4319);
   U1160 : MUX2_X1 port map( A => n916, B => DATAIN(7), S => n45, Z => n4320);
   U1161 : MUX2_X1 port map( A => n917, B => DATAIN(8), S => n44, Z => n4321);
   U1162 : MUX2_X1 port map( A => n918, B => DATAIN(9), S => n44, Z => n4322);
   U1163 : MUX2_X1 port map( A => n919, B => DATAIN(10), S => n44, Z => n4323);
   U1164 : MUX2_X1 port map( A => n920, B => DATAIN(11), S => n44, Z => n4324);
   U1165 : MUX2_X1 port map( A => n921, B => DATAIN(12), S => n44, Z => n4325);
   U1166 : MUX2_X1 port map( A => n922, B => DATAIN(13), S => n44, Z => n4326);
   U1167 : MUX2_X1 port map( A => n923, B => DATAIN(14), S => n44, Z => n4327);
   U1168 : MUX2_X1 port map( A => n924, B => DATAIN(15), S => n44, Z => n4328);
   U1169 : MUX2_X1 port map( A => n925, B => DATAIN(16), S => n44, Z => n4329);
   U1170 : MUX2_X1 port map( A => n926, B => DATAIN(17), S => n44, Z => n4330);
   U1171 : MUX2_X1 port map( A => n927, B => DATAIN(18), S => n44, Z => n4331);
   U1172 : MUX2_X1 port map( A => n928, B => DATAIN(19), S => n44, Z => n4332);
   U1173 : MUX2_X1 port map( A => n929, B => DATAIN(20), S => n43, Z => n4333);
   U1174 : MUX2_X1 port map( A => n930, B => DATAIN(21), S => n43, Z => n4334);
   U1175 : MUX2_X1 port map( A => n931, B => DATAIN(22), S => n43, Z => n4335);
   U1176 : MUX2_X1 port map( A => n932, B => DATAIN(23), S => n43, Z => n4336);
   U1177 : MUX2_X1 port map( A => n933, B => DATAIN(24), S => n43, Z => n4337);
   U1178 : MUX2_X1 port map( A => n934, B => DATAIN(25), S => n43, Z => n4338);
   U1179 : MUX2_X1 port map( A => n935, B => DATAIN(26), S => n43, Z => n4339);
   U1180 : MUX2_X1 port map( A => n936, B => DATAIN(27), S => n43, Z => n4340);
   U1181 : MUX2_X1 port map( A => n937, B => DATAIN(28), S => n43, Z => n4341);
   U1182 : MUX2_X1 port map( A => n938, B => DATAIN(29), S => n43, Z => n4342);
   U1183 : MUX2_X1 port map( A => n939, B => DATAIN(30), S => n43, Z => n4343);
   U1184 : MUX2_X1 port map( A => n940, B => DATAIN(31), S => n43, Z => n4344);
   U1185 : AND2_X1 port map( A1 => n841, A2 => n570, ZN => n909);
   U1186 : MUX2_X1 port map( A => n2501, B => DATAIN(31), S => n48, Z => n3558)
                           ;
   U1187 : MUX2_X1 port map( A => n2522, B => DATAIN(30), S => n48, Z => n3557)
                           ;
   U1188 : MUX2_X1 port map( A => n2543, B => DATAIN(29), S => n48, Z => n3556)
                           ;
   U1189 : MUX2_X1 port map( A => n2564, B => DATAIN(28), S => n48, Z => n3555)
                           ;
   U1190 : MUX2_X1 port map( A => n2585, B => DATAIN(27), S => n48, Z => n3554)
                           ;
   U1191 : MUX2_X1 port map( A => n2606, B => DATAIN(26), S => n48, Z => n3553)
                           ;
   U1192 : MUX2_X1 port map( A => n2627, B => DATAIN(25), S => n48, Z => n3552)
                           ;
   U1193 : MUX2_X1 port map( A => n2648, B => DATAIN(24), S => n48, Z => n3551)
                           ;
   U1194 : MUX2_X1 port map( A => n2669, B => DATAIN(23), S => n47, Z => n3550)
                           ;
   U1195 : MUX2_X1 port map( A => n2690, B => DATAIN(22), S => n47, Z => n3549)
                           ;
   U1196 : MUX2_X1 port map( A => n2711, B => DATAIN(21), S => n47, Z => n3548)
                           ;
   U1197 : MUX2_X1 port map( A => n2732, B => DATAIN(20), S => n47, Z => n3547)
                           ;
   U1198 : MUX2_X1 port map( A => n2753, B => DATAIN(19), S => n47, Z => n3546)
                           ;
   U1199 : MUX2_X1 port map( A => n2774, B => DATAIN(18), S => n47, Z => n3545)
                           ;
   U1200 : MUX2_X1 port map( A => n2795, B => DATAIN(17), S => n47, Z => n3544)
                           ;
   U1201 : MUX2_X1 port map( A => n2816, B => DATAIN(16), S => n47, Z => n3543)
                           ;
   U1202 : MUX2_X1 port map( A => n2837, B => DATAIN(15), S => n47, Z => n3542)
                           ;
   U1203 : MUX2_X1 port map( A => n2858, B => DATAIN(14), S => n47, Z => n3541)
                           ;
   U1204 : MUX2_X1 port map( A => n2879, B => DATAIN(13), S => n47, Z => n3540)
                           ;
   U1205 : MUX2_X1 port map( A => n2900, B => DATAIN(12), S => n47, Z => n3539)
                           ;
   U1206 : MUX2_X1 port map( A => n2921, B => DATAIN(11), S => n46, Z => n3538)
                           ;
   U1207 : MUX2_X1 port map( A => n2942, B => DATAIN(10), S => n46, Z => n3537)
                           ;
   U1208 : MUX2_X1 port map( A => n2963, B => DATAIN(9), S => n46, Z => n3536);
   U1209 : MUX2_X1 port map( A => n3560, B => DATAIN(8), S => n46, Z => n3535);
   U1210 : MUX2_X1 port map( A => n3581, B => DATAIN(7), S => n46, Z => n3534);
   U1211 : MUX2_X1 port map( A => n3602, B => DATAIN(6), S => n46, Z => n3533);
   U1212 : MUX2_X1 port map( A => n3623, B => DATAIN(5), S => n46, Z => n3532);
   U1213 : MUX2_X1 port map( A => n3644, B => DATAIN(4), S => n46, Z => n3531);
   U1214 : MUX2_X1 port map( A => n3665, B => DATAIN(3), S => n46, Z => n3530);
   U1215 : MUX2_X1 port map( A => n3686, B => DATAIN(2), S => n46, Z => n3529);
   U1216 : MUX2_X1 port map( A => n3707, B => DATAIN(1), S => n46, Z => n3528);
   U1217 : MUX2_X1 port map( A => n3728, B => DATAIN(0), S => n46, Z => n3527);
   U1218 : AND2_X1 port map( A1 => n705, A2 => n604, ZN => n941);
   U1219 : MUX2_X1 port map( A => n2500, B => DATAIN(31), S => n51, Z => n3526)
                           ;
   U1220 : MUX2_X1 port map( A => n2521, B => DATAIN(30), S => n51, Z => n3525)
                           ;
   U1221 : MUX2_X1 port map( A => n2542, B => DATAIN(29), S => n51, Z => n3524)
                           ;
   U1222 : MUX2_X1 port map( A => n2563, B => DATAIN(28), S => n51, Z => n3523)
                           ;
   U1223 : MUX2_X1 port map( A => n2584, B => DATAIN(27), S => n51, Z => n3522)
                           ;
   U1224 : MUX2_X1 port map( A => n2605, B => DATAIN(26), S => n51, Z => n3521)
                           ;
   U1225 : MUX2_X1 port map( A => n2626, B => DATAIN(25), S => n51, Z => n3520)
                           ;
   U1226 : MUX2_X1 port map( A => n2647, B => DATAIN(24), S => n51, Z => n3519)
                           ;
   U1227 : MUX2_X1 port map( A => n2668, B => DATAIN(23), S => n50, Z => n3518)
                           ;
   U1228 : MUX2_X1 port map( A => n2689, B => DATAIN(22), S => n50, Z => n3517)
                           ;
   U1229 : MUX2_X1 port map( A => n2710, B => DATAIN(21), S => n50, Z => n3516)
                           ;
   U1230 : MUX2_X1 port map( A => n2731, B => DATAIN(20), S => n50, Z => n3515)
                           ;
   U1231 : MUX2_X1 port map( A => n2752, B => DATAIN(19), S => n50, Z => n3514)
                           ;
   U1232 : MUX2_X1 port map( A => n2773, B => DATAIN(18), S => n50, Z => n3513)
                           ;
   U1233 : MUX2_X1 port map( A => n2794, B => DATAIN(17), S => n50, Z => n3512)
                           ;
   U1234 : MUX2_X1 port map( A => n2815, B => DATAIN(16), S => n50, Z => n3511)
                           ;
   U1235 : MUX2_X1 port map( A => n2836, B => DATAIN(15), S => n50, Z => n3510)
                           ;
   U1236 : MUX2_X1 port map( A => n2857, B => DATAIN(14), S => n50, Z => n3509)
                           ;
   U1237 : MUX2_X1 port map( A => n2878, B => DATAIN(13), S => n50, Z => n3508)
                           ;
   U1238 : MUX2_X1 port map( A => n2899, B => DATAIN(12), S => n50, Z => n3507)
                           ;
   U1239 : MUX2_X1 port map( A => n2920, B => DATAIN(11), S => n49, Z => n3506)
                           ;
   U1240 : MUX2_X1 port map( A => n2941, B => DATAIN(10), S => n49, Z => n3505)
                           ;
   U1241 : MUX2_X1 port map( A => n2962, B => DATAIN(9), S => n49, Z => n3504);
   U1242 : MUX2_X1 port map( A => n3559, B => DATAIN(8), S => n49, Z => n3503);
   U1243 : MUX2_X1 port map( A => n3580, B => DATAIN(7), S => n49, Z => n3502);
   U1244 : MUX2_X1 port map( A => n3601, B => DATAIN(6), S => n49, Z => n3501);
   U1245 : MUX2_X1 port map( A => n3622, B => DATAIN(5), S => n49, Z => n3500);
   U1246 : MUX2_X1 port map( A => n3643, B => DATAIN(4), S => n49, Z => n3499);
   U1247 : MUX2_X1 port map( A => n3664, B => DATAIN(3), S => n49, Z => n3498);
   U1248 : MUX2_X1 port map( A => n3685, B => DATAIN(2), S => n49, Z => n3497);
   U1249 : MUX2_X1 port map( A => n3706, B => DATAIN(1), S => n49, Z => n3496);
   U1250 : MUX2_X1 port map( A => n3727, B => DATAIN(0), S => n49, Z => n3495);
   U1251 : AND2_X1 port map( A1 => n739, A2 => n604, ZN => n942);
   U1252 : MUX2_X1 port map( A => n2499, B => DATAIN(31), S => n54, Z => n3494)
                           ;
   U1253 : MUX2_X1 port map( A => n2520, B => DATAIN(30), S => n54, Z => n3493)
                           ;
   U1254 : MUX2_X1 port map( A => n2541, B => DATAIN(29), S => n54, Z => n3492)
                           ;
   U1255 : MUX2_X1 port map( A => n2562, B => DATAIN(28), S => n54, Z => n3491)
                           ;
   U1256 : MUX2_X1 port map( A => n2583, B => DATAIN(27), S => n54, Z => n3490)
                           ;
   U1257 : MUX2_X1 port map( A => n2604, B => DATAIN(26), S => n54, Z => n3489)
                           ;
   U1258 : MUX2_X1 port map( A => n2625, B => DATAIN(25), S => n54, Z => n3488)
                           ;
   U1259 : MUX2_X1 port map( A => n2646, B => DATAIN(24), S => n54, Z => n3487)
                           ;
   U1260 : MUX2_X1 port map( A => n2667, B => DATAIN(23), S => n53, Z => n3486)
                           ;
   U1261 : MUX2_X1 port map( A => n2688, B => DATAIN(22), S => n53, Z => n3485)
                           ;
   U1262 : MUX2_X1 port map( A => n2709, B => DATAIN(21), S => n53, Z => n3484)
                           ;
   U1263 : MUX2_X1 port map( A => n2730, B => DATAIN(20), S => n53, Z => n3483)
                           ;
   U1264 : MUX2_X1 port map( A => n2751, B => DATAIN(19), S => n53, Z => n3482)
                           ;
   U1265 : MUX2_X1 port map( A => n2772, B => DATAIN(18), S => n53, Z => n3481)
                           ;
   U1266 : MUX2_X1 port map( A => n2793, B => DATAIN(17), S => n53, Z => n3480)
                           ;
   U1267 : MUX2_X1 port map( A => n2814, B => DATAIN(16), S => n53, Z => n3479)
                           ;
   U1268 : MUX2_X1 port map( A => n2835, B => DATAIN(15), S => n53, Z => n3478)
                           ;
   U1269 : MUX2_X1 port map( A => n2856, B => DATAIN(14), S => n53, Z => n3477)
                           ;
   U1270 : MUX2_X1 port map( A => n2877, B => DATAIN(13), S => n53, Z => n3476)
                           ;
   U1271 : MUX2_X1 port map( A => n2898, B => DATAIN(12), S => n53, Z => n3475)
                           ;
   U1272 : MUX2_X1 port map( A => n2919, B => DATAIN(11), S => n52, Z => n3474)
                           ;
   U1273 : MUX2_X1 port map( A => n2940, B => DATAIN(10), S => n52, Z => n3473)
                           ;
   U1274 : MUX2_X1 port map( A => n2961, B => DATAIN(9), S => n52, Z => n3472);
   U1275 : MUX2_X1 port map( A => n2982, B => DATAIN(8), S => n52, Z => n3471);
   U1276 : MUX2_X1 port map( A => n3579, B => DATAIN(7), S => n52, Z => n3470);
   U1277 : MUX2_X1 port map( A => n3600, B => DATAIN(6), S => n52, Z => n3469);
   U1278 : MUX2_X1 port map( A => n3621, B => DATAIN(5), S => n52, Z => n3468);
   U1279 : MUX2_X1 port map( A => n3642, B => DATAIN(4), S => n52, Z => n3467);
   U1280 : MUX2_X1 port map( A => n3663, B => DATAIN(3), S => n52, Z => n3466);
   U1281 : MUX2_X1 port map( A => n3684, B => DATAIN(2), S => n52, Z => n3465);
   U1282 : MUX2_X1 port map( A => n3705, B => DATAIN(1), S => n52, Z => n3464);
   U1283 : MUX2_X1 port map( A => n3726, B => DATAIN(0), S => n52, Z => n3463);
   U1284 : AND2_X1 port map( A1 => n773, A2 => n604, ZN => n943);
   U1285 : MUX2_X1 port map( A => n2498, B => DATAIN(31), S => n57, Z => n3462)
                           ;
   U1286 : MUX2_X1 port map( A => n2519, B => DATAIN(30), S => n57, Z => n3461)
                           ;
   U1287 : MUX2_X1 port map( A => n2540, B => DATAIN(29), S => n57, Z => n3460)
                           ;
   U1288 : MUX2_X1 port map( A => n2561, B => DATAIN(28), S => n57, Z => n3459)
                           ;
   U1289 : MUX2_X1 port map( A => n2582, B => DATAIN(27), S => n57, Z => n3458)
                           ;
   U1290 : MUX2_X1 port map( A => n2603, B => DATAIN(26), S => n57, Z => n3457)
                           ;
   U1291 : MUX2_X1 port map( A => n2624, B => DATAIN(25), S => n57, Z => n3456)
                           ;
   U1292 : MUX2_X1 port map( A => n2645, B => DATAIN(24), S => n57, Z => n3455)
                           ;
   U1293 : MUX2_X1 port map( A => n2666, B => DATAIN(23), S => n56, Z => n3454)
                           ;
   U1294 : MUX2_X1 port map( A => n2687, B => DATAIN(22), S => n56, Z => n3453)
                           ;
   U1295 : MUX2_X1 port map( A => n2708, B => DATAIN(21), S => n56, Z => n3452)
                           ;
   U1296 : MUX2_X1 port map( A => n2729, B => DATAIN(20), S => n56, Z => n3451)
                           ;
   U1297 : MUX2_X1 port map( A => n2750, B => DATAIN(19), S => n56, Z => n3450)
                           ;
   U1298 : MUX2_X1 port map( A => n2771, B => DATAIN(18), S => n56, Z => n3449)
                           ;
   U1299 : MUX2_X1 port map( A => n2792, B => DATAIN(17), S => n56, Z => n3448)
                           ;
   U1300 : MUX2_X1 port map( A => n2813, B => DATAIN(16), S => n56, Z => n3447)
                           ;
   U1301 : MUX2_X1 port map( A => n2834, B => DATAIN(15), S => n56, Z => n3446)
                           ;
   U1302 : MUX2_X1 port map( A => n2855, B => DATAIN(14), S => n56, Z => n3445)
                           ;
   U1303 : MUX2_X1 port map( A => n2876, B => DATAIN(13), S => n56, Z => n3444)
                           ;
   U1304 : MUX2_X1 port map( A => n2897, B => DATAIN(12), S => n56, Z => n3443)
                           ;
   U1305 : MUX2_X1 port map( A => n2918, B => DATAIN(11), S => n55, Z => n3442)
                           ;
   U1306 : MUX2_X1 port map( A => n2939, B => DATAIN(10), S => n55, Z => n3441)
                           ;
   U1307 : MUX2_X1 port map( A => n2960, B => DATAIN(9), S => n55, Z => n3440);
   U1308 : MUX2_X1 port map( A => n2981, B => DATAIN(8), S => n55, Z => n3439);
   U1309 : MUX2_X1 port map( A => n3578, B => DATAIN(7), S => n55, Z => n3438);
   U1310 : MUX2_X1 port map( A => n3599, B => DATAIN(6), S => n55, Z => n3437);
   U1311 : MUX2_X1 port map( A => n3620, B => DATAIN(5), S => n55, Z => n3436);
   U1312 : MUX2_X1 port map( A => n3641, B => DATAIN(4), S => n55, Z => n3435);
   U1313 : MUX2_X1 port map( A => n3662, B => DATAIN(3), S => n55, Z => n3434);
   U1314 : MUX2_X1 port map( A => n3683, B => DATAIN(2), S => n55, Z => n3433);
   U1315 : MUX2_X1 port map( A => n3704, B => DATAIN(1), S => n55, Z => n3432);
   U1316 : MUX2_X1 port map( A => n3725, B => DATAIN(0), S => n55, Z => n3431);
   U1317 : AND2_X1 port map( A1 => n807, A2 => n604, ZN => n944);
   U1318 : AND3_X1 port map( A1 => n945, A2 => n946, A3 => n947, ZN => n604);
   U1319 : MUX2_X1 port map( A => n2497, B => DATAIN(31), S => n60, Z => n3430)
                           ;
   U1320 : MUX2_X1 port map( A => n2518, B => DATAIN(30), S => n60, Z => n3429)
                           ;
   U1321 : MUX2_X1 port map( A => n2539, B => DATAIN(29), S => n60, Z => n3428)
                           ;
   U1322 : MUX2_X1 port map( A => n2560, B => DATAIN(28), S => n60, Z => n3427)
                           ;
   U1323 : MUX2_X1 port map( A => n2581, B => DATAIN(27), S => n60, Z => n3426)
                           ;
   U1324 : MUX2_X1 port map( A => n2602, B => DATAIN(26), S => n60, Z => n3425)
                           ;
   U1325 : MUX2_X1 port map( A => n2623, B => DATAIN(25), S => n60, Z => n3424)
                           ;
   U1326 : MUX2_X1 port map( A => n2644, B => DATAIN(24), S => n60, Z => n3423)
                           ;
   U1327 : MUX2_X1 port map( A => n2665, B => DATAIN(23), S => n59, Z => n3422)
                           ;
   U1328 : MUX2_X1 port map( A => n2686, B => DATAIN(22), S => n59, Z => n3421)
                           ;
   U1329 : MUX2_X1 port map( A => n2707, B => DATAIN(21), S => n59, Z => n3420)
                           ;
   U1330 : MUX2_X1 port map( A => n2728, B => DATAIN(20), S => n59, Z => n3419)
                           ;
   U1331 : MUX2_X1 port map( A => n2749, B => DATAIN(19), S => n59, Z => n3418)
                           ;
   U1332 : MUX2_X1 port map( A => n2770, B => DATAIN(18), S => n59, Z => n3417)
                           ;
   U1333 : MUX2_X1 port map( A => n2791, B => DATAIN(17), S => n59, Z => n3416)
                           ;
   U1334 : MUX2_X1 port map( A => n2812, B => DATAIN(16), S => n59, Z => n3415)
                           ;
   U1335 : MUX2_X1 port map( A => n2833, B => DATAIN(15), S => n59, Z => n3414)
                           ;
   U1336 : MUX2_X1 port map( A => n2854, B => DATAIN(14), S => n59, Z => n3413)
                           ;
   U1337 : MUX2_X1 port map( A => n2875, B => DATAIN(13), S => n59, Z => n3412)
                           ;
   U1338 : MUX2_X1 port map( A => n2896, B => DATAIN(12), S => n59, Z => n3411)
                           ;
   U1339 : MUX2_X1 port map( A => n2917, B => DATAIN(11), S => n58, Z => n3410)
                           ;
   U1340 : MUX2_X1 port map( A => n2938, B => DATAIN(10), S => n58, Z => n3409)
                           ;
   U1341 : MUX2_X1 port map( A => n2959, B => DATAIN(9), S => n58, Z => n3408);
   U1342 : MUX2_X1 port map( A => n2980, B => DATAIN(8), S => n58, Z => n3407);
   U1343 : MUX2_X1 port map( A => n3577, B => DATAIN(7), S => n58, Z => n3406);
   U1344 : MUX2_X1 port map( A => n3598, B => DATAIN(6), S => n58, Z => n3405);
   U1345 : MUX2_X1 port map( A => n3619, B => DATAIN(5), S => n58, Z => n3404);
   U1346 : MUX2_X1 port map( A => n3640, B => DATAIN(4), S => n58, Z => n3403);
   U1347 : MUX2_X1 port map( A => n3661, B => DATAIN(3), S => n58, Z => n3402);
   U1348 : MUX2_X1 port map( A => n3682, B => DATAIN(2), S => n58, Z => n3401);
   U1349 : MUX2_X1 port map( A => n3703, B => DATAIN(1), S => n58, Z => n3400);
   U1350 : MUX2_X1 port map( A => n3724, B => DATAIN(0), S => n58, Z => n3399);
   U1351 : AND2_X1 port map( A1 => n705, A2 => n467, ZN => n948);
   U1352 : MUX2_X1 port map( A => n2496, B => DATAIN(31), S => n63, Z => n3398)
                           ;
   U1353 : MUX2_X1 port map( A => n2517, B => DATAIN(30), S => n63, Z => n3397)
                           ;
   U1354 : MUX2_X1 port map( A => n2538, B => DATAIN(29), S => n63, Z => n3396)
                           ;
   U1355 : MUX2_X1 port map( A => n2559, B => DATAIN(28), S => n63, Z => n3395)
                           ;
   U1356 : MUX2_X1 port map( A => n2580, B => DATAIN(27), S => n63, Z => n3394)
                           ;
   U1357 : MUX2_X1 port map( A => n2601, B => DATAIN(26), S => n63, Z => n3393)
                           ;
   U1358 : MUX2_X1 port map( A => n2622, B => DATAIN(25), S => n63, Z => n3392)
                           ;
   U1359 : MUX2_X1 port map( A => n2643, B => DATAIN(24), S => n63, Z => n3391)
                           ;
   U1360 : MUX2_X1 port map( A => n2664, B => DATAIN(23), S => n62, Z => n3390)
                           ;
   U1361 : MUX2_X1 port map( A => n2685, B => DATAIN(22), S => n62, Z => n3389)
                           ;
   U1362 : MUX2_X1 port map( A => n2706, B => DATAIN(21), S => n62, Z => n3388)
                           ;
   U1363 : MUX2_X1 port map( A => n2727, B => DATAIN(20), S => n62, Z => n3387)
                           ;
   U1364 : MUX2_X1 port map( A => n2748, B => DATAIN(19), S => n62, Z => n3386)
                           ;
   U1365 : MUX2_X1 port map( A => n2769, B => DATAIN(18), S => n62, Z => n3385)
                           ;
   U1366 : MUX2_X1 port map( A => n2790, B => DATAIN(17), S => n62, Z => n3384)
                           ;
   U1367 : MUX2_X1 port map( A => n2811, B => DATAIN(16), S => n62, Z => n3383)
                           ;
   U1368 : MUX2_X1 port map( A => n2832, B => DATAIN(15), S => n62, Z => n3382)
                           ;
   U1369 : MUX2_X1 port map( A => n2853, B => DATAIN(14), S => n62, Z => n3381)
                           ;
   U1370 : MUX2_X1 port map( A => n2874, B => DATAIN(13), S => n62, Z => n3380)
                           ;
   U1371 : MUX2_X1 port map( A => n2895, B => DATAIN(12), S => n62, Z => n3379)
                           ;
   U1372 : MUX2_X1 port map( A => n2916, B => DATAIN(11), S => n61, Z => n3378)
                           ;
   U1373 : MUX2_X1 port map( A => n2937, B => DATAIN(10), S => n61, Z => n3377)
                           ;
   U1374 : MUX2_X1 port map( A => n2958, B => DATAIN(9), S => n61, Z => n3376);
   U1375 : MUX2_X1 port map( A => n2979, B => DATAIN(8), S => n61, Z => n3375);
   U1376 : MUX2_X1 port map( A => n3576, B => DATAIN(7), S => n61, Z => n3374);
   U1377 : MUX2_X1 port map( A => n3597, B => DATAIN(6), S => n61, Z => n3373);
   U1378 : MUX2_X1 port map( A => n3618, B => DATAIN(5), S => n61, Z => n3372);
   U1379 : MUX2_X1 port map( A => n3639, B => DATAIN(4), S => n61, Z => n3371);
   U1380 : MUX2_X1 port map( A => n3660, B => DATAIN(3), S => n61, Z => n3370);
   U1381 : MUX2_X1 port map( A => n3681, B => DATAIN(2), S => n61, Z => n3369);
   U1382 : MUX2_X1 port map( A => n3702, B => DATAIN(1), S => n61, Z => n3368);
   U1383 : MUX2_X1 port map( A => n3723, B => DATAIN(0), S => n61, Z => n3367);
   U1384 : AND2_X1 port map( A1 => n739, A2 => n467, ZN => n949);
   U1385 : MUX2_X1 port map( A => n2493, B => DATAIN(31), S => n66, Z => n3366)
                           ;
   U1386 : MUX2_X1 port map( A => n2514, B => DATAIN(30), S => n66, Z => n3365)
                           ;
   U1387 : MUX2_X1 port map( A => n2535, B => DATAIN(29), S => n66, Z => n3364)
                           ;
   U1388 : MUX2_X1 port map( A => n2556, B => DATAIN(28), S => n66, Z => n3363)
                           ;
   U1389 : MUX2_X1 port map( A => n2577, B => DATAIN(27), S => n66, Z => n3362)
                           ;
   U1390 : MUX2_X1 port map( A => n2598, B => DATAIN(26), S => n66, Z => n3361)
                           ;
   U1391 : MUX2_X1 port map( A => n2619, B => DATAIN(25), S => n66, Z => n3360)
                           ;
   U1392 : MUX2_X1 port map( A => n2640, B => DATAIN(24), S => n66, Z => n3359)
                           ;
   U1393 : MUX2_X1 port map( A => n2661, B => DATAIN(23), S => n65, Z => n3358)
                           ;
   U1394 : MUX2_X1 port map( A => n2682, B => DATAIN(22), S => n65, Z => n3357)
                           ;
   U1395 : MUX2_X1 port map( A => n2703, B => DATAIN(21), S => n65, Z => n3356)
                           ;
   U1396 : MUX2_X1 port map( A => n2724, B => DATAIN(20), S => n65, Z => n3355)
                           ;
   U1397 : MUX2_X1 port map( A => n2745, B => DATAIN(19), S => n65, Z => n3354)
                           ;
   U1398 : MUX2_X1 port map( A => n2766, B => DATAIN(18), S => n65, Z => n3353)
                           ;
   U1399 : MUX2_X1 port map( A => n2787, B => DATAIN(17), S => n65, Z => n3352)
                           ;
   U1400 : MUX2_X1 port map( A => n2808, B => DATAIN(16), S => n65, Z => n3351)
                           ;
   U1401 : MUX2_X1 port map( A => n2829, B => DATAIN(15), S => n65, Z => n3350)
                           ;
   U1402 : MUX2_X1 port map( A => n2850, B => DATAIN(14), S => n65, Z => n3349)
                           ;
   U1403 : MUX2_X1 port map( A => n2871, B => DATAIN(13), S => n65, Z => n3348)
                           ;
   U1404 : MUX2_X1 port map( A => n2892, B => DATAIN(12), S => n65, Z => n3347)
                           ;
   U1405 : MUX2_X1 port map( A => n2913, B => DATAIN(11), S => n64, Z => n3346)
                           ;
   U1406 : MUX2_X1 port map( A => n2934, B => DATAIN(10), S => n64, Z => n3345)
                           ;
   U1407 : MUX2_X1 port map( A => n2955, B => DATAIN(9), S => n64, Z => n3344);
   U1408 : MUX2_X1 port map( A => n2976, B => DATAIN(8), S => n64, Z => n3343);
   U1409 : MUX2_X1 port map( A => n3573, B => DATAIN(7), S => n64, Z => n3342);
   U1410 : MUX2_X1 port map( A => n3594, B => DATAIN(6), S => n64, Z => n3341);
   U1411 : MUX2_X1 port map( A => n3615, B => DATAIN(5), S => n64, Z => n3340);
   U1412 : MUX2_X1 port map( A => n3636, B => DATAIN(4), S => n64, Z => n3339);
   U1413 : MUX2_X1 port map( A => n3657, B => DATAIN(3), S => n64, Z => n3338);
   U1414 : MUX2_X1 port map( A => n3678, B => DATAIN(2), S => n64, Z => n3337);
   U1415 : MUX2_X1 port map( A => n3699, B => DATAIN(1), S => n64, Z => n3336);
   U1416 : MUX2_X1 port map( A => n3720, B => DATAIN(0), S => n64, Z => n3335);
   U1417 : AND2_X1 port map( A1 => n773, A2 => n467, ZN => n950);
   U1418 : MUX2_X1 port map( A => n2492, B => DATAIN(31), S => n69, Z => n3334)
                           ;
   U1419 : MUX2_X1 port map( A => n2513, B => DATAIN(30), S => n69, Z => n3333)
                           ;
   U1420 : MUX2_X1 port map( A => n2534, B => DATAIN(29), S => n69, Z => n3332)
                           ;
   U1421 : MUX2_X1 port map( A => n2555, B => DATAIN(28), S => n69, Z => n3331)
                           ;
   U1422 : MUX2_X1 port map( A => n2576, B => DATAIN(27), S => n69, Z => n3330)
                           ;
   U1423 : MUX2_X1 port map( A => n2597, B => DATAIN(26), S => n69, Z => n3329)
                           ;
   U1424 : MUX2_X1 port map( A => n2618, B => DATAIN(25), S => n69, Z => n3328)
                           ;
   U1425 : MUX2_X1 port map( A => n2639, B => DATAIN(24), S => n69, Z => n3327)
                           ;
   U1426 : MUX2_X1 port map( A => n2660, B => DATAIN(23), S => n68, Z => n3326)
                           ;
   U1427 : MUX2_X1 port map( A => n2681, B => DATAIN(22), S => n68, Z => n3325)
                           ;
   U1428 : MUX2_X1 port map( A => n2702, B => DATAIN(21), S => n68, Z => n3324)
                           ;
   U1429 : MUX2_X1 port map( A => n2723, B => DATAIN(20), S => n68, Z => n3323)
                           ;
   U1430 : MUX2_X1 port map( A => n2744, B => DATAIN(19), S => n68, Z => n3322)
                           ;
   U1431 : MUX2_X1 port map( A => n2765, B => DATAIN(18), S => n68, Z => n3321)
                           ;
   U1432 : MUX2_X1 port map( A => n2786, B => DATAIN(17), S => n68, Z => n3320)
                           ;
   U1433 : MUX2_X1 port map( A => n2807, B => DATAIN(16), S => n68, Z => n3319)
                           ;
   U1434 : MUX2_X1 port map( A => n2828, B => DATAIN(15), S => n68, Z => n3318)
                           ;
   U1435 : MUX2_X1 port map( A => n2849, B => DATAIN(14), S => n68, Z => n3317)
                           ;
   U1436 : MUX2_X1 port map( A => n2870, B => DATAIN(13), S => n68, Z => n3316)
                           ;
   U1437 : MUX2_X1 port map( A => n2891, B => DATAIN(12), S => n68, Z => n3315)
                           ;
   U1438 : MUX2_X1 port map( A => n2912, B => DATAIN(11), S => n67, Z => n3314)
                           ;
   U1439 : MUX2_X1 port map( A => n2933, B => DATAIN(10), S => n67, Z => n3313)
                           ;
   U1440 : MUX2_X1 port map( A => n2954, B => DATAIN(9), S => n67, Z => n3312);
   U1441 : MUX2_X1 port map( A => n2975, B => DATAIN(8), S => n67, Z => n3311);
   U1442 : MUX2_X1 port map( A => n3572, B => DATAIN(7), S => n67, Z => n3310);
   U1443 : MUX2_X1 port map( A => n3593, B => DATAIN(6), S => n67, Z => n3309);
   U1444 : MUX2_X1 port map( A => n3614, B => DATAIN(5), S => n67, Z => n3308);
   U1445 : MUX2_X1 port map( A => n3635, B => DATAIN(4), S => n67, Z => n3307);
   U1446 : MUX2_X1 port map( A => n3656, B => DATAIN(3), S => n67, Z => n3306);
   U1447 : MUX2_X1 port map( A => n3677, B => DATAIN(2), S => n67, Z => n3305);
   U1448 : MUX2_X1 port map( A => n3698, B => DATAIN(1), S => n67, Z => n3304);
   U1449 : MUX2_X1 port map( A => n3719, B => DATAIN(0), S => n67, Z => n3303);
   U1450 : AND2_X1 port map( A1 => n807, A2 => n467, ZN => n951);
   U1451 : AND3_X1 port map( A1 => n947, A2 => n946, A3 => ADD_WR(3), ZN => 
                           n467);
   U1452 : INV_X1 port map( A => ADD_WR(4), ZN => n946);
   U1453 : MUX2_X1 port map( A => n2509, B => DATAIN(31), S => n72, Z => n3302)
                           ;
   U1454 : MUX2_X1 port map( A => n2530, B => DATAIN(30), S => n72, Z => n3301)
                           ;
   U1455 : MUX2_X1 port map( A => n2551, B => DATAIN(29), S => n72, Z => n3300)
                           ;
   U1456 : MUX2_X1 port map( A => n2572, B => DATAIN(28), S => n72, Z => n3299)
                           ;
   U1457 : MUX2_X1 port map( A => n2593, B => DATAIN(27), S => n72, Z => n3298)
                           ;
   U1458 : MUX2_X1 port map( A => n2614, B => DATAIN(26), S => n72, Z => n3297)
                           ;
   U1459 : MUX2_X1 port map( A => n2635, B => DATAIN(25), S => n72, Z => n3296)
                           ;
   U1460 : MUX2_X1 port map( A => n2656, B => DATAIN(24), S => n72, Z => n3295)
                           ;
   U1461 : MUX2_X1 port map( A => n2677, B => DATAIN(23), S => n71, Z => n3294)
                           ;
   U1462 : MUX2_X1 port map( A => n2698, B => DATAIN(22), S => n71, Z => n3293)
                           ;
   U1463 : MUX2_X1 port map( A => n2719, B => DATAIN(21), S => n71, Z => n3292)
                           ;
   U1464 : MUX2_X1 port map( A => n2740, B => DATAIN(20), S => n71, Z => n3291)
                           ;
   U1465 : MUX2_X1 port map( A => n2761, B => DATAIN(19), S => n71, Z => n3290)
                           ;
   U1466 : MUX2_X1 port map( A => n2782, B => DATAIN(18), S => n71, Z => n3289)
                           ;
   U1467 : MUX2_X1 port map( A => n2803, B => DATAIN(17), S => n71, Z => n3288)
                           ;
   U1468 : MUX2_X1 port map( A => n2824, B => DATAIN(16), S => n71, Z => n3287)
                           ;
   U1469 : MUX2_X1 port map( A => n2845, B => DATAIN(15), S => n71, Z => n3286)
                           ;
   U1470 : MUX2_X1 port map( A => n2866, B => DATAIN(14), S => n71, Z => n3285)
                           ;
   U1471 : MUX2_X1 port map( A => n2887, B => DATAIN(13), S => n71, Z => n3284)
                           ;
   U1472 : MUX2_X1 port map( A => n2908, B => DATAIN(12), S => n71, Z => n3283)
                           ;
   U1473 : MUX2_X1 port map( A => n2929, B => DATAIN(11), S => n70, Z => n3282)
                           ;
   U1474 : MUX2_X1 port map( A => n2950, B => DATAIN(10), S => n70, Z => n3281)
                           ;
   U1475 : MUX2_X1 port map( A => n2971, B => DATAIN(9), S => n70, Z => n3280);
   U1476 : MUX2_X1 port map( A => n3568, B => DATAIN(8), S => n70, Z => n3279);
   U1477 : MUX2_X1 port map( A => n3589, B => DATAIN(7), S => n70, Z => n3278);
   U1478 : MUX2_X1 port map( A => n3610, B => DATAIN(6), S => n70, Z => n3277);
   U1479 : MUX2_X1 port map( A => n3631, B => DATAIN(5), S => n70, Z => n3276);
   U1480 : MUX2_X1 port map( A => n3652, B => DATAIN(4), S => n70, Z => n3275);
   U1481 : MUX2_X1 port map( A => n3673, B => DATAIN(3), S => n70, Z => n3274);
   U1482 : MUX2_X1 port map( A => n3694, B => DATAIN(2), S => n70, Z => n3273);
   U1483 : MUX2_X1 port map( A => n3715, B => DATAIN(1), S => n70, Z => n3272);
   U1484 : MUX2_X1 port map( A => n3736, B => DATAIN(0), S => n70, Z => n3271);
   U1485 : AND2_X1 port map( A1 => n841, A2 => n705, ZN => n952);
   U1486 : AND3_X1 port map( A1 => n953, A2 => n954, A3 => ADD_WR(1), ZN => 
                           n705);
   U1487 : MUX2_X1 port map( A => n2508, B => DATAIN(31), S => n75, Z => n3270)
                           ;
   U1488 : MUX2_X1 port map( A => n2529, B => DATAIN(30), S => n75, Z => n3269)
                           ;
   U1489 : MUX2_X1 port map( A => n2550, B => DATAIN(29), S => n75, Z => n3268)
                           ;
   U1490 : MUX2_X1 port map( A => n2571, B => DATAIN(28), S => n75, Z => n3267)
                           ;
   U1491 : MUX2_X1 port map( A => n2592, B => DATAIN(27), S => n75, Z => n3266)
                           ;
   U1492 : MUX2_X1 port map( A => n2613, B => DATAIN(26), S => n75, Z => n3265)
                           ;
   U1493 : MUX2_X1 port map( A => n2634, B => DATAIN(25), S => n75, Z => n3264)
                           ;
   U1494 : MUX2_X1 port map( A => n2655, B => DATAIN(24), S => n75, Z => n3263)
                           ;
   U1495 : MUX2_X1 port map( A => n2676, B => DATAIN(23), S => n74, Z => n3262)
                           ;
   U1496 : MUX2_X1 port map( A => n2697, B => DATAIN(22), S => n74, Z => n3261)
                           ;
   U1497 : MUX2_X1 port map( A => n2718, B => DATAIN(21), S => n74, Z => n3260)
                           ;
   U1498 : MUX2_X1 port map( A => n2739, B => DATAIN(20), S => n74, Z => n3259)
                           ;
   U1499 : MUX2_X1 port map( A => n2760, B => DATAIN(19), S => n74, Z => n3258)
                           ;
   U1500 : MUX2_X1 port map( A => n2781, B => DATAIN(18), S => n74, Z => n3257)
                           ;
   U1501 : MUX2_X1 port map( A => n2802, B => DATAIN(17), S => n74, Z => n3256)
                           ;
   U1502 : MUX2_X1 port map( A => n2823, B => DATAIN(16), S => n74, Z => n3255)
                           ;
   U1503 : MUX2_X1 port map( A => n2844, B => DATAIN(15), S => n74, Z => n3254)
                           ;
   U1504 : MUX2_X1 port map( A => n2865, B => DATAIN(14), S => n74, Z => n3253)
                           ;
   U1505 : MUX2_X1 port map( A => n2886, B => DATAIN(13), S => n74, Z => n3252)
                           ;
   U1506 : MUX2_X1 port map( A => n2907, B => DATAIN(12), S => n74, Z => n3251)
                           ;
   U1507 : MUX2_X1 port map( A => n2928, B => DATAIN(11), S => n73, Z => n3250)
                           ;
   U1508 : MUX2_X1 port map( A => n2949, B => DATAIN(10), S => n73, Z => n3249)
                           ;
   U1509 : MUX2_X1 port map( A => n2970, B => DATAIN(9), S => n73, Z => n3248);
   U1510 : MUX2_X1 port map( A => n3567, B => DATAIN(8), S => n73, Z => n3247);
   U1511 : MUX2_X1 port map( A => n3588, B => DATAIN(7), S => n73, Z => n3246);
   U1512 : MUX2_X1 port map( A => n3609, B => DATAIN(6), S => n73, Z => n3245);
   U1513 : MUX2_X1 port map( A => n3630, B => DATAIN(5), S => n73, Z => n3244);
   U1514 : MUX2_X1 port map( A => n3651, B => DATAIN(4), S => n73, Z => n3243);
   U1515 : MUX2_X1 port map( A => n3672, B => DATAIN(3), S => n73, Z => n3242);
   U1516 : MUX2_X1 port map( A => n3693, B => DATAIN(2), S => n73, Z => n3241);
   U1517 : MUX2_X1 port map( A => n3714, B => DATAIN(1), S => n73, Z => n3240);
   U1518 : MUX2_X1 port map( A => n3735, B => DATAIN(0), S => n73, Z => n3239);
   U1519 : AND2_X1 port map( A1 => n841, A2 => n739, ZN => n955);
   U1520 : AND3_X1 port map( A1 => ADD_WR(0), A2 => n954, A3 => ADD_WR(1), ZN 
                           => n739);
   U1521 : MUX2_X1 port map( A => n2506, B => DATAIN(31), S => n78, Z => n3238)
                           ;
   U1522 : MUX2_X1 port map( A => n2527, B => DATAIN(30), S => n78, Z => n3237)
                           ;
   U1523 : MUX2_X1 port map( A => n2548, B => DATAIN(29), S => n78, Z => n3236)
                           ;
   U1524 : MUX2_X1 port map( A => n2569, B => DATAIN(28), S => n78, Z => n3235)
                           ;
   U1525 : MUX2_X1 port map( A => n2590, B => DATAIN(27), S => n78, Z => n3234)
                           ;
   U1526 : MUX2_X1 port map( A => n2611, B => DATAIN(26), S => n78, Z => n3233)
                           ;
   U1527 : MUX2_X1 port map( A => n2632, B => DATAIN(25), S => n78, Z => n3232)
                           ;
   U1528 : MUX2_X1 port map( A => n2653, B => DATAIN(24), S => n78, Z => n3231)
                           ;
   U1529 : MUX2_X1 port map( A => n2674, B => DATAIN(23), S => n77, Z => n3230)
                           ;
   U1530 : MUX2_X1 port map( A => n2695, B => DATAIN(22), S => n77, Z => n3229)
                           ;
   U1531 : MUX2_X1 port map( A => n2716, B => DATAIN(21), S => n77, Z => n3228)
                           ;
   U1532 : MUX2_X1 port map( A => n2737, B => DATAIN(20), S => n77, Z => n3227)
                           ;
   U1533 : MUX2_X1 port map( A => n2758, B => DATAIN(19), S => n77, Z => n3226)
                           ;
   U1534 : MUX2_X1 port map( A => n2779, B => DATAIN(18), S => n77, Z => n3225)
                           ;
   U1535 : MUX2_X1 port map( A => n2800, B => DATAIN(17), S => n77, Z => n3224)
                           ;
   U1536 : MUX2_X1 port map( A => n2821, B => DATAIN(16), S => n77, Z => n3223)
                           ;
   U1537 : MUX2_X1 port map( A => n2842, B => DATAIN(15), S => n77, Z => n3222)
                           ;
   U1538 : MUX2_X1 port map( A => n2863, B => DATAIN(14), S => n77, Z => n3221)
                           ;
   U1539 : MUX2_X1 port map( A => n2884, B => DATAIN(13), S => n77, Z => n3220)
                           ;
   U1540 : MUX2_X1 port map( A => n2905, B => DATAIN(12), S => n77, Z => n3219)
                           ;
   U1541 : MUX2_X1 port map( A => n2926, B => DATAIN(11), S => n76, Z => n3218)
                           ;
   U1542 : MUX2_X1 port map( A => n2947, B => DATAIN(10), S => n76, Z => n3217)
                           ;
   U1543 : MUX2_X1 port map( A => n2968, B => DATAIN(9), S => n76, Z => n3216);
   U1544 : MUX2_X1 port map( A => n3565, B => DATAIN(8), S => n76, Z => n3215);
   U1545 : MUX2_X1 port map( A => n3586, B => DATAIN(7), S => n76, Z => n3214);
   U1546 : MUX2_X1 port map( A => n3607, B => DATAIN(6), S => n76, Z => n3213);
   U1547 : MUX2_X1 port map( A => n3628, B => DATAIN(5), S => n76, Z => n3212);
   U1548 : MUX2_X1 port map( A => n3649, B => DATAIN(4), S => n76, Z => n3211);
   U1549 : MUX2_X1 port map( A => n3670, B => DATAIN(3), S => n76, Z => n3210);
   U1550 : MUX2_X1 port map( A => n3691, B => DATAIN(2), S => n76, Z => n3209);
   U1551 : MUX2_X1 port map( A => n3712, B => DATAIN(1), S => n76, Z => n3208);
   U1552 : MUX2_X1 port map( A => n3733, B => DATAIN(0), S => n76, Z => n3207);
   U1553 : AND2_X1 port map( A1 => n841, A2 => n773, ZN => n956);
   U1554 : AND3_X1 port map( A1 => ADD_WR(2), A2 => n953, A3 => ADD_WR(1), ZN 
                           => n773);
   U1555 : MUX2_X1 port map( A => n2505, B => DATAIN(31), S => n81, Z => n3206)
                           ;
   U1556 : MUX2_X1 port map( A => n2526, B => DATAIN(30), S => n81, Z => n3205)
                           ;
   U1557 : MUX2_X1 port map( A => n2547, B => DATAIN(29), S => n81, Z => n3204)
                           ;
   U1558 : MUX2_X1 port map( A => n2568, B => DATAIN(28), S => n81, Z => n3203)
                           ;
   U1559 : MUX2_X1 port map( A => n2589, B => DATAIN(27), S => n81, Z => n3202)
                           ;
   U1560 : MUX2_X1 port map( A => n2610, B => DATAIN(26), S => n81, Z => n3201)
                           ;
   U1561 : MUX2_X1 port map( A => n2631, B => DATAIN(25), S => n81, Z => n3200)
                           ;
   U1562 : MUX2_X1 port map( A => n2652, B => DATAIN(24), S => n81, Z => n3199)
                           ;
   U1563 : MUX2_X1 port map( A => n2673, B => DATAIN(23), S => n80, Z => n3198)
                           ;
   U1564 : MUX2_X1 port map( A => n2694, B => DATAIN(22), S => n80, Z => n3197)
                           ;
   U1565 : MUX2_X1 port map( A => n2715, B => DATAIN(21), S => n80, Z => n3196)
                           ;
   U1566 : MUX2_X1 port map( A => n2736, B => DATAIN(20), S => n80, Z => n3195)
                           ;
   U1567 : MUX2_X1 port map( A => n2757, B => DATAIN(19), S => n80, Z => n3194)
                           ;
   U1568 : MUX2_X1 port map( A => n2778, B => DATAIN(18), S => n80, Z => n3193)
                           ;
   U1569 : MUX2_X1 port map( A => n2799, B => DATAIN(17), S => n80, Z => n3192)
                           ;
   U1570 : MUX2_X1 port map( A => n2820, B => DATAIN(16), S => n80, Z => n3191)
                           ;
   U1571 : MUX2_X1 port map( A => n2841, B => DATAIN(15), S => n80, Z => n3190)
                           ;
   U1572 : MUX2_X1 port map( A => n2862, B => DATAIN(14), S => n80, Z => n3189)
                           ;
   U1573 : MUX2_X1 port map( A => n2883, B => DATAIN(13), S => n80, Z => n3188)
                           ;
   U1574 : MUX2_X1 port map( A => n2904, B => DATAIN(12), S => n80, Z => n3187)
                           ;
   U1575 : MUX2_X1 port map( A => n2925, B => DATAIN(11), S => n79, Z => n3186)
                           ;
   U1576 : MUX2_X1 port map( A => n2946, B => DATAIN(10), S => n79, Z => n3185)
                           ;
   U1577 : MUX2_X1 port map( A => n2967, B => DATAIN(9), S => n79, Z => n3184);
   U1578 : MUX2_X1 port map( A => n3564, B => DATAIN(8), S => n79, Z => n3183);
   U1579 : MUX2_X1 port map( A => n3585, B => DATAIN(7), S => n79, Z => n3182);
   U1580 : MUX2_X1 port map( A => n3606, B => DATAIN(6), S => n79, Z => n3181);
   U1581 : MUX2_X1 port map( A => n3627, B => DATAIN(5), S => n79, Z => n3180);
   U1582 : MUX2_X1 port map( A => n3648, B => DATAIN(4), S => n79, Z => n3179);
   U1583 : MUX2_X1 port map( A => n3669, B => DATAIN(3), S => n79, Z => n3178);
   U1584 : MUX2_X1 port map( A => n3690, B => DATAIN(2), S => n79, Z => n3177);
   U1585 : MUX2_X1 port map( A => n3711, B => DATAIN(1), S => n79, Z => n3176);
   U1586 : MUX2_X1 port map( A => n3732, B => DATAIN(0), S => n79, Z => n3175);
   U1587 : AND2_X1 port map( A1 => n841, A2 => n807, ZN => n957);
   U1588 : AND3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => ADD_WR(1),
                           ZN => n807);
   U1589 : AND3_X1 port map( A1 => n947, A2 => n945, A3 => ADD_WR(4), ZN => 
                           n841);
   U1590 : INV_X1 port map( A => ADD_WR(3), ZN => n945);
   U1591 : MUX2_X1 port map( A => n2503, B => DATAIN(31), S => n84, Z => n3174)
                           ;
   U1592 : MUX2_X1 port map( A => n2524, B => DATAIN(30), S => n84, Z => n3173)
                           ;
   U1593 : MUX2_X1 port map( A => n2545, B => DATAIN(29), S => n84, Z => n3172)
                           ;
   U1594 : MUX2_X1 port map( A => n2566, B => DATAIN(28), S => n84, Z => n3171)
                           ;
   U1595 : MUX2_X1 port map( A => n2587, B => DATAIN(27), S => n84, Z => n3170)
                           ;
   U1596 : MUX2_X1 port map( A => n2608, B => DATAIN(26), S => n84, Z => n3169)
                           ;
   U1597 : MUX2_X1 port map( A => n2629, B => DATAIN(25), S => n84, Z => n3168)
                           ;
   U1598 : MUX2_X1 port map( A => n2650, B => DATAIN(24), S => n84, Z => n3167)
                           ;
   U1599 : MUX2_X1 port map( A => n2671, B => DATAIN(23), S => n83, Z => n3166)
                           ;
   U1600 : MUX2_X1 port map( A => n2692, B => DATAIN(22), S => n83, Z => n3165)
                           ;
   U1601 : MUX2_X1 port map( A => n2713, B => DATAIN(21), S => n83, Z => n3164)
                           ;
   U1602 : MUX2_X1 port map( A => n2734, B => DATAIN(20), S => n83, Z => n3163)
                           ;
   U1603 : MUX2_X1 port map( A => n2755, B => DATAIN(19), S => n83, Z => n3162)
                           ;
   U1604 : MUX2_X1 port map( A => n2776, B => DATAIN(18), S => n83, Z => n3161)
                           ;
   U1605 : MUX2_X1 port map( A => n2797, B => DATAIN(17), S => n83, Z => n3160)
                           ;
   U1606 : MUX2_X1 port map( A => n2818, B => DATAIN(16), S => n83, Z => n3159)
                           ;
   U1607 : MUX2_X1 port map( A => n2839, B => DATAIN(15), S => n83, Z => n3158)
                           ;
   U1608 : MUX2_X1 port map( A => n2860, B => DATAIN(14), S => n83, Z => n3157)
                           ;
   U1609 : MUX2_X1 port map( A => n2881, B => DATAIN(13), S => n83, Z => n3156)
                           ;
   U1610 : MUX2_X1 port map( A => n2902, B => DATAIN(12), S => n83, Z => n3155)
                           ;
   U1611 : MUX2_X1 port map( A => n2923, B => DATAIN(11), S => n82, Z => n3154)
                           ;
   U1612 : MUX2_X1 port map( A => n2944, B => DATAIN(10), S => n82, Z => n3153)
                           ;
   U1613 : MUX2_X1 port map( A => n2965, B => DATAIN(9), S => n82, Z => n3152);
   U1614 : MUX2_X1 port map( A => n3562, B => DATAIN(8), S => n82, Z => n3151);
   U1615 : MUX2_X1 port map( A => n3583, B => DATAIN(7), S => n82, Z => n3150);
   U1616 : MUX2_X1 port map( A => n3604, B => DATAIN(6), S => n82, Z => n3149);
   U1617 : MUX2_X1 port map( A => n3625, B => DATAIN(5), S => n82, Z => n3148);
   U1618 : MUX2_X1 port map( A => n3646, B => DATAIN(4), S => n82, Z => n3147);
   U1619 : MUX2_X1 port map( A => n3667, B => DATAIN(3), S => n82, Z => n3146);
   U1620 : MUX2_X1 port map( A => n3688, B => DATAIN(2), S => n82, Z => n3145);
   U1621 : MUX2_X1 port map( A => n3709, B => DATAIN(1), S => n82, Z => n3144);
   U1622 : MUX2_X1 port map( A => n3730, B => DATAIN(0), S => n82, Z => n3143);
   U1623 : AND2_X1 port map( A1 => n704, A2 => n468, ZN => n958);
   U1624 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => ADD_WR(0),
                           ZN => n468);
   U1625 : MUX2_X1 port map( A => n2502, B => DATAIN(31), S => n87, Z => n3142)
                           ;
   U1626 : MUX2_X1 port map( A => n2523, B => DATAIN(30), S => n87, Z => n3141)
                           ;
   U1627 : MUX2_X1 port map( A => n2544, B => DATAIN(29), S => n87, Z => n3140)
                           ;
   U1628 : MUX2_X1 port map( A => n2565, B => DATAIN(28), S => n87, Z => n3139)
                           ;
   U1629 : MUX2_X1 port map( A => n2586, B => DATAIN(27), S => n87, Z => n3138)
                           ;
   U1630 : MUX2_X1 port map( A => n2607, B => DATAIN(26), S => n87, Z => n3137)
                           ;
   U1631 : MUX2_X1 port map( A => n2628, B => DATAIN(25), S => n87, Z => n3136)
                           ;
   U1632 : MUX2_X1 port map( A => n2649, B => DATAIN(24), S => n87, Z => n3135)
                           ;
   U1633 : MUX2_X1 port map( A => n2670, B => DATAIN(23), S => n86, Z => n3134)
                           ;
   U1634 : MUX2_X1 port map( A => n2691, B => DATAIN(22), S => n86, Z => n3133)
                           ;
   U1635 : MUX2_X1 port map( A => n2712, B => DATAIN(21), S => n86, Z => n3132)
                           ;
   U1636 : MUX2_X1 port map( A => n2733, B => DATAIN(20), S => n86, Z => n3131)
                           ;
   U1637 : MUX2_X1 port map( A => n2754, B => DATAIN(19), S => n86, Z => n3130)
                           ;
   U1638 : MUX2_X1 port map( A => n2775, B => DATAIN(18), S => n86, Z => n3129)
                           ;
   U1639 : MUX2_X1 port map( A => n2796, B => DATAIN(17), S => n86, Z => n3128)
                           ;
   U1640 : MUX2_X1 port map( A => n2817, B => DATAIN(16), S => n86, Z => n3127)
                           ;
   U1641 : MUX2_X1 port map( A => n2838, B => DATAIN(15), S => n86, Z => n3126)
                           ;
   U1642 : MUX2_X1 port map( A => n2859, B => DATAIN(14), S => n86, Z => n3125)
                           ;
   U1643 : MUX2_X1 port map( A => n2880, B => DATAIN(13), S => n86, Z => n3124)
                           ;
   U1644 : MUX2_X1 port map( A => n2901, B => DATAIN(12), S => n86, Z => n3123)
                           ;
   U1645 : MUX2_X1 port map( A => n2922, B => DATAIN(11), S => n85, Z => n3122)
                           ;
   U1646 : MUX2_X1 port map( A => n2943, B => DATAIN(10), S => n85, Z => n3121)
                           ;
   U1647 : MUX2_X1 port map( A => n2964, B => DATAIN(9), S => n85, Z => n3120);
   U1648 : MUX2_X1 port map( A => n3561, B => DATAIN(8), S => n85, Z => n3119);
   U1649 : MUX2_X1 port map( A => n3582, B => DATAIN(7), S => n85, Z => n3118);
   U1650 : MUX2_X1 port map( A => n3603, B => DATAIN(6), S => n85, Z => n3117);
   U1651 : MUX2_X1 port map( A => n3624, B => DATAIN(5), S => n85, Z => n3116);
   U1652 : MUX2_X1 port map( A => n3645, B => DATAIN(4), S => n85, Z => n3115);
   U1653 : MUX2_X1 port map( A => n3666, B => DATAIN(3), S => n85, Z => n3114);
   U1654 : MUX2_X1 port map( A => n3687, B => DATAIN(2), S => n85, Z => n3113);
   U1655 : MUX2_X1 port map( A => n3708, B => DATAIN(1), S => n85, Z => n3112);
   U1656 : MUX2_X1 port map( A => n3729, B => DATAIN(0), S => n85, Z => n3111);
   U1657 : AND2_X1 port map( A1 => n704, A2 => n502, ZN => n959);
   U1658 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => n953, ZN 
                           => n502);
   U1659 : MUX2_X1 port map( A => n3832, B => DATAIN(31), S => n90, Z => n3110)
                           ;
   U1660 : MUX2_X1 port map( A => n3831, B => DATAIN(30), S => n90, Z => n3109)
                           ;
   U1661 : MUX2_X1 port map( A => n3830, B => DATAIN(29), S => n90, Z => n3108)
                           ;
   U1662 : MUX2_X1 port map( A => n3829, B => DATAIN(28), S => n90, Z => n3107)
                           ;
   U1663 : MUX2_X1 port map( A => n3828, B => DATAIN(27), S => n90, Z => n3106)
                           ;
   U1664 : MUX2_X1 port map( A => n3827, B => DATAIN(26), S => n90, Z => n3105)
                           ;
   U1665 : MUX2_X1 port map( A => n3826, B => DATAIN(25), S => n90, Z => n3104)
                           ;
   U1666 : MUX2_X1 port map( A => n3825, B => DATAIN(24), S => n90, Z => n3103)
                           ;
   U1667 : MUX2_X1 port map( A => n3824, B => DATAIN(23), S => n89, Z => n3102)
                           ;
   U1668 : MUX2_X1 port map( A => n3823, B => DATAIN(22), S => n89, Z => n3101)
                           ;
   U1669 : MUX2_X1 port map( A => n3822, B => DATAIN(21), S => n89, Z => n3100)
                           ;
   U1670 : MUX2_X1 port map( A => n3821, B => DATAIN(20), S => n89, Z => n3099)
                           ;
   U1671 : MUX2_X1 port map( A => n3820, B => DATAIN(19), S => n89, Z => n3098)
                           ;
   U1672 : MUX2_X1 port map( A => n3819, B => DATAIN(18), S => n89, Z => n3097)
                           ;
   U1673 : MUX2_X1 port map( A => n3818, B => DATAIN(17), S => n89, Z => n3096)
                           ;
   U1674 : MUX2_X1 port map( A => n3817, B => DATAIN(16), S => n89, Z => n3095)
                           ;
   U1675 : MUX2_X1 port map( A => n3816, B => DATAIN(15), S => n89, Z => n3094)
                           ;
   U1676 : MUX2_X1 port map( A => n3815, B => DATAIN(14), S => n89, Z => n3093)
                           ;
   U1677 : MUX2_X1 port map( A => n3814, B => DATAIN(13), S => n89, Z => n3092)
                           ;
   U1678 : MUX2_X1 port map( A => n3813, B => DATAIN(12), S => n89, Z => n3091)
                           ;
   U1679 : MUX2_X1 port map( A => n3812, B => DATAIN(11), S => n88, Z => n3090)
                           ;
   U1680 : MUX2_X1 port map( A => n3811, B => DATAIN(10), S => n88, Z => n3089)
                           ;
   U1681 : MUX2_X1 port map( A => n3810, B => DATAIN(9), S => n88, Z => n3088);
   U1682 : MUX2_X1 port map( A => n3809, B => DATAIN(8), S => n88, Z => n3087);
   U1683 : MUX2_X1 port map( A => n3808, B => DATAIN(7), S => n88, Z => n3086);
   U1684 : MUX2_X1 port map( A => n3807, B => DATAIN(6), S => n88, Z => n3085);
   U1685 : MUX2_X1 port map( A => n3806, B => DATAIN(5), S => n88, Z => n3084);
   U1686 : MUX2_X1 port map( A => n3805, B => DATAIN(4), S => n88, Z => n3083);
   U1687 : MUX2_X1 port map( A => n3804, B => DATAIN(3), S => n88, Z => n3082);
   U1688 : MUX2_X1 port map( A => n3803, B => DATAIN(2), S => n88, Z => n3081);
   U1689 : MUX2_X1 port map( A => n3802, B => DATAIN(1), S => n88, Z => n3080);
   U1690 : MUX2_X1 port map( A => n3801, B => DATAIN(0), S => n88, Z => n3079);
   U1691 : AND2_X1 port map( A1 => n704, A2 => n536, ZN => n960);
   U1692 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n954, ZN 
                           => n536);
   U1693 : MUX2_X1 port map( A => n3800, B => DATAIN(31), S => n93, Z => n3078)
                           ;
   U1694 : MUX2_X1 port map( A => n3799, B => DATAIN(30), S => n93, Z => n3077)
                           ;
   U1695 : MUX2_X1 port map( A => n3798, B => DATAIN(29), S => n93, Z => n3076)
                           ;
   U1696 : MUX2_X1 port map( A => n3797, B => DATAIN(28), S => n93, Z => n3075)
                           ;
   U1697 : MUX2_X1 port map( A => n3796, B => DATAIN(27), S => n93, Z => n3074)
                           ;
   U1698 : MUX2_X1 port map( A => n3795, B => DATAIN(26), S => n93, Z => n3073)
                           ;
   U1699 : MUX2_X1 port map( A => n3794, B => DATAIN(25), S => n93, Z => n3072)
                           ;
   U1700 : MUX2_X1 port map( A => n3793, B => DATAIN(24), S => n93, Z => n3071)
                           ;
   U1701 : MUX2_X1 port map( A => n3792, B => DATAIN(23), S => n92, Z => n3070)
                           ;
   U1702 : MUX2_X1 port map( A => n3791, B => DATAIN(22), S => n92, Z => n3069)
                           ;
   U1703 : MUX2_X1 port map( A => n3790, B => DATAIN(21), S => n92, Z => n3068)
                           ;
   U1704 : MUX2_X1 port map( A => n3789, B => DATAIN(20), S => n92, Z => n3067)
                           ;
   U1705 : MUX2_X1 port map( A => n3788, B => DATAIN(19), S => n92, Z => n3066)
                           ;
   U1706 : MUX2_X1 port map( A => n3787, B => DATAIN(18), S => n92, Z => n3065)
                           ;
   U1707 : MUX2_X1 port map( A => n3786, B => DATAIN(17), S => n92, Z => n3064)
                           ;
   U1708 : MUX2_X1 port map( A => n3785, B => DATAIN(16), S => n92, Z => n3063)
                           ;
   U1709 : MUX2_X1 port map( A => n3784, B => DATAIN(15), S => n92, Z => n3062)
                           ;
   U1710 : MUX2_X1 port map( A => n3783, B => DATAIN(14), S => n92, Z => n3061)
                           ;
   U1711 : MUX2_X1 port map( A => n3782, B => DATAIN(13), S => n92, Z => n3060)
                           ;
   U1712 : MUX2_X1 port map( A => n3781, B => DATAIN(12), S => n92, Z => n3059)
                           ;
   U1713 : MUX2_X1 port map( A => n3780, B => DATAIN(11), S => n91, Z => n3058)
                           ;
   U1714 : MUX2_X1 port map( A => n3779, B => DATAIN(10), S => n91, Z => n3057)
                           ;
   U1715 : MUX2_X1 port map( A => n3778, B => DATAIN(9), S => n91, Z => n3056);
   U1716 : MUX2_X1 port map( A => n3777, B => DATAIN(8), S => n91, Z => n3055);
   U1717 : MUX2_X1 port map( A => n3776, B => DATAIN(7), S => n91, Z => n3054);
   U1718 : MUX2_X1 port map( A => n3775, B => DATAIN(6), S => n91, Z => n3053);
   U1719 : MUX2_X1 port map( A => n3774, B => DATAIN(5), S => n91, Z => n3052);
   U1720 : MUX2_X1 port map( A => n3773, B => DATAIN(4), S => n91, Z => n3051);
   U1721 : MUX2_X1 port map( A => n3772, B => DATAIN(3), S => n91, Z => n3050);
   U1722 : MUX2_X1 port map( A => n3771, B => DATAIN(2), S => n91, Z => n3049);
   U1723 : MUX2_X1 port map( A => n3770, B => DATAIN(1), S => n91, Z => n3048);
   U1724 : MUX2_X1 port map( A => n3769, B => DATAIN(0), S => n91, Z => n3047);
   U1725 : AND2_X1 port map( A1 => n704, A2 => n570, ZN => n961);
   U1726 : NOR3_X1 port map( A1 => n953, A2 => ADD_WR(1), A3 => n954, ZN => 
                           n570);
   U1727 : INV_X1 port map( A => ADD_WR(2), ZN => n954);
   U1728 : AND3_X1 port map( A1 => ADD_WR(3), A2 => n947, A3 => ADD_WR(4), ZN 
                           => n704);
   U1729 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n947);
   U1730 : OAI222_X1 port map( A1 => n298, A2 => n96, B1 => n963, B2 => n99, C1
                           => n3716, C2 => n102, ZN => n3046);
   U1731 : NOR4_X1 port map( A1 => n966, A2 => n967, A3 => n968, A4 => n969, ZN
                           => n963);
   U1732 : OAI221_X1 port map( B1 => n3833, B2 => n105, C1 => n971, C2 => n108,
                           A => n973, ZN => n969);
   U1733 : AOI22_X1 port map( A1 => n111, A2 => n3730, B1 => n114, B2 => n673, 
                           ZN => n973);
   U1734 : OAI221_X1 port map( B1 => n976, B2 => n117, C1 => n3737, C2 => n120,
                           A => n979, ZN => n968);
   U1735 : AOI22_X1 port map( A1 => n123, A2 => n774, B1 => n126, B2 => n3729, 
                           ZN => n979);
   U1736 : OAI211_X1 port map( C1 => n3734, C2 => n129, A => n983, B => n984, 
                           ZN => n967);
   U1737 : AOI221_X1 port map( B1 => n132, B2 => n908, C1 => n135, C2 => n3735,
                           A => n987, ZN => n984);
   U1738 : OAI22_X1 port map( A1 => n3731, A2 => n138, B1 => n989, B2 => n141, 
                           ZN => n987);
   U1739 : AOI22_X1 port map( A1 => n144, A2 => n3736, B1 => n147, B2 => n808, 
                           ZN => n983);
   U1740 : NAND4_X1 port map( A1 => n993, A2 => n994, A3 => n995, A4 => n996, 
                           ZN => n966);
   U1741 : AOI221_X1 port map( B1 => n150, B2 => n3719, C1 => n153, C2 => n3720
                           , A => n999, ZN => n996);
   U1742 : OAI22_X1 port map( A1 => n3718, A2 => n156, B1 => n3717, B2 => n159,
                           ZN => n999);
   U1743 : AOI221_X1 port map( B1 => n162, B2 => n3723, C1 => n165, C2 => n3724
                           , A => n1004, ZN => n995);
   U1744 : OAI22_X1 port map( A1 => n3722, A2 => n168, B1 => n3721, B2 => n171,
                           ZN => n1004);
   U1745 : AOI221_X1 port map( B1 => n174, B2 => n605, C1 => n177, C2 => n638, 
                           A => n1009, ZN => n994);
   U1746 : OAI22_X1 port map( A1 => n1010, A2 => n180, B1 => n1012, B2 => n183,
                           ZN => n1009);
   U1747 : AOI221_X1 port map( B1 => n186, B2 => n571, C1 => n189, C2 => n3769,
                           A => n1016, ZN => n993);
   U1748 : OAI22_X1 port map( A1 => n1017, A2 => n192, B1 => n1019, B2 => n195,
                           ZN => n1016);
   U1749 : OAI222_X1 port map( A1 => n299, A2 => n96, B1 => n1021, B2 => n99, 
                           C1 => n3695, C2 => n102, ZN => n3045);
   U1750 : NOR4_X1 port map( A1 => n1022, A2 => n1023, A3 => n1024, A4 => n1025
                           , ZN => n1021);
   U1751 : OAI221_X1 port map( B1 => n3834, B2 => n105, C1 => n1026, C2 => n108
                           , A => n1027, ZN => n1025);
   U1752 : AOI22_X1 port map( A1 => n111, A2 => n3709, B1 => n114, B2 => n674, 
                           ZN => n1027);
   U1753 : OAI221_X1 port map( B1 => n1028, B2 => n117, C1 => n3738, C2 => n120
                           , A => n1029, ZN => n1024);
   U1754 : AOI22_X1 port map( A1 => n123, A2 => n776, B1 => n126, B2 => n3708, 
                           ZN => n1029);
   U1755 : OAI211_X1 port map( C1 => n3713, C2 => n129, A => n1030, B => n1031,
                           ZN => n1023);
   U1756 : AOI221_X1 port map( B1 => n132, B2 => n910, C1 => n135, C2 => n3714,
                           A => n1032, ZN => n1031);
   U1757 : OAI22_X1 port map( A1 => n3710, A2 => n138, B1 => n1033, B2 => n141,
                           ZN => n1032);
   U1758 : AOI22_X1 port map( A1 => n144, A2 => n3715, B1 => n147, B2 => n810, 
                           ZN => n1030);
   U1759 : NAND4_X1 port map( A1 => n1034, A2 => n1035, A3 => n1036, A4 => 
                           n1037, ZN => n1022);
   U1760 : AOI221_X1 port map( B1 => n150, B2 => n3698, C1 => n153, C2 => n3699
                           , A => n1038, ZN => n1037);
   U1761 : OAI22_X1 port map( A1 => n3697, A2 => n156, B1 => n3696, B2 => n159,
                           ZN => n1038);
   U1762 : AOI221_X1 port map( B1 => n162, B2 => n3702, C1 => n165, C2 => n3703
                           , A => n1039, ZN => n1036);
   U1763 : OAI22_X1 port map( A1 => n3701, A2 => n168, B1 => n3700, B2 => n171,
                           ZN => n1039);
   U1764 : AOI221_X1 port map( B1 => n174, B2 => n607, C1 => n177, C2 => n640, 
                           A => n1040, ZN => n1035);
   U1765 : OAI22_X1 port map( A1 => n1041, A2 => n180, B1 => n1042, B2 => n183,
                           ZN => n1040);
   U1766 : AOI221_X1 port map( B1 => n186, B2 => n573, C1 => n189, C2 => n3770,
                           A => n1043, ZN => n1034);
   U1767 : OAI22_X1 port map( A1 => n1044, A2 => n192, B1 => n1045, B2 => n195,
                           ZN => n1043);
   U1768 : OAI222_X1 port map( A1 => n300, A2 => n96, B1 => n1046, B2 => n99, 
                           C1 => n3674, C2 => n102, ZN => n3044);
   U1769 : NOR4_X1 port map( A1 => n1047, A2 => n1048, A3 => n1049, A4 => n1050
                           , ZN => n1046);
   U1770 : OAI221_X1 port map( B1 => n3835, B2 => n105, C1 => n1051, C2 => n108
                           , A => n1052, ZN => n1050);
   U1771 : AOI22_X1 port map( A1 => n111, A2 => n3688, B1 => n114, B2 => n675, 
                           ZN => n1052);
   U1772 : OAI221_X1 port map( B1 => n1053, B2 => n117, C1 => n3739, C2 => n120
                           , A => n1054, ZN => n1049);
   U1773 : AOI22_X1 port map( A1 => n123, A2 => n777, B1 => n126, B2 => n3687, 
                           ZN => n1054);
   U1774 : OAI211_X1 port map( C1 => n3692, C2 => n129, A => n1055, B => n1056,
                           ZN => n1048);
   U1775 : AOI221_X1 port map( B1 => n132, B2 => n911, C1 => n135, C2 => n3693,
                           A => n1057, ZN => n1056);
   U1776 : OAI22_X1 port map( A1 => n3689, A2 => n138, B1 => n1058, B2 => n141,
                           ZN => n1057);
   U1777 : AOI22_X1 port map( A1 => n144, A2 => n3694, B1 => n147, B2 => n811, 
                           ZN => n1055);
   U1778 : NAND4_X1 port map( A1 => n1059, A2 => n1060, A3 => n1061, A4 => 
                           n1062, ZN => n1047);
   U1779 : AOI221_X1 port map( B1 => n150, B2 => n3677, C1 => n153, C2 => n3678
                           , A => n1063, ZN => n1062);
   U1780 : OAI22_X1 port map( A1 => n3676, A2 => n156, B1 => n3675, B2 => n159,
                           ZN => n1063);
   U1781 : AOI221_X1 port map( B1 => n162, B2 => n3681, C1 => n165, C2 => n3682
                           , A => n1064, ZN => n1061);
   U1782 : OAI22_X1 port map( A1 => n3680, A2 => n168, B1 => n3679, B2 => n171,
                           ZN => n1064);
   U1783 : AOI221_X1 port map( B1 => n174, B2 => n608, C1 => n177, C2 => n641, 
                           A => n1065, ZN => n1060);
   U1784 : OAI22_X1 port map( A1 => n1066, A2 => n180, B1 => n1067, B2 => n183,
                           ZN => n1065);
   U1785 : AOI221_X1 port map( B1 => n186, B2 => n574, C1 => n189, C2 => n3771,
                           A => n1068, ZN => n1059);
   U1786 : OAI22_X1 port map( A1 => n1069, A2 => n192, B1 => n1070, B2 => n195,
                           ZN => n1068);
   U1787 : OAI222_X1 port map( A1 => n301, A2 => n96, B1 => n1071, B2 => n99, 
                           C1 => n3653, C2 => n102, ZN => n3043);
   U1788 : NOR4_X1 port map( A1 => n1072, A2 => n1073, A3 => n1074, A4 => n1075
                           , ZN => n1071);
   U1789 : OAI221_X1 port map( B1 => n3836, B2 => n105, C1 => n1076, C2 => n108
                           , A => n1077, ZN => n1075);
   U1790 : AOI22_X1 port map( A1 => n111, A2 => n3667, B1 => n114, B2 => n676, 
                           ZN => n1077);
   U1791 : OAI221_X1 port map( B1 => n1078, B2 => n117, C1 => n3740, C2 => n120
                           , A => n1079, ZN => n1074);
   U1792 : AOI22_X1 port map( A1 => n123, A2 => n778, B1 => n126, B2 => n3666, 
                           ZN => n1079);
   U1793 : OAI211_X1 port map( C1 => n3671, C2 => n129, A => n1080, B => n1081,
                           ZN => n1073);
   U1794 : AOI221_X1 port map( B1 => n132, B2 => n912, C1 => n135, C2 => n3672,
                           A => n1082, ZN => n1081);
   U1795 : OAI22_X1 port map( A1 => n3668, A2 => n138, B1 => n1083, B2 => n141,
                           ZN => n1082);
   U1796 : AOI22_X1 port map( A1 => n144, A2 => n3673, B1 => n147, B2 => n812, 
                           ZN => n1080);
   U1797 : NAND4_X1 port map( A1 => n1084, A2 => n1085, A3 => n1086, A4 => 
                           n1087, ZN => n1072);
   U1798 : AOI221_X1 port map( B1 => n150, B2 => n3656, C1 => n153, C2 => n3657
                           , A => n1088, ZN => n1087);
   U1799 : OAI22_X1 port map( A1 => n3655, A2 => n156, B1 => n3654, B2 => n159,
                           ZN => n1088);
   U1800 : AOI221_X1 port map( B1 => n162, B2 => n3660, C1 => n165, C2 => n3661
                           , A => n1089, ZN => n1086);
   U1801 : OAI22_X1 port map( A1 => n3659, A2 => n168, B1 => n3658, B2 => n171,
                           ZN => n1089);
   U1802 : AOI221_X1 port map( B1 => n174, B2 => n609, C1 => n177, C2 => n642, 
                           A => n1090, ZN => n1085);
   U1803 : OAI22_X1 port map( A1 => n1091, A2 => n180, B1 => n1092, B2 => n183,
                           ZN => n1090);
   U1804 : AOI221_X1 port map( B1 => n186, B2 => n575, C1 => n189, C2 => n3772,
                           A => n1093, ZN => n1084);
   U1805 : OAI22_X1 port map( A1 => n1094, A2 => n192, B1 => n1095, B2 => n195,
                           ZN => n1093);
   U1806 : OAI222_X1 port map( A1 => n302, A2 => n96, B1 => n1096, B2 => n99, 
                           C1 => n3632, C2 => n102, ZN => n3042);
   U1807 : NOR4_X1 port map( A1 => n1097, A2 => n1098, A3 => n1099, A4 => n1100
                           , ZN => n1096);
   U1808 : OAI221_X1 port map( B1 => n3837, B2 => n105, C1 => n1101, C2 => n108
                           , A => n1102, ZN => n1100);
   U1809 : AOI22_X1 port map( A1 => n111, A2 => n3646, B1 => n114, B2 => n677, 
                           ZN => n1102);
   U1810 : OAI221_X1 port map( B1 => n1103, B2 => n117, C1 => n3741, C2 => n120
                           , A => n1104, ZN => n1099);
   U1811 : AOI22_X1 port map( A1 => n123, A2 => n779, B1 => n126, B2 => n3645, 
                           ZN => n1104);
   U1812 : OAI211_X1 port map( C1 => n3650, C2 => n129, A => n1105, B => n1106,
                           ZN => n1098);
   U1813 : AOI221_X1 port map( B1 => n132, B2 => n913, C1 => n135, C2 => n3651,
                           A => n1107, ZN => n1106);
   U1814 : OAI22_X1 port map( A1 => n3647, A2 => n138, B1 => n1108, B2 => n141,
                           ZN => n1107);
   U1815 : AOI22_X1 port map( A1 => n144, A2 => n3652, B1 => n147, B2 => n813, 
                           ZN => n1105);
   U1816 : NAND4_X1 port map( A1 => n1109, A2 => n1110, A3 => n1111, A4 => 
                           n1112, ZN => n1097);
   U1817 : AOI221_X1 port map( B1 => n150, B2 => n3635, C1 => n153, C2 => n3636
                           , A => n1113, ZN => n1112);
   U1818 : OAI22_X1 port map( A1 => n3634, A2 => n156, B1 => n3633, B2 => n159,
                           ZN => n1113);
   U1819 : AOI221_X1 port map( B1 => n162, B2 => n3639, C1 => n165, C2 => n3640
                           , A => n1114, ZN => n1111);
   U1820 : OAI22_X1 port map( A1 => n3638, A2 => n168, B1 => n3637, B2 => n171,
                           ZN => n1114);
   U1821 : AOI221_X1 port map( B1 => n174, B2 => n610, C1 => n177, C2 => n643, 
                           A => n1115, ZN => n1110);
   U1822 : OAI22_X1 port map( A1 => n1116, A2 => n180, B1 => n1117, B2 => n183,
                           ZN => n1115);
   U1823 : AOI221_X1 port map( B1 => n186, B2 => n576, C1 => n189, C2 => n3773,
                           A => n1118, ZN => n1109);
   U1824 : OAI22_X1 port map( A1 => n1119, A2 => n192, B1 => n1120, B2 => n195,
                           ZN => n1118);
   U1825 : OAI222_X1 port map( A1 => n303, A2 => n96, B1 => n1121, B2 => n99, 
                           C1 => n3611, C2 => n102, ZN => n3041);
   U1826 : NOR4_X1 port map( A1 => n1122, A2 => n1123, A3 => n1124, A4 => n1125
                           , ZN => n1121);
   U1827 : OAI221_X1 port map( B1 => n3838, B2 => n105, C1 => n1126, C2 => n108
                           , A => n1127, ZN => n1125);
   U1828 : AOI22_X1 port map( A1 => n111, A2 => n3625, B1 => n114, B2 => n678, 
                           ZN => n1127);
   U1829 : OAI221_X1 port map( B1 => n1128, B2 => n117, C1 => n3742, C2 => n120
                           , A => n1129, ZN => n1124);
   U1830 : AOI22_X1 port map( A1 => n123, A2 => n780, B1 => n126, B2 => n3624, 
                           ZN => n1129);
   U1831 : OAI211_X1 port map( C1 => n3629, C2 => n129, A => n1130, B => n1131,
                           ZN => n1123);
   U1832 : AOI221_X1 port map( B1 => n132, B2 => n914, C1 => n135, C2 => n3630,
                           A => n1132, ZN => n1131);
   U1833 : OAI22_X1 port map( A1 => n3626, A2 => n138, B1 => n1133, B2 => n141,
                           ZN => n1132);
   U1834 : AOI22_X1 port map( A1 => n144, A2 => n3631, B1 => n147, B2 => n814, 
                           ZN => n1130);
   U1835 : NAND4_X1 port map( A1 => n1134, A2 => n1135, A3 => n1136, A4 => 
                           n1137, ZN => n1122);
   U1836 : AOI221_X1 port map( B1 => n150, B2 => n3614, C1 => n153, C2 => n3615
                           , A => n1138, ZN => n1137);
   U1837 : OAI22_X1 port map( A1 => n3613, A2 => n156, B1 => n3612, B2 => n159,
                           ZN => n1138);
   U1838 : AOI221_X1 port map( B1 => n162, B2 => n3618, C1 => n165, C2 => n3619
                           , A => n1139, ZN => n1136);
   U1839 : OAI22_X1 port map( A1 => n3617, A2 => n168, B1 => n3616, B2 => n171,
                           ZN => n1139);
   U1840 : AOI221_X1 port map( B1 => n174, B2 => n611, C1 => n177, C2 => n644, 
                           A => n1140, ZN => n1135);
   U1841 : OAI22_X1 port map( A1 => n1141, A2 => n180, B1 => n1142, B2 => n183,
                           ZN => n1140);
   U1842 : AOI221_X1 port map( B1 => n186, B2 => n577, C1 => n189, C2 => n3774,
                           A => n1143, ZN => n1134);
   U1843 : OAI22_X1 port map( A1 => n1144, A2 => n192, B1 => n1145, B2 => n195,
                           ZN => n1143);
   U1844 : OAI222_X1 port map( A1 => n304, A2 => n96, B1 => n1146, B2 => n99, 
                           C1 => n3590, C2 => n102, ZN => n3040);
   U1845 : NOR4_X1 port map( A1 => n1147, A2 => n1148, A3 => n1149, A4 => n1150
                           , ZN => n1146);
   U1846 : OAI221_X1 port map( B1 => n3839, B2 => n105, C1 => n1151, C2 => n108
                           , A => n1152, ZN => n1150);
   U1847 : AOI22_X1 port map( A1 => n111, A2 => n3604, B1 => n114, B2 => n679, 
                           ZN => n1152);
   U1848 : OAI221_X1 port map( B1 => n1153, B2 => n117, C1 => n3743, C2 => n120
                           , A => n1154, ZN => n1149);
   U1849 : AOI22_X1 port map( A1 => n123, A2 => n781, B1 => n126, B2 => n3603, 
                           ZN => n1154);
   U1850 : OAI211_X1 port map( C1 => n3608, C2 => n129, A => n1155, B => n1156,
                           ZN => n1148);
   U1851 : AOI221_X1 port map( B1 => n132, B2 => n915, C1 => n135, C2 => n3609,
                           A => n1157, ZN => n1156);
   U1852 : OAI22_X1 port map( A1 => n3605, A2 => n138, B1 => n1158, B2 => n141,
                           ZN => n1157);
   U1853 : AOI22_X1 port map( A1 => n144, A2 => n3610, B1 => n147, B2 => n815, 
                           ZN => n1155);
   U1854 : NAND4_X1 port map( A1 => n1159, A2 => n1160, A3 => n1161, A4 => 
                           n1162, ZN => n1147);
   U1855 : AOI221_X1 port map( B1 => n150, B2 => n3593, C1 => n153, C2 => n3594
                           , A => n1163, ZN => n1162);
   U1856 : OAI22_X1 port map( A1 => n3592, A2 => n156, B1 => n3591, B2 => n159,
                           ZN => n1163);
   U1857 : AOI221_X1 port map( B1 => n162, B2 => n3597, C1 => n165, C2 => n3598
                           , A => n1164, ZN => n1161);
   U1858 : OAI22_X1 port map( A1 => n3596, A2 => n168, B1 => n3595, B2 => n171,
                           ZN => n1164);
   U1859 : AOI221_X1 port map( B1 => n174, B2 => n612, C1 => n177, C2 => n645, 
                           A => n1165, ZN => n1160);
   U1860 : OAI22_X1 port map( A1 => n1166, A2 => n180, B1 => n1167, B2 => n183,
                           ZN => n1165);
   U1861 : AOI221_X1 port map( B1 => n186, B2 => n578, C1 => n189, C2 => n3775,
                           A => n1168, ZN => n1159);
   U1862 : OAI22_X1 port map( A1 => n1169, A2 => n192, B1 => n1170, B2 => n195,
                           ZN => n1168);
   U1863 : OAI222_X1 port map( A1 => n305, A2 => n96, B1 => n1171, B2 => n99, 
                           C1 => n3569, C2 => n102, ZN => n3039);
   U1864 : NOR4_X1 port map( A1 => n1172, A2 => n1173, A3 => n1174, A4 => n1175
                           , ZN => n1171);
   U1865 : OAI221_X1 port map( B1 => n3840, B2 => n105, C1 => n1176, C2 => n108
                           , A => n1177, ZN => n1175);
   U1866 : AOI22_X1 port map( A1 => n111, A2 => n3583, B1 => n114, B2 => n680, 
                           ZN => n1177);
   U1867 : OAI221_X1 port map( B1 => n1178, B2 => n117, C1 => n3744, C2 => n120
                           , A => n1179, ZN => n1174);
   U1868 : AOI22_X1 port map( A1 => n123, A2 => n782, B1 => n126, B2 => n3582, 
                           ZN => n1179);
   U1869 : OAI211_X1 port map( C1 => n3587, C2 => n129, A => n1180, B => n1181,
                           ZN => n1173);
   U1870 : AOI221_X1 port map( B1 => n132, B2 => n916, C1 => n135, C2 => n3588,
                           A => n1182, ZN => n1181);
   U1871 : OAI22_X1 port map( A1 => n3584, A2 => n138, B1 => n1183, B2 => n141,
                           ZN => n1182);
   U1872 : AOI22_X1 port map( A1 => n144, A2 => n3589, B1 => n147, B2 => n816, 
                           ZN => n1180);
   U1873 : NAND4_X1 port map( A1 => n1184, A2 => n1185, A3 => n1186, A4 => 
                           n1187, ZN => n1172);
   U1874 : AOI221_X1 port map( B1 => n150, B2 => n3572, C1 => n153, C2 => n3573
                           , A => n1188, ZN => n1187);
   U1875 : OAI22_X1 port map( A1 => n3571, A2 => n156, B1 => n3570, B2 => n159,
                           ZN => n1188);
   U1876 : AOI221_X1 port map( B1 => n162, B2 => n3576, C1 => n165, C2 => n3577
                           , A => n1189, ZN => n1186);
   U1877 : OAI22_X1 port map( A1 => n3575, A2 => n168, B1 => n3574, B2 => n171,
                           ZN => n1189);
   U1878 : AOI221_X1 port map( B1 => n174, B2 => n613, C1 => n177, C2 => n646, 
                           A => n1190, ZN => n1185);
   U1879 : OAI22_X1 port map( A1 => n1191, A2 => n180, B1 => n1192, B2 => n183,
                           ZN => n1190);
   U1880 : AOI221_X1 port map( B1 => n186, B2 => n579, C1 => n189, C2 => n3776,
                           A => n1193, ZN => n1184);
   U1881 : OAI22_X1 port map( A1 => n1194, A2 => n192, B1 => n1195, B2 => n195,
                           ZN => n1193);
   U1882 : OAI222_X1 port map( A1 => n306, A2 => n95, B1 => n1196, B2 => n98, 
                           C1 => n2972, C2 => n102, ZN => n3038);
   U1883 : NOR4_X1 port map( A1 => n1197, A2 => n1198, A3 => n1199, A4 => n1200
                           , ZN => n1196);
   U1884 : OAI221_X1 port map( B1 => n3841, B2 => n104, C1 => n1201, C2 => n107
                           , A => n1202, ZN => n1200);
   U1885 : AOI22_X1 port map( A1 => n110, A2 => n3562, B1 => n113, B2 => n681, 
                           ZN => n1202);
   U1886 : OAI221_X1 port map( B1 => n1203, B2 => n116, C1 => n3745, C2 => n119
                           , A => n1204, ZN => n1199);
   U1887 : AOI22_X1 port map( A1 => n122, A2 => n783, B1 => n125, B2 => n3561, 
                           ZN => n1204);
   U1888 : OAI211_X1 port map( C1 => n3566, C2 => n128, A => n1205, B => n1206,
                           ZN => n1198);
   U1889 : AOI221_X1 port map( B1 => n131, B2 => n917, C1 => n134, C2 => n3567,
                           A => n1207, ZN => n1206);
   U1890 : OAI22_X1 port map( A1 => n3563, A2 => n137, B1 => n1208, B2 => n140,
                           ZN => n1207);
   U1891 : AOI22_X1 port map( A1 => n143, A2 => n3568, B1 => n146, B2 => n817, 
                           ZN => n1205);
   U1892 : NAND4_X1 port map( A1 => n1209, A2 => n1210, A3 => n1211, A4 => 
                           n1212, ZN => n1197);
   U1893 : AOI221_X1 port map( B1 => n149, B2 => n2975, C1 => n152, C2 => n2976
                           , A => n1213, ZN => n1212);
   U1894 : OAI22_X1 port map( A1 => n2974, A2 => n155, B1 => n2973, B2 => n158,
                           ZN => n1213);
   U1895 : AOI221_X1 port map( B1 => n161, B2 => n2979, C1 => n164, C2 => n2980
                           , A => n1214, ZN => n1211);
   U1896 : OAI22_X1 port map( A1 => n2978, A2 => n167, B1 => n2977, B2 => n170,
                           ZN => n1214);
   U1897 : AOI221_X1 port map( B1 => n173, B2 => n614, C1 => n176, C2 => n647, 
                           A => n1215, ZN => n1210);
   U1898 : OAI22_X1 port map( A1 => n1216, A2 => n179, B1 => n1217, B2 => n182,
                           ZN => n1215);
   U1899 : AOI221_X1 port map( B1 => n185, B2 => n580, C1 => n188, C2 => n3777,
                           A => n1218, ZN => n1209);
   U1900 : OAI22_X1 port map( A1 => n1219, A2 => n191, B1 => n1220, B2 => n194,
                           ZN => n1218);
   U1901 : OAI222_X1 port map( A1 => n307, A2 => n95, B1 => n1221, B2 => n98, 
                           C1 => n2951, C2 => n102, ZN => n3037);
   U1902 : NOR4_X1 port map( A1 => n1222, A2 => n1223, A3 => n1224, A4 => n1225
                           , ZN => n1221);
   U1903 : OAI221_X1 port map( B1 => n3842, B2 => n104, C1 => n1226, C2 => n107
                           , A => n1227, ZN => n1225);
   U1904 : AOI22_X1 port map( A1 => n110, A2 => n2965, B1 => n113, B2 => n682, 
                           ZN => n1227);
   U1905 : OAI221_X1 port map( B1 => n1228, B2 => n116, C1 => n3746, C2 => n119
                           , A => n1229, ZN => n1224);
   U1906 : AOI22_X1 port map( A1 => n122, A2 => n784, B1 => n125, B2 => n2964, 
                           ZN => n1229);
   U1907 : OAI211_X1 port map( C1 => n2969, C2 => n128, A => n1230, B => n1231,
                           ZN => n1223);
   U1908 : AOI221_X1 port map( B1 => n131, B2 => n918, C1 => n134, C2 => n2970,
                           A => n1232, ZN => n1231);
   U1909 : OAI22_X1 port map( A1 => n2966, A2 => n137, B1 => n1233, B2 => n140,
                           ZN => n1232);
   U1910 : AOI22_X1 port map( A1 => n143, A2 => n2971, B1 => n146, B2 => n818, 
                           ZN => n1230);
   U1911 : NAND4_X1 port map( A1 => n1234, A2 => n1235, A3 => n1236, A4 => 
                           n1237, ZN => n1222);
   U1912 : AOI221_X1 port map( B1 => n149, B2 => n2954, C1 => n152, C2 => n2955
                           , A => n1238, ZN => n1237);
   U1913 : OAI22_X1 port map( A1 => n2953, A2 => n155, B1 => n2952, B2 => n158,
                           ZN => n1238);
   U1914 : AOI221_X1 port map( B1 => n161, B2 => n2958, C1 => n164, C2 => n2959
                           , A => n1239, ZN => n1236);
   U1915 : OAI22_X1 port map( A1 => n2957, A2 => n167, B1 => n2956, B2 => n170,
                           ZN => n1239);
   U1916 : AOI221_X1 port map( B1 => n173, B2 => n615, C1 => n176, C2 => n648, 
                           A => n1240, ZN => n1235);
   U1917 : OAI22_X1 port map( A1 => n1241, A2 => n179, B1 => n1242, B2 => n182,
                           ZN => n1240);
   U1918 : AOI221_X1 port map( B1 => n185, B2 => n581, C1 => n188, C2 => n3778,
                           A => n1243, ZN => n1234);
   U1919 : OAI22_X1 port map( A1 => n1244, A2 => n191, B1 => n1245, B2 => n194,
                           ZN => n1243);
   U1920 : OAI222_X1 port map( A1 => n308, A2 => n95, B1 => n1246, B2 => n98, 
                           C1 => n2930, C2 => n101, ZN => n3036);
   U1921 : NOR4_X1 port map( A1 => n1247, A2 => n1248, A3 => n1249, A4 => n1250
                           , ZN => n1246);
   U1922 : OAI221_X1 port map( B1 => n3843, B2 => n104, C1 => n1251, C2 => n107
                           , A => n1252, ZN => n1250);
   U1923 : AOI22_X1 port map( A1 => n110, A2 => n2944, B1 => n113, B2 => n683, 
                           ZN => n1252);
   U1924 : OAI221_X1 port map( B1 => n1253, B2 => n116, C1 => n3747, C2 => n119
                           , A => n1254, ZN => n1249);
   U1925 : AOI22_X1 port map( A1 => n122, A2 => n785, B1 => n125, B2 => n2943, 
                           ZN => n1254);
   U1926 : OAI211_X1 port map( C1 => n2948, C2 => n128, A => n1255, B => n1256,
                           ZN => n1248);
   U1927 : AOI221_X1 port map( B1 => n131, B2 => n919, C1 => n134, C2 => n2949,
                           A => n1257, ZN => n1256);
   U1928 : OAI22_X1 port map( A1 => n2945, A2 => n137, B1 => n1258, B2 => n140,
                           ZN => n1257);
   U1929 : AOI22_X1 port map( A1 => n143, A2 => n2950, B1 => n146, B2 => n819, 
                           ZN => n1255);
   U1930 : NAND4_X1 port map( A1 => n1259, A2 => n1260, A3 => n1261, A4 => 
                           n1262, ZN => n1247);
   U1931 : AOI221_X1 port map( B1 => n149, B2 => n2933, C1 => n152, C2 => n2934
                           , A => n1263, ZN => n1262);
   U1932 : OAI22_X1 port map( A1 => n2932, A2 => n155, B1 => n2931, B2 => n158,
                           ZN => n1263);
   U1933 : AOI221_X1 port map( B1 => n161, B2 => n2937, C1 => n164, C2 => n2938
                           , A => n1264, ZN => n1261);
   U1934 : OAI22_X1 port map( A1 => n2936, A2 => n167, B1 => n2935, B2 => n170,
                           ZN => n1264);
   U1935 : AOI221_X1 port map( B1 => n173, B2 => n616, C1 => n176, C2 => n649, 
                           A => n1265, ZN => n1260);
   U1936 : OAI22_X1 port map( A1 => n1266, A2 => n179, B1 => n1267, B2 => n182,
                           ZN => n1265);
   U1937 : AOI221_X1 port map( B1 => n185, B2 => n582, C1 => n188, C2 => n3779,
                           A => n1268, ZN => n1259);
   U1938 : OAI22_X1 port map( A1 => n1269, A2 => n191, B1 => n1270, B2 => n194,
                           ZN => n1268);
   U1939 : OAI222_X1 port map( A1 => n309, A2 => n95, B1 => n1271, B2 => n98, 
                           C1 => n2909, C2 => n101, ZN => n3035);
   U1940 : NOR4_X1 port map( A1 => n1272, A2 => n1273, A3 => n1274, A4 => n1275
                           , ZN => n1271);
   U1941 : OAI221_X1 port map( B1 => n3844, B2 => n104, C1 => n1276, C2 => n107
                           , A => n1277, ZN => n1275);
   U1942 : AOI22_X1 port map( A1 => n110, A2 => n2923, B1 => n113, B2 => n684, 
                           ZN => n1277);
   U1943 : OAI221_X1 port map( B1 => n1278, B2 => n116, C1 => n3748, C2 => n119
                           , A => n1279, ZN => n1274);
   U1944 : AOI22_X1 port map( A1 => n122, A2 => n786, B1 => n125, B2 => n2922, 
                           ZN => n1279);
   U1945 : OAI211_X1 port map( C1 => n2927, C2 => n128, A => n1280, B => n1281,
                           ZN => n1273);
   U1946 : AOI221_X1 port map( B1 => n131, B2 => n920, C1 => n134, C2 => n2928,
                           A => n1282, ZN => n1281);
   U1947 : OAI22_X1 port map( A1 => n2924, A2 => n137, B1 => n1283, B2 => n140,
                           ZN => n1282);
   U1948 : AOI22_X1 port map( A1 => n143, A2 => n2929, B1 => n146, B2 => n820, 
                           ZN => n1280);
   U1949 : NAND4_X1 port map( A1 => n1284, A2 => n1285, A3 => n1286, A4 => 
                           n1287, ZN => n1272);
   U1950 : AOI221_X1 port map( B1 => n149, B2 => n2912, C1 => n152, C2 => n2913
                           , A => n1288, ZN => n1287);
   U1951 : OAI22_X1 port map( A1 => n2911, A2 => n155, B1 => n2910, B2 => n158,
                           ZN => n1288);
   U1952 : AOI221_X1 port map( B1 => n161, B2 => n2916, C1 => n164, C2 => n2917
                           , A => n1289, ZN => n1286);
   U1953 : OAI22_X1 port map( A1 => n2915, A2 => n167, B1 => n2914, B2 => n170,
                           ZN => n1289);
   U1954 : AOI221_X1 port map( B1 => n173, B2 => n617, C1 => n176, C2 => n650, 
                           A => n1290, ZN => n1285);
   U1955 : OAI22_X1 port map( A1 => n1291, A2 => n179, B1 => n1292, B2 => n182,
                           ZN => n1290);
   U1956 : AOI221_X1 port map( B1 => n185, B2 => n583, C1 => n188, C2 => n3780,
                           A => n1293, ZN => n1284);
   U1957 : OAI22_X1 port map( A1 => n1294, A2 => n191, B1 => n1295, B2 => n194,
                           ZN => n1293);
   U1958 : OAI222_X1 port map( A1 => n310, A2 => n95, B1 => n1296, B2 => n98, 
                           C1 => n2888, C2 => n101, ZN => n3034);
   U1959 : NOR4_X1 port map( A1 => n1297, A2 => n1298, A3 => n1299, A4 => n1300
                           , ZN => n1296);
   U1960 : OAI221_X1 port map( B1 => n3845, B2 => n104, C1 => n1301, C2 => n107
                           , A => n1302, ZN => n1300);
   U1961 : AOI22_X1 port map( A1 => n110, A2 => n2902, B1 => n113, B2 => n685, 
                           ZN => n1302);
   U1962 : OAI221_X1 port map( B1 => n1303, B2 => n116, C1 => n3749, C2 => n119
                           , A => n1304, ZN => n1299);
   U1963 : AOI22_X1 port map( A1 => n122, A2 => n787, B1 => n125, B2 => n2901, 
                           ZN => n1304);
   U1964 : OAI211_X1 port map( C1 => n2906, C2 => n128, A => n1305, B => n1306,
                           ZN => n1298);
   U1965 : AOI221_X1 port map( B1 => n131, B2 => n921, C1 => n134, C2 => n2907,
                           A => n1307, ZN => n1306);
   U1966 : OAI22_X1 port map( A1 => n2903, A2 => n137, B1 => n1308, B2 => n140,
                           ZN => n1307);
   U1967 : AOI22_X1 port map( A1 => n143, A2 => n2908, B1 => n146, B2 => n821, 
                           ZN => n1305);
   U1968 : NAND4_X1 port map( A1 => n1309, A2 => n1310, A3 => n1311, A4 => 
                           n1312, ZN => n1297);
   U1969 : AOI221_X1 port map( B1 => n149, B2 => n2891, C1 => n152, C2 => n2892
                           , A => n1313, ZN => n1312);
   U1970 : OAI22_X1 port map( A1 => n2890, A2 => n155, B1 => n2889, B2 => n158,
                           ZN => n1313);
   U1971 : AOI221_X1 port map( B1 => n161, B2 => n2895, C1 => n164, C2 => n2896
                           , A => n1314, ZN => n1311);
   U1972 : OAI22_X1 port map( A1 => n2894, A2 => n167, B1 => n2893, B2 => n170,
                           ZN => n1314);
   U1973 : AOI221_X1 port map( B1 => n173, B2 => n618, C1 => n176, C2 => n651, 
                           A => n1315, ZN => n1310);
   U1974 : OAI22_X1 port map( A1 => n1316, A2 => n179, B1 => n1317, B2 => n182,
                           ZN => n1315);
   U1975 : AOI221_X1 port map( B1 => n185, B2 => n584, C1 => n188, C2 => n3781,
                           A => n1318, ZN => n1309);
   U1976 : OAI22_X1 port map( A1 => n1319, A2 => n191, B1 => n1320, B2 => n194,
                           ZN => n1318);
   U1977 : OAI222_X1 port map( A1 => n311, A2 => n95, B1 => n1321, B2 => n98, 
                           C1 => n2867, C2 => n101, ZN => n3033);
   U1978 : NOR4_X1 port map( A1 => n1322, A2 => n1323, A3 => n1324, A4 => n1325
                           , ZN => n1321);
   U1979 : OAI221_X1 port map( B1 => n3846, B2 => n104, C1 => n1326, C2 => n107
                           , A => n1327, ZN => n1325);
   U1980 : AOI22_X1 port map( A1 => n110, A2 => n2881, B1 => n113, B2 => n686, 
                           ZN => n1327);
   U1981 : OAI221_X1 port map( B1 => n1328, B2 => n116, C1 => n3750, C2 => n119
                           , A => n1329, ZN => n1324);
   U1982 : AOI22_X1 port map( A1 => n122, A2 => n788, B1 => n125, B2 => n2880, 
                           ZN => n1329);
   U1983 : OAI211_X1 port map( C1 => n2885, C2 => n128, A => n1330, B => n1331,
                           ZN => n1323);
   U1984 : AOI221_X1 port map( B1 => n131, B2 => n922, C1 => n134, C2 => n2886,
                           A => n1332, ZN => n1331);
   U1985 : OAI22_X1 port map( A1 => n2882, A2 => n137, B1 => n1333, B2 => n140,
                           ZN => n1332);
   U1986 : AOI22_X1 port map( A1 => n143, A2 => n2887, B1 => n146, B2 => n822, 
                           ZN => n1330);
   U1987 : NAND4_X1 port map( A1 => n1334, A2 => n1335, A3 => n1336, A4 => 
                           n1337, ZN => n1322);
   U1988 : AOI221_X1 port map( B1 => n149, B2 => n2870, C1 => n152, C2 => n2871
                           , A => n1338, ZN => n1337);
   U1989 : OAI22_X1 port map( A1 => n2869, A2 => n155, B1 => n2868, B2 => n158,
                           ZN => n1338);
   U1990 : AOI221_X1 port map( B1 => n161, B2 => n2874, C1 => n164, C2 => n2875
                           , A => n1339, ZN => n1336);
   U1991 : OAI22_X1 port map( A1 => n2873, A2 => n167, B1 => n2872, B2 => n170,
                           ZN => n1339);
   U1992 : AOI221_X1 port map( B1 => n173, B2 => n619, C1 => n176, C2 => n652, 
                           A => n1340, ZN => n1335);
   U1993 : OAI22_X1 port map( A1 => n1341, A2 => n179, B1 => n1342, B2 => n182,
                           ZN => n1340);
   U1994 : AOI221_X1 port map( B1 => n185, B2 => n585, C1 => n188, C2 => n3782,
                           A => n1343, ZN => n1334);
   U1995 : OAI22_X1 port map( A1 => n1344, A2 => n191, B1 => n1345, B2 => n194,
                           ZN => n1343);
   U1996 : OAI222_X1 port map( A1 => n312, A2 => n95, B1 => n1346, B2 => n98, 
                           C1 => n2846, C2 => n101, ZN => n3032);
   U1997 : NOR4_X1 port map( A1 => n1347, A2 => n1348, A3 => n1349, A4 => n1350
                           , ZN => n1346);
   U1998 : OAI221_X1 port map( B1 => n3847, B2 => n104, C1 => n1351, C2 => n107
                           , A => n1352, ZN => n1350);
   U1999 : AOI22_X1 port map( A1 => n110, A2 => n2860, B1 => n113, B2 => n687, 
                           ZN => n1352);
   U2000 : OAI221_X1 port map( B1 => n1353, B2 => n116, C1 => n3751, C2 => n119
                           , A => n1354, ZN => n1349);
   U2001 : AOI22_X1 port map( A1 => n122, A2 => n789, B1 => n125, B2 => n2859, 
                           ZN => n1354);
   U2002 : OAI211_X1 port map( C1 => n2864, C2 => n128, A => n1355, B => n1356,
                           ZN => n1348);
   U2003 : AOI221_X1 port map( B1 => n131, B2 => n923, C1 => n134, C2 => n2865,
                           A => n1357, ZN => n1356);
   U2004 : OAI22_X1 port map( A1 => n2861, A2 => n137, B1 => n1358, B2 => n140,
                           ZN => n1357);
   U2005 : AOI22_X1 port map( A1 => n143, A2 => n2866, B1 => n146, B2 => n823, 
                           ZN => n1355);
   U2006 : NAND4_X1 port map( A1 => n1359, A2 => n1360, A3 => n1361, A4 => 
                           n1362, ZN => n1347);
   U2007 : AOI221_X1 port map( B1 => n149, B2 => n2849, C1 => n152, C2 => n2850
                           , A => n1363, ZN => n1362);
   U2008 : OAI22_X1 port map( A1 => n2848, A2 => n155, B1 => n2847, B2 => n158,
                           ZN => n1363);
   U2009 : AOI221_X1 port map( B1 => n161, B2 => n2853, C1 => n164, C2 => n2854
                           , A => n1364, ZN => n1361);
   U2010 : OAI22_X1 port map( A1 => n2852, A2 => n167, B1 => n2851, B2 => n170,
                           ZN => n1364);
   U2011 : AOI221_X1 port map( B1 => n173, B2 => n620, C1 => n176, C2 => n653, 
                           A => n1365, ZN => n1360);
   U2012 : OAI22_X1 port map( A1 => n1366, A2 => n179, B1 => n1367, B2 => n182,
                           ZN => n1365);
   U2013 : AOI221_X1 port map( B1 => n185, B2 => n586, C1 => n188, C2 => n3783,
                           A => n1368, ZN => n1359);
   U2014 : OAI22_X1 port map( A1 => n1369, A2 => n191, B1 => n1370, B2 => n194,
                           ZN => n1368);
   U2015 : OAI222_X1 port map( A1 => n313, A2 => n95, B1 => n1371, B2 => n98, 
                           C1 => n2825, C2 => n101, ZN => n3031);
   U2016 : NOR4_X1 port map( A1 => n1372, A2 => n1373, A3 => n1374, A4 => n1375
                           , ZN => n1371);
   U2017 : OAI221_X1 port map( B1 => n3848, B2 => n104, C1 => n1376, C2 => n107
                           , A => n1377, ZN => n1375);
   U2018 : AOI22_X1 port map( A1 => n110, A2 => n2839, B1 => n113, B2 => n688, 
                           ZN => n1377);
   U2019 : OAI221_X1 port map( B1 => n1378, B2 => n116, C1 => n3752, C2 => n119
                           , A => n1379, ZN => n1374);
   U2020 : AOI22_X1 port map( A1 => n122, A2 => n790, B1 => n125, B2 => n2838, 
                           ZN => n1379);
   U2021 : OAI211_X1 port map( C1 => n2843, C2 => n128, A => n1380, B => n1381,
                           ZN => n1373);
   U2022 : AOI221_X1 port map( B1 => n131, B2 => n924, C1 => n134, C2 => n2844,
                           A => n1382, ZN => n1381);
   U2023 : OAI22_X1 port map( A1 => n2840, A2 => n137, B1 => n1383, B2 => n140,
                           ZN => n1382);
   U2024 : AOI22_X1 port map( A1 => n143, A2 => n2845, B1 => n146, B2 => n824, 
                           ZN => n1380);
   U2025 : NAND4_X1 port map( A1 => n1384, A2 => n1385, A3 => n1386, A4 => 
                           n1387, ZN => n1372);
   U2026 : AOI221_X1 port map( B1 => n149, B2 => n2828, C1 => n152, C2 => n2829
                           , A => n1388, ZN => n1387);
   U2027 : OAI22_X1 port map( A1 => n2827, A2 => n155, B1 => n2826, B2 => n158,
                           ZN => n1388);
   U2028 : AOI221_X1 port map( B1 => n161, B2 => n2832, C1 => n164, C2 => n2833
                           , A => n1389, ZN => n1386);
   U2029 : OAI22_X1 port map( A1 => n2831, A2 => n167, B1 => n2830, B2 => n170,
                           ZN => n1389);
   U2030 : AOI221_X1 port map( B1 => n173, B2 => n621, C1 => n176, C2 => n654, 
                           A => n1390, ZN => n1385);
   U2031 : OAI22_X1 port map( A1 => n1391, A2 => n179, B1 => n1392, B2 => n182,
                           ZN => n1390);
   U2032 : AOI221_X1 port map( B1 => n185, B2 => n587, C1 => n188, C2 => n3784,
                           A => n1393, ZN => n1384);
   U2033 : OAI22_X1 port map( A1 => n1394, A2 => n191, B1 => n1395, B2 => n194,
                           ZN => n1393);
   U2034 : OAI222_X1 port map( A1 => n314, A2 => n95, B1 => n1396, B2 => n98, 
                           C1 => n2804, C2 => n101, ZN => n3030);
   U2035 : NOR4_X1 port map( A1 => n1397, A2 => n1398, A3 => n1399, A4 => n1400
                           , ZN => n1396);
   U2036 : OAI221_X1 port map( B1 => n3849, B2 => n104, C1 => n1401, C2 => n107
                           , A => n1402, ZN => n1400);
   U2037 : AOI22_X1 port map( A1 => n110, A2 => n2818, B1 => n113, B2 => n689, 
                           ZN => n1402);
   U2038 : OAI221_X1 port map( B1 => n1403, B2 => n116, C1 => n3753, C2 => n119
                           , A => n1404, ZN => n1399);
   U2039 : AOI22_X1 port map( A1 => n122, A2 => n791, B1 => n125, B2 => n2817, 
                           ZN => n1404);
   U2040 : OAI211_X1 port map( C1 => n2822, C2 => n128, A => n1405, B => n1406,
                           ZN => n1398);
   U2041 : AOI221_X1 port map( B1 => n131, B2 => n925, C1 => n134, C2 => n2823,
                           A => n1407, ZN => n1406);
   U2042 : OAI22_X1 port map( A1 => n2819, A2 => n137, B1 => n1408, B2 => n140,
                           ZN => n1407);
   U2043 : AOI22_X1 port map( A1 => n143, A2 => n2824, B1 => n146, B2 => n825, 
                           ZN => n1405);
   U2044 : NAND4_X1 port map( A1 => n1409, A2 => n1410, A3 => n1411, A4 => 
                           n1412, ZN => n1397);
   U2045 : AOI221_X1 port map( B1 => n149, B2 => n2807, C1 => n152, C2 => n2808
                           , A => n1413, ZN => n1412);
   U2046 : OAI22_X1 port map( A1 => n2806, A2 => n155, B1 => n2805, B2 => n158,
                           ZN => n1413);
   U2047 : AOI221_X1 port map( B1 => n161, B2 => n2811, C1 => n164, C2 => n2812
                           , A => n1414, ZN => n1411);
   U2048 : OAI22_X1 port map( A1 => n2810, A2 => n167, B1 => n2809, B2 => n170,
                           ZN => n1414);
   U2049 : AOI221_X1 port map( B1 => n173, B2 => n622, C1 => n176, C2 => n655, 
                           A => n1415, ZN => n1410);
   U2050 : OAI22_X1 port map( A1 => n1416, A2 => n179, B1 => n1417, B2 => n182,
                           ZN => n1415);
   U2051 : AOI221_X1 port map( B1 => n185, B2 => n588, C1 => n188, C2 => n3785,
                           A => n1418, ZN => n1409);
   U2052 : OAI22_X1 port map( A1 => n1419, A2 => n191, B1 => n1420, B2 => n194,
                           ZN => n1418);
   U2053 : OAI222_X1 port map( A1 => n315, A2 => n95, B1 => n1421, B2 => n98, 
                           C1 => n2783, C2 => n101, ZN => n3029);
   U2054 : NOR4_X1 port map( A1 => n1422, A2 => n1423, A3 => n1424, A4 => n1425
                           , ZN => n1421);
   U2055 : OAI221_X1 port map( B1 => n3850, B2 => n104, C1 => n1426, C2 => n107
                           , A => n1427, ZN => n1425);
   U2056 : AOI22_X1 port map( A1 => n110, A2 => n2797, B1 => n113, B2 => n690, 
                           ZN => n1427);
   U2057 : OAI221_X1 port map( B1 => n1428, B2 => n116, C1 => n3754, C2 => n119
                           , A => n1429, ZN => n1424);
   U2058 : AOI22_X1 port map( A1 => n122, A2 => n792, B1 => n125, B2 => n2796, 
                           ZN => n1429);
   U2059 : OAI211_X1 port map( C1 => n2801, C2 => n128, A => n1430, B => n1431,
                           ZN => n1423);
   U2060 : AOI221_X1 port map( B1 => n131, B2 => n926, C1 => n134, C2 => n2802,
                           A => n1432, ZN => n1431);
   U2061 : OAI22_X1 port map( A1 => n2798, A2 => n137, B1 => n1433, B2 => n140,
                           ZN => n1432);
   U2062 : AOI22_X1 port map( A1 => n143, A2 => n2803, B1 => n146, B2 => n826, 
                           ZN => n1430);
   U2063 : NAND4_X1 port map( A1 => n1434, A2 => n1435, A3 => n1436, A4 => 
                           n1437, ZN => n1422);
   U2064 : AOI221_X1 port map( B1 => n149, B2 => n2786, C1 => n152, C2 => n2787
                           , A => n1438, ZN => n1437);
   U2065 : OAI22_X1 port map( A1 => n2785, A2 => n155, B1 => n2784, B2 => n158,
                           ZN => n1438);
   U2066 : AOI221_X1 port map( B1 => n161, B2 => n2790, C1 => n164, C2 => n2791
                           , A => n1439, ZN => n1436);
   U2067 : OAI22_X1 port map( A1 => n2789, A2 => n167, B1 => n2788, B2 => n170,
                           ZN => n1439);
   U2068 : AOI221_X1 port map( B1 => n173, B2 => n623, C1 => n176, C2 => n656, 
                           A => n1440, ZN => n1435);
   U2069 : OAI22_X1 port map( A1 => n1441, A2 => n179, B1 => n1442, B2 => n182,
                           ZN => n1440);
   U2070 : AOI221_X1 port map( B1 => n185, B2 => n589, C1 => n188, C2 => n3786,
                           A => n1443, ZN => n1434);
   U2071 : OAI22_X1 port map( A1 => n1444, A2 => n191, B1 => n1445, B2 => n194,
                           ZN => n1443);
   U2072 : OAI222_X1 port map( A1 => n316, A2 => n95, B1 => n1446, B2 => n98, 
                           C1 => n2762, C2 => n101, ZN => n3028);
   U2073 : NOR4_X1 port map( A1 => n1447, A2 => n1448, A3 => n1449, A4 => n1450
                           , ZN => n1446);
   U2074 : OAI221_X1 port map( B1 => n3851, B2 => n104, C1 => n1451, C2 => n107
                           , A => n1452, ZN => n1450);
   U2075 : AOI22_X1 port map( A1 => n110, A2 => n2776, B1 => n113, B2 => n691, 
                           ZN => n1452);
   U2076 : OAI221_X1 port map( B1 => n1453, B2 => n116, C1 => n3755, C2 => n119
                           , A => n1454, ZN => n1449);
   U2077 : AOI22_X1 port map( A1 => n122, A2 => n793, B1 => n125, B2 => n2775, 
                           ZN => n1454);
   U2078 : OAI211_X1 port map( C1 => n2780, C2 => n128, A => n1455, B => n1456,
                           ZN => n1448);
   U2079 : AOI221_X1 port map( B1 => n131, B2 => n927, C1 => n134, C2 => n2781,
                           A => n1457, ZN => n1456);
   U2080 : OAI22_X1 port map( A1 => n2777, A2 => n137, B1 => n1458, B2 => n140,
                           ZN => n1457);
   U2081 : AOI22_X1 port map( A1 => n143, A2 => n2782, B1 => n146, B2 => n827, 
                           ZN => n1455);
   U2082 : NAND4_X1 port map( A1 => n1459, A2 => n1460, A3 => n1461, A4 => 
                           n1462, ZN => n1447);
   U2083 : AOI221_X1 port map( B1 => n149, B2 => n2765, C1 => n152, C2 => n2766
                           , A => n1463, ZN => n1462);
   U2084 : OAI22_X1 port map( A1 => n2764, A2 => n155, B1 => n2763, B2 => n158,
                           ZN => n1463);
   U2085 : AOI221_X1 port map( B1 => n161, B2 => n2769, C1 => n164, C2 => n2770
                           , A => n1464, ZN => n1461);
   U2086 : OAI22_X1 port map( A1 => n2768, A2 => n167, B1 => n2767, B2 => n170,
                           ZN => n1464);
   U2087 : AOI221_X1 port map( B1 => n173, B2 => n624, C1 => n176, C2 => n657, 
                           A => n1465, ZN => n1460);
   U2088 : OAI22_X1 port map( A1 => n1466, A2 => n179, B1 => n1467, B2 => n182,
                           ZN => n1465);
   U2089 : AOI221_X1 port map( B1 => n185, B2 => n590, C1 => n188, C2 => n3787,
                           A => n1468, ZN => n1459);
   U2090 : OAI22_X1 port map( A1 => n1469, A2 => n191, B1 => n1470, B2 => n194,
                           ZN => n1468);
   U2091 : OAI222_X1 port map( A1 => n317, A2 => n95, B1 => n1471, B2 => n98, 
                           C1 => n2741, C2 => n101, ZN => n3027);
   U2092 : NOR4_X1 port map( A1 => n1472, A2 => n1473, A3 => n1474, A4 => n1475
                           , ZN => n1471);
   U2093 : OAI221_X1 port map( B1 => n3852, B2 => n104, C1 => n1476, C2 => n107
                           , A => n1477, ZN => n1475);
   U2094 : AOI22_X1 port map( A1 => n110, A2 => n2755, B1 => n113, B2 => n692, 
                           ZN => n1477);
   U2095 : OAI221_X1 port map( B1 => n1478, B2 => n116, C1 => n3756, C2 => n119
                           , A => n1479, ZN => n1474);
   U2096 : AOI22_X1 port map( A1 => n122, A2 => n794, B1 => n125, B2 => n2754, 
                           ZN => n1479);
   U2097 : OAI211_X1 port map( C1 => n2759, C2 => n128, A => n1480, B => n1481,
                           ZN => n1473);
   U2098 : AOI221_X1 port map( B1 => n131, B2 => n928, C1 => n134, C2 => n2760,
                           A => n1482, ZN => n1481);
   U2099 : OAI22_X1 port map( A1 => n2756, A2 => n137, B1 => n1483, B2 => n140,
                           ZN => n1482);
   U2100 : AOI22_X1 port map( A1 => n143, A2 => n2761, B1 => n146, B2 => n828, 
                           ZN => n1480);
   U2101 : NAND4_X1 port map( A1 => n1484, A2 => n1485, A3 => n1486, A4 => 
                           n1487, ZN => n1472);
   U2102 : AOI221_X1 port map( B1 => n149, B2 => n2744, C1 => n152, C2 => n2745
                           , A => n1488, ZN => n1487);
   U2103 : OAI22_X1 port map( A1 => n2743, A2 => n155, B1 => n2742, B2 => n158,
                           ZN => n1488);
   U2104 : AOI221_X1 port map( B1 => n161, B2 => n2748, C1 => n164, C2 => n2749
                           , A => n1489, ZN => n1486);
   U2105 : OAI22_X1 port map( A1 => n2747, A2 => n167, B1 => n2746, B2 => n170,
                           ZN => n1489);
   U2106 : AOI221_X1 port map( B1 => n173, B2 => n625, C1 => n176, C2 => n658, 
                           A => n1490, ZN => n1485);
   U2107 : OAI22_X1 port map( A1 => n1491, A2 => n179, B1 => n1492, B2 => n182,
                           ZN => n1490);
   U2108 : AOI221_X1 port map( B1 => n185, B2 => n591, C1 => n188, C2 => n3788,
                           A => n1493, ZN => n1484);
   U2109 : OAI22_X1 port map( A1 => n1494, A2 => n191, B1 => n1495, B2 => n194,
                           ZN => n1493);
   U2110 : OAI222_X1 port map( A1 => n318, A2 => n94, B1 => n1496, B2 => n97, 
                           C1 => n2720, C2 => n101, ZN => n3026);
   U2111 : NOR4_X1 port map( A1 => n1497, A2 => n1498, A3 => n1499, A4 => n1500
                           , ZN => n1496);
   U2112 : OAI221_X1 port map( B1 => n3853, B2 => n103, C1 => n1501, C2 => n106
                           , A => n1502, ZN => n1500);
   U2113 : AOI22_X1 port map( A1 => n109, A2 => n2734, B1 => n112, B2 => n693, 
                           ZN => n1502);
   U2114 : OAI221_X1 port map( B1 => n1503, B2 => n115, C1 => n3757, C2 => n118
                           , A => n1504, ZN => n1499);
   U2115 : AOI22_X1 port map( A1 => n121, A2 => n795, B1 => n124, B2 => n2733, 
                           ZN => n1504);
   U2116 : OAI211_X1 port map( C1 => n2738, C2 => n127, A => n1505, B => n1506,
                           ZN => n1498);
   U2117 : AOI221_X1 port map( B1 => n130, B2 => n929, C1 => n133, C2 => n2739,
                           A => n1507, ZN => n1506);
   U2118 : OAI22_X1 port map( A1 => n2735, A2 => n136, B1 => n1508, B2 => n139,
                           ZN => n1507);
   U2119 : AOI22_X1 port map( A1 => n142, A2 => n2740, B1 => n145, B2 => n829, 
                           ZN => n1505);
   U2120 : NAND4_X1 port map( A1 => n1509, A2 => n1510, A3 => n1511, A4 => 
                           n1512, ZN => n1497);
   U2121 : AOI221_X1 port map( B1 => n148, B2 => n2723, C1 => n151, C2 => n2724
                           , A => n1513, ZN => n1512);
   U2122 : OAI22_X1 port map( A1 => n2722, A2 => n154, B1 => n2721, B2 => n157,
                           ZN => n1513);
   U2123 : AOI221_X1 port map( B1 => n160, B2 => n2727, C1 => n163, C2 => n2728
                           , A => n1514, ZN => n1511);
   U2124 : OAI22_X1 port map( A1 => n2726, A2 => n166, B1 => n2725, B2 => n169,
                           ZN => n1514);
   U2125 : AOI221_X1 port map( B1 => n172, B2 => n626, C1 => n175, C2 => n659, 
                           A => n1515, ZN => n1510);
   U2126 : OAI22_X1 port map( A1 => n1516, A2 => n178, B1 => n1517, B2 => n181,
                           ZN => n1515);
   U2127 : AOI221_X1 port map( B1 => n184, B2 => n592, C1 => n187, C2 => n3789,
                           A => n1518, ZN => n1509);
   U2128 : OAI22_X1 port map( A1 => n1519, A2 => n190, B1 => n1520, B2 => n193,
                           ZN => n1518);
   U2129 : OAI222_X1 port map( A1 => n319, A2 => n94, B1 => n1521, B2 => n97, 
                           C1 => n2699, C2 => n101, ZN => n3025);
   U2130 : NOR4_X1 port map( A1 => n1522, A2 => n1523, A3 => n1524, A4 => n1525
                           , ZN => n1521);
   U2131 : OAI221_X1 port map( B1 => n3854, B2 => n103, C1 => n1526, C2 => n106
                           , A => n1527, ZN => n1525);
   U2132 : AOI22_X1 port map( A1 => n109, A2 => n2713, B1 => n112, B2 => n694, 
                           ZN => n1527);
   U2133 : OAI221_X1 port map( B1 => n1528, B2 => n115, C1 => n3758, C2 => n118
                           , A => n1529, ZN => n1524);
   U2134 : AOI22_X1 port map( A1 => n121, A2 => n796, B1 => n124, B2 => n2712, 
                           ZN => n1529);
   U2135 : OAI211_X1 port map( C1 => n2717, C2 => n127, A => n1530, B => n1531,
                           ZN => n1523);
   U2136 : AOI221_X1 port map( B1 => n130, B2 => n930, C1 => n133, C2 => n2718,
                           A => n1532, ZN => n1531);
   U2137 : OAI22_X1 port map( A1 => n2714, A2 => n136, B1 => n1533, B2 => n139,
                           ZN => n1532);
   U2138 : AOI22_X1 port map( A1 => n142, A2 => n2719, B1 => n145, B2 => n830, 
                           ZN => n1530);
   U2139 : NAND4_X1 port map( A1 => n1534, A2 => n1535, A3 => n1536, A4 => 
                           n1537, ZN => n1522);
   U2140 : AOI221_X1 port map( B1 => n148, B2 => n2702, C1 => n151, C2 => n2703
                           , A => n1538, ZN => n1537);
   U2141 : OAI22_X1 port map( A1 => n2701, A2 => n154, B1 => n2700, B2 => n157,
                           ZN => n1538);
   U2142 : AOI221_X1 port map( B1 => n160, B2 => n2706, C1 => n163, C2 => n2707
                           , A => n1539, ZN => n1536);
   U2143 : OAI22_X1 port map( A1 => n2705, A2 => n166, B1 => n2704, B2 => n169,
                           ZN => n1539);
   U2144 : AOI221_X1 port map( B1 => n172, B2 => n627, C1 => n175, C2 => n660, 
                           A => n1540, ZN => n1535);
   U2145 : OAI22_X1 port map( A1 => n1541, A2 => n178, B1 => n1542, B2 => n181,
                           ZN => n1540);
   U2146 : AOI221_X1 port map( B1 => n184, B2 => n593, C1 => n187, C2 => n3790,
                           A => n1543, ZN => n1534);
   U2147 : OAI22_X1 port map( A1 => n1544, A2 => n190, B1 => n1545, B2 => n193,
                           ZN => n1543);
   U2148 : OAI222_X1 port map( A1 => n320, A2 => n94, B1 => n1546, B2 => n97, 
                           C1 => n2678, C2 => n100, ZN => n3024);
   U2149 : NOR4_X1 port map( A1 => n1547, A2 => n1548, A3 => n1549, A4 => n1550
                           , ZN => n1546);
   U2150 : OAI221_X1 port map( B1 => n3855, B2 => n103, C1 => n1551, C2 => n106
                           , A => n1552, ZN => n1550);
   U2151 : AOI22_X1 port map( A1 => n109, A2 => n2692, B1 => n112, B2 => n695, 
                           ZN => n1552);
   U2152 : OAI221_X1 port map( B1 => n1553, B2 => n115, C1 => n3759, C2 => n118
                           , A => n1554, ZN => n1549);
   U2153 : AOI22_X1 port map( A1 => n121, A2 => n797, B1 => n124, B2 => n2691, 
                           ZN => n1554);
   U2154 : OAI211_X1 port map( C1 => n2696, C2 => n127, A => n1555, B => n1556,
                           ZN => n1548);
   U2155 : AOI221_X1 port map( B1 => n130, B2 => n931, C1 => n133, C2 => n2697,
                           A => n1557, ZN => n1556);
   U2156 : OAI22_X1 port map( A1 => n2693, A2 => n136, B1 => n1558, B2 => n139,
                           ZN => n1557);
   U2157 : AOI22_X1 port map( A1 => n142, A2 => n2698, B1 => n145, B2 => n831, 
                           ZN => n1555);
   U2158 : NAND4_X1 port map( A1 => n1559, A2 => n1560, A3 => n1561, A4 => 
                           n1562, ZN => n1547);
   U2159 : AOI221_X1 port map( B1 => n148, B2 => n2681, C1 => n151, C2 => n2682
                           , A => n1563, ZN => n1562);
   U2160 : OAI22_X1 port map( A1 => n2680, A2 => n154, B1 => n2679, B2 => n157,
                           ZN => n1563);
   U2161 : AOI221_X1 port map( B1 => n160, B2 => n2685, C1 => n163, C2 => n2686
                           , A => n1564, ZN => n1561);
   U2162 : OAI22_X1 port map( A1 => n2684, A2 => n166, B1 => n2683, B2 => n169,
                           ZN => n1564);
   U2163 : AOI221_X1 port map( B1 => n172, B2 => n628, C1 => n175, C2 => n661, 
                           A => n1565, ZN => n1560);
   U2164 : OAI22_X1 port map( A1 => n1566, A2 => n178, B1 => n1567, B2 => n181,
                           ZN => n1565);
   U2165 : AOI221_X1 port map( B1 => n184, B2 => n594, C1 => n187, C2 => n3791,
                           A => n1568, ZN => n1559);
   U2166 : OAI22_X1 port map( A1 => n1569, A2 => n190, B1 => n1570, B2 => n193,
                           ZN => n1568);
   U2167 : OAI222_X1 port map( A1 => n321, A2 => n94, B1 => n1571, B2 => n97, 
                           C1 => n2657, C2 => n100, ZN => n3023);
   U2168 : NOR4_X1 port map( A1 => n1572, A2 => n1573, A3 => n1574, A4 => n1575
                           , ZN => n1571);
   U2169 : OAI221_X1 port map( B1 => n3856, B2 => n103, C1 => n1576, C2 => n106
                           , A => n1577, ZN => n1575);
   U2170 : AOI22_X1 port map( A1 => n109, A2 => n2671, B1 => n112, B2 => n696, 
                           ZN => n1577);
   U2171 : OAI221_X1 port map( B1 => n1578, B2 => n115, C1 => n3760, C2 => n118
                           , A => n1579, ZN => n1574);
   U2172 : AOI22_X1 port map( A1 => n121, A2 => n798, B1 => n124, B2 => n2670, 
                           ZN => n1579);
   U2173 : OAI211_X1 port map( C1 => n2675, C2 => n127, A => n1580, B => n1581,
                           ZN => n1573);
   U2174 : AOI221_X1 port map( B1 => n130, B2 => n932, C1 => n133, C2 => n2676,
                           A => n1582, ZN => n1581);
   U2175 : OAI22_X1 port map( A1 => n2672, A2 => n136, B1 => n1583, B2 => n139,
                           ZN => n1582);
   U2176 : AOI22_X1 port map( A1 => n142, A2 => n2677, B1 => n145, B2 => n832, 
                           ZN => n1580);
   U2177 : NAND4_X1 port map( A1 => n1584, A2 => n1585, A3 => n1586, A4 => 
                           n1587, ZN => n1572);
   U2178 : AOI221_X1 port map( B1 => n148, B2 => n2660, C1 => n151, C2 => n2661
                           , A => n1588, ZN => n1587);
   U2179 : OAI22_X1 port map( A1 => n2659, A2 => n154, B1 => n2658, B2 => n157,
                           ZN => n1588);
   U2180 : AOI221_X1 port map( B1 => n160, B2 => n2664, C1 => n163, C2 => n2665
                           , A => n1589, ZN => n1586);
   U2181 : OAI22_X1 port map( A1 => n2663, A2 => n166, B1 => n2662, B2 => n169,
                           ZN => n1589);
   U2182 : AOI221_X1 port map( B1 => n172, B2 => n629, C1 => n175, C2 => n662, 
                           A => n1590, ZN => n1585);
   U2183 : OAI22_X1 port map( A1 => n1591, A2 => n178, B1 => n1592, B2 => n181,
                           ZN => n1590);
   U2184 : AOI221_X1 port map( B1 => n184, B2 => n595, C1 => n187, C2 => n3792,
                           A => n1593, ZN => n1584);
   U2185 : OAI22_X1 port map( A1 => n1594, A2 => n190, B1 => n1595, B2 => n193,
                           ZN => n1593);
   U2186 : OAI222_X1 port map( A1 => n322, A2 => n94, B1 => n1596, B2 => n97, 
                           C1 => n2636, C2 => n100, ZN => n3022);
   U2187 : NOR4_X1 port map( A1 => n1597, A2 => n1598, A3 => n1599, A4 => n1600
                           , ZN => n1596);
   U2188 : OAI221_X1 port map( B1 => n3857, B2 => n103, C1 => n1601, C2 => n106
                           , A => n1602, ZN => n1600);
   U2189 : AOI22_X1 port map( A1 => n109, A2 => n2650, B1 => n112, B2 => n697, 
                           ZN => n1602);
   U2190 : OAI221_X1 port map( B1 => n1603, B2 => n115, C1 => n3761, C2 => n118
                           , A => n1604, ZN => n1599);
   U2191 : AOI22_X1 port map( A1 => n121, A2 => n799, B1 => n124, B2 => n2649, 
                           ZN => n1604);
   U2192 : OAI211_X1 port map( C1 => n2654, C2 => n127, A => n1605, B => n1606,
                           ZN => n1598);
   U2193 : AOI221_X1 port map( B1 => n130, B2 => n933, C1 => n133, C2 => n2655,
                           A => n1607, ZN => n1606);
   U2194 : OAI22_X1 port map( A1 => n2651, A2 => n136, B1 => n1608, B2 => n139,
                           ZN => n1607);
   U2195 : AOI22_X1 port map( A1 => n142, A2 => n2656, B1 => n145, B2 => n833, 
                           ZN => n1605);
   U2196 : NAND4_X1 port map( A1 => n1609, A2 => n1610, A3 => n1611, A4 => 
                           n1612, ZN => n1597);
   U2197 : AOI221_X1 port map( B1 => n148, B2 => n2639, C1 => n151, C2 => n2640
                           , A => n1613, ZN => n1612);
   U2198 : OAI22_X1 port map( A1 => n2638, A2 => n154, B1 => n2637, B2 => n157,
                           ZN => n1613);
   U2199 : AOI221_X1 port map( B1 => n160, B2 => n2643, C1 => n163, C2 => n2644
                           , A => n1614, ZN => n1611);
   U2200 : OAI22_X1 port map( A1 => n2642, A2 => n166, B1 => n2641, B2 => n169,
                           ZN => n1614);
   U2201 : AOI221_X1 port map( B1 => n172, B2 => n630, C1 => n175, C2 => n663, 
                           A => n1615, ZN => n1610);
   U2202 : OAI22_X1 port map( A1 => n1616, A2 => n178, B1 => n1617, B2 => n181,
                           ZN => n1615);
   U2203 : AOI221_X1 port map( B1 => n184, B2 => n596, C1 => n187, C2 => n3793,
                           A => n1618, ZN => n1609);
   U2204 : OAI22_X1 port map( A1 => n1619, A2 => n190, B1 => n1620, B2 => n193,
                           ZN => n1618);
   U2205 : OAI222_X1 port map( A1 => n323, A2 => n94, B1 => n1621, B2 => n97, 
                           C1 => n2615, C2 => n100, ZN => n3021);
   U2206 : NOR4_X1 port map( A1 => n1622, A2 => n1623, A3 => n1624, A4 => n1625
                           , ZN => n1621);
   U2207 : OAI221_X1 port map( B1 => n3858, B2 => n103, C1 => n1626, C2 => n106
                           , A => n1627, ZN => n1625);
   U2208 : AOI22_X1 port map( A1 => n109, A2 => n2629, B1 => n112, B2 => n698, 
                           ZN => n1627);
   U2209 : OAI221_X1 port map( B1 => n1628, B2 => n115, C1 => n3762, C2 => n118
                           , A => n1629, ZN => n1624);
   U2210 : AOI22_X1 port map( A1 => n121, A2 => n800, B1 => n124, B2 => n2628, 
                           ZN => n1629);
   U2211 : OAI211_X1 port map( C1 => n2633, C2 => n127, A => n1630, B => n1631,
                           ZN => n1623);
   U2212 : AOI221_X1 port map( B1 => n130, B2 => n934, C1 => n133, C2 => n2634,
                           A => n1632, ZN => n1631);
   U2213 : OAI22_X1 port map( A1 => n2630, A2 => n136, B1 => n1633, B2 => n139,
                           ZN => n1632);
   U2214 : AOI22_X1 port map( A1 => n142, A2 => n2635, B1 => n145, B2 => n834, 
                           ZN => n1630);
   U2215 : NAND4_X1 port map( A1 => n1634, A2 => n1635, A3 => n1636, A4 => 
                           n1637, ZN => n1622);
   U2216 : AOI221_X1 port map( B1 => n148, B2 => n2618, C1 => n151, C2 => n2619
                           , A => n1638, ZN => n1637);
   U2217 : OAI22_X1 port map( A1 => n2617, A2 => n154, B1 => n2616, B2 => n157,
                           ZN => n1638);
   U2218 : AOI221_X1 port map( B1 => n160, B2 => n2622, C1 => n163, C2 => n2623
                           , A => n1639, ZN => n1636);
   U2219 : OAI22_X1 port map( A1 => n2621, A2 => n166, B1 => n2620, B2 => n169,
                           ZN => n1639);
   U2220 : AOI221_X1 port map( B1 => n172, B2 => n631, C1 => n175, C2 => n664, 
                           A => n1640, ZN => n1635);
   U2221 : OAI22_X1 port map( A1 => n1641, A2 => n178, B1 => n1642, B2 => n181,
                           ZN => n1640);
   U2222 : AOI221_X1 port map( B1 => n184, B2 => n597, C1 => n187, C2 => n3794,
                           A => n1643, ZN => n1634);
   U2223 : OAI22_X1 port map( A1 => n1644, A2 => n190, B1 => n1645, B2 => n193,
                           ZN => n1643);
   U2224 : OAI222_X1 port map( A1 => n324, A2 => n94, B1 => n1646, B2 => n97, 
                           C1 => n2594, C2 => n100, ZN => n3020);
   U2225 : NOR4_X1 port map( A1 => n1647, A2 => n1648, A3 => n1649, A4 => n1650
                           , ZN => n1646);
   U2226 : OAI221_X1 port map( B1 => n3859, B2 => n103, C1 => n1651, C2 => n106
                           , A => n1652, ZN => n1650);
   U2227 : AOI22_X1 port map( A1 => n109, A2 => n2608, B1 => n112, B2 => n699, 
                           ZN => n1652);
   U2228 : OAI221_X1 port map( B1 => n1653, B2 => n115, C1 => n3763, C2 => n118
                           , A => n1654, ZN => n1649);
   U2229 : AOI22_X1 port map( A1 => n121, A2 => n801, B1 => n124, B2 => n2607, 
                           ZN => n1654);
   U2230 : OAI211_X1 port map( C1 => n2612, C2 => n127, A => n1655, B => n1656,
                           ZN => n1648);
   U2231 : AOI221_X1 port map( B1 => n130, B2 => n935, C1 => n133, C2 => n2613,
                           A => n1657, ZN => n1656);
   U2232 : OAI22_X1 port map( A1 => n2609, A2 => n136, B1 => n1658, B2 => n139,
                           ZN => n1657);
   U2233 : AOI22_X1 port map( A1 => n142, A2 => n2614, B1 => n145, B2 => n835, 
                           ZN => n1655);
   U2234 : NAND4_X1 port map( A1 => n1659, A2 => n1660, A3 => n1661, A4 => 
                           n1662, ZN => n1647);
   U2235 : AOI221_X1 port map( B1 => n148, B2 => n2597, C1 => n151, C2 => n2598
                           , A => n1663, ZN => n1662);
   U2236 : OAI22_X1 port map( A1 => n2596, A2 => n154, B1 => n2595, B2 => n157,
                           ZN => n1663);
   U2237 : AOI221_X1 port map( B1 => n160, B2 => n2601, C1 => n163, C2 => n2602
                           , A => n1664, ZN => n1661);
   U2238 : OAI22_X1 port map( A1 => n2600, A2 => n166, B1 => n2599, B2 => n169,
                           ZN => n1664);
   U2239 : AOI221_X1 port map( B1 => n172, B2 => n632, C1 => n175, C2 => n665, 
                           A => n1665, ZN => n1660);
   U2240 : OAI22_X1 port map( A1 => n1666, A2 => n178, B1 => n1667, B2 => n181,
                           ZN => n1665);
   U2241 : AOI221_X1 port map( B1 => n184, B2 => n598, C1 => n187, C2 => n3795,
                           A => n1668, ZN => n1659);
   U2242 : OAI22_X1 port map( A1 => n1669, A2 => n190, B1 => n1670, B2 => n193,
                           ZN => n1668);
   U2243 : OAI222_X1 port map( A1 => n325, A2 => n94, B1 => n1671, B2 => n97, 
                           C1 => n2573, C2 => n100, ZN => n3019);
   U2244 : NOR4_X1 port map( A1 => n1672, A2 => n1673, A3 => n1674, A4 => n1675
                           , ZN => n1671);
   U2245 : OAI221_X1 port map( B1 => n3860, B2 => n103, C1 => n1676, C2 => n106
                           , A => n1677, ZN => n1675);
   U2246 : AOI22_X1 port map( A1 => n109, A2 => n2587, B1 => n112, B2 => n700, 
                           ZN => n1677);
   U2247 : OAI221_X1 port map( B1 => n1678, B2 => n115, C1 => n3764, C2 => n118
                           , A => n1679, ZN => n1674);
   U2248 : AOI22_X1 port map( A1 => n121, A2 => n802, B1 => n124, B2 => n2586, 
                           ZN => n1679);
   U2249 : OAI211_X1 port map( C1 => n2591, C2 => n127, A => n1680, B => n1681,
                           ZN => n1673);
   U2250 : AOI221_X1 port map( B1 => n130, B2 => n936, C1 => n133, C2 => n2592,
                           A => n1682, ZN => n1681);
   U2251 : OAI22_X1 port map( A1 => n2588, A2 => n136, B1 => n1683, B2 => n139,
                           ZN => n1682);
   U2252 : AOI22_X1 port map( A1 => n142, A2 => n2593, B1 => n145, B2 => n836, 
                           ZN => n1680);
   U2253 : NAND4_X1 port map( A1 => n1684, A2 => n1685, A3 => n1686, A4 => 
                           n1687, ZN => n1672);
   U2254 : AOI221_X1 port map( B1 => n148, B2 => n2576, C1 => n151, C2 => n2577
                           , A => n1688, ZN => n1687);
   U2255 : OAI22_X1 port map( A1 => n2575, A2 => n154, B1 => n2574, B2 => n157,
                           ZN => n1688);
   U2256 : AOI221_X1 port map( B1 => n160, B2 => n2580, C1 => n163, C2 => n2581
                           , A => n1689, ZN => n1686);
   U2257 : OAI22_X1 port map( A1 => n2579, A2 => n166, B1 => n2578, B2 => n169,
                           ZN => n1689);
   U2258 : AOI221_X1 port map( B1 => n172, B2 => n633, C1 => n175, C2 => n666, 
                           A => n1690, ZN => n1685);
   U2259 : OAI22_X1 port map( A1 => n1691, A2 => n178, B1 => n1692, B2 => n181,
                           ZN => n1690);
   U2260 : AOI221_X1 port map( B1 => n184, B2 => n599, C1 => n187, C2 => n3796,
                           A => n1693, ZN => n1684);
   U2261 : OAI22_X1 port map( A1 => n1694, A2 => n190, B1 => n1695, B2 => n193,
                           ZN => n1693);
   U2262 : OAI222_X1 port map( A1 => n326, A2 => n94, B1 => n1696, B2 => n97, 
                           C1 => n2552, C2 => n100, ZN => n3018);
   U2263 : NOR4_X1 port map( A1 => n1697, A2 => n1698, A3 => n1699, A4 => n1700
                           , ZN => n1696);
   U2264 : OAI221_X1 port map( B1 => n3861, B2 => n103, C1 => n1701, C2 => n106
                           , A => n1702, ZN => n1700);
   U2265 : AOI22_X1 port map( A1 => n109, A2 => n2566, B1 => n112, B2 => n701, 
                           ZN => n1702);
   U2266 : OAI221_X1 port map( B1 => n1703, B2 => n115, C1 => n3765, C2 => n118
                           , A => n1704, ZN => n1699);
   U2267 : AOI22_X1 port map( A1 => n121, A2 => n803, B1 => n124, B2 => n2565, 
                           ZN => n1704);
   U2268 : OAI211_X1 port map( C1 => n2570, C2 => n127, A => n1705, B => n1706,
                           ZN => n1698);
   U2269 : AOI221_X1 port map( B1 => n130, B2 => n937, C1 => n133, C2 => n2571,
                           A => n1707, ZN => n1706);
   U2270 : OAI22_X1 port map( A1 => n2567, A2 => n136, B1 => n1708, B2 => n139,
                           ZN => n1707);
   U2271 : AOI22_X1 port map( A1 => n142, A2 => n2572, B1 => n145, B2 => n837, 
                           ZN => n1705);
   U2272 : NAND4_X1 port map( A1 => n1709, A2 => n1710, A3 => n1711, A4 => 
                           n1712, ZN => n1697);
   U2273 : AOI221_X1 port map( B1 => n148, B2 => n2555, C1 => n151, C2 => n2556
                           , A => n1713, ZN => n1712);
   U2274 : OAI22_X1 port map( A1 => n2554, A2 => n154, B1 => n2553, B2 => n157,
                           ZN => n1713);
   U2275 : AOI221_X1 port map( B1 => n160, B2 => n2559, C1 => n163, C2 => n2560
                           , A => n1714, ZN => n1711);
   U2276 : OAI22_X1 port map( A1 => n2558, A2 => n166, B1 => n2557, B2 => n169,
                           ZN => n1714);
   U2277 : AOI221_X1 port map( B1 => n172, B2 => n634, C1 => n175, C2 => n667, 
                           A => n1715, ZN => n1710);
   U2278 : OAI22_X1 port map( A1 => n1716, A2 => n178, B1 => n1717, B2 => n181,
                           ZN => n1715);
   U2279 : AOI221_X1 port map( B1 => n184, B2 => n600, C1 => n187, C2 => n3797,
                           A => n1718, ZN => n1709);
   U2280 : OAI22_X1 port map( A1 => n1719, A2 => n190, B1 => n1720, B2 => n193,
                           ZN => n1718);
   U2281 : OAI222_X1 port map( A1 => n327, A2 => n94, B1 => n1721, B2 => n97, 
                           C1 => n2531, C2 => n100, ZN => n3017);
   U2282 : NOR4_X1 port map( A1 => n1722, A2 => n1723, A3 => n1724, A4 => n1725
                           , ZN => n1721);
   U2283 : OAI221_X1 port map( B1 => n3862, B2 => n103, C1 => n1726, C2 => n106
                           , A => n1727, ZN => n1725);
   U2284 : AOI22_X1 port map( A1 => n109, A2 => n2545, B1 => n112, B2 => n702, 
                           ZN => n1727);
   U2285 : OAI221_X1 port map( B1 => n1728, B2 => n115, C1 => n3766, C2 => n118
                           , A => n1729, ZN => n1724);
   U2286 : AOI22_X1 port map( A1 => n121, A2 => n804, B1 => n124, B2 => n2544, 
                           ZN => n1729);
   U2287 : OAI211_X1 port map( C1 => n2549, C2 => n127, A => n1730, B => n1731,
                           ZN => n1723);
   U2288 : AOI221_X1 port map( B1 => n130, B2 => n938, C1 => n133, C2 => n2550,
                           A => n1732, ZN => n1731);
   U2289 : OAI22_X1 port map( A1 => n2546, A2 => n136, B1 => n1733, B2 => n139,
                           ZN => n1732);
   U2290 : AOI22_X1 port map( A1 => n142, A2 => n2551, B1 => n145, B2 => n838, 
                           ZN => n1730);
   U2291 : NAND4_X1 port map( A1 => n1734, A2 => n1735, A3 => n1736, A4 => 
                           n1737, ZN => n1722);
   U2292 : AOI221_X1 port map( B1 => n148, B2 => n2534, C1 => n151, C2 => n2535
                           , A => n1738, ZN => n1737);
   U2293 : OAI22_X1 port map( A1 => n2533, A2 => n154, B1 => n2532, B2 => n157,
                           ZN => n1738);
   U2294 : AOI221_X1 port map( B1 => n160, B2 => n2538, C1 => n163, C2 => n2539
                           , A => n1739, ZN => n1736);
   U2295 : OAI22_X1 port map( A1 => n2537, A2 => n166, B1 => n2536, B2 => n169,
                           ZN => n1739);
   U2296 : AOI221_X1 port map( B1 => n172, B2 => n635, C1 => n175, C2 => n668, 
                           A => n1740, ZN => n1735);
   U2297 : OAI22_X1 port map( A1 => n1741, A2 => n178, B1 => n1742, B2 => n181,
                           ZN => n1740);
   U2298 : AOI221_X1 port map( B1 => n184, B2 => n601, C1 => n187, C2 => n3798,
                           A => n1743, ZN => n1734);
   U2299 : OAI22_X1 port map( A1 => n1744, A2 => n190, B1 => n1745, B2 => n193,
                           ZN => n1743);
   U2300 : OAI222_X1 port map( A1 => n328, A2 => n94, B1 => n1746, B2 => n97, 
                           C1 => n2510, C2 => n100, ZN => n3016);
   U2301 : NOR4_X1 port map( A1 => n1747, A2 => n1748, A3 => n1749, A4 => n1750
                           , ZN => n1746);
   U2302 : OAI221_X1 port map( B1 => n3863, B2 => n103, C1 => n1751, C2 => n106
                           , A => n1752, ZN => n1750);
   U2303 : AOI22_X1 port map( A1 => n109, A2 => n2524, B1 => n112, B2 => n703, 
                           ZN => n1752);
   U2304 : OAI221_X1 port map( B1 => n1753, B2 => n115, C1 => n3767, C2 => n118
                           , A => n1754, ZN => n1749);
   U2305 : AOI22_X1 port map( A1 => n121, A2 => n805, B1 => n124, B2 => n2523, 
                           ZN => n1754);
   U2306 : OAI211_X1 port map( C1 => n2528, C2 => n127, A => n1755, B => n1756,
                           ZN => n1748);
   U2307 : AOI221_X1 port map( B1 => n130, B2 => n939, C1 => n133, C2 => n2529,
                           A => n1757, ZN => n1756);
   U2308 : OAI22_X1 port map( A1 => n2525, A2 => n136, B1 => n1758, B2 => n139,
                           ZN => n1757);
   U2309 : AOI22_X1 port map( A1 => n142, A2 => n2530, B1 => n145, B2 => n839, 
                           ZN => n1755);
   U2310 : NAND4_X1 port map( A1 => n1759, A2 => n1760, A3 => n1761, A4 => 
                           n1762, ZN => n1747);
   U2311 : AOI221_X1 port map( B1 => n148, B2 => n2513, C1 => n151, C2 => n2514
                           , A => n1763, ZN => n1762);
   U2312 : OAI22_X1 port map( A1 => n2512, A2 => n154, B1 => n2511, B2 => n157,
                           ZN => n1763);
   U2313 : AOI221_X1 port map( B1 => n160, B2 => n2517, C1 => n163, C2 => n2518
                           , A => n1764, ZN => n1761);
   U2314 : OAI22_X1 port map( A1 => n2516, A2 => n166, B1 => n2515, B2 => n169,
                           ZN => n1764);
   U2315 : AOI221_X1 port map( B1 => n172, B2 => n636, C1 => n175, C2 => n669, 
                           A => n1765, ZN => n1760);
   U2316 : OAI22_X1 port map( A1 => n1766, A2 => n178, B1 => n1767, B2 => n181,
                           ZN => n1765);
   U2317 : AOI221_X1 port map( B1 => n184, B2 => n602, C1 => n187, C2 => n3799,
                           A => n1768, ZN => n1759);
   U2318 : OAI22_X1 port map( A1 => n1769, A2 => n190, B1 => n1770, B2 => n193,
                           ZN => n1768);
   U2319 : OAI222_X1 port map( A1 => n329, A2 => n94, B1 => n1771, B2 => n97, 
                           C1 => n2489, C2 => n100, ZN => n3015);
   U2320 : NAND2_X1 port map( A1 => n100, A2 => n1772, ZN => n964);
   U2321 : NOR4_X1 port map( A1 => n1773, A2 => n1774, A3 => n1775, A4 => n1776
                           , ZN => n1771);
   U2322 : OAI221_X1 port map( B1 => n3864, B2 => n103, C1 => n1777, C2 => n106
                           , A => n1778, ZN => n1776);
   U2323 : AOI22_X1 port map( A1 => n109, A2 => n2503, B1 => n112, B2 => n671, 
                           ZN => n1778);
   U2324 : AND2_X1 port map( A1 => n1779, A2 => n1780, ZN => n975);
   U2325 : AND2_X1 port map( A1 => n1779, A2 => n1781, ZN => n974);
   U2326 : NAND2_X1 port map( A1 => n1782, A2 => n1783, ZN => n972);
   U2327 : NAND2_X1 port map( A1 => n1784, A2 => n1780, ZN => n970);
   U2328 : OAI221_X1 port map( B1 => n1785, B2 => n115, C1 => n3768, C2 => n118
                           , A => n1786, ZN => n1775);
   U2329 : AOI22_X1 port map( A1 => n121, A2 => n806, B1 => n124, B2 => n2502, 
                           ZN => n1786);
   U2330 : AND2_X1 port map( A1 => n1784, A2 => n1781, ZN => n981);
   U2331 : AND2_X1 port map( A1 => n1784, A2 => n1783, ZN => n980);
   U2332 : NAND2_X1 port map( A1 => n1779, A2 => n1783, ZN => n978);
   U2333 : NAND2_X1 port map( A1 => n1779, A2 => n1787, ZN => n977);
   U2334 : NOR3_X1 port map( A1 => n1788, A2 => ADD_RS2(0), A3 => n1789, ZN => 
                           n1779);
   U2335 : OAI211_X1 port map( C1 => n2507, C2 => n127, A => n1790, B => n1791,
                           ZN => n1774);
   U2336 : AOI221_X1 port map( B1 => n130, B2 => n940, C1 => n133, C2 => n2508,
                           A => n1792, ZN => n1791);
   U2337 : OAI22_X1 port map( A1 => n2504, A2 => n136, B1 => n1793, B2 => n139,
                           ZN => n1792);
   U2338 : NAND2_X1 port map( A1 => n1794, A2 => n1783, ZN => n990);
   U2339 : NAND2_X1 port map( A1 => n1794, A2 => n1787, ZN => n988);
   U2340 : AND2_X1 port map( A1 => n1782, A2 => n1780, ZN => n986);
   U2341 : AND2_X1 port map( A1 => n1782, A2 => n1787, ZN => n985);
   U2342 : AOI22_X1 port map( A1 => n142, A2 => n2509, B1 => n145, B2 => n840, 
                           ZN => n1790);
   U2343 : AND2_X1 port map( A1 => n1794, A2 => n1781, ZN => n992);
   U2344 : AND2_X1 port map( A1 => n1794, A2 => n1780, ZN => n991);
   U2345 : NOR3_X1 port map( A1 => ADD_RS2(0), A2 => ADD_RS2(3), A3 => n1788, 
                           ZN => n1794);
   U2346 : NAND2_X1 port map( A1 => n1782, A2 => n1781, ZN => n982);
   U2347 : NOR3_X1 port map( A1 => n1795, A2 => ADD_RS2(3), A3 => n1788, ZN => 
                           n1782);
   U2348 : NAND4_X1 port map( A1 => n1796, A2 => n1797, A3 => n1798, A4 => 
                           n1799, ZN => n1773);
   U2349 : AOI221_X1 port map( B1 => n148, B2 => n2492, C1 => n151, C2 => n2493
                           , A => n1800, ZN => n1799);
   U2350 : OAI22_X1 port map( A1 => n2491, A2 => n154, B1 => n2490, B2 => n157,
                           ZN => n1800);
   U2351 : NAND2_X1 port map( A1 => n1787, A2 => n1801, ZN => n1001);
   U2352 : NAND2_X1 port map( A1 => n1787, A2 => n1802, ZN => n1000);
   U2353 : AND2_X1 port map( A1 => n1801, A2 => n1783, ZN => n998);
   U2354 : AND2_X1 port map( A1 => n1783, A2 => n1802, ZN => n997);
   U2355 : AOI221_X1 port map( B1 => n160, B2 => n2496, C1 => n163, C2 => n2497
                           , A => n1803, ZN => n1798);
   U2356 : OAI22_X1 port map( A1 => n2495, A2 => n166, B1 => n2494, B2 => n169,
                           ZN => n1803);
   U2357 : NAND2_X1 port map( A1 => n1781, A2 => n1801, ZN => n1006);
   U2358 : NAND2_X1 port map( A1 => n1781, A2 => n1802, ZN => n1005);
   U2359 : AND2_X1 port map( A1 => n1780, A2 => n1801, ZN => n1003);
   U2360 : NOR3_X1 port map( A1 => ADD_RS2(0), A2 => ADD_RS2(4), A3 => n1789, 
                           ZN => n1801);
   U2361 : AND2_X1 port map( A1 => n1780, A2 => n1802, ZN => n1002);
   U2362 : NOR3_X1 port map( A1 => n1795, A2 => ADD_RS2(4), A3 => n1789, ZN => 
                           n1802);
   U2363 : AOI221_X1 port map( B1 => n172, B2 => n637, C1 => n175, C2 => n670, 
                           A => n1804, ZN => n1797);
   U2364 : OAI22_X1 port map( A1 => n1805, A2 => n178, B1 => n1806, B2 => n181,
                           ZN => n1804);
   U2365 : NAND2_X1 port map( A1 => n1807, A2 => n1783, ZN => n1013);
   U2366 : NAND2_X1 port map( A1 => n1808, A2 => n1783, ZN => n1011);
   U2367 : NOR2_X1 port map( A1 => n1809, A2 => n1810, ZN => n1783);
   U2368 : AND2_X1 port map( A1 => n1807, A2 => n1787, ZN => n1008);
   U2369 : AND2_X1 port map( A1 => n1808, A2 => n1787, ZN => n1007);
   U2370 : AOI221_X1 port map( B1 => n184, B2 => n603, C1 => n187, C2 => n3800,
                           A => n1811, ZN => n1796);
   U2371 : OAI22_X1 port map( A1 => n1812, A2 => n190, B1 => n1813, B2 => n193,
                           ZN => n1811);
   U2372 : NAND2_X1 port map( A1 => n1807, A2 => n1780, ZN => n1020);
   U2373 : NAND2_X1 port map( A1 => n1808, A2 => n1780, ZN => n1018);
   U2374 : NOR2_X1 port map( A1 => n1810, A2 => ADD_RS2(2), ZN => n1780);
   U2375 : NOR3_X1 port map( A1 => ADD_RS2(3), A2 => ADD_RS2(4), A3 => 
                           ADD_RS2(0), ZN => n1808);
   U2376 : AND2_X1 port map( A1 => n1784, A2 => n1787, ZN => n1015);
   U2377 : NOR2_X1 port map( A1 => n1809, A2 => ADD_RS2(1), ZN => n1787);
   U2378 : INV_X1 port map( A => ADD_RS2(2), ZN => n1809);
   U2379 : NOR3_X1 port map( A1 => n1788, A2 => n1795, A3 => n1789, ZN => n1784
                           );
   U2380 : INV_X1 port map( A => ADD_RS2(3), ZN => n1789);
   U2381 : INV_X1 port map( A => ADD_RS2(4), ZN => n1788);
   U2382 : AND2_X1 port map( A1 => n1807, A2 => n1781, ZN => n1014);
   U2383 : NOR2_X1 port map( A1 => ADD_RS2(1), A2 => ADD_RS2(2), ZN => n1781);
   U2384 : NOR3_X1 port map( A1 => ADD_RS2(3), A2 => ADD_RS2(4), A3 => n1795, 
                           ZN => n1807);
   U2385 : INV_X1 port map( A => ADD_RS2(0), ZN => n1795);
   U2386 : NAND2_X1 port map( A1 => n1814, A2 => n100, ZN => n962);
   U2387 : AND3_X1 port map( A1 => RD2, A2 => ENABLE, A3 => n419, ZN => n965);
   U2388 : INV_X1 port map( A => n1772, ZN => n1814);
   U2389 : NAND4_X1 port map( A1 => n1815, A2 => n1816, A3 => n1817, A4 => 
                           n1818, ZN => n1772);
   U2390 : NOR3_X1 port map( A1 => n1819, A2 => n1820, A3 => n1821, ZN => n1818
                           );
   U2391 : XNOR2_X1 port map( A => ADD_WR(1), B => n1810, ZN => n1821);
   U2392 : INV_X1 port map( A => ADD_RS2(1), ZN => n1810);
   U2393 : XNOR2_X1 port map( A => n953, B => ADD_RS2(0), ZN => n1819);
   U2394 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS2(3), ZN => n1817);
   U2395 : XNOR2_X1 port map( A => ADD_WR(4), B => ADD_RS2(4), ZN => n1816);
   U2396 : XNOR2_X1 port map( A => ADD_RS2(2), B => ADD_WR(2), ZN => n1815);
   U2397 : OAI222_X1 port map( A1 => n329, A2 => n198, B1 => n1823, B2 => n201,
                           C1 => n2488, C2 => n204, ZN => n3014);
   U2398 : NOR4_X1 port map( A1 => n1826, A2 => n1827, A3 => n1828, A4 => n1829
                           , ZN => n1823);
   U2399 : OAI221_X1 port map( B1 => n3864, B2 => n207, C1 => n1777, C2 => n210
                           , A => n1832, ZN => n1829);
   U2400 : AOI22_X1 port map( A1 => n213, A2 => n2503, B1 => n216, B2 => n671, 
                           ZN => n1832);
   U2401 : OAI221_X1 port map( B1 => n1785, B2 => n219, C1 => n3768, C2 => n222
                           , A => n1837, ZN => n1828);
   U2402 : AOI22_X1 port map( A1 => n225, A2 => n806, B1 => n228, B2 => n2502, 
                           ZN => n1837);
   U2403 : OAI211_X1 port map( C1 => n2507, C2 => n231, A => n1841, B => n1842,
                           ZN => n1827);
   U2404 : AOI221_X1 port map( B1 => n234, B2 => n940, C1 => n237, C2 => n2508,
                           A => n1845, ZN => n1842);
   U2405 : OAI22_X1 port map( A1 => n2504, A2 => n240, B1 => n1793, B2 => n243,
                           ZN => n1845);
   U2406 : AOI22_X1 port map( A1 => n246, A2 => n2509, B1 => n249, B2 => n840, 
                           ZN => n1841);
   U2407 : NAND4_X1 port map( A1 => n1850, A2 => n1851, A3 => n1852, A4 => 
                           n1853, ZN => n1826);
   U2408 : AOI221_X1 port map( B1 => n252, B2 => n2492, C1 => n255, C2 => n2493
                           , A => n1856, ZN => n1853);
   U2409 : OAI22_X1 port map( A1 => n2491, A2 => n258, B1 => n2490, B2 => n261,
                           ZN => n1856);
   U2410 : AOI221_X1 port map( B1 => n264, B2 => n2496, C1 => n267, C2 => n2497
                           , A => n1861, ZN => n1852);
   U2411 : OAI22_X1 port map( A1 => n2495, A2 => n270, B1 => n2494, B2 => n273,
                           ZN => n1861);
   U2412 : AOI221_X1 port map( B1 => n276, B2 => n637, C1 => n279, C2 => n670, 
                           A => n1866, ZN => n1851);
   U2413 : OAI22_X1 port map( A1 => n1805, A2 => n282, B1 => n1806, B2 => n285,
                           ZN => n1866);
   U2414 : AOI221_X1 port map( B1 => n288, B2 => n603, C1 => n291, C2 => n3800,
                           A => n1871, ZN => n1850);
   U2415 : OAI22_X1 port map( A1 => n1812, A2 => n294, B1 => n1813, B2 => n297,
                           ZN => n1871);
   U2416 : OAI222_X1 port map( A1 => n328, A2 => n198, B1 => n1874, B2 => n201,
                           C1 => n2487, C2 => n204, ZN => n3013);
   U2417 : NOR4_X1 port map( A1 => n1875, A2 => n1876, A3 => n1877, A4 => n1878
                           , ZN => n1874);
   U2418 : OAI221_X1 port map( B1 => n3863, B2 => n207, C1 => n1751, C2 => n210
                           , A => n1879, ZN => n1878);
   U2419 : AOI22_X1 port map( A1 => n213, A2 => n2524, B1 => n216, B2 => n703, 
                           ZN => n1879);
   U2420 : OAI221_X1 port map( B1 => n1753, B2 => n219, C1 => n3767, C2 => n222
                           , A => n1880, ZN => n1877);
   U2421 : AOI22_X1 port map( A1 => n225, A2 => n805, B1 => n228, B2 => n2523, 
                           ZN => n1880);
   U2422 : OAI211_X1 port map( C1 => n2528, C2 => n231, A => n1881, B => n1882,
                           ZN => n1876);
   U2423 : AOI221_X1 port map( B1 => n234, B2 => n939, C1 => n237, C2 => n2529,
                           A => n1883, ZN => n1882);
   U2424 : OAI22_X1 port map( A1 => n2525, A2 => n240, B1 => n1758, B2 => n243,
                           ZN => n1883);
   U2425 : AOI22_X1 port map( A1 => n246, A2 => n2530, B1 => n249, B2 => n839, 
                           ZN => n1881);
   U2426 : NAND4_X1 port map( A1 => n1884, A2 => n1885, A3 => n1886, A4 => 
                           n1887, ZN => n1875);
   U2427 : AOI221_X1 port map( B1 => n252, B2 => n2513, C1 => n255, C2 => n2514
                           , A => n1888, ZN => n1887);
   U2428 : OAI22_X1 port map( A1 => n2512, A2 => n258, B1 => n2511, B2 => n261,
                           ZN => n1888);
   U2429 : AOI221_X1 port map( B1 => n264, B2 => n2517, C1 => n267, C2 => n2518
                           , A => n1889, ZN => n1886);
   U2430 : OAI22_X1 port map( A1 => n2516, A2 => n270, B1 => n2515, B2 => n273,
                           ZN => n1889);
   U2431 : AOI221_X1 port map( B1 => n276, B2 => n636, C1 => n279, C2 => n669, 
                           A => n1890, ZN => n1885);
   U2432 : OAI22_X1 port map( A1 => n1766, A2 => n282, B1 => n1767, B2 => n285,
                           ZN => n1890);
   U2433 : AOI221_X1 port map( B1 => n288, B2 => n602, C1 => n291, C2 => n3799,
                           A => n1891, ZN => n1884);
   U2434 : OAI22_X1 port map( A1 => n1769, A2 => n294, B1 => n1770, B2 => n297,
                           ZN => n1891);
   U2435 : OAI222_X1 port map( A1 => n327, A2 => n198, B1 => n1892, B2 => n201,
                           C1 => n2486, C2 => n204, ZN => n3012);
   U2436 : NOR4_X1 port map( A1 => n1893, A2 => n1894, A3 => n1895, A4 => n1896
                           , ZN => n1892);
   U2437 : OAI221_X1 port map( B1 => n3862, B2 => n207, C1 => n1726, C2 => n210
                           , A => n1897, ZN => n1896);
   U2438 : AOI22_X1 port map( A1 => n213, A2 => n2545, B1 => n216, B2 => n702, 
                           ZN => n1897);
   U2439 : OAI221_X1 port map( B1 => n1728, B2 => n219, C1 => n3766, C2 => n222
                           , A => n1898, ZN => n1895);
   U2440 : AOI22_X1 port map( A1 => n225, A2 => n804, B1 => n228, B2 => n2544, 
                           ZN => n1898);
   U2441 : OAI211_X1 port map( C1 => n2549, C2 => n231, A => n1899, B => n1900,
                           ZN => n1894);
   U2442 : AOI221_X1 port map( B1 => n234, B2 => n938, C1 => n237, C2 => n2550,
                           A => n1901, ZN => n1900);
   U2443 : OAI22_X1 port map( A1 => n2546, A2 => n240, B1 => n1733, B2 => n243,
                           ZN => n1901);
   U2444 : AOI22_X1 port map( A1 => n246, A2 => n2551, B1 => n249, B2 => n838, 
                           ZN => n1899);
   U2445 : NAND4_X1 port map( A1 => n1902, A2 => n1903, A3 => n1904, A4 => 
                           n1905, ZN => n1893);
   U2446 : AOI221_X1 port map( B1 => n252, B2 => n2534, C1 => n255, C2 => n2535
                           , A => n1906, ZN => n1905);
   U2447 : OAI22_X1 port map( A1 => n2533, A2 => n258, B1 => n2532, B2 => n261,
                           ZN => n1906);
   U2448 : AOI221_X1 port map( B1 => n264, B2 => n2538, C1 => n267, C2 => n2539
                           , A => n1907, ZN => n1904);
   U2449 : OAI22_X1 port map( A1 => n2537, A2 => n270, B1 => n2536, B2 => n273,
                           ZN => n1907);
   U2450 : AOI221_X1 port map( B1 => n276, B2 => n635, C1 => n279, C2 => n668, 
                           A => n1908, ZN => n1903);
   U2451 : OAI22_X1 port map( A1 => n1741, A2 => n282, B1 => n1742, B2 => n285,
                           ZN => n1908);
   U2452 : AOI221_X1 port map( B1 => n288, B2 => n601, C1 => n291, C2 => n3798,
                           A => n1909, ZN => n1902);
   U2453 : OAI22_X1 port map( A1 => n1744, A2 => n294, B1 => n1745, B2 => n297,
                           ZN => n1909);
   U2454 : OAI222_X1 port map( A1 => n326, A2 => n198, B1 => n1910, B2 => n201,
                           C1 => n2485, C2 => n204, ZN => n3011);
   U2455 : NOR4_X1 port map( A1 => n1911, A2 => n1912, A3 => n1913, A4 => n1914
                           , ZN => n1910);
   U2456 : OAI221_X1 port map( B1 => n3861, B2 => n207, C1 => n1701, C2 => n210
                           , A => n1915, ZN => n1914);
   U2457 : AOI22_X1 port map( A1 => n213, A2 => n2566, B1 => n216, B2 => n701, 
                           ZN => n1915);
   U2458 : OAI221_X1 port map( B1 => n1703, B2 => n219, C1 => n3765, C2 => n222
                           , A => n1916, ZN => n1913);
   U2459 : AOI22_X1 port map( A1 => n225, A2 => n803, B1 => n228, B2 => n2565, 
                           ZN => n1916);
   U2460 : OAI211_X1 port map( C1 => n2570, C2 => n231, A => n1917, B => n1918,
                           ZN => n1912);
   U2461 : AOI221_X1 port map( B1 => n234, B2 => n937, C1 => n237, C2 => n2571,
                           A => n1919, ZN => n1918);
   U2462 : OAI22_X1 port map( A1 => n2567, A2 => n240, B1 => n1708, B2 => n243,
                           ZN => n1919);
   U2463 : AOI22_X1 port map( A1 => n246, A2 => n2572, B1 => n249, B2 => n837, 
                           ZN => n1917);
   U2464 : NAND4_X1 port map( A1 => n1920, A2 => n1921, A3 => n1922, A4 => 
                           n1923, ZN => n1911);
   U2465 : AOI221_X1 port map( B1 => n252, B2 => n2555, C1 => n255, C2 => n2556
                           , A => n1924, ZN => n1923);
   U2466 : OAI22_X1 port map( A1 => n2554, A2 => n258, B1 => n2553, B2 => n261,
                           ZN => n1924);
   U2467 : AOI221_X1 port map( B1 => n264, B2 => n2559, C1 => n267, C2 => n2560
                           , A => n1925, ZN => n1922);
   U2468 : OAI22_X1 port map( A1 => n2558, A2 => n270, B1 => n2557, B2 => n273,
                           ZN => n1925);
   U2469 : AOI221_X1 port map( B1 => n276, B2 => n634, C1 => n279, C2 => n667, 
                           A => n1926, ZN => n1921);
   U2470 : OAI22_X1 port map( A1 => n1716, A2 => n282, B1 => n1717, B2 => n285,
                           ZN => n1926);
   U2471 : AOI221_X1 port map( B1 => n288, B2 => n600, C1 => n291, C2 => n3797,
                           A => n1927, ZN => n1920);
   U2472 : OAI22_X1 port map( A1 => n1719, A2 => n294, B1 => n1720, B2 => n297,
                           ZN => n1927);
   U2473 : OAI222_X1 port map( A1 => n325, A2 => n198, B1 => n1928, B2 => n201,
                           C1 => n2484, C2 => n204, ZN => n3010);
   U2474 : NOR4_X1 port map( A1 => n1929, A2 => n1930, A3 => n1931, A4 => n1932
                           , ZN => n1928);
   U2475 : OAI221_X1 port map( B1 => n3860, B2 => n207, C1 => n1676, C2 => n210
                           , A => n1933, ZN => n1932);
   U2476 : AOI22_X1 port map( A1 => n213, A2 => n2587, B1 => n216, B2 => n700, 
                           ZN => n1933);
   U2477 : OAI221_X1 port map( B1 => n1678, B2 => n219, C1 => n3764, C2 => n222
                           , A => n1934, ZN => n1931);
   U2478 : AOI22_X1 port map( A1 => n225, A2 => n802, B1 => n228, B2 => n2586, 
                           ZN => n1934);
   U2479 : OAI211_X1 port map( C1 => n2591, C2 => n231, A => n1935, B => n1936,
                           ZN => n1930);
   U2480 : AOI221_X1 port map( B1 => n234, B2 => n936, C1 => n237, C2 => n2592,
                           A => n1937, ZN => n1936);
   U2481 : OAI22_X1 port map( A1 => n2588, A2 => n240, B1 => n1683, B2 => n243,
                           ZN => n1937);
   U2482 : AOI22_X1 port map( A1 => n246, A2 => n2593, B1 => n249, B2 => n836, 
                           ZN => n1935);
   U2483 : NAND4_X1 port map( A1 => n1938, A2 => n1939, A3 => n1940, A4 => 
                           n1941, ZN => n1929);
   U2484 : AOI221_X1 port map( B1 => n252, B2 => n2576, C1 => n255, C2 => n2577
                           , A => n1942, ZN => n1941);
   U2485 : OAI22_X1 port map( A1 => n2575, A2 => n258, B1 => n2574, B2 => n261,
                           ZN => n1942);
   U2486 : AOI221_X1 port map( B1 => n264, B2 => n2580, C1 => n267, C2 => n2581
                           , A => n1943, ZN => n1940);
   U2487 : OAI22_X1 port map( A1 => n2579, A2 => n270, B1 => n2578, B2 => n273,
                           ZN => n1943);
   U2488 : AOI221_X1 port map( B1 => n276, B2 => n633, C1 => n279, C2 => n666, 
                           A => n1944, ZN => n1939);
   U2489 : OAI22_X1 port map( A1 => n1691, A2 => n282, B1 => n1692, B2 => n285,
                           ZN => n1944);
   U2490 : AOI221_X1 port map( B1 => n288, B2 => n599, C1 => n291, C2 => n3796,
                           A => n1945, ZN => n1938);
   U2491 : OAI22_X1 port map( A1 => n1694, A2 => n294, B1 => n1695, B2 => n297,
                           ZN => n1945);
   U2492 : OAI222_X1 port map( A1 => n324, A2 => n198, B1 => n1946, B2 => n201,
                           C1 => n2483, C2 => n204, ZN => n3009);
   U2493 : NOR4_X1 port map( A1 => n1947, A2 => n1948, A3 => n1949, A4 => n1950
                           , ZN => n1946);
   U2494 : OAI221_X1 port map( B1 => n3859, B2 => n207, C1 => n1651, C2 => n210
                           , A => n1951, ZN => n1950);
   U2495 : AOI22_X1 port map( A1 => n213, A2 => n2608, B1 => n216, B2 => n699, 
                           ZN => n1951);
   U2496 : OAI221_X1 port map( B1 => n1653, B2 => n219, C1 => n3763, C2 => n222
                           , A => n1952, ZN => n1949);
   U2497 : AOI22_X1 port map( A1 => n225, A2 => n801, B1 => n228, B2 => n2607, 
                           ZN => n1952);
   U2498 : OAI211_X1 port map( C1 => n2612, C2 => n231, A => n1953, B => n1954,
                           ZN => n1948);
   U2499 : AOI221_X1 port map( B1 => n234, B2 => n935, C1 => n237, C2 => n2613,
                           A => n1955, ZN => n1954);
   U2500 : OAI22_X1 port map( A1 => n2609, A2 => n240, B1 => n1658, B2 => n243,
                           ZN => n1955);
   U2501 : AOI22_X1 port map( A1 => n246, A2 => n2614, B1 => n249, B2 => n835, 
                           ZN => n1953);
   U2502 : NAND4_X1 port map( A1 => n1956, A2 => n1957, A3 => n1958, A4 => 
                           n1959, ZN => n1947);
   U2503 : AOI221_X1 port map( B1 => n252, B2 => n2597, C1 => n255, C2 => n2598
                           , A => n1960, ZN => n1959);
   U2504 : OAI22_X1 port map( A1 => n2596, A2 => n258, B1 => n2595, B2 => n261,
                           ZN => n1960);
   U2505 : AOI221_X1 port map( B1 => n264, B2 => n2601, C1 => n267, C2 => n2602
                           , A => n1961, ZN => n1958);
   U2506 : OAI22_X1 port map( A1 => n2600, A2 => n270, B1 => n2599, B2 => n273,
                           ZN => n1961);
   U2507 : AOI221_X1 port map( B1 => n276, B2 => n632, C1 => n279, C2 => n665, 
                           A => n1962, ZN => n1957);
   U2508 : OAI22_X1 port map( A1 => n1666, A2 => n282, B1 => n1667, B2 => n285,
                           ZN => n1962);
   U2509 : AOI221_X1 port map( B1 => n288, B2 => n598, C1 => n291, C2 => n3795,
                           A => n1963, ZN => n1956);
   U2510 : OAI22_X1 port map( A1 => n1669, A2 => n294, B1 => n1670, B2 => n297,
                           ZN => n1963);
   U2511 : OAI222_X1 port map( A1 => n323, A2 => n198, B1 => n1964, B2 => n201,
                           C1 => n2482, C2 => n204, ZN => n3008);
   U2512 : NOR4_X1 port map( A1 => n1965, A2 => n1966, A3 => n1967, A4 => n1968
                           , ZN => n1964);
   U2513 : OAI221_X1 port map( B1 => n3858, B2 => n207, C1 => n1626, C2 => n210
                           , A => n1969, ZN => n1968);
   U2514 : AOI22_X1 port map( A1 => n213, A2 => n2629, B1 => n216, B2 => n698, 
                           ZN => n1969);
   U2515 : OAI221_X1 port map( B1 => n1628, B2 => n219, C1 => n3762, C2 => n222
                           , A => n1970, ZN => n1967);
   U2516 : AOI22_X1 port map( A1 => n225, A2 => n800, B1 => n228, B2 => n2628, 
                           ZN => n1970);
   U2517 : OAI211_X1 port map( C1 => n2633, C2 => n231, A => n1971, B => n1972,
                           ZN => n1966);
   U2518 : AOI221_X1 port map( B1 => n234, B2 => n934, C1 => n237, C2 => n2634,
                           A => n1973, ZN => n1972);
   U2519 : OAI22_X1 port map( A1 => n2630, A2 => n240, B1 => n1633, B2 => n243,
                           ZN => n1973);
   U2520 : AOI22_X1 port map( A1 => n246, A2 => n2635, B1 => n249, B2 => n834, 
                           ZN => n1971);
   U2521 : NAND4_X1 port map( A1 => n1974, A2 => n1975, A3 => n1976, A4 => 
                           n1977, ZN => n1965);
   U2522 : AOI221_X1 port map( B1 => n252, B2 => n2618, C1 => n255, C2 => n2619
                           , A => n1978, ZN => n1977);
   U2523 : OAI22_X1 port map( A1 => n2617, A2 => n258, B1 => n2616, B2 => n261,
                           ZN => n1978);
   U2524 : AOI221_X1 port map( B1 => n264, B2 => n2622, C1 => n267, C2 => n2623
                           , A => n1979, ZN => n1976);
   U2525 : OAI22_X1 port map( A1 => n2621, A2 => n270, B1 => n2620, B2 => n273,
                           ZN => n1979);
   U2526 : AOI221_X1 port map( B1 => n276, B2 => n631, C1 => n279, C2 => n664, 
                           A => n1980, ZN => n1975);
   U2527 : OAI22_X1 port map( A1 => n1641, A2 => n282, B1 => n1642, B2 => n285,
                           ZN => n1980);
   U2528 : AOI221_X1 port map( B1 => n288, B2 => n597, C1 => n291, C2 => n3794,
                           A => n1981, ZN => n1974);
   U2529 : OAI22_X1 port map( A1 => n1644, A2 => n294, B1 => n1645, B2 => n297,
                           ZN => n1981);
   U2530 : OAI222_X1 port map( A1 => n322, A2 => n198, B1 => n1982, B2 => n201,
                           C1 => n2481, C2 => n204, ZN => n3007);
   U2531 : NOR4_X1 port map( A1 => n1983, A2 => n1984, A3 => n1985, A4 => n1986
                           , ZN => n1982);
   U2532 : OAI221_X1 port map( B1 => n3857, B2 => n207, C1 => n1601, C2 => n210
                           , A => n1987, ZN => n1986);
   U2533 : AOI22_X1 port map( A1 => n213, A2 => n2650, B1 => n216, B2 => n697, 
                           ZN => n1987);
   U2534 : OAI221_X1 port map( B1 => n1603, B2 => n219, C1 => n3761, C2 => n222
                           , A => n1988, ZN => n1985);
   U2535 : AOI22_X1 port map( A1 => n225, A2 => n799, B1 => n228, B2 => n2649, 
                           ZN => n1988);
   U2536 : OAI211_X1 port map( C1 => n2654, C2 => n231, A => n1989, B => n1990,
                           ZN => n1984);
   U2537 : AOI221_X1 port map( B1 => n234, B2 => n933, C1 => n237, C2 => n2655,
                           A => n1991, ZN => n1990);
   U2538 : OAI22_X1 port map( A1 => n2651, A2 => n240, B1 => n1608, B2 => n243,
                           ZN => n1991);
   U2539 : AOI22_X1 port map( A1 => n246, A2 => n2656, B1 => n249, B2 => n833, 
                           ZN => n1989);
   U2540 : NAND4_X1 port map( A1 => n1992, A2 => n1993, A3 => n1994, A4 => 
                           n1995, ZN => n1983);
   U2541 : AOI221_X1 port map( B1 => n252, B2 => n2639, C1 => n255, C2 => n2640
                           , A => n1996, ZN => n1995);
   U2542 : OAI22_X1 port map( A1 => n2638, A2 => n258, B1 => n2637, B2 => n261,
                           ZN => n1996);
   U2543 : AOI221_X1 port map( B1 => n264, B2 => n2643, C1 => n267, C2 => n2644
                           , A => n1997, ZN => n1994);
   U2544 : OAI22_X1 port map( A1 => n2642, A2 => n270, B1 => n2641, B2 => n273,
                           ZN => n1997);
   U2545 : AOI221_X1 port map( B1 => n276, B2 => n630, C1 => n279, C2 => n663, 
                           A => n1998, ZN => n1993);
   U2546 : OAI22_X1 port map( A1 => n1616, A2 => n282, B1 => n1617, B2 => n285,
                           ZN => n1998);
   U2547 : AOI221_X1 port map( B1 => n288, B2 => n596, C1 => n291, C2 => n3793,
                           A => n1999, ZN => n1992);
   U2548 : OAI22_X1 port map( A1 => n1619, A2 => n294, B1 => n1620, B2 => n297,
                           ZN => n1999);
   U2549 : OAI222_X1 port map( A1 => n321, A2 => n197, B1 => n2000, B2 => n200,
                           C1 => n2480, C2 => n204, ZN => n3006);
   U2550 : NOR4_X1 port map( A1 => n2001, A2 => n2002, A3 => n2003, A4 => n2004
                           , ZN => n2000);
   U2551 : OAI221_X1 port map( B1 => n3856, B2 => n206, C1 => n1576, C2 => n209
                           , A => n2005, ZN => n2004);
   U2552 : AOI22_X1 port map( A1 => n212, A2 => n2671, B1 => n215, B2 => n696, 
                           ZN => n2005);
   U2553 : OAI221_X1 port map( B1 => n1578, B2 => n218, C1 => n3760, C2 => n221
                           , A => n2006, ZN => n2003);
   U2554 : AOI22_X1 port map( A1 => n224, A2 => n798, B1 => n227, B2 => n2670, 
                           ZN => n2006);
   U2555 : OAI211_X1 port map( C1 => n2675, C2 => n230, A => n2007, B => n2008,
                           ZN => n2002);
   U2556 : AOI221_X1 port map( B1 => n233, B2 => n932, C1 => n236, C2 => n2676,
                           A => n2009, ZN => n2008);
   U2557 : OAI22_X1 port map( A1 => n2672, A2 => n239, B1 => n1583, B2 => n242,
                           ZN => n2009);
   U2558 : AOI22_X1 port map( A1 => n245, A2 => n2677, B1 => n248, B2 => n832, 
                           ZN => n2007);
   U2559 : NAND4_X1 port map( A1 => n2010, A2 => n2011, A3 => n2012, A4 => 
                           n2013, ZN => n2001);
   U2560 : AOI221_X1 port map( B1 => n251, B2 => n2660, C1 => n254, C2 => n2661
                           , A => n2014, ZN => n2013);
   U2561 : OAI22_X1 port map( A1 => n2659, A2 => n257, B1 => n2658, B2 => n260,
                           ZN => n2014);
   U2562 : AOI221_X1 port map( B1 => n263, B2 => n2664, C1 => n266, C2 => n2665
                           , A => n2015, ZN => n2012);
   U2563 : OAI22_X1 port map( A1 => n2663, A2 => n269, B1 => n2662, B2 => n272,
                           ZN => n2015);
   U2564 : AOI221_X1 port map( B1 => n275, B2 => n629, C1 => n278, C2 => n662, 
                           A => n2016, ZN => n2011);
   U2565 : OAI22_X1 port map( A1 => n1591, A2 => n281, B1 => n1592, B2 => n284,
                           ZN => n2016);
   U2566 : AOI221_X1 port map( B1 => n287, B2 => n595, C1 => n290, C2 => n3792,
                           A => n2017, ZN => n2010);
   U2567 : OAI22_X1 port map( A1 => n1594, A2 => n293, B1 => n1595, B2 => n296,
                           ZN => n2017);
   U2568 : OAI222_X1 port map( A1 => n320, A2 => n197, B1 => n2018, B2 => n200,
                           C1 => n2479, C2 => n204, ZN => n3005);
   U2569 : NOR4_X1 port map( A1 => n2019, A2 => n2020, A3 => n2021, A4 => n2022
                           , ZN => n2018);
   U2570 : OAI221_X1 port map( B1 => n3855, B2 => n206, C1 => n1551, C2 => n209
                           , A => n2023, ZN => n2022);
   U2571 : AOI22_X1 port map( A1 => n212, A2 => n2692, B1 => n215, B2 => n695, 
                           ZN => n2023);
   U2572 : OAI221_X1 port map( B1 => n1553, B2 => n218, C1 => n3759, C2 => n221
                           , A => n2024, ZN => n2021);
   U2573 : AOI22_X1 port map( A1 => n224, A2 => n797, B1 => n227, B2 => n2691, 
                           ZN => n2024);
   U2574 : OAI211_X1 port map( C1 => n2696, C2 => n230, A => n2025, B => n2026,
                           ZN => n2020);
   U2575 : AOI221_X1 port map( B1 => n233, B2 => n931, C1 => n236, C2 => n2697,
                           A => n2027, ZN => n2026);
   U2576 : OAI22_X1 port map( A1 => n2693, A2 => n239, B1 => n1558, B2 => n242,
                           ZN => n2027);
   U2577 : AOI22_X1 port map( A1 => n245, A2 => n2698, B1 => n248, B2 => n831, 
                           ZN => n2025);
   U2578 : NAND4_X1 port map( A1 => n2028, A2 => n2029, A3 => n2030, A4 => 
                           n2031, ZN => n2019);
   U2579 : AOI221_X1 port map( B1 => n251, B2 => n2681, C1 => n254, C2 => n2682
                           , A => n2032, ZN => n2031);
   U2580 : OAI22_X1 port map( A1 => n2680, A2 => n257, B1 => n2679, B2 => n260,
                           ZN => n2032);
   U2581 : AOI221_X1 port map( B1 => n263, B2 => n2685, C1 => n266, C2 => n2686
                           , A => n2033, ZN => n2030);
   U2582 : OAI22_X1 port map( A1 => n2684, A2 => n269, B1 => n2683, B2 => n272,
                           ZN => n2033);
   U2583 : AOI221_X1 port map( B1 => n275, B2 => n628, C1 => n278, C2 => n661, 
                           A => n2034, ZN => n2029);
   U2584 : OAI22_X1 port map( A1 => n1566, A2 => n281, B1 => n1567, B2 => n284,
                           ZN => n2034);
   U2585 : AOI221_X1 port map( B1 => n287, B2 => n594, C1 => n290, C2 => n3791,
                           A => n2035, ZN => n2028);
   U2586 : OAI22_X1 port map( A1 => n1569, A2 => n293, B1 => n1570, B2 => n296,
                           ZN => n2035);
   U2587 : OAI222_X1 port map( A1 => n319, A2 => n197, B1 => n2036, B2 => n200,
                           C1 => n2478, C2 => n203, ZN => n3004);
   U2588 : NOR4_X1 port map( A1 => n2037, A2 => n2038, A3 => n2039, A4 => n2040
                           , ZN => n2036);
   U2589 : OAI221_X1 port map( B1 => n3854, B2 => n206, C1 => n1526, C2 => n209
                           , A => n2041, ZN => n2040);
   U2590 : AOI22_X1 port map( A1 => n212, A2 => n2713, B1 => n215, B2 => n694, 
                           ZN => n2041);
   U2591 : OAI221_X1 port map( B1 => n1528, B2 => n218, C1 => n3758, C2 => n221
                           , A => n2042, ZN => n2039);
   U2592 : AOI22_X1 port map( A1 => n224, A2 => n796, B1 => n227, B2 => n2712, 
                           ZN => n2042);
   U2593 : OAI211_X1 port map( C1 => n2717, C2 => n230, A => n2043, B => n2044,
                           ZN => n2038);
   U2594 : AOI221_X1 port map( B1 => n233, B2 => n930, C1 => n236, C2 => n2718,
                           A => n2045, ZN => n2044);
   U2595 : OAI22_X1 port map( A1 => n2714, A2 => n239, B1 => n1533, B2 => n242,
                           ZN => n2045);
   U2596 : AOI22_X1 port map( A1 => n245, A2 => n2719, B1 => n248, B2 => n830, 
                           ZN => n2043);
   U2597 : NAND4_X1 port map( A1 => n2046, A2 => n2047, A3 => n2048, A4 => 
                           n2049, ZN => n2037);
   U2598 : AOI221_X1 port map( B1 => n251, B2 => n2702, C1 => n254, C2 => n2703
                           , A => n2050, ZN => n2049);
   U2599 : OAI22_X1 port map( A1 => n2701, A2 => n257, B1 => n2700, B2 => n260,
                           ZN => n2050);
   U2600 : AOI221_X1 port map( B1 => n263, B2 => n2706, C1 => n266, C2 => n2707
                           , A => n2051, ZN => n2048);
   U2601 : OAI22_X1 port map( A1 => n2705, A2 => n269, B1 => n2704, B2 => n272,
                           ZN => n2051);
   U2602 : AOI221_X1 port map( B1 => n275, B2 => n627, C1 => n278, C2 => n660, 
                           A => n2052, ZN => n2047);
   U2603 : OAI22_X1 port map( A1 => n1541, A2 => n281, B1 => n1542, B2 => n284,
                           ZN => n2052);
   U2604 : AOI221_X1 port map( B1 => n287, B2 => n593, C1 => n290, C2 => n3790,
                           A => n2053, ZN => n2046);
   U2605 : OAI22_X1 port map( A1 => n1544, A2 => n293, B1 => n1545, B2 => n296,
                           ZN => n2053);
   U2606 : OAI222_X1 port map( A1 => n318, A2 => n197, B1 => n2054, B2 => n200,
                           C1 => n2477, C2 => n203, ZN => n3003);
   U2607 : NOR4_X1 port map( A1 => n2055, A2 => n2056, A3 => n2057, A4 => n2058
                           , ZN => n2054);
   U2608 : OAI221_X1 port map( B1 => n3853, B2 => n206, C1 => n1501, C2 => n209
                           , A => n2059, ZN => n2058);
   U2609 : AOI22_X1 port map( A1 => n212, A2 => n2734, B1 => n215, B2 => n693, 
                           ZN => n2059);
   U2610 : OAI221_X1 port map( B1 => n1503, B2 => n218, C1 => n3757, C2 => n221
                           , A => n2060, ZN => n2057);
   U2611 : AOI22_X1 port map( A1 => n224, A2 => n795, B1 => n227, B2 => n2733, 
                           ZN => n2060);
   U2612 : OAI211_X1 port map( C1 => n2738, C2 => n230, A => n2061, B => n2062,
                           ZN => n2056);
   U2613 : AOI221_X1 port map( B1 => n233, B2 => n929, C1 => n236, C2 => n2739,
                           A => n2063, ZN => n2062);
   U2614 : OAI22_X1 port map( A1 => n2735, A2 => n239, B1 => n1508, B2 => n242,
                           ZN => n2063);
   U2615 : AOI22_X1 port map( A1 => n245, A2 => n2740, B1 => n248, B2 => n829, 
                           ZN => n2061);
   U2616 : NAND4_X1 port map( A1 => n2064, A2 => n2065, A3 => n2066, A4 => 
                           n2067, ZN => n2055);
   U2617 : AOI221_X1 port map( B1 => n251, B2 => n2723, C1 => n254, C2 => n2724
                           , A => n2068, ZN => n2067);
   U2618 : OAI22_X1 port map( A1 => n2722, A2 => n257, B1 => n2721, B2 => n260,
                           ZN => n2068);
   U2619 : AOI221_X1 port map( B1 => n263, B2 => n2727, C1 => n266, C2 => n2728
                           , A => n2069, ZN => n2066);
   U2620 : OAI22_X1 port map( A1 => n2726, A2 => n269, B1 => n2725, B2 => n272,
                           ZN => n2069);
   U2621 : AOI221_X1 port map( B1 => n275, B2 => n626, C1 => n278, C2 => n659, 
                           A => n2070, ZN => n2065);
   U2622 : OAI22_X1 port map( A1 => n1516, A2 => n281, B1 => n1517, B2 => n284,
                           ZN => n2070);
   U2623 : AOI221_X1 port map( B1 => n287, B2 => n592, C1 => n290, C2 => n3789,
                           A => n2071, ZN => n2064);
   U2624 : OAI22_X1 port map( A1 => n1519, A2 => n293, B1 => n1520, B2 => n296,
                           ZN => n2071);
   U2625 : OAI222_X1 port map( A1 => n317, A2 => n197, B1 => n2072, B2 => n200,
                           C1 => n2476, C2 => n203, ZN => n3002);
   U2626 : NOR4_X1 port map( A1 => n2073, A2 => n2074, A3 => n2075, A4 => n2076
                           , ZN => n2072);
   U2627 : OAI221_X1 port map( B1 => n3852, B2 => n206, C1 => n1476, C2 => n209
                           , A => n2077, ZN => n2076);
   U2628 : AOI22_X1 port map( A1 => n212, A2 => n2755, B1 => n215, B2 => n692, 
                           ZN => n2077);
   U2629 : OAI221_X1 port map( B1 => n1478, B2 => n218, C1 => n3756, C2 => n221
                           , A => n2078, ZN => n2075);
   U2630 : AOI22_X1 port map( A1 => n224, A2 => n794, B1 => n227, B2 => n2754, 
                           ZN => n2078);
   U2631 : OAI211_X1 port map( C1 => n2759, C2 => n230, A => n2079, B => n2080,
                           ZN => n2074);
   U2632 : AOI221_X1 port map( B1 => n233, B2 => n928, C1 => n236, C2 => n2760,
                           A => n2081, ZN => n2080);
   U2633 : OAI22_X1 port map( A1 => n2756, A2 => n239, B1 => n1483, B2 => n242,
                           ZN => n2081);
   U2634 : AOI22_X1 port map( A1 => n245, A2 => n2761, B1 => n248, B2 => n828, 
                           ZN => n2079);
   U2635 : NAND4_X1 port map( A1 => n2082, A2 => n2083, A3 => n2084, A4 => 
                           n2085, ZN => n2073);
   U2636 : AOI221_X1 port map( B1 => n251, B2 => n2744, C1 => n254, C2 => n2745
                           , A => n2086, ZN => n2085);
   U2637 : OAI22_X1 port map( A1 => n2743, A2 => n257, B1 => n2742, B2 => n260,
                           ZN => n2086);
   U2638 : AOI221_X1 port map( B1 => n263, B2 => n2748, C1 => n266, C2 => n2749
                           , A => n2087, ZN => n2084);
   U2639 : OAI22_X1 port map( A1 => n2747, A2 => n269, B1 => n2746, B2 => n272,
                           ZN => n2087);
   U2640 : AOI221_X1 port map( B1 => n275, B2 => n625, C1 => n278, C2 => n658, 
                           A => n2088, ZN => n2083);
   U2641 : OAI22_X1 port map( A1 => n1491, A2 => n281, B1 => n1492, B2 => n284,
                           ZN => n2088);
   U2642 : AOI221_X1 port map( B1 => n287, B2 => n591, C1 => n290, C2 => n3788,
                           A => n2089, ZN => n2082);
   U2643 : OAI22_X1 port map( A1 => n1494, A2 => n293, B1 => n1495, B2 => n296,
                           ZN => n2089);
   U2644 : OAI222_X1 port map( A1 => n316, A2 => n197, B1 => n2090, B2 => n200,
                           C1 => n2475, C2 => n203, ZN => n3001);
   U2645 : NOR4_X1 port map( A1 => n2091, A2 => n2092, A3 => n2093, A4 => n2094
                           , ZN => n2090);
   U2646 : OAI221_X1 port map( B1 => n3851, B2 => n206, C1 => n1451, C2 => n209
                           , A => n2095, ZN => n2094);
   U2647 : AOI22_X1 port map( A1 => n212, A2 => n2776, B1 => n215, B2 => n691, 
                           ZN => n2095);
   U2648 : OAI221_X1 port map( B1 => n1453, B2 => n218, C1 => n3755, C2 => n221
                           , A => n2096, ZN => n2093);
   U2649 : AOI22_X1 port map( A1 => n224, A2 => n793, B1 => n227, B2 => n2775, 
                           ZN => n2096);
   U2650 : OAI211_X1 port map( C1 => n2780, C2 => n230, A => n2097, B => n2098,
                           ZN => n2092);
   U2651 : AOI221_X1 port map( B1 => n233, B2 => n927, C1 => n236, C2 => n2781,
                           A => n2099, ZN => n2098);
   U2652 : OAI22_X1 port map( A1 => n2777, A2 => n239, B1 => n1458, B2 => n242,
                           ZN => n2099);
   U2653 : AOI22_X1 port map( A1 => n245, A2 => n2782, B1 => n248, B2 => n827, 
                           ZN => n2097);
   U2654 : NAND4_X1 port map( A1 => n2100, A2 => n2101, A3 => n2102, A4 => 
                           n2103, ZN => n2091);
   U2655 : AOI221_X1 port map( B1 => n251, B2 => n2765, C1 => n254, C2 => n2766
                           , A => n2104, ZN => n2103);
   U2656 : OAI22_X1 port map( A1 => n2764, A2 => n257, B1 => n2763, B2 => n260,
                           ZN => n2104);
   U2657 : AOI221_X1 port map( B1 => n263, B2 => n2769, C1 => n266, C2 => n2770
                           , A => n2105, ZN => n2102);
   U2658 : OAI22_X1 port map( A1 => n2768, A2 => n269, B1 => n2767, B2 => n272,
                           ZN => n2105);
   U2659 : AOI221_X1 port map( B1 => n275, B2 => n624, C1 => n278, C2 => n657, 
                           A => n2106, ZN => n2101);
   U2660 : OAI22_X1 port map( A1 => n1466, A2 => n281, B1 => n1467, B2 => n284,
                           ZN => n2106);
   U2661 : AOI221_X1 port map( B1 => n287, B2 => n590, C1 => n290, C2 => n3787,
                           A => n2107, ZN => n2100);
   U2662 : OAI22_X1 port map( A1 => n1469, A2 => n293, B1 => n1470, B2 => n296,
                           ZN => n2107);
   U2663 : OAI222_X1 port map( A1 => n315, A2 => n197, B1 => n2108, B2 => n200,
                           C1 => n2474, C2 => n203, ZN => n3000);
   U2664 : NOR4_X1 port map( A1 => n2109, A2 => n2110, A3 => n2111, A4 => n2112
                           , ZN => n2108);
   U2665 : OAI221_X1 port map( B1 => n3850, B2 => n206, C1 => n1426, C2 => n209
                           , A => n2113, ZN => n2112);
   U2666 : AOI22_X1 port map( A1 => n212, A2 => n2797, B1 => n215, B2 => n690, 
                           ZN => n2113);
   U2667 : OAI221_X1 port map( B1 => n1428, B2 => n218, C1 => n3754, C2 => n221
                           , A => n2114, ZN => n2111);
   U2668 : AOI22_X1 port map( A1 => n224, A2 => n792, B1 => n227, B2 => n2796, 
                           ZN => n2114);
   U2669 : OAI211_X1 port map( C1 => n2801, C2 => n230, A => n2115, B => n2116,
                           ZN => n2110);
   U2670 : AOI221_X1 port map( B1 => n233, B2 => n926, C1 => n236, C2 => n2802,
                           A => n2117, ZN => n2116);
   U2671 : OAI22_X1 port map( A1 => n2798, A2 => n239, B1 => n1433, B2 => n242,
                           ZN => n2117);
   U2672 : AOI22_X1 port map( A1 => n245, A2 => n2803, B1 => n248, B2 => n826, 
                           ZN => n2115);
   U2673 : NAND4_X1 port map( A1 => n2118, A2 => n2119, A3 => n2120, A4 => 
                           n2121, ZN => n2109);
   U2674 : AOI221_X1 port map( B1 => n251, B2 => n2786, C1 => n254, C2 => n2787
                           , A => n2122, ZN => n2121);
   U2675 : OAI22_X1 port map( A1 => n2785, A2 => n257, B1 => n2784, B2 => n260,
                           ZN => n2122);
   U2676 : AOI221_X1 port map( B1 => n263, B2 => n2790, C1 => n266, C2 => n2791
                           , A => n2123, ZN => n2120);
   U2677 : OAI22_X1 port map( A1 => n2789, A2 => n269, B1 => n2788, B2 => n272,
                           ZN => n2123);
   U2678 : AOI221_X1 port map( B1 => n275, B2 => n623, C1 => n278, C2 => n656, 
                           A => n2124, ZN => n2119);
   U2679 : OAI22_X1 port map( A1 => n1441, A2 => n281, B1 => n1442, B2 => n284,
                           ZN => n2124);
   U2680 : AOI221_X1 port map( B1 => n287, B2 => n589, C1 => n290, C2 => n3786,
                           A => n2125, ZN => n2118);
   U2681 : OAI22_X1 port map( A1 => n1444, A2 => n293, B1 => n1445, B2 => n296,
                           ZN => n2125);
   U2682 : OAI222_X1 port map( A1 => n314, A2 => n197, B1 => n2126, B2 => n200,
                           C1 => n2473, C2 => n203, ZN => n2999);
   U2683 : NOR4_X1 port map( A1 => n2127, A2 => n2128, A3 => n2129, A4 => n2130
                           , ZN => n2126);
   U2684 : OAI221_X1 port map( B1 => n3849, B2 => n206, C1 => n1401, C2 => n209
                           , A => n2131, ZN => n2130);
   U2685 : AOI22_X1 port map( A1 => n212, A2 => n2818, B1 => n215, B2 => n689, 
                           ZN => n2131);
   U2686 : OAI221_X1 port map( B1 => n1403, B2 => n218, C1 => n3753, C2 => n221
                           , A => n2132, ZN => n2129);
   U2687 : AOI22_X1 port map( A1 => n224, A2 => n791, B1 => n227, B2 => n2817, 
                           ZN => n2132);
   U2688 : OAI211_X1 port map( C1 => n2822, C2 => n230, A => n2133, B => n2134,
                           ZN => n2128);
   U2689 : AOI221_X1 port map( B1 => n233, B2 => n925, C1 => n236, C2 => n2823,
                           A => n2135, ZN => n2134);
   U2690 : OAI22_X1 port map( A1 => n2819, A2 => n239, B1 => n1408, B2 => n242,
                           ZN => n2135);
   U2691 : AOI22_X1 port map( A1 => n245, A2 => n2824, B1 => n248, B2 => n825, 
                           ZN => n2133);
   U2692 : NAND4_X1 port map( A1 => n2136, A2 => n2137, A3 => n2138, A4 => 
                           n2139, ZN => n2127);
   U2693 : AOI221_X1 port map( B1 => n251, B2 => n2807, C1 => n254, C2 => n2808
                           , A => n2140, ZN => n2139);
   U2694 : OAI22_X1 port map( A1 => n2806, A2 => n257, B1 => n2805, B2 => n260,
                           ZN => n2140);
   U2695 : AOI221_X1 port map( B1 => n263, B2 => n2811, C1 => n266, C2 => n2812
                           , A => n2141, ZN => n2138);
   U2696 : OAI22_X1 port map( A1 => n2810, A2 => n269, B1 => n2809, B2 => n272,
                           ZN => n2141);
   U2697 : AOI221_X1 port map( B1 => n275, B2 => n622, C1 => n278, C2 => n655, 
                           A => n2142, ZN => n2137);
   U2698 : OAI22_X1 port map( A1 => n1416, A2 => n281, B1 => n1417, B2 => n284,
                           ZN => n2142);
   U2699 : AOI221_X1 port map( B1 => n287, B2 => n588, C1 => n290, C2 => n3785,
                           A => n2143, ZN => n2136);
   U2700 : OAI22_X1 port map( A1 => n1419, A2 => n293, B1 => n1420, B2 => n296,
                           ZN => n2143);
   U2701 : OAI222_X1 port map( A1 => n313, A2 => n197, B1 => n2144, B2 => n200,
                           C1 => n2472, C2 => n203, ZN => n2998);
   U2702 : NOR4_X1 port map( A1 => n2145, A2 => n2146, A3 => n2147, A4 => n2148
                           , ZN => n2144);
   U2703 : OAI221_X1 port map( B1 => n3848, B2 => n206, C1 => n1376, C2 => n209
                           , A => n2149, ZN => n2148);
   U2704 : AOI22_X1 port map( A1 => n212, A2 => n2839, B1 => n215, B2 => n688, 
                           ZN => n2149);
   U2705 : OAI221_X1 port map( B1 => n1378, B2 => n218, C1 => n3752, C2 => n221
                           , A => n2150, ZN => n2147);
   U2706 : AOI22_X1 port map( A1 => n224, A2 => n790, B1 => n227, B2 => n2838, 
                           ZN => n2150);
   U2707 : OAI211_X1 port map( C1 => n2843, C2 => n230, A => n2151, B => n2152,
                           ZN => n2146);
   U2708 : AOI221_X1 port map( B1 => n233, B2 => n924, C1 => n236, C2 => n2844,
                           A => n2153, ZN => n2152);
   U2709 : OAI22_X1 port map( A1 => n2840, A2 => n239, B1 => n1383, B2 => n242,
                           ZN => n2153);
   U2710 : AOI22_X1 port map( A1 => n245, A2 => n2845, B1 => n248, B2 => n824, 
                           ZN => n2151);
   U2711 : NAND4_X1 port map( A1 => n2154, A2 => n2155, A3 => n2156, A4 => 
                           n2157, ZN => n2145);
   U2712 : AOI221_X1 port map( B1 => n251, B2 => n2828, C1 => n254, C2 => n2829
                           , A => n2158, ZN => n2157);
   U2713 : OAI22_X1 port map( A1 => n2827, A2 => n257, B1 => n2826, B2 => n260,
                           ZN => n2158);
   U2714 : AOI221_X1 port map( B1 => n263, B2 => n2832, C1 => n266, C2 => n2833
                           , A => n2159, ZN => n2156);
   U2715 : OAI22_X1 port map( A1 => n2831, A2 => n269, B1 => n2830, B2 => n272,
                           ZN => n2159);
   U2716 : AOI221_X1 port map( B1 => n275, B2 => n621, C1 => n278, C2 => n654, 
                           A => n2160, ZN => n2155);
   U2717 : OAI22_X1 port map( A1 => n1391, A2 => n281, B1 => n1392, B2 => n284,
                           ZN => n2160);
   U2718 : AOI221_X1 port map( B1 => n287, B2 => n587, C1 => n290, C2 => n3784,
                           A => n2161, ZN => n2154);
   U2719 : OAI22_X1 port map( A1 => n1394, A2 => n293, B1 => n1395, B2 => n296,
                           ZN => n2161);
   U2720 : OAI222_X1 port map( A1 => n312, A2 => n197, B1 => n2162, B2 => n200,
                           C1 => n2471, C2 => n203, ZN => n2997);
   U2721 : NOR4_X1 port map( A1 => n2163, A2 => n2164, A3 => n2165, A4 => n2166
                           , ZN => n2162);
   U2722 : OAI221_X1 port map( B1 => n3847, B2 => n206, C1 => n1351, C2 => n209
                           , A => n2167, ZN => n2166);
   U2723 : AOI22_X1 port map( A1 => n212, A2 => n2860, B1 => n215, B2 => n687, 
                           ZN => n2167);
   U2724 : OAI221_X1 port map( B1 => n1353, B2 => n218, C1 => n3751, C2 => n221
                           , A => n2168, ZN => n2165);
   U2725 : AOI22_X1 port map( A1 => n224, A2 => n789, B1 => n227, B2 => n2859, 
                           ZN => n2168);
   U2726 : OAI211_X1 port map( C1 => n2864, C2 => n230, A => n2169, B => n2170,
                           ZN => n2164);
   U2727 : AOI221_X1 port map( B1 => n233, B2 => n923, C1 => n236, C2 => n2865,
                           A => n2171, ZN => n2170);
   U2728 : OAI22_X1 port map( A1 => n2861, A2 => n239, B1 => n1358, B2 => n242,
                           ZN => n2171);
   U2729 : AOI22_X1 port map( A1 => n245, A2 => n2866, B1 => n248, B2 => n823, 
                           ZN => n2169);
   U2730 : NAND4_X1 port map( A1 => n2172, A2 => n2173, A3 => n2174, A4 => 
                           n2175, ZN => n2163);
   U2731 : AOI221_X1 port map( B1 => n251, B2 => n2849, C1 => n254, C2 => n2850
                           , A => n2176, ZN => n2175);
   U2732 : OAI22_X1 port map( A1 => n2848, A2 => n257, B1 => n2847, B2 => n260,
                           ZN => n2176);
   U2733 : AOI221_X1 port map( B1 => n263, B2 => n2853, C1 => n266, C2 => n2854
                           , A => n2177, ZN => n2174);
   U2734 : OAI22_X1 port map( A1 => n2852, A2 => n269, B1 => n2851, B2 => n272,
                           ZN => n2177);
   U2735 : AOI221_X1 port map( B1 => n275, B2 => n620, C1 => n278, C2 => n653, 
                           A => n2178, ZN => n2173);
   U2736 : OAI22_X1 port map( A1 => n1366, A2 => n281, B1 => n1367, B2 => n284,
                           ZN => n2178);
   U2737 : AOI221_X1 port map( B1 => n287, B2 => n586, C1 => n290, C2 => n3783,
                           A => n2179, ZN => n2172);
   U2738 : OAI22_X1 port map( A1 => n1369, A2 => n293, B1 => n1370, B2 => n296,
                           ZN => n2179);
   U2739 : OAI222_X1 port map( A1 => n311, A2 => n197, B1 => n2180, B2 => n200,
                           C1 => n2470, C2 => n203, ZN => n2996);
   U2740 : NOR4_X1 port map( A1 => n2181, A2 => n2182, A3 => n2183, A4 => n2184
                           , ZN => n2180);
   U2741 : OAI221_X1 port map( B1 => n3846, B2 => n206, C1 => n1326, C2 => n209
                           , A => n2185, ZN => n2184);
   U2742 : AOI22_X1 port map( A1 => n212, A2 => n2881, B1 => n215, B2 => n686, 
                           ZN => n2185);
   U2743 : OAI221_X1 port map( B1 => n1328, B2 => n218, C1 => n3750, C2 => n221
                           , A => n2186, ZN => n2183);
   U2744 : AOI22_X1 port map( A1 => n224, A2 => n788, B1 => n227, B2 => n2880, 
                           ZN => n2186);
   U2745 : OAI211_X1 port map( C1 => n2885, C2 => n230, A => n2187, B => n2188,
                           ZN => n2182);
   U2746 : AOI221_X1 port map( B1 => n233, B2 => n922, C1 => n236, C2 => n2886,
                           A => n2189, ZN => n2188);
   U2747 : OAI22_X1 port map( A1 => n2882, A2 => n239, B1 => n1333, B2 => n242,
                           ZN => n2189);
   U2748 : AOI22_X1 port map( A1 => n245, A2 => n2887, B1 => n248, B2 => n822, 
                           ZN => n2187);
   U2749 : NAND4_X1 port map( A1 => n2190, A2 => n2191, A3 => n2192, A4 => 
                           n2193, ZN => n2181);
   U2750 : AOI221_X1 port map( B1 => n251, B2 => n2870, C1 => n254, C2 => n2871
                           , A => n2194, ZN => n2193);
   U2751 : OAI22_X1 port map( A1 => n2869, A2 => n257, B1 => n2868, B2 => n260,
                           ZN => n2194);
   U2752 : AOI221_X1 port map( B1 => n263, B2 => n2874, C1 => n266, C2 => n2875
                           , A => n2195, ZN => n2192);
   U2753 : OAI22_X1 port map( A1 => n2873, A2 => n269, B1 => n2872, B2 => n272,
                           ZN => n2195);
   U2754 : AOI221_X1 port map( B1 => n275, B2 => n619, C1 => n278, C2 => n652, 
                           A => n2196, ZN => n2191);
   U2755 : OAI22_X1 port map( A1 => n1341, A2 => n281, B1 => n1342, B2 => n284,
                           ZN => n2196);
   U2756 : AOI221_X1 port map( B1 => n287, B2 => n585, C1 => n290, C2 => n3782,
                           A => n2197, ZN => n2190);
   U2757 : OAI22_X1 port map( A1 => n1344, A2 => n293, B1 => n1345, B2 => n296,
                           ZN => n2197);
   U2758 : OAI222_X1 port map( A1 => n310, A2 => n197, B1 => n2198, B2 => n200,
                           C1 => n2469, C2 => n203, ZN => n2995);
   U2759 : NOR4_X1 port map( A1 => n2199, A2 => n2200, A3 => n2201, A4 => n2202
                           , ZN => n2198);
   U2760 : OAI221_X1 port map( B1 => n3845, B2 => n206, C1 => n1301, C2 => n209
                           , A => n2203, ZN => n2202);
   U2761 : AOI22_X1 port map( A1 => n212, A2 => n2902, B1 => n215, B2 => n685, 
                           ZN => n2203);
   U2762 : OAI221_X1 port map( B1 => n1303, B2 => n218, C1 => n3749, C2 => n221
                           , A => n2204, ZN => n2201);
   U2763 : AOI22_X1 port map( A1 => n224, A2 => n787, B1 => n227, B2 => n2901, 
                           ZN => n2204);
   U2764 : OAI211_X1 port map( C1 => n2906, C2 => n230, A => n2205, B => n2206,
                           ZN => n2200);
   U2765 : AOI221_X1 port map( B1 => n233, B2 => n921, C1 => n236, C2 => n2907,
                           A => n2207, ZN => n2206);
   U2766 : OAI22_X1 port map( A1 => n2903, A2 => n239, B1 => n1308, B2 => n242,
                           ZN => n2207);
   U2767 : AOI22_X1 port map( A1 => n245, A2 => n2908, B1 => n248, B2 => n821, 
                           ZN => n2205);
   U2768 : NAND4_X1 port map( A1 => n2208, A2 => n2209, A3 => n2210, A4 => 
                           n2211, ZN => n2199);
   U2769 : AOI221_X1 port map( B1 => n251, B2 => n2891, C1 => n254, C2 => n2892
                           , A => n2212, ZN => n2211);
   U2770 : OAI22_X1 port map( A1 => n2890, A2 => n257, B1 => n2889, B2 => n260,
                           ZN => n2212);
   U2771 : AOI221_X1 port map( B1 => n263, B2 => n2895, C1 => n266, C2 => n2896
                           , A => n2213, ZN => n2210);
   U2772 : OAI22_X1 port map( A1 => n2894, A2 => n269, B1 => n2893, B2 => n272,
                           ZN => n2213);
   U2773 : AOI221_X1 port map( B1 => n275, B2 => n618, C1 => n278, C2 => n651, 
                           A => n2214, ZN => n2209);
   U2774 : OAI22_X1 port map( A1 => n1316, A2 => n281, B1 => n1317, B2 => n284,
                           ZN => n2214);
   U2775 : AOI221_X1 port map( B1 => n287, B2 => n584, C1 => n290, C2 => n3781,
                           A => n2215, ZN => n2208);
   U2776 : OAI22_X1 port map( A1 => n1319, A2 => n293, B1 => n1320, B2 => n296,
                           ZN => n2215);
   U2777 : OAI222_X1 port map( A1 => n309, A2 => n196, B1 => n2216, B2 => n199,
                           C1 => n2468, C2 => n203, ZN => n2994);
   U2778 : NOR4_X1 port map( A1 => n2217, A2 => n2218, A3 => n2219, A4 => n2220
                           , ZN => n2216);
   U2779 : OAI221_X1 port map( B1 => n3844, B2 => n205, C1 => n1276, C2 => n208
                           , A => n2221, ZN => n2220);
   U2780 : AOI22_X1 port map( A1 => n211, A2 => n2923, B1 => n214, B2 => n684, 
                           ZN => n2221);
   U2781 : OAI221_X1 port map( B1 => n1278, B2 => n217, C1 => n3748, C2 => n220
                           , A => n2222, ZN => n2219);
   U2782 : AOI22_X1 port map( A1 => n223, A2 => n786, B1 => n226, B2 => n2922, 
                           ZN => n2222);
   U2783 : OAI211_X1 port map( C1 => n2927, C2 => n229, A => n2223, B => n2224,
                           ZN => n2218);
   U2784 : AOI221_X1 port map( B1 => n232, B2 => n920, C1 => n235, C2 => n2928,
                           A => n2225, ZN => n2224);
   U2785 : OAI22_X1 port map( A1 => n2924, A2 => n238, B1 => n1283, B2 => n241,
                           ZN => n2225);
   U2786 : AOI22_X1 port map( A1 => n244, A2 => n2929, B1 => n247, B2 => n820, 
                           ZN => n2223);
   U2787 : NAND4_X1 port map( A1 => n2226, A2 => n2227, A3 => n2228, A4 => 
                           n2229, ZN => n2217);
   U2788 : AOI221_X1 port map( B1 => n250, B2 => n2912, C1 => n253, C2 => n2913
                           , A => n2230, ZN => n2229);
   U2789 : OAI22_X1 port map( A1 => n2911, A2 => n256, B1 => n2910, B2 => n259,
                           ZN => n2230);
   U2790 : AOI221_X1 port map( B1 => n262, B2 => n2916, C1 => n265, C2 => n2917
                           , A => n2231, ZN => n2228);
   U2791 : OAI22_X1 port map( A1 => n2915, A2 => n268, B1 => n2914, B2 => n271,
                           ZN => n2231);
   U2792 : AOI221_X1 port map( B1 => n274, B2 => n617, C1 => n277, C2 => n650, 
                           A => n2232, ZN => n2227);
   U2793 : OAI22_X1 port map( A1 => n1291, A2 => n280, B1 => n1292, B2 => n283,
                           ZN => n2232);
   U2794 : AOI221_X1 port map( B1 => n286, B2 => n583, C1 => n289, C2 => n3780,
                           A => n2233, ZN => n2226);
   U2795 : OAI22_X1 port map( A1 => n1294, A2 => n292, B1 => n1295, B2 => n295,
                           ZN => n2233);
   U2796 : OAI222_X1 port map( A1 => n308, A2 => n196, B1 => n2234, B2 => n199,
                           C1 => n2467, C2 => n203, ZN => n2993);
   U2797 : NOR4_X1 port map( A1 => n2235, A2 => n2236, A3 => n2237, A4 => n2238
                           , ZN => n2234);
   U2798 : OAI221_X1 port map( B1 => n3843, B2 => n205, C1 => n1251, C2 => n208
                           , A => n2239, ZN => n2238);
   U2799 : AOI22_X1 port map( A1 => n211, A2 => n2944, B1 => n214, B2 => n683, 
                           ZN => n2239);
   U2800 : OAI221_X1 port map( B1 => n1253, B2 => n217, C1 => n3747, C2 => n220
                           , A => n2240, ZN => n2237);
   U2801 : AOI22_X1 port map( A1 => n223, A2 => n785, B1 => n226, B2 => n2943, 
                           ZN => n2240);
   U2802 : OAI211_X1 port map( C1 => n2948, C2 => n229, A => n2241, B => n2242,
                           ZN => n2236);
   U2803 : AOI221_X1 port map( B1 => n232, B2 => n919, C1 => n235, C2 => n2949,
                           A => n2243, ZN => n2242);
   U2804 : OAI22_X1 port map( A1 => n2945, A2 => n238, B1 => n1258, B2 => n241,
                           ZN => n2243);
   U2805 : AOI22_X1 port map( A1 => n244, A2 => n2950, B1 => n247, B2 => n819, 
                           ZN => n2241);
   U2806 : NAND4_X1 port map( A1 => n2244, A2 => n2245, A3 => n2246, A4 => 
                           n2247, ZN => n2235);
   U2807 : AOI221_X1 port map( B1 => n250, B2 => n2933, C1 => n253, C2 => n2934
                           , A => n2248, ZN => n2247);
   U2808 : OAI22_X1 port map( A1 => n2932, A2 => n256, B1 => n2931, B2 => n259,
                           ZN => n2248);
   U2809 : AOI221_X1 port map( B1 => n262, B2 => n2937, C1 => n265, C2 => n2938
                           , A => n2249, ZN => n2246);
   U2810 : OAI22_X1 port map( A1 => n2936, A2 => n268, B1 => n2935, B2 => n271,
                           ZN => n2249);
   U2811 : AOI221_X1 port map( B1 => n274, B2 => n616, C1 => n277, C2 => n649, 
                           A => n2250, ZN => n2245);
   U2812 : OAI22_X1 port map( A1 => n1266, A2 => n280, B1 => n1267, B2 => n283,
                           ZN => n2250);
   U2813 : AOI221_X1 port map( B1 => n286, B2 => n582, C1 => n289, C2 => n3779,
                           A => n2251, ZN => n2244);
   U2814 : OAI22_X1 port map( A1 => n1269, A2 => n292, B1 => n1270, B2 => n295,
                           ZN => n2251);
   U2815 : OAI222_X1 port map( A1 => n307, A2 => n196, B1 => n2252, B2 => n199,
                           C1 => n2466, C2 => n202, ZN => n2992);
   U2816 : NOR4_X1 port map( A1 => n2253, A2 => n2254, A3 => n2255, A4 => n2256
                           , ZN => n2252);
   U2817 : OAI221_X1 port map( B1 => n3842, B2 => n205, C1 => n1226, C2 => n208
                           , A => n2257, ZN => n2256);
   U2818 : AOI22_X1 port map( A1 => n211, A2 => n2965, B1 => n214, B2 => n682, 
                           ZN => n2257);
   U2819 : OAI221_X1 port map( B1 => n1228, B2 => n217, C1 => n3746, C2 => n220
                           , A => n2258, ZN => n2255);
   U2820 : AOI22_X1 port map( A1 => n223, A2 => n784, B1 => n226, B2 => n2964, 
                           ZN => n2258);
   U2821 : OAI211_X1 port map( C1 => n2969, C2 => n229, A => n2259, B => n2260,
                           ZN => n2254);
   U2822 : AOI221_X1 port map( B1 => n232, B2 => n918, C1 => n235, C2 => n2970,
                           A => n2261, ZN => n2260);
   U2823 : OAI22_X1 port map( A1 => n2966, A2 => n238, B1 => n1233, B2 => n241,
                           ZN => n2261);
   U2824 : AOI22_X1 port map( A1 => n244, A2 => n2971, B1 => n247, B2 => n818, 
                           ZN => n2259);
   U2825 : NAND4_X1 port map( A1 => n2262, A2 => n2263, A3 => n2264, A4 => 
                           n2265, ZN => n2253);
   U2826 : AOI221_X1 port map( B1 => n250, B2 => n2954, C1 => n253, C2 => n2955
                           , A => n2266, ZN => n2265);
   U2827 : OAI22_X1 port map( A1 => n2953, A2 => n256, B1 => n2952, B2 => n259,
                           ZN => n2266);
   U2828 : AOI221_X1 port map( B1 => n262, B2 => n2958, C1 => n265, C2 => n2959
                           , A => n2267, ZN => n2264);
   U2829 : OAI22_X1 port map( A1 => n2957, A2 => n268, B1 => n2956, B2 => n271,
                           ZN => n2267);
   U2830 : AOI221_X1 port map( B1 => n274, B2 => n615, C1 => n277, C2 => n648, 
                           A => n2268, ZN => n2263);
   U2831 : OAI22_X1 port map( A1 => n1241, A2 => n280, B1 => n1242, B2 => n283,
                           ZN => n2268);
   U2832 : AOI221_X1 port map( B1 => n286, B2 => n581, C1 => n289, C2 => n3778,
                           A => n2269, ZN => n2262);
   U2833 : OAI22_X1 port map( A1 => n1244, A2 => n292, B1 => n1245, B2 => n295,
                           ZN => n2269);
   U2834 : OAI222_X1 port map( A1 => n306, A2 => n196, B1 => n2270, B2 => n199,
                           C1 => n2465, C2 => n202, ZN => n2991);
   U2835 : NOR4_X1 port map( A1 => n2271, A2 => n2272, A3 => n2273, A4 => n2274
                           , ZN => n2270);
   U2836 : OAI221_X1 port map( B1 => n3841, B2 => n205, C1 => n1201, C2 => n208
                           , A => n2275, ZN => n2274);
   U2837 : AOI22_X1 port map( A1 => n211, A2 => n3562, B1 => n214, B2 => n681, 
                           ZN => n2275);
   U2838 : OAI221_X1 port map( B1 => n1203, B2 => n217, C1 => n3745, C2 => n220
                           , A => n2276, ZN => n2273);
   U2839 : AOI22_X1 port map( A1 => n223, A2 => n783, B1 => n226, B2 => n3561, 
                           ZN => n2276);
   U2840 : OAI211_X1 port map( C1 => n3566, C2 => n229, A => n2277, B => n2278,
                           ZN => n2272);
   U2841 : AOI221_X1 port map( B1 => n232, B2 => n917, C1 => n235, C2 => n3567,
                           A => n2279, ZN => n2278);
   U2842 : OAI22_X1 port map( A1 => n3563, A2 => n238, B1 => n1208, B2 => n241,
                           ZN => n2279);
   U2843 : AOI22_X1 port map( A1 => n244, A2 => n3568, B1 => n247, B2 => n817, 
                           ZN => n2277);
   U2844 : NAND4_X1 port map( A1 => n2280, A2 => n2281, A3 => n2282, A4 => 
                           n2283, ZN => n2271);
   U2845 : AOI221_X1 port map( B1 => n250, B2 => n2975, C1 => n253, C2 => n2976
                           , A => n2284, ZN => n2283);
   U2846 : OAI22_X1 port map( A1 => n2974, A2 => n256, B1 => n2973, B2 => n259,
                           ZN => n2284);
   U2847 : AOI221_X1 port map( B1 => n262, B2 => n2979, C1 => n265, C2 => n2980
                           , A => n2285, ZN => n2282);
   U2848 : OAI22_X1 port map( A1 => n2978, A2 => n268, B1 => n2977, B2 => n271,
                           ZN => n2285);
   U2849 : AOI221_X1 port map( B1 => n274, B2 => n614, C1 => n277, C2 => n647, 
                           A => n2286, ZN => n2281);
   U2850 : OAI22_X1 port map( A1 => n1216, A2 => n280, B1 => n1217, B2 => n283,
                           ZN => n2286);
   U2851 : AOI221_X1 port map( B1 => n286, B2 => n580, C1 => n289, C2 => n3777,
                           A => n2287, ZN => n2280);
   U2852 : OAI22_X1 port map( A1 => n1219, A2 => n292, B1 => n1220, B2 => n295,
                           ZN => n2287);
   U2853 : OAI222_X1 port map( A1 => n305, A2 => n196, B1 => n2288, B2 => n199,
                           C1 => n2464, C2 => n202, ZN => n2990);
   U2854 : NOR4_X1 port map( A1 => n2289, A2 => n2290, A3 => n2291, A4 => n2292
                           , ZN => n2288);
   U2855 : OAI221_X1 port map( B1 => n3840, B2 => n205, C1 => n1176, C2 => n208
                           , A => n2293, ZN => n2292);
   U2856 : AOI22_X1 port map( A1 => n211, A2 => n3583, B1 => n214, B2 => n680, 
                           ZN => n2293);
   U2857 : OAI221_X1 port map( B1 => n1178, B2 => n217, C1 => n3744, C2 => n220
                           , A => n2294, ZN => n2291);
   U2858 : AOI22_X1 port map( A1 => n223, A2 => n782, B1 => n226, B2 => n3582, 
                           ZN => n2294);
   U2859 : OAI211_X1 port map( C1 => n3587, C2 => n229, A => n2295, B => n2296,
                           ZN => n2290);
   U2860 : AOI221_X1 port map( B1 => n232, B2 => n916, C1 => n235, C2 => n3588,
                           A => n2297, ZN => n2296);
   U2861 : OAI22_X1 port map( A1 => n3584, A2 => n238, B1 => n1183, B2 => n241,
                           ZN => n2297);
   U2862 : AOI22_X1 port map( A1 => n244, A2 => n3589, B1 => n247, B2 => n816, 
                           ZN => n2295);
   U2863 : NAND4_X1 port map( A1 => n2298, A2 => n2299, A3 => n2300, A4 => 
                           n2301, ZN => n2289);
   U2864 : AOI221_X1 port map( B1 => n250, B2 => n3572, C1 => n253, C2 => n3573
                           , A => n2302, ZN => n2301);
   U2865 : OAI22_X1 port map( A1 => n3571, A2 => n256, B1 => n3570, B2 => n259,
                           ZN => n2302);
   U2866 : AOI221_X1 port map( B1 => n262, B2 => n3576, C1 => n265, C2 => n3577
                           , A => n2303, ZN => n2300);
   U2867 : OAI22_X1 port map( A1 => n3575, A2 => n268, B1 => n3574, B2 => n271,
                           ZN => n2303);
   U2868 : AOI221_X1 port map( B1 => n274, B2 => n613, C1 => n277, C2 => n646, 
                           A => n2304, ZN => n2299);
   U2869 : OAI22_X1 port map( A1 => n1191, A2 => n280, B1 => n1192, B2 => n283,
                           ZN => n2304);
   U2870 : AOI221_X1 port map( B1 => n286, B2 => n579, C1 => n289, C2 => n3776,
                           A => n2305, ZN => n2298);
   U2871 : OAI22_X1 port map( A1 => n1194, A2 => n292, B1 => n1195, B2 => n295,
                           ZN => n2305);
   U2872 : OAI222_X1 port map( A1 => n304, A2 => n196, B1 => n2306, B2 => n199,
                           C1 => n2463, C2 => n202, ZN => n2989);
   U2873 : NOR4_X1 port map( A1 => n2307, A2 => n2308, A3 => n2309, A4 => n2310
                           , ZN => n2306);
   U2874 : OAI221_X1 port map( B1 => n3839, B2 => n205, C1 => n1151, C2 => n208
                           , A => n2311, ZN => n2310);
   U2875 : AOI22_X1 port map( A1 => n211, A2 => n3604, B1 => n214, B2 => n679, 
                           ZN => n2311);
   U2876 : OAI221_X1 port map( B1 => n1153, B2 => n217, C1 => n3743, C2 => n220
                           , A => n2312, ZN => n2309);
   U2877 : AOI22_X1 port map( A1 => n223, A2 => n781, B1 => n226, B2 => n3603, 
                           ZN => n2312);
   U2878 : OAI211_X1 port map( C1 => n3608, C2 => n229, A => n2313, B => n2314,
                           ZN => n2308);
   U2879 : AOI221_X1 port map( B1 => n232, B2 => n915, C1 => n235, C2 => n3609,
                           A => n2315, ZN => n2314);
   U2880 : OAI22_X1 port map( A1 => n3605, A2 => n238, B1 => n1158, B2 => n241,
                           ZN => n2315);
   U2881 : AOI22_X1 port map( A1 => n244, A2 => n3610, B1 => n247, B2 => n815, 
                           ZN => n2313);
   U2882 : NAND4_X1 port map( A1 => n2316, A2 => n2317, A3 => n2318, A4 => 
                           n2319, ZN => n2307);
   U2883 : AOI221_X1 port map( B1 => n250, B2 => n3593, C1 => n253, C2 => n3594
                           , A => n2320, ZN => n2319);
   U2884 : OAI22_X1 port map( A1 => n3592, A2 => n256, B1 => n3591, B2 => n259,
                           ZN => n2320);
   U2885 : AOI221_X1 port map( B1 => n262, B2 => n3597, C1 => n265, C2 => n3598
                           , A => n2321, ZN => n2318);
   U2886 : OAI22_X1 port map( A1 => n3596, A2 => n268, B1 => n3595, B2 => n271,
                           ZN => n2321);
   U2887 : AOI221_X1 port map( B1 => n274, B2 => n612, C1 => n277, C2 => n645, 
                           A => n2322, ZN => n2317);
   U2888 : OAI22_X1 port map( A1 => n1166, A2 => n280, B1 => n1167, B2 => n283,
                           ZN => n2322);
   U2889 : AOI221_X1 port map( B1 => n286, B2 => n578, C1 => n289, C2 => n3775,
                           A => n2323, ZN => n2316);
   U2890 : OAI22_X1 port map( A1 => n1169, A2 => n292, B1 => n1170, B2 => n295,
                           ZN => n2323);
   U2891 : OAI222_X1 port map( A1 => n303, A2 => n196, B1 => n2324, B2 => n199,
                           C1 => n2462, C2 => n202, ZN => n2988);
   U2892 : NOR4_X1 port map( A1 => n2325, A2 => n2326, A3 => n2327, A4 => n2328
                           , ZN => n2324);
   U2893 : OAI221_X1 port map( B1 => n3838, B2 => n205, C1 => n1126, C2 => n208
                           , A => n2329, ZN => n2328);
   U2894 : AOI22_X1 port map( A1 => n211, A2 => n3625, B1 => n214, B2 => n678, 
                           ZN => n2329);
   U2895 : OAI221_X1 port map( B1 => n1128, B2 => n217, C1 => n3742, C2 => n220
                           , A => n2330, ZN => n2327);
   U2896 : AOI22_X1 port map( A1 => n223, A2 => n780, B1 => n226, B2 => n3624, 
                           ZN => n2330);
   U2897 : OAI211_X1 port map( C1 => n3629, C2 => n229, A => n2331, B => n2332,
                           ZN => n2326);
   U2898 : AOI221_X1 port map( B1 => n232, B2 => n914, C1 => n235, C2 => n3630,
                           A => n2333, ZN => n2332);
   U2899 : OAI22_X1 port map( A1 => n3626, A2 => n238, B1 => n1133, B2 => n241,
                           ZN => n2333);
   U2900 : AOI22_X1 port map( A1 => n244, A2 => n3631, B1 => n247, B2 => n814, 
                           ZN => n2331);
   U2901 : NAND4_X1 port map( A1 => n2334, A2 => n2335, A3 => n2336, A4 => 
                           n2337, ZN => n2325);
   U2902 : AOI221_X1 port map( B1 => n250, B2 => n3614, C1 => n253, C2 => n3615
                           , A => n2338, ZN => n2337);
   U2903 : OAI22_X1 port map( A1 => n3613, A2 => n256, B1 => n3612, B2 => n259,
                           ZN => n2338);
   U2904 : AOI221_X1 port map( B1 => n262, B2 => n3618, C1 => n265, C2 => n3619
                           , A => n2339, ZN => n2336);
   U2905 : OAI22_X1 port map( A1 => n3617, A2 => n268, B1 => n3616, B2 => n271,
                           ZN => n2339);
   U2906 : AOI221_X1 port map( B1 => n274, B2 => n611, C1 => n277, C2 => n644, 
                           A => n2340, ZN => n2335);
   U2907 : OAI22_X1 port map( A1 => n1141, A2 => n280, B1 => n1142, B2 => n283,
                           ZN => n2340);
   U2908 : AOI221_X1 port map( B1 => n286, B2 => n577, C1 => n289, C2 => n3774,
                           A => n2341, ZN => n2334);
   U2909 : OAI22_X1 port map( A1 => n1144, A2 => n292, B1 => n1145, B2 => n295,
                           ZN => n2341);
   U2910 : OAI222_X1 port map( A1 => n302, A2 => n196, B1 => n2342, B2 => n199,
                           C1 => n2461, C2 => n202, ZN => n2987);
   U2911 : NOR4_X1 port map( A1 => n2343, A2 => n2344, A3 => n2345, A4 => n2346
                           , ZN => n2342);
   U2912 : OAI221_X1 port map( B1 => n3837, B2 => n205, C1 => n1101, C2 => n208
                           , A => n2347, ZN => n2346);
   U2913 : AOI22_X1 port map( A1 => n211, A2 => n3646, B1 => n214, B2 => n677, 
                           ZN => n2347);
   U2914 : OAI221_X1 port map( B1 => n1103, B2 => n217, C1 => n3741, C2 => n220
                           , A => n2348, ZN => n2345);
   U2915 : AOI22_X1 port map( A1 => n223, A2 => n779, B1 => n226, B2 => n3645, 
                           ZN => n2348);
   U2916 : OAI211_X1 port map( C1 => n3650, C2 => n229, A => n2349, B => n2350,
                           ZN => n2344);
   U2917 : AOI221_X1 port map( B1 => n232, B2 => n913, C1 => n235, C2 => n3651,
                           A => n2351, ZN => n2350);
   U2918 : OAI22_X1 port map( A1 => n3647, A2 => n238, B1 => n1108, B2 => n241,
                           ZN => n2351);
   U2919 : AOI22_X1 port map( A1 => n244, A2 => n3652, B1 => n247, B2 => n813, 
                           ZN => n2349);
   U2920 : NAND4_X1 port map( A1 => n2352, A2 => n2353, A3 => n2354, A4 => 
                           n2355, ZN => n2343);
   U2921 : AOI221_X1 port map( B1 => n250, B2 => n3635, C1 => n253, C2 => n3636
                           , A => n2356, ZN => n2355);
   U2922 : OAI22_X1 port map( A1 => n3634, A2 => n256, B1 => n3633, B2 => n259,
                           ZN => n2356);
   U2923 : AOI221_X1 port map( B1 => n262, B2 => n3639, C1 => n265, C2 => n3640
                           , A => n2357, ZN => n2354);
   U2924 : OAI22_X1 port map( A1 => n3638, A2 => n268, B1 => n3637, B2 => n271,
                           ZN => n2357);
   U2925 : AOI221_X1 port map( B1 => n274, B2 => n610, C1 => n277, C2 => n643, 
                           A => n2358, ZN => n2353);
   U2926 : OAI22_X1 port map( A1 => n1116, A2 => n280, B1 => n1117, B2 => n283,
                           ZN => n2358);
   U2927 : AOI221_X1 port map( B1 => n286, B2 => n576, C1 => n289, C2 => n3773,
                           A => n2359, ZN => n2352);
   U2928 : OAI22_X1 port map( A1 => n1119, A2 => n292, B1 => n1120, B2 => n295,
                           ZN => n2359);
   U2929 : OAI222_X1 port map( A1 => n301, A2 => n196, B1 => n2360, B2 => n199,
                           C1 => n2460, C2 => n202, ZN => n2986);
   U2930 : NOR4_X1 port map( A1 => n2361, A2 => n2362, A3 => n2363, A4 => n2364
                           , ZN => n2360);
   U2931 : OAI221_X1 port map( B1 => n3836, B2 => n205, C1 => n1076, C2 => n208
                           , A => n2365, ZN => n2364);
   U2932 : AOI22_X1 port map( A1 => n211, A2 => n3667, B1 => n214, B2 => n676, 
                           ZN => n2365);
   U2933 : OAI221_X1 port map( B1 => n1078, B2 => n217, C1 => n3740, C2 => n220
                           , A => n2366, ZN => n2363);
   U2934 : AOI22_X1 port map( A1 => n223, A2 => n778, B1 => n226, B2 => n3666, 
                           ZN => n2366);
   U2935 : OAI211_X1 port map( C1 => n3671, C2 => n229, A => n2367, B => n2368,
                           ZN => n2362);
   U2936 : AOI221_X1 port map( B1 => n232, B2 => n912, C1 => n235, C2 => n3672,
                           A => n2369, ZN => n2368);
   U2937 : OAI22_X1 port map( A1 => n3668, A2 => n238, B1 => n1083, B2 => n241,
                           ZN => n2369);
   U2938 : AOI22_X1 port map( A1 => n244, A2 => n3673, B1 => n247, B2 => n812, 
                           ZN => n2367);
   U2939 : NAND4_X1 port map( A1 => n2370, A2 => n2371, A3 => n2372, A4 => 
                           n2373, ZN => n2361);
   U2940 : AOI221_X1 port map( B1 => n250, B2 => n3656, C1 => n253, C2 => n3657
                           , A => n2374, ZN => n2373);
   U2941 : OAI22_X1 port map( A1 => n3655, A2 => n256, B1 => n3654, B2 => n259,
                           ZN => n2374);
   U2942 : AOI221_X1 port map( B1 => n262, B2 => n3660, C1 => n265, C2 => n3661
                           , A => n2375, ZN => n2372);
   U2943 : OAI22_X1 port map( A1 => n3659, A2 => n268, B1 => n3658, B2 => n271,
                           ZN => n2375);
   U2944 : AOI221_X1 port map( B1 => n274, B2 => n609, C1 => n277, C2 => n642, 
                           A => n2376, ZN => n2371);
   U2945 : OAI22_X1 port map( A1 => n1091, A2 => n280, B1 => n1092, B2 => n283,
                           ZN => n2376);
   U2946 : AOI221_X1 port map( B1 => n286, B2 => n575, C1 => n289, C2 => n3772,
                           A => n2377, ZN => n2370);
   U2947 : OAI22_X1 port map( A1 => n1094, A2 => n292, B1 => n1095, B2 => n295,
                           ZN => n2377);
   U2948 : OAI222_X1 port map( A1 => n300, A2 => n196, B1 => n2378, B2 => n199,
                           C1 => n2459, C2 => n202, ZN => n2985);
   U2949 : NOR4_X1 port map( A1 => n2379, A2 => n2380, A3 => n2381, A4 => n2382
                           , ZN => n2378);
   U2950 : OAI221_X1 port map( B1 => n3835, B2 => n205, C1 => n1051, C2 => n208
                           , A => n2383, ZN => n2382);
   U2951 : AOI22_X1 port map( A1 => n211, A2 => n3688, B1 => n214, B2 => n675, 
                           ZN => n2383);
   U2952 : OAI221_X1 port map( B1 => n1053, B2 => n217, C1 => n3739, C2 => n220
                           , A => n2384, ZN => n2381);
   U2953 : AOI22_X1 port map( A1 => n223, A2 => n777, B1 => n226, B2 => n3687, 
                           ZN => n2384);
   U2954 : OAI211_X1 port map( C1 => n3692, C2 => n229, A => n2385, B => n2386,
                           ZN => n2380);
   U2955 : AOI221_X1 port map( B1 => n232, B2 => n911, C1 => n235, C2 => n3693,
                           A => n2387, ZN => n2386);
   U2956 : OAI22_X1 port map( A1 => n3689, A2 => n238, B1 => n1058, B2 => n241,
                           ZN => n2387);
   U2957 : AOI22_X1 port map( A1 => n244, A2 => n3694, B1 => n247, B2 => n811, 
                           ZN => n2385);
   U2958 : NAND4_X1 port map( A1 => n2388, A2 => n2389, A3 => n2390, A4 => 
                           n2391, ZN => n2379);
   U2959 : AOI221_X1 port map( B1 => n250, B2 => n3677, C1 => n253, C2 => n3678
                           , A => n2392, ZN => n2391);
   U2960 : OAI22_X1 port map( A1 => n3676, A2 => n256, B1 => n3675, B2 => n259,
                           ZN => n2392);
   U2961 : AOI221_X1 port map( B1 => n262, B2 => n3681, C1 => n265, C2 => n3682
                           , A => n2393, ZN => n2390);
   U2962 : OAI22_X1 port map( A1 => n3680, A2 => n268, B1 => n3679, B2 => n271,
                           ZN => n2393);
   U2963 : AOI221_X1 port map( B1 => n274, B2 => n608, C1 => n277, C2 => n641, 
                           A => n2394, ZN => n2389);
   U2964 : OAI22_X1 port map( A1 => n1066, A2 => n280, B1 => n1067, B2 => n283,
                           ZN => n2394);
   U2965 : AOI221_X1 port map( B1 => n286, B2 => n574, C1 => n289, C2 => n3771,
                           A => n2395, ZN => n2388);
   U2966 : OAI22_X1 port map( A1 => n1069, A2 => n292, B1 => n1070, B2 => n295,
                           ZN => n2395);
   U2967 : OAI222_X1 port map( A1 => n299, A2 => n196, B1 => n2396, B2 => n199,
                           C1 => n2458, C2 => n202, ZN => n2984);
   U2968 : NOR4_X1 port map( A1 => n2397, A2 => n2398, A3 => n2399, A4 => n2400
                           , ZN => n2396);
   U2969 : OAI221_X1 port map( B1 => n3834, B2 => n205, C1 => n1026, C2 => n208
                           , A => n2401, ZN => n2400);
   U2970 : AOI22_X1 port map( A1 => n211, A2 => n3709, B1 => n214, B2 => n674, 
                           ZN => n2401);
   U2971 : OAI221_X1 port map( B1 => n1028, B2 => n217, C1 => n3738, C2 => n220
                           , A => n2402, ZN => n2399);
   U2972 : AOI22_X1 port map( A1 => n223, A2 => n776, B1 => n226, B2 => n3708, 
                           ZN => n2402);
   U2973 : OAI211_X1 port map( C1 => n3713, C2 => n229, A => n2403, B => n2404,
                           ZN => n2398);
   U2974 : AOI221_X1 port map( B1 => n232, B2 => n910, C1 => n235, C2 => n3714,
                           A => n2405, ZN => n2404);
   U2975 : OAI22_X1 port map( A1 => n3710, A2 => n238, B1 => n1033, B2 => n241,
                           ZN => n2405);
   U2976 : AOI22_X1 port map( A1 => n244, A2 => n3715, B1 => n247, B2 => n810, 
                           ZN => n2403);
   U2977 : NAND4_X1 port map( A1 => n2406, A2 => n2407, A3 => n2408, A4 => 
                           n2409, ZN => n2397);
   U2978 : AOI221_X1 port map( B1 => n250, B2 => n3698, C1 => n253, C2 => n3699
                           , A => n2410, ZN => n2409);
   U2979 : OAI22_X1 port map( A1 => n3697, A2 => n256, B1 => n3696, B2 => n259,
                           ZN => n2410);
   U2980 : AOI221_X1 port map( B1 => n262, B2 => n3702, C1 => n265, C2 => n3703
                           , A => n2411, ZN => n2408);
   U2981 : OAI22_X1 port map( A1 => n3701, A2 => n268, B1 => n3700, B2 => n271,
                           ZN => n2411);
   U2982 : AOI221_X1 port map( B1 => n274, B2 => n607, C1 => n277, C2 => n640, 
                           A => n2412, ZN => n2407);
   U2983 : OAI22_X1 port map( A1 => n1041, A2 => n280, B1 => n1042, B2 => n283,
                           ZN => n2412);
   U2984 : AOI221_X1 port map( B1 => n286, B2 => n573, C1 => n289, C2 => n3770,
                           A => n2413, ZN => n2406);
   U2985 : OAI22_X1 port map( A1 => n1044, A2 => n292, B1 => n1045, B2 => n295,
                           ZN => n2413);
   U2986 : OAI222_X1 port map( A1 => n298, A2 => n196, B1 => n2414, B2 => n199,
                           C1 => n2457, C2 => n202, ZN => n2983);
   U2987 : NAND2_X1 port map( A1 => n202, A2 => n2415, ZN => n1824);
   U2988 : NOR4_X1 port map( A1 => n2416, A2 => n2417, A3 => n2418, A4 => n2419
                           , ZN => n2414);
   U2989 : OAI221_X1 port map( B1 => n3833, B2 => n205, C1 => n971, C2 => n208,
                           A => n2420, ZN => n2419);
   U2990 : AOI22_X1 port map( A1 => n211, A2 => n3730, B1 => n214, B2 => n673, 
                           ZN => n2420);
   U2991 : AND2_X1 port map( A1 => n2421, A2 => n2422, ZN => n1834);
   U2992 : AND2_X1 port map( A1 => n2421, A2 => n2423, ZN => n1833);
   U2993 : NAND2_X1 port map( A1 => n2424, A2 => n2425, ZN => n1831);
   U2994 : NAND2_X1 port map( A1 => n2426, A2 => n2422, ZN => n1830);
   U2995 : OAI221_X1 port map( B1 => n976, B2 => n217, C1 => n3737, C2 => n220,
                           A => n2427, ZN => n2418);
   U2996 : AOI22_X1 port map( A1 => n223, A2 => n774, B1 => n226, B2 => n3729, 
                           ZN => n2427);
   U2997 : AND2_X1 port map( A1 => n2426, A2 => n2423, ZN => n1839);
   U2998 : AND2_X1 port map( A1 => n2426, A2 => n2425, ZN => n1838);
   U2999 : NAND2_X1 port map( A1 => n2421, A2 => n2425, ZN => n1836);
   U3000 : NAND2_X1 port map( A1 => n2421, A2 => n2428, ZN => n1835);
   U3001 : NOR3_X1 port map( A1 => n2429, A2 => ADD_RS1(0), A3 => n2430, ZN => 
                           n2421);
   U3002 : OAI211_X1 port map( C1 => n3734, C2 => n229, A => n2431, B => n2432,
                           ZN => n2417);
   U3003 : AOI221_X1 port map( B1 => n232, B2 => n908, C1 => n235, C2 => n3735,
                           A => n2433, ZN => n2432);
   U3004 : OAI22_X1 port map( A1 => n3731, A2 => n238, B1 => n989, B2 => n241, 
                           ZN => n2433);
   U3005 : NAND2_X1 port map( A1 => n2434, A2 => n2425, ZN => n1847);
   U3006 : NAND2_X1 port map( A1 => n2434, A2 => n2428, ZN => n1846);
   U3007 : AND2_X1 port map( A1 => n2424, A2 => n2422, ZN => n1844);
   U3008 : AND2_X1 port map( A1 => n2424, A2 => n2428, ZN => n1843);
   U3009 : AOI22_X1 port map( A1 => n244, A2 => n3736, B1 => n247, B2 => n808, 
                           ZN => n2431);
   U3010 : AND2_X1 port map( A1 => n2434, A2 => n2423, ZN => n1849);
   U3011 : AND2_X1 port map( A1 => n2434, A2 => n2422, ZN => n1848);
   U3012 : NOR3_X1 port map( A1 => ADD_RS1(0), A2 => ADD_RS1(3), A3 => n2429, 
                           ZN => n2434);
   U3013 : NAND2_X1 port map( A1 => n2424, A2 => n2423, ZN => n1840);
   U3014 : NOR3_X1 port map( A1 => n2435, A2 => ADD_RS1(3), A3 => n2429, ZN => 
                           n2424);
   U3015 : NAND4_X1 port map( A1 => n2436, A2 => n2437, A3 => n2438, A4 => 
                           n2439, ZN => n2416);
   U3016 : AOI221_X1 port map( B1 => n250, B2 => n3719, C1 => n253, C2 => n3720
                           , A => n2440, ZN => n2439);
   U3017 : OAI22_X1 port map( A1 => n3718, A2 => n256, B1 => n3717, B2 => n259,
                           ZN => n2440);
   U3018 : NAND2_X1 port map( A1 => n2428, A2 => n2441, ZN => n1858);
   U3019 : NAND2_X1 port map( A1 => n2428, A2 => n2442, ZN => n1857);
   U3020 : AND2_X1 port map( A1 => n2441, A2 => n2425, ZN => n1855);
   U3021 : AND2_X1 port map( A1 => n2425, A2 => n2442, ZN => n1854);
   U3022 : AOI221_X1 port map( B1 => n262, B2 => n3723, C1 => n265, C2 => n3724
                           , A => n2443, ZN => n2438);
   U3023 : OAI22_X1 port map( A1 => n3722, A2 => n268, B1 => n3721, B2 => n271,
                           ZN => n2443);
   U3024 : NAND2_X1 port map( A1 => n2423, A2 => n2441, ZN => n1863);
   U3025 : NAND2_X1 port map( A1 => n2423, A2 => n2442, ZN => n1862);
   U3026 : AND2_X1 port map( A1 => n2422, A2 => n2441, ZN => n1860);
   U3027 : NOR3_X1 port map( A1 => ADD_RS1(0), A2 => ADD_RS1(4), A3 => n2430, 
                           ZN => n2441);
   U3028 : AND2_X1 port map( A1 => n2422, A2 => n2442, ZN => n1859);
   U3029 : NOR3_X1 port map( A1 => n2435, A2 => ADD_RS1(4), A3 => n2430, ZN => 
                           n2442);
   U3030 : AOI221_X1 port map( B1 => n274, B2 => n605, C1 => n277, C2 => n638, 
                           A => n2444, ZN => n2437);
   U3031 : OAI22_X1 port map( A1 => n1010, A2 => n280, B1 => n1012, B2 => n283,
                           ZN => n2444);
   U3032 : NAND2_X1 port map( A1 => n2445, A2 => n2425, ZN => n1868);
   U3033 : NAND2_X1 port map( A1 => n2446, A2 => n2425, ZN => n1867);
   U3034 : NOR2_X1 port map( A1 => n2447, A2 => n2448, ZN => n2425);
   U3035 : AND2_X1 port map( A1 => n2445, A2 => n2428, ZN => n1865);
   U3036 : AND2_X1 port map( A1 => n2446, A2 => n2428, ZN => n1864);
   U3037 : AOI221_X1 port map( B1 => n286, B2 => n571, C1 => n289, C2 => n3769,
                           A => n2449, ZN => n2436);
   U3038 : OAI22_X1 port map( A1 => n1017, A2 => n292, B1 => n1019, B2 => n295,
                           ZN => n2449);
   U3039 : NAND2_X1 port map( A1 => n2445, A2 => n2422, ZN => n1873);
   U3040 : NAND2_X1 port map( A1 => n2446, A2 => n2422, ZN => n1872);
   U3041 : NOR2_X1 port map( A1 => n2448, A2 => ADD_RS1(2), ZN => n2422);
   U3042 : NOR3_X1 port map( A1 => ADD_RS1(3), A2 => ADD_RS1(4), A3 => 
                           ADD_RS1(0), ZN => n2446);
   U3043 : AND2_X1 port map( A1 => n2426, A2 => n2428, ZN => n1870);
   U3044 : NOR2_X1 port map( A1 => n2447, A2 => ADD_RS1(1), ZN => n2428);
   U3045 : INV_X1 port map( A => ADD_RS1(2), ZN => n2447);
   U3046 : NOR3_X1 port map( A1 => n2429, A2 => n2435, A3 => n2430, ZN => n2426
                           );
   U3047 : INV_X1 port map( A => ADD_RS1(3), ZN => n2430);
   U3048 : INV_X1 port map( A => ADD_RS1(4), ZN => n2429);
   U3049 : AND2_X1 port map( A1 => n2445, A2 => n2423, ZN => n1869);
   U3050 : NOR2_X1 port map( A1 => ADD_RS1(1), A2 => ADD_RS1(2), ZN => n2423);
   U3051 : NOR3_X1 port map( A1 => ADD_RS1(3), A2 => ADD_RS1(4), A3 => n2435, 
                           ZN => n2445);
   U3052 : INV_X1 port map( A => ADD_RS1(0), ZN => n2435);
   U3053 : NAND2_X1 port map( A1 => n2450, A2 => n202, ZN => n1822);
   U3054 : AND3_X1 port map( A1 => n419, A2 => ENABLE, A3 => RD1, ZN => n1825);
   U3055 : INV_X1 port map( A => n2415, ZN => n2450);
   U3056 : NAND4_X1 port map( A1 => n2451, A2 => n2452, A3 => n2453, A4 => 
                           n2454, ZN => n2415);
   U3057 : NOR3_X1 port map( A1 => n2455, A2 => n1820, A3 => n2456, ZN => n2454
                           );
   U3058 : XNOR2_X1 port map( A => ADD_WR(1), B => n2448, ZN => n2456);
   U3059 : INV_X1 port map( A => ADD_RS1(1), ZN => n2448);
   U3060 : INV_X1 port map( A => WR, ZN => n1820);
   U3061 : XNOR2_X1 port map( A => n953, B => ADD_RS1(0), ZN => n2455);
   U3062 : INV_X1 port map( A => ADD_WR(0), ZN => n953);
   U3063 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS1(3), ZN => n2453);
   U3064 : XNOR2_X1 port map( A => ADD_WR(4), B => ADD_RS1(4), ZN => n2452);
   U3065 : XNOR2_X1 port map( A => ADD_RS1(2), B => ADD_WR(2), ZN => n2451);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_0 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_0;

architecture SYN_bhv of regn_N5_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15 : 
      std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n15, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n10);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n14, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n9);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n13, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n8);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n12, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n7);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n11, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n6);
   U2 : OAI21_X1 port map( B1 => n6, B2 => EN, A => n1, ZN => n11);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n1);
   U4 : OAI21_X1 port map( B1 => n7, B2 => EN, A => n2, ZN => n12);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n8, B2 => EN, A => n3, ZN => n13);
   U7 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n9, B2 => EN, A => n4, ZN => n14);
   U9 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n4);
   U10 : OAI21_X1 port map( B1 => n10, B2 => EN, A => n5, ZN => n15);
   U11 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n5);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity instruction_decomposition is

   port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype : in
         std_logic;  ADD_RS1, ADD_RS2, ADD_WR : out std_logic_vector (4 downto 
         0);  IMM : out std_logic_vector (31 downto 0));

end instruction_decomposition;

architecture SYN_bhv of instruction_decomposition is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal IMM_24_port, IMM_23_port, IMM_22_port, IMM_21_port, IMM_20_port, 
      IMM_19_port, IMM_18_port, IMM_17_port, IMM_16_port, IMM_15_port, 
      IMM_14_port, IMM_13_port, IMM_12_port, IMM_11_port, IMM_10_port, 
      IMM_9_port, IMM_8_port, IMM_7_port, IMM_6_port, IMM_5_port, IMM_4_port, 
      IMM_3_port, IMM_2_port, IMM_1_port, IMM_0_port, n21, n22, n23, n24, n25, 
      n26, n27, n28, n29, n30, n31, n32, n1, n2, IMM_31_port, n4, n5, n6, n7, 
      n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20 : std_logic
      ;

begin
   IMM <= ( IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, 
      IMM_31_port, IMM_31_port, IMM_24_port, IMM_23_port, IMM_22_port, 
      IMM_21_port, IMM_20_port, IMM_19_port, IMM_18_port, IMM_17_port, 
      IMM_16_port, IMM_15_port, IMM_14_port, IMM_13_port, IMM_12_port, 
      IMM_11_port, IMM_10_port, IMM_9_port, IMM_8_port, IMM_7_port, IMM_6_port,
      IMM_5_port, IMM_4_port, IMM_3_port, IMM_2_port, IMM_1_port, IMM_0_port );
   
   U72 : NAND3_X1 port map( A1 => INST_IN(29), A2 => INST_IN(27), A3 => 
                           INST_IN(31), ZN => n31);
   U73 : NAND3_X1 port map( A1 => INST_IN(26), A2 => Itype, A3 => n32, ZN => 
                           n30);
   U2 : INV_X1 port map( A => Rtype, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n28, A2 => Jtype, ZN => n24);
   U4 : INV_X1 port map( A => n27, ZN => n2);
   U5 : OAI21_X1 port map( B1 => Itype, B2 => Jtype, A => n4, ZN => n27);
   U6 : NOR2_X1 port map( A1 => Rtype, A2 => Itype, ZN => n28);
   U7 : NOR2_X1 port map( A1 => n28, A2 => n10, ZN => ADD_RS1(0));
   U8 : NOR2_X1 port map( A1 => n1, A2 => n15, ZN => ADD_RS2(0));
   U9 : NOR2_X1 port map( A1 => n28, A2 => n7, ZN => ADD_RS1(3));
   U10 : NOR2_X1 port map( A1 => n1, A2 => n12, ZN => ADD_RS2(3));
   U11 : NOR2_X1 port map( A1 => n1, A2 => n11, ZN => ADD_RS2(4));
   U12 : NOR2_X1 port map( A1 => n28, A2 => n8, ZN => ADD_RS1(2));
   U13 : NOR2_X1 port map( A1 => n1, A2 => n13, ZN => ADD_RS2(2));
   U14 : OR2_X1 port map( A1 => n26, A2 => n16, ZN => n25);
   U15 : NOR2_X1 port map( A1 => n28, A2 => n9, ZN => ADD_RS1(1));
   U16 : NOR2_X1 port map( A1 => n1, A2 => n14, ZN => ADD_RS2(1));
   U17 : NAND2_X1 port map( A1 => Itype, A2 => n4, ZN => n26);
   U18 : INV_X1 port map( A => Itype, ZN => n5);
   U19 : AND2_X1 port map( A1 => INST_IN(0), A2 => n2, ZN => IMM_0_port);
   U20 : AND2_X1 port map( A1 => INST_IN(1), A2 => n2, ZN => IMM_1_port);
   U21 : AND2_X1 port map( A1 => INST_IN(2), A2 => n2, ZN => IMM_2_port);
   U22 : AND2_X1 port map( A1 => INST_IN(3), A2 => n2, ZN => IMM_3_port);
   U23 : AND2_X1 port map( A1 => INST_IN(4), A2 => n2, ZN => IMM_4_port);
   U24 : AND2_X1 port map( A1 => INST_IN(5), A2 => n2, ZN => IMM_5_port);
   U25 : AND2_X1 port map( A1 => INST_IN(6), A2 => n2, ZN => IMM_6_port);
   U26 : AND2_X1 port map( A1 => INST_IN(7), A2 => n2, ZN => IMM_7_port);
   U27 : AND2_X1 port map( A1 => INST_IN(8), A2 => n2, ZN => IMM_8_port);
   U28 : AND2_X1 port map( A1 => INST_IN(9), A2 => n2, ZN => IMM_9_port);
   U29 : AND2_X1 port map( A1 => INST_IN(10), A2 => n2, ZN => IMM_10_port);
   U30 : NOR2_X1 port map( A1 => n27, A2 => n20, ZN => IMM_11_port);
   U31 : NOR2_X1 port map( A1 => n27, A2 => n19, ZN => IMM_12_port);
   U32 : NOR2_X1 port map( A1 => n27, A2 => n18, ZN => IMM_13_port);
   U33 : NOR2_X1 port map( A1 => n27, A2 => n17, ZN => IMM_14_port);
   U34 : NOR2_X1 port map( A1 => n27, A2 => n16, ZN => IMM_15_port);
   U35 : OAI21_X1 port map( B1 => n24, B2 => n15, A => n25, ZN => IMM_16_port);
   U36 : OAI21_X1 port map( B1 => n24, B2 => n14, A => n25, ZN => IMM_17_port);
   U37 : OAI21_X1 port map( B1 => n24, B2 => n13, A => n25, ZN => IMM_18_port);
   U38 : OAI21_X1 port map( B1 => n24, B2 => n12, A => n25, ZN => IMM_19_port);
   U39 : OAI21_X1 port map( B1 => n24, B2 => n11, A => n25, ZN => IMM_20_port);
   U40 : OAI21_X1 port map( B1 => n24, B2 => n10, A => n25, ZN => IMM_21_port);
   U41 : OAI21_X1 port map( B1 => n24, B2 => n9, A => n25, ZN => IMM_22_port);
   U42 : OAI21_X1 port map( B1 => n24, B2 => n8, A => n25, ZN => IMM_23_port);
   U43 : OAI21_X1 port map( B1 => n24, B2 => n7, A => n25, ZN => IMM_24_port);
   U44 : OAI221_X1 port map( B1 => n26, B2 => n15, C1 => n20, C2 => n4, A => 
                           n24, ZN => ADD_WR(0));
   U45 : OAI221_X1 port map( B1 => n26, B2 => n14, C1 => n19, C2 => n4, A => 
                           n24, ZN => ADD_WR(1));
   U46 : OAI221_X1 port map( B1 => n26, B2 => n13, C1 => n18, C2 => n4, A => 
                           n24, ZN => ADD_WR(2));
   U47 : OAI221_X1 port map( B1 => n26, B2 => n12, C1 => n17, C2 => n4, A => 
                           n24, ZN => ADD_WR(3));
   U48 : OAI221_X1 port map( B1 => n26, B2 => n11, C1 => n16, C2 => n4, A => 
                           n24, ZN => ADD_WR(4));
   U49 : NOR2_X1 port map( A1 => n28, A2 => n6, ZN => ADD_RS1(4));
   U50 : INV_X1 port map( A => INST_IN(25), ZN => n6);
   U51 : INV_X1 port map( A => n21, ZN => IMM_31_port);
   U52 : OAI21_X1 port map( B1 => n22, B2 => n23, A => n4, ZN => n21);
   U53 : AND3_X1 port map( A1 => Jtype, A2 => n5, A3 => INST_IN(25), ZN => n22)
                           ;
   U54 : NOR2_X1 port map( A1 => n16, A2 => n5, ZN => n23);
   U55 : INV_X1 port map( A => n29, ZN => n1);
   U56 : OAI21_X1 port map( B1 => n30, B2 => n31, A => n4, ZN => n29);
   U57 : INV_X1 port map( A => INST_IN(15), ZN => n16);
   U58 : INV_X1 port map( A => INST_IN(16), ZN => n15);
   U59 : INV_X1 port map( A => INST_IN(17), ZN => n14);
   U60 : INV_X1 port map( A => INST_IN(19), ZN => n12);
   U61 : INV_X1 port map( A => INST_IN(18), ZN => n13);
   U62 : INV_X1 port map( A => INST_IN(20), ZN => n11);
   U63 : NOR2_X1 port map( A1 => INST_IN(30), A2 => INST_IN(28), ZN => n32);
   U64 : INV_X1 port map( A => INST_IN(21), ZN => n10);
   U65 : INV_X1 port map( A => INST_IN(22), ZN => n9);
   U66 : INV_X1 port map( A => INST_IN(24), ZN => n7);
   U67 : INV_X1 port map( A => INST_IN(23), ZN => n8);
   U68 : INV_X1 port map( A => INST_IN(11), ZN => n20);
   U69 : INV_X1 port map( A => INST_IN(12), ZN => n19);
   U70 : INV_X1 port map( A => INST_IN(13), ZN => n18);
   U71 : INV_X1 port map( A => INST_IN(14), ZN => n17);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity instruction_type is

   port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype : 
         out std_logic);

end instruction_type;

architecture SYN_bhv of instruction_type is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n1, n2, n3, n4, n5, 
      n6, n7, n8 : std_logic;

begin
   
   U21 : OAI33_X1 port map( A1 => n5, A2 => INST_IN(29), A3 => n2, B1 => n4, B2
                           => INST_IN(30), B3 => INST_IN(26), ZN => n17);
   U1 : NOR2_X1 port map( A1 => n9, A2 => n10, ZN => Rtype);
   U2 : OAI22_X1 port map( A1 => n10, A2 => n5, B1 => n7, B2 => n4, ZN => n16);
   U3 : NOR2_X1 port map( A1 => n9, A2 => n6, ZN => Jtype);
   U4 : NAND4_X1 port map( A1 => n5, A2 => n4, A3 => n3, A4 => n1, ZN => n9);
   U5 : NAND2_X1 port map( A1 => n6, A2 => n8, ZN => n10);
   U6 : INV_X1 port map( A => n14, ZN => n7);
   U7 : INV_X1 port map( A => n18, ZN => n2);
   U8 : OAI221_X1 port map( B1 => n7, B2 => INST_IN(30), C1 => n3, C2 => 
                           INST_IN(26), A => n10, ZN => n18);
   U9 : OAI211_X1 port map( C1 => INST_IN(31), C2 => n11, A => n12, B => n13, 
                           ZN => Itype);
   U10 : NAND4_X1 port map( A1 => INST_IN(29), A2 => INST_IN(28), A3 => n14, A4
                           => n1, ZN => n13);
   U11 : NAND4_X1 port map( A1 => INST_IN(31), A2 => INST_IN(27), A3 => n15, A4
                           => INST_IN(26), ZN => n12);
   U12 : AOI21_X1 port map( B1 => INST_IN(30), B2 => n16, A => n17, ZN => n11);
   U13 : NOR2_X1 port map( A1 => n8, A2 => INST_IN(27), ZN => n14);
   U14 : NOR2_X1 port map( A1 => INST_IN(30), A2 => INST_IN(28), ZN => n15);
   U15 : INV_X1 port map( A => INST_IN(30), ZN => n3);
   U16 : INV_X1 port map( A => INST_IN(28), ZN => n5);
   U17 : INV_X1 port map( A => INST_IN(29), ZN => n4);
   U18 : INV_X1 port map( A => INST_IN(26), ZN => n8);
   U19 : INV_X1 port map( A => INST_IN(31), ZN => n1);
   U20 : INV_X1 port map( A => INST_IN(27), ZN => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_0 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_0;

architecture SYN_bhv of regn_N32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, DOUT_27_port,
      DOUT_26_port, DOUT_24_port, DOUT_23_port, DOUT_22_port, DOUT_21_port, 
      DOUT_20_port, DOUT_18_port, DOUT_17_port, DOUT_16_port, DOUT_14_port, 
      DOUT_13_port, DOUT_12_port, n51, n52, DOUT_7_port, DOUT_6_port, 
      DOUT_5_port, DOUT_4_port, DOUT_3_port, DOUT_2_port, DOUT_1_port, 
      DOUT_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n53, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n9, DOUT_19_port, n11, n12
      , n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, 
      n27, n28, n29, n30, n31, n32, DOUT_8_port, DOUT_9_port, DOUT_10_port, 
      DOUT_11_port, DOUT_15_port, n49, DOUT_25_port, n_1922, n_1923, n_1924, 
      n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, 
      n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941 : 
      std_logic;

begin
   DOUT <= ( DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, 
      DOUT_27_port, DOUT_26_port, DOUT_25_port, DOUT_24_port, DOUT_23_port, 
      DOUT_22_port, DOUT_21_port, DOUT_20_port, DOUT_19_port, DOUT_18_port, 
      DOUT_17_port, DOUT_16_port, DOUT_15_port, DOUT_14_port, DOUT_13_port, 
      DOUT_12_port, DOUT_11_port, DOUT_10_port, DOUT_9_port, DOUT_8_port, 
      DOUT_7_port, DOUT_6_port, DOUT_5_port, DOUT_4_port, DOUT_3_port, 
      DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n96, CK => CLK, RN => n32, Q => 
                           DOUT_31_port, QN => n_1922);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n95, CK => CLK, RN => n32, Q => 
                           DOUT_30_port, QN => n_1923);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n94, CK => CLK, RN => n32, Q => 
                           DOUT_29_port, QN => n_1924);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n93, CK => CLK, RN => n32, Q => 
                           DOUT_28_port, QN => n_1925);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n92, CK => CLK, RN => n32, Q => 
                           DOUT_27_port, QN => n_1926);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n91, CK => CLK, RN => n32, Q => 
                           DOUT_26_port, QN => n_1927);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n90, CK => CLK, RN => n32, Q => 
                           DOUT_25_port, QN => n_1928);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n89, CK => CLK, RN => n32, Q => 
                           DOUT_24_port, QN => n_1929);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n88, CK => CLK, RN => n31, Q => 
                           DOUT_23_port, QN => n_1930);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n87, CK => CLK, RN => n31, Q => 
                           DOUT_22_port, QN => n_1931);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n86, CK => CLK, RN => n31, Q => 
                           DOUT_21_port, QN => n_1932);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n85, CK => CLK, RN => n31, Q => 
                           DOUT_20_port, QN => n53);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n83, CK => CLK, RN => n31, Q => 
                           DOUT_18_port, QN => n_1933);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n82, CK => CLK, RN => n31, Q => 
                           DOUT_17_port, QN => n_1934);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n81, CK => CLK, RN => n31, Q => 
                           DOUT_16_port, QN => n_1935);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n80, CK => CLK, RN => n31, Q => 
                           DOUT_15_port, QN => n_1936);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n79, CK => CLK, RN => n31, Q => 
                           DOUT_14_port, QN => n_1937);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n78, CK => CLK, RN => n31, Q => 
                           DOUT_13_port, QN => n_1938);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n77, CK => CLK, RN => n31, Q => 
                           DOUT_12_port, QN => n_1939);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n76, CK => CLK, RN => n30, Q => 
                           DOUT_11_port, QN => n_1940);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n75, CK => CLK, RN => n30, Q => n9
                           , QN => n43);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n74, CK => CLK, RN => n30, Q => n51
                           , QN => n42);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n73, CK => CLK, RN => n30, Q => n52
                           , QN => n41);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n72, CK => CLK, RN => n30, Q => 
                           DOUT_7_port, QN => n40);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n71, CK => CLK, RN => n30, Q => 
                           DOUT_6_port, QN => n39);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n70, CK => CLK, RN => n30, Q => 
                           DOUT_5_port, QN => n38);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n69, CK => CLK, RN => n30, Q => 
                           DOUT_4_port, QN => n37);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n68, CK => CLK, RN => n30, Q => 
                           DOUT_3_port, QN => n36);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n67, CK => CLK, RN => n30, Q => 
                           DOUT_2_port, QN => n35);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n66, CK => CLK, RN => n30, Q => 
                           DOUT_1_port, QN => n34);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n65, CK => CLK, RN => n30, Q => 
                           DOUT_0_port, QN => n33);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n84, CK => CLK, RN => n31, Q => 
                           DOUT_19_port, QN => n_1941);
   U2 : INV_X1 port map( A => EN, ZN => n11);
   U3 : INV_X1 port map( A => n43, ZN => DOUT_10_port);
   U4 : MUX2_X1 port map( A => DIN(28), B => DOUT_28_port, S => n11, Z => n93);
   U5 : MUX2_X1 port map( A => DIN(25), B => DOUT_25_port, S => n11, Z => n90);
   U6 : NAND2_X1 port map( A1 => DOUT_15_port, A2 => n12, ZN => n13);
   U7 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n14);
   U8 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => n80);
   U9 : INV_X1 port map( A => EN, ZN => n12);
   U10 : BUF_X1 port map( A => RST, Z => n30);
   U11 : BUF_X1 port map( A => RST, Z => n31);
   U12 : BUF_X1 port map( A => RST, Z => n32);
   U13 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n8);
   U14 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n7);
   U15 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n6);
   U16 : OAI21_X1 port map( B1 => n35, B2 => EN, A => n3, ZN => n67);
   U17 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n3);
   U18 : OAI21_X1 port map( B1 => n34, B2 => EN, A => n2, ZN => n66);
   U19 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n2);
   U20 : OAI21_X1 port map( B1 => n33, B2 => EN, A => n1, ZN => n65);
   U21 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n1);
   U22 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n4);
   U23 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n5);
   U24 : INV_X1 port map( A => EN, ZN => n27);
   U25 : INV_X1 port map( A => EN, ZN => n18);
   U26 : INV_X1 port map( A => EN, ZN => n21);
   U27 : OAI21_X1 port map( B1 => n37, B2 => EN, A => n5, ZN => n69);
   U28 : OAI21_X1 port map( B1 => n38, B2 => EN, A => n6, ZN => n70);
   U29 : OAI21_X1 port map( B1 => n40, B2 => EN, A => n8, ZN => n72);
   U30 : NAND2_X1 port map( A1 => DIN(29), A2 => n15, ZN => n16);
   U31 : NAND2_X1 port map( A1 => DOUT_29_port, A2 => n18, ZN => n17);
   U32 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => n94);
   U33 : INV_X1 port map( A => n18, ZN => n15);
   U34 : OAI21_X1 port map( B1 => n39, B2 => EN, A => n7, ZN => n71);
   U35 : NAND2_X1 port map( A1 => DIN(31), A2 => n24, ZN => n19);
   U36 : NAND2_X1 port map( A1 => DOUT_31_port, A2 => n21, ZN => n20);
   U37 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => n96);
   U38 : OAI21_X1 port map( B1 => n36, B2 => EN, A => n4, ZN => n68);
   U39 : NAND2_X1 port map( A1 => DIN(27), A2 => n15, ZN => n22);
   U40 : NAND2_X1 port map( A1 => DOUT_27_port, A2 => n12, ZN => n23);
   U41 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => n92);
   U42 : NAND2_X1 port map( A1 => DIN(23), A2 => n24, ZN => n25);
   U43 : NAND2_X1 port map( A1 => DOUT_23_port, A2 => n27, ZN => n26);
   U44 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => n88);
   U45 : INV_X1 port map( A => n27, ZN => n24);
   U46 : NAND2_X1 port map( A1 => DIN(19), A2 => n24, ZN => n28);
   U47 : NAND2_X1 port map( A1 => DOUT_19_port, A2 => n12, ZN => n29);
   U48 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => n84);
   U49 : INV_X1 port map( A => n41, ZN => DOUT_8_port);
   U50 : MUX2_X1 port map( A => n52, B => DIN(8), S => EN, Z => n73);
   U51 : INV_X1 port map( A => n42, ZN => DOUT_9_port);
   U52 : MUX2_X1 port map( A => n51, B => DIN(9), S => EN, Z => n74);
   U53 : MUX2_X1 port map( A => n9, B => DIN(10), S => EN, Z => n75);
   U54 : MUX2_X1 port map( A => DOUT_11_port, B => DIN(11), S => EN, Z => n76);
   U55 : MUX2_X1 port map( A => DOUT_12_port, B => DIN(12), S => EN, Z => n77);
   U56 : MUX2_X1 port map( A => DOUT_13_port, B => DIN(13), S => EN, Z => n78);
   U57 : MUX2_X1 port map( A => DOUT_14_port, B => DIN(14), S => EN, Z => n79);
   U58 : MUX2_X1 port map( A => DOUT_16_port, B => DIN(16), S => EN, Z => n81);
   U59 : MUX2_X1 port map( A => DOUT_17_port, B => DIN(17), S => EN, Z => n82);
   U60 : MUX2_X1 port map( A => DOUT_18_port, B => DIN(18), S => EN, Z => n83);
   U61 : INV_X1 port map( A => n53, ZN => n49);
   U62 : MUX2_X1 port map( A => n49, B => DIN(20), S => EN, Z => n85);
   U63 : MUX2_X1 port map( A => DOUT_21_port, B => DIN(21), S => EN, Z => n86);
   U64 : MUX2_X1 port map( A => DOUT_22_port, B => DIN(22), S => EN, Z => n87);
   U65 : MUX2_X1 port map( A => DOUT_24_port, B => DIN(24), S => EN, Z => n89);
   U66 : MUX2_X1 port map( A => DOUT_26_port, B => DIN(26), S => EN, Z => n91);
   U67 : MUX2_X1 port map( A => DOUT_30_port, B => DIN(30), S => EN, Z => n95);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_0;

architecture SYN_bhv of mux21_NBIT32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n43, n54, n65, n1, n2, n3, n4, n5, n6, n7, 
      n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B(19), A2 => n16, ZN => n5);
   U2 : NAND2_X1 port map( A1 => B(15), A2 => n16, ZN => n8);
   U3 : INV_X1 port map( A => n17, ZN => n16);
   U4 : INV_X1 port map( A => n19, ZN => n15);
   U5 : NAND2_X1 port map( A1 => A(23), A2 => n19, ZN => n9);
   U6 : NAND2_X1 port map( A1 => A(31), A2 => n18, ZN => n1);
   U7 : NAND2_X1 port map( A1 => B(31), A2 => n15, ZN => n2);
   U8 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => Z(31));
   U9 : NAND2_X1 port map( A1 => B(23), A2 => n16, ZN => n10);
   U10 : NAND2_X1 port map( A1 => A(19), A2 => n3, ZN => n4);
   U11 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Z(19));
   U12 : INV_X1 port map( A => n16, ZN => n3);
   U13 : NAND2_X1 port map( A1 => A(15), A2 => n6, ZN => n7);
   U14 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => Z(15));
   U15 : INV_X1 port map( A => n16, ZN => n6);
   U16 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Z(23));
   U17 : AOI22_X1 port map( A1 => A(7), A2 => n19, B1 => B(7), B2 => n15, ZN =>
                           n36);
   U18 : INV_X1 port map( A => n37, ZN => Z(6));
   U19 : AOI22_X1 port map( A1 => A(6), A2 => n19, B1 => B(6), B2 => n15, ZN =>
                           n37);
   U20 : INV_X1 port map( A => n38, ZN => Z(5));
   U21 : AOI22_X1 port map( A1 => A(5), A2 => n18, B1 => B(5), B2 => n15, ZN =>
                           n38);
   U22 : INV_X1 port map( A => n43, ZN => Z(2));
   U23 : AOI22_X1 port map( A1 => A(2), A2 => n17, B1 => B(2), B2 => n15, ZN =>
                           n43);
   U24 : INV_X1 port map( A => n54, ZN => Z(1));
   U25 : AOI22_X1 port map( A1 => A(1), A2 => n18, B1 => B(1), B2 => n15, ZN =>
                           n54);
   U26 : INV_X1 port map( A => n65, ZN => Z(0));
   U27 : AOI22_X1 port map( A1 => A(0), A2 => n19, B1 => B(0), B2 => n15, ZN =>
                           n65);
   U28 : INV_X1 port map( A => n40, ZN => Z(3));
   U29 : AOI22_X1 port map( A1 => A(3), A2 => n17, B1 => B(3), B2 => n15, ZN =>
                           n40);
   U30 : INV_X1 port map( A => n39, ZN => Z(4));
   U31 : AOI22_X1 port map( A1 => A(4), A2 => n18, B1 => B(4), B2 => n15, ZN =>
                           n39);
   U32 : NAND2_X1 port map( A1 => A(27), A2 => n18, ZN => n11);
   U33 : NAND2_X1 port map( A1 => B(27), A2 => n15, ZN => n12);
   U34 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => Z(27));
   U35 : NAND2_X1 port map( A1 => A(25), A2 => n17, ZN => n13);
   U36 : NAND2_X1 port map( A1 => B(25), A2 => n16, ZN => n14);
   U37 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => Z(25));
   U38 : INV_X1 port map( A => n36, ZN => Z(7));
   U39 : INV_X1 port map( A => S, ZN => n17);
   U40 : INV_X1 port map( A => S, ZN => n18);
   U41 : INV_X1 port map( A => S, ZN => n19);
   U42 : MUX2_X1 port map( A => A(8), B => B(8), S => n16, Z => Z(8));
   U43 : MUX2_X1 port map( A => A(9), B => B(9), S => n16, Z => Z(9));
   U44 : MUX2_X1 port map( A => A(10), B => B(10), S => n16, Z => Z(10));
   U45 : MUX2_X1 port map( A => A(11), B => B(11), S => n16, Z => Z(11));
   U46 : MUX2_X1 port map( A => A(12), B => B(12), S => n16, Z => Z(12));
   U47 : MUX2_X1 port map( A => A(13), B => B(13), S => n16, Z => Z(13));
   U48 : MUX2_X1 port map( A => A(14), B => B(14), S => n16, Z => Z(14));
   U49 : MUX2_X1 port map( A => A(16), B => B(16), S => n16, Z => Z(16));
   U50 : MUX2_X1 port map( A => A(17), B => B(17), S => n16, Z => Z(17));
   U51 : MUX2_X1 port map( A => A(18), B => B(18), S => n16, Z => Z(18));
   U52 : MUX2_X1 port map( A => A(20), B => B(20), S => n16, Z => Z(20));
   U53 : MUX2_X1 port map( A => A(21), B => B(21), S => n16, Z => Z(21));
   U54 : MUX2_X1 port map( A => A(22), B => B(22), S => n16, Z => Z(22));
   U55 : MUX2_X1 port map( A => A(24), B => B(24), S => n16, Z => Z(24));
   U56 : MUX2_X1 port map( A => A(26), B => B(26), S => n15, Z => Z(26));
   U57 : MUX2_X1 port map( A => A(28), B => B(28), S => n15, Z => Z(28));
   U58 : MUX2_X1 port map( A => A(29), B => B(29), S => n15, Z => Z(29));
   U59 : MUX2_X1 port map( A => A(30), B => B(30), S => n15, Z => Z(30));

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HazardDetection is

   port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : in std_logic_vector (4
         downto 0);  DRAM_R : in std_logic;  INS_IN, PC_IN : in 
         std_logic_vector (31 downto 0);  Bubble : out std_logic;  HDU_INS_OUT,
         HDU_PC_OUT, HDU_NPC_OUT : out std_logic_vector (31 downto 0));

end HazardDetection;

architecture SYN_arch of HazardDetection is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component HazardDetection_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n7, n8, n11, n1, n2, n3, n4, n5, n6, n9, n10, n12, n13, n14, n15, n16
      , n_1942 : std_logic;

begin
   HDU_INS_OUT <= ( INS_IN(31), INS_IN(30), INS_IN(29), INS_IN(28), INS_IN(27),
      INS_IN(26), INS_IN(25), INS_IN(24), INS_IN(23), INS_IN(22), INS_IN(21), 
      INS_IN(20), INS_IN(19), INS_IN(18), INS_IN(17), INS_IN(16), INS_IN(15), 
      INS_IN(14), INS_IN(13), INS_IN(12), INS_IN(11), INS_IN(10), INS_IN(9), 
      INS_IN(8), INS_IN(7), INS_IN(6), INS_IN(5), INS_IN(4), INS_IN(3), 
      INS_IN(2), INS_IN(1), INS_IN(0) );
   HDU_NPC_OUT <= ( PC_IN(31), PC_IN(30), PC_IN(29), PC_IN(28), PC_IN(27), 
      PC_IN(26), PC_IN(25), PC_IN(24), PC_IN(23), PC_IN(22), PC_IN(21), 
      PC_IN(20), PC_IN(19), PC_IN(18), PC_IN(17), PC_IN(16), PC_IN(15), 
      PC_IN(14), PC_IN(13), PC_IN(12), PC_IN(11), PC_IN(10), PC_IN(9), PC_IN(8)
      , PC_IN(7), PC_IN(6), PC_IN(5), PC_IN(4), PC_IN(3), PC_IN(2), PC_IN(1), 
      PC_IN(0) );
   
   n7 <= '0';
   n8 <= '1';
   n11 <= '0';
   sub_25 : HazardDetection_DW01_sub_0 port map( A(31) => PC_IN(31), A(30) => 
                           PC_IN(30), A(29) => PC_IN(29), A(28) => PC_IN(28), 
                           A(27) => PC_IN(27), A(26) => PC_IN(26), A(25) => 
                           PC_IN(25), A(24) => PC_IN(24), A(23) => PC_IN(23), 
                           A(22) => PC_IN(22), A(21) => PC_IN(21), A(20) => 
                           PC_IN(20), A(19) => PC_IN(19), A(18) => PC_IN(18), 
                           A(17) => PC_IN(17), A(16) => PC_IN(16), A(15) => 
                           PC_IN(15), A(14) => PC_IN(14), A(13) => PC_IN(13), 
                           A(12) => PC_IN(12), A(11) => PC_IN(11), A(10) => 
                           PC_IN(10), A(9) => PC_IN(9), A(8) => PC_IN(8), A(7) 
                           => PC_IN(7), A(6) => PC_IN(6), A(5) => PC_IN(5), 
                           A(4) => PC_IN(4), A(3) => PC_IN(3), A(2) => PC_IN(2)
                           , A(1) => PC_IN(1), A(0) => PC_IN(0), B(31) => n7, 
                           B(30) => n7, B(29) => n7, B(28) => n7, B(27) => n7, 
                           B(26) => n7, B(25) => n7, B(24) => n7, B(23) => n7, 
                           B(22) => n7, B(21) => n7, B(20) => n7, B(19) => n7, 
                           B(18) => n7, B(17) => n7, B(16) => n7, B(15) => n7, 
                           B(14) => n7, B(13) => n7, B(12) => n7, B(11) => n7, 
                           B(10) => n7, B(9) => n7, B(8) => n7, B(7) => n7, 
                           B(6) => n7, B(5) => n7, B(4) => n7, B(3) => n7, B(2)
                           => n8, B(1) => n7, B(0) => n7, CI => n11, DIFF(31) 
                           => HDU_PC_OUT(31), DIFF(30) => HDU_PC_OUT(30), 
                           DIFF(29) => HDU_PC_OUT(29), DIFF(28) => 
                           HDU_PC_OUT(28), DIFF(27) => HDU_PC_OUT(27), DIFF(26)
                           => HDU_PC_OUT(26), DIFF(25) => HDU_PC_OUT(25), 
                           DIFF(24) => HDU_PC_OUT(24), DIFF(23) => 
                           HDU_PC_OUT(23), DIFF(22) => HDU_PC_OUT(22), DIFF(21)
                           => HDU_PC_OUT(21), DIFF(20) => HDU_PC_OUT(20), 
                           DIFF(19) => HDU_PC_OUT(19), DIFF(18) => 
                           HDU_PC_OUT(18), DIFF(17) => HDU_PC_OUT(17), DIFF(16)
                           => HDU_PC_OUT(16), DIFF(15) => HDU_PC_OUT(15), 
                           DIFF(14) => HDU_PC_OUT(14), DIFF(13) => 
                           HDU_PC_OUT(13), DIFF(12) => HDU_PC_OUT(12), DIFF(11)
                           => HDU_PC_OUT(11), DIFF(10) => HDU_PC_OUT(10), 
                           DIFF(9) => HDU_PC_OUT(9), DIFF(8) => HDU_PC_OUT(8), 
                           DIFF(7) => HDU_PC_OUT(7), DIFF(6) => HDU_PC_OUT(6), 
                           DIFF(5) => HDU_PC_OUT(5), DIFF(4) => HDU_PC_OUT(4), 
                           DIFF(3) => HDU_PC_OUT(3), DIFF(2) => HDU_PC_OUT(2), 
                           DIFF(1) => HDU_PC_OUT(1), DIFF(0) => HDU_PC_OUT(0), 
                           CO => n_1942);
   U4 : AND3_X1 port map( A1 => DRAM_R, A2 => n1, A3 => RST, ZN => Bubble);
   U5 : OAI33_X1 port map( A1 => n2, A2 => n3, A3 => n4, B1 => n5, B2 => n6, B3
                           => n9, ZN => n1);
   U6 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RS2(4), Z => n9);
   U8 : XOR2_X1 port map( A => ADD_WR(2), B => ADD_RS2(2), Z => n6);
   U9 : NAND3_X1 port map( A1 => n10, A2 => n12, A3 => n13, ZN => n5);
   U11 : XNOR2_X1 port map( A => ADD_WR(0), B => ADD_RS2(0), ZN => n13);
   U12 : XNOR2_X1 port map( A => ADD_WR(1), B => ADD_RS2(1), ZN => n12);
   U13 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS2(3), ZN => n10);
   U14 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RS1(4), Z => n4);
   U15 : XOR2_X1 port map( A => ADD_WR(2), B => ADD_RS1(2), Z => n3);
   U16 : NAND3_X1 port map( A1 => n14, A2 => n15, A3 => n16, ZN => n2);
   U17 : XNOR2_X1 port map( A => ADD_WR(0), B => ADD_RS1(0), ZN => n16);
   U18 : XNOR2_X1 port map( A => ADD_WR(1), B => ADD_RS1(1), ZN => n15);
   U19 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS1(3), ZN => n14);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Writeback is

   port( WB_MUX_SEL : in std_logic;  DATA_IN, ALU_RES_IN : in std_logic_vector 
         (31 downto 0);  ADD_WR_IN : in std_logic_vector (4 downto 0);  
         DATA_OUT : out std_logic_vector (31 downto 0);  ADD_WR_OUT : out 
         std_logic_vector (4 downto 0));

end Writeback;

architecture SYN_struct of Writeback is

   component mux21_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;

begin
   ADD_WR_OUT <= ( ADD_WR_IN(4), ADD_WR_IN(3), ADD_WR_IN(2), ADD_WR_IN(1), 
      ADD_WR_IN(0) );
   
   WBmux : mux21_NBIT32_2 port map( A(31) => DATA_IN(31), A(30) => DATA_IN(30),
                           A(29) => DATA_IN(29), A(28) => DATA_IN(28), A(27) =>
                           DATA_IN(27), A(26) => DATA_IN(26), A(25) => 
                           DATA_IN(25), A(24) => DATA_IN(24), A(23) => 
                           DATA_IN(23), A(22) => DATA_IN(22), A(21) => 
                           DATA_IN(21), A(20) => DATA_IN(20), A(19) => 
                           DATA_IN(19), A(18) => DATA_IN(18), A(17) => 
                           DATA_IN(17), A(16) => DATA_IN(16), A(15) => 
                           DATA_IN(15), A(14) => DATA_IN(14), A(13) => 
                           DATA_IN(13), A(12) => DATA_IN(12), A(11) => 
                           DATA_IN(11), A(10) => DATA_IN(10), A(9) => 
                           DATA_IN(9), A(8) => DATA_IN(8), A(7) => DATA_IN(7), 
                           A(6) => DATA_IN(6), A(5) => DATA_IN(5), A(4) => 
                           DATA_IN(4), A(3) => DATA_IN(3), A(2) => DATA_IN(2), 
                           A(1) => DATA_IN(1), A(0) => DATA_IN(0), B(31) => 
                           ALU_RES_IN(31), B(30) => ALU_RES_IN(30), B(29) => 
                           ALU_RES_IN(29), B(28) => ALU_RES_IN(28), B(27) => 
                           ALU_RES_IN(27), B(26) => ALU_RES_IN(26), B(25) => 
                           ALU_RES_IN(25), B(24) => ALU_RES_IN(24), B(23) => 
                           ALU_RES_IN(23), B(22) => ALU_RES_IN(22), B(21) => 
                           ALU_RES_IN(21), B(20) => ALU_RES_IN(20), B(19) => 
                           ALU_RES_IN(19), B(18) => ALU_RES_IN(18), B(17) => 
                           ALU_RES_IN(17), B(16) => ALU_RES_IN(16), B(15) => 
                           ALU_RES_IN(15), B(14) => ALU_RES_IN(14), B(13) => 
                           ALU_RES_IN(13), B(12) => ALU_RES_IN(12), B(11) => 
                           ALU_RES_IN(11), B(10) => ALU_RES_IN(10), B(9) => 
                           ALU_RES_IN(9), B(8) => ALU_RES_IN(8), B(7) => 
                           ALU_RES_IN(7), B(6) => ALU_RES_IN(6), B(5) => 
                           ALU_RES_IN(5), B(4) => ALU_RES_IN(4), B(3) => 
                           ALU_RES_IN(3), B(2) => ALU_RES_IN(2), B(1) => 
                           ALU_RES_IN(1), B(0) => ALU_RES_IN(0), S => 
                           WB_MUX_SEL, Z(31) => DATA_OUT(31), Z(30) => 
                           DATA_OUT(30), Z(29) => DATA_OUT(29), Z(28) => 
                           DATA_OUT(28), Z(27) => DATA_OUT(27), Z(26) => 
                           DATA_OUT(26), Z(25) => DATA_OUT(25), Z(24) => 
                           DATA_OUT(24), Z(23) => DATA_OUT(23), Z(22) => 
                           DATA_OUT(22), Z(21) => DATA_OUT(21), Z(20) => 
                           DATA_OUT(20), Z(19) => DATA_OUT(19), Z(18) => 
                           DATA_OUT(18), Z(17) => DATA_OUT(17), Z(16) => 
                           DATA_OUT(16), Z(15) => DATA_OUT(15), Z(14) => 
                           DATA_OUT(14), Z(13) => DATA_OUT(13), Z(12) => 
                           DATA_OUT(12), Z(11) => DATA_OUT(11), Z(10) => 
                           DATA_OUT(10), Z(9) => DATA_OUT(9), Z(8) => 
                           DATA_OUT(8), Z(7) => DATA_OUT(7), Z(6) => 
                           DATA_OUT(6), Z(5) => DATA_OUT(5), Z(4) => 
                           DATA_OUT(4), Z(3) => DATA_OUT(3), Z(2) => 
                           DATA_OUT(2), Z(1) => DATA_OUT(1), Z(0) => 
                           DATA_OUT(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Memory is

   port( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, DRAM_EN_IN : in std_logic; 
         PC_SEL : in std_logic_vector (1 downto 0);  NPC_IN, NPC_ABS, NPC_REL, 
         ALU_RES_IN, B_IN : in std_logic_vector (31 downto 0);  ADD_WR_IN : in 
         std_logic_vector (4 downto 0);  DRAM_DATA_IN : in std_logic_vector (31
         downto 0);  PC_OUT : out std_logic_vector (31 downto 0);  DRAM_EN_OUT,
         DRAM_R_OUT, DRAM_W_OUT : out std_logic;  DRAM_ADDR_OUT, DRAM_DATA_OUT,
         DATA_OUT, ALU_RES_OUT, OP_MEM : out std_logic_vector (31 downto 0);  
         ADD_WR_MEM, ADD_WR_OUT : out std_logic_vector (4 downto 0));

end Memory;

architecture SYN_struct of Memory is

   component mux41_NBIT32_2
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component regn_N32_1
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N5_1
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N32_2
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port : std_logic;

begin
   DRAM_EN_OUT <= DRAM_EN_IN;
   DRAM_R_OUT <= DRAM_R_IN;
   DRAM_W_OUT <= DRAM_W_IN;
   DRAM_ADDR_OUT <= ( ALU_RES_IN(31), ALU_RES_IN(30), ALU_RES_IN(29), 
      ALU_RES_IN(28), ALU_RES_IN(27), ALU_RES_IN(26), ALU_RES_IN(25), 
      ALU_RES_IN(24), ALU_RES_IN(23), ALU_RES_IN(22), ALU_RES_IN(21), 
      ALU_RES_IN(20), ALU_RES_IN(19), ALU_RES_IN(18), ALU_RES_IN(17), 
      ALU_RES_IN(16), ALU_RES_IN(15), ALU_RES_IN(14), ALU_RES_IN(13), 
      ALU_RES_IN(12), ALU_RES_IN(11), ALU_RES_IN(10), ALU_RES_IN(9), 
      ALU_RES_IN(8), ALU_RES_IN(7), ALU_RES_IN(6), ALU_RES_IN(5), ALU_RES_IN(4)
      , ALU_RES_IN(3), ALU_RES_IN(2), ALU_RES_IN(1), ALU_RES_IN(0) );
   DRAM_DATA_OUT <= ( B_IN(31), B_IN(30), B_IN(29), B_IN(28), B_IN(27), 
      B_IN(26), B_IN(25), B_IN(24), B_IN(23), B_IN(22), B_IN(21), B_IN(20), 
      B_IN(19), B_IN(18), B_IN(17), B_IN(16), B_IN(15), B_IN(14), B_IN(13), 
      B_IN(12), B_IN(11), B_IN(10), B_IN(9), B_IN(8), B_IN(7), B_IN(6), B_IN(5)
      , B_IN(4), B_IN(3), B_IN(2), B_IN(1), B_IN(0) );
   OP_MEM <= ( ALU_RES_IN(31), ALU_RES_IN(30), ALU_RES_IN(29), ALU_RES_IN(28), 
      ALU_RES_IN(27), ALU_RES_IN(26), ALU_RES_IN(25), ALU_RES_IN(24), 
      ALU_RES_IN(23), ALU_RES_IN(22), ALU_RES_IN(21), ALU_RES_IN(20), 
      ALU_RES_IN(19), ALU_RES_IN(18), ALU_RES_IN(17), ALU_RES_IN(16), 
      ALU_RES_IN(15), ALU_RES_IN(14), ALU_RES_IN(13), ALU_RES_IN(12), 
      ALU_RES_IN(11), ALU_RES_IN(10), ALU_RES_IN(9), ALU_RES_IN(8), 
      ALU_RES_IN(7), ALU_RES_IN(6), ALU_RES_IN(5), ALU_RES_IN(4), ALU_RES_IN(3)
      , ALU_RES_IN(2), ALU_RES_IN(1), ALU_RES_IN(0) );
   ADD_WR_MEM <= ( ADD_WR_IN(4), ADD_WR_IN(3), ADD_WR_IN(2), ADD_WR_IN(1), 
      ADD_WR_IN(0) );
   
   X_Logic0_port <= '0';
   LMD : regn_N32_2 port map( DIN(31) => DRAM_DATA_IN(31), DIN(30) => 
                           DRAM_DATA_IN(30), DIN(29) => DRAM_DATA_IN(29), 
                           DIN(28) => DRAM_DATA_IN(28), DIN(27) => 
                           DRAM_DATA_IN(27), DIN(26) => DRAM_DATA_IN(26), 
                           DIN(25) => DRAM_DATA_IN(25), DIN(24) => 
                           DRAM_DATA_IN(24), DIN(23) => DRAM_DATA_IN(23), 
                           DIN(22) => DRAM_DATA_IN(22), DIN(21) => 
                           DRAM_DATA_IN(21), DIN(20) => DRAM_DATA_IN(20), 
                           DIN(19) => DRAM_DATA_IN(19), DIN(18) => 
                           DRAM_DATA_IN(18), DIN(17) => DRAM_DATA_IN(17), 
                           DIN(16) => DRAM_DATA_IN(16), DIN(15) => 
                           DRAM_DATA_IN(15), DIN(14) => DRAM_DATA_IN(14), 
                           DIN(13) => DRAM_DATA_IN(13), DIN(12) => 
                           DRAM_DATA_IN(12), DIN(11) => DRAM_DATA_IN(11), 
                           DIN(10) => DRAM_DATA_IN(10), DIN(9) => 
                           DRAM_DATA_IN(9), DIN(8) => DRAM_DATA_IN(8), DIN(7) 
                           => DRAM_DATA_IN(7), DIN(6) => DRAM_DATA_IN(6), 
                           DIN(5) => DRAM_DATA_IN(5), DIN(4) => DRAM_DATA_IN(4)
                           , DIN(3) => DRAM_DATA_IN(3), DIN(2) => 
                           DRAM_DATA_IN(2), DIN(1) => DRAM_DATA_IN(1), DIN(0) 
                           => DRAM_DATA_IN(0), CLK => CLK, EN => MEM_EN_IN, RST
                           => RST, DOUT(31) => DATA_OUT(31), DOUT(30) => 
                           DATA_OUT(30), DOUT(29) => DATA_OUT(29), DOUT(28) => 
                           DATA_OUT(28), DOUT(27) => DATA_OUT(27), DOUT(26) => 
                           DATA_OUT(26), DOUT(25) => DATA_OUT(25), DOUT(24) => 
                           DATA_OUT(24), DOUT(23) => DATA_OUT(23), DOUT(22) => 
                           DATA_OUT(22), DOUT(21) => DATA_OUT(21), DOUT(20) => 
                           DATA_OUT(20), DOUT(19) => DATA_OUT(19), DOUT(18) => 
                           DATA_OUT(18), DOUT(17) => DATA_OUT(17), DOUT(16) => 
                           DATA_OUT(16), DOUT(15) => DATA_OUT(15), DOUT(14) => 
                           DATA_OUT(14), DOUT(13) => DATA_OUT(13), DOUT(12) => 
                           DATA_OUT(12), DOUT(11) => DATA_OUT(11), DOUT(10) => 
                           DATA_OUT(10), DOUT(9) => DATA_OUT(9), DOUT(8) => 
                           DATA_OUT(8), DOUT(7) => DATA_OUT(7), DOUT(6) => 
                           DATA_OUT(6), DOUT(5) => DATA_OUT(5), DOUT(4) => 
                           DATA_OUT(4), DOUT(3) => DATA_OUT(3), DOUT(2) => 
                           DATA_OUT(2), DOUT(1) => DATA_OUT(1), DOUT(0) => 
                           DATA_OUT(0));
   reg0 : regn_N5_1 port map( DIN(4) => ADD_WR_IN(4), DIN(3) => ADD_WR_IN(3), 
                           DIN(2) => ADD_WR_IN(2), DIN(1) => ADD_WR_IN(1), 
                           DIN(0) => ADD_WR_IN(0), CLK => CLK, EN => MEM_EN_IN,
                           RST => RST, DOUT(4) => ADD_WR_OUT(4), DOUT(3) => 
                           ADD_WR_OUT(3), DOUT(2) => ADD_WR_OUT(2), DOUT(1) => 
                           ADD_WR_OUT(1), DOUT(0) => ADD_WR_OUT(0));
   reg1 : regn_N32_1 port map( DIN(31) => ALU_RES_IN(31), DIN(30) => 
                           ALU_RES_IN(30), DIN(29) => ALU_RES_IN(29), DIN(28) 
                           => ALU_RES_IN(28), DIN(27) => ALU_RES_IN(27), 
                           DIN(26) => ALU_RES_IN(26), DIN(25) => ALU_RES_IN(25)
                           , DIN(24) => ALU_RES_IN(24), DIN(23) => 
                           ALU_RES_IN(23), DIN(22) => ALU_RES_IN(22), DIN(21) 
                           => ALU_RES_IN(21), DIN(20) => ALU_RES_IN(20), 
                           DIN(19) => ALU_RES_IN(19), DIN(18) => ALU_RES_IN(18)
                           , DIN(17) => ALU_RES_IN(17), DIN(16) => 
                           ALU_RES_IN(16), DIN(15) => ALU_RES_IN(15), DIN(14) 
                           => ALU_RES_IN(14), DIN(13) => ALU_RES_IN(13), 
                           DIN(12) => ALU_RES_IN(12), DIN(11) => ALU_RES_IN(11)
                           , DIN(10) => ALU_RES_IN(10), DIN(9) => ALU_RES_IN(9)
                           , DIN(8) => ALU_RES_IN(8), DIN(7) => ALU_RES_IN(7), 
                           DIN(6) => ALU_RES_IN(6), DIN(5) => ALU_RES_IN(5), 
                           DIN(4) => ALU_RES_IN(4), DIN(3) => ALU_RES_IN(3), 
                           DIN(2) => ALU_RES_IN(2), DIN(1) => ALU_RES_IN(1), 
                           DIN(0) => ALU_RES_IN(0), CLK => CLK, EN => MEM_EN_IN
                           , RST => RST, DOUT(31) => ALU_RES_OUT(31), DOUT(30) 
                           => ALU_RES_OUT(30), DOUT(29) => ALU_RES_OUT(29), 
                           DOUT(28) => ALU_RES_OUT(28), DOUT(27) => 
                           ALU_RES_OUT(27), DOUT(26) => ALU_RES_OUT(26), 
                           DOUT(25) => ALU_RES_OUT(25), DOUT(24) => 
                           ALU_RES_OUT(24), DOUT(23) => ALU_RES_OUT(23), 
                           DOUT(22) => ALU_RES_OUT(22), DOUT(21) => 
                           ALU_RES_OUT(21), DOUT(20) => ALU_RES_OUT(20), 
                           DOUT(19) => ALU_RES_OUT(19), DOUT(18) => 
                           ALU_RES_OUT(18), DOUT(17) => ALU_RES_OUT(17), 
                           DOUT(16) => ALU_RES_OUT(16), DOUT(15) => 
                           ALU_RES_OUT(15), DOUT(14) => ALU_RES_OUT(14), 
                           DOUT(13) => ALU_RES_OUT(13), DOUT(12) => 
                           ALU_RES_OUT(12), DOUT(11) => ALU_RES_OUT(11), 
                           DOUT(10) => ALU_RES_OUT(10), DOUT(9) => 
                           ALU_RES_OUT(9), DOUT(8) => ALU_RES_OUT(8), DOUT(7) 
                           => ALU_RES_OUT(7), DOUT(6) => ALU_RES_OUT(6), 
                           DOUT(5) => ALU_RES_OUT(5), DOUT(4) => ALU_RES_OUT(4)
                           , DOUT(3) => ALU_RES_OUT(3), DOUT(2) => 
                           ALU_RES_OUT(2), DOUT(1) => ALU_RES_OUT(1), DOUT(0) 
                           => ALU_RES_OUT(0));
   PCsel : mux41_NBIT32_2 port map( A(31) => NPC_IN(31), A(30) => NPC_IN(30), 
                           A(29) => NPC_IN(29), A(28) => NPC_IN(28), A(27) => 
                           NPC_IN(27), A(26) => NPC_IN(26), A(25) => NPC_IN(25)
                           , A(24) => NPC_IN(24), A(23) => NPC_IN(23), A(22) =>
                           NPC_IN(22), A(21) => NPC_IN(21), A(20) => NPC_IN(20)
                           , A(19) => NPC_IN(19), A(18) => NPC_IN(18), A(17) =>
                           NPC_IN(17), A(16) => NPC_IN(16), A(15) => NPC_IN(15)
                           , A(14) => NPC_IN(14), A(13) => NPC_IN(13), A(12) =>
                           NPC_IN(12), A(11) => NPC_IN(11), A(10) => NPC_IN(10)
                           , A(9) => NPC_IN(9), A(8) => NPC_IN(8), A(7) => 
                           NPC_IN(7), A(6) => NPC_IN(6), A(5) => NPC_IN(5), 
                           A(4) => NPC_IN(4), A(3) => NPC_IN(3), A(2) => 
                           NPC_IN(2), A(1) => NPC_IN(1), A(0) => NPC_IN(0), 
                           B(31) => NPC_REL(31), B(30) => NPC_REL(30), B(29) =>
                           NPC_REL(29), B(28) => NPC_REL(28), B(27) => 
                           NPC_REL(27), B(26) => NPC_REL(26), B(25) => 
                           NPC_REL(25), B(24) => NPC_REL(24), B(23) => 
                           NPC_REL(23), B(22) => NPC_REL(22), B(21) => 
                           NPC_REL(21), B(20) => NPC_REL(20), B(19) => 
                           NPC_REL(19), B(18) => NPC_REL(18), B(17) => 
                           NPC_REL(17), B(16) => NPC_REL(16), B(15) => 
                           NPC_REL(15), B(14) => NPC_REL(14), B(13) => 
                           NPC_REL(13), B(12) => NPC_REL(12), B(11) => 
                           NPC_REL(11), B(10) => NPC_REL(10), B(9) => 
                           NPC_REL(9), B(8) => NPC_REL(8), B(7) => NPC_REL(7), 
                           B(6) => NPC_REL(6), B(5) => NPC_REL(5), B(4) => 
                           NPC_REL(4), B(3) => NPC_REL(3), B(2) => NPC_REL(2), 
                           B(1) => NPC_REL(1), B(0) => NPC_REL(0), C(31) => 
                           NPC_ABS(31), C(30) => NPC_ABS(30), C(29) => 
                           NPC_ABS(29), C(28) => NPC_ABS(28), C(27) => 
                           NPC_ABS(27), C(26) => NPC_ABS(26), C(25) => 
                           NPC_ABS(25), C(24) => NPC_ABS(24), C(23) => 
                           NPC_ABS(23), C(22) => NPC_ABS(22), C(21) => 
                           NPC_ABS(21), C(20) => NPC_ABS(20), C(19) => 
                           NPC_ABS(19), C(18) => NPC_ABS(18), C(17) => 
                           NPC_ABS(17), C(16) => NPC_ABS(16), C(15) => 
                           NPC_ABS(15), C(14) => NPC_ABS(14), C(13) => 
                           NPC_ABS(13), C(12) => NPC_ABS(12), C(11) => 
                           NPC_ABS(11), C(10) => NPC_ABS(10), C(9) => 
                           NPC_ABS(9), C(8) => NPC_ABS(8), C(7) => NPC_ABS(7), 
                           C(6) => NPC_ABS(6), C(5) => NPC_ABS(5), C(4) => 
                           NPC_ABS(4), C(3) => NPC_ABS(3), C(2) => NPC_ABS(2), 
                           C(1) => NPC_ABS(1), C(0) => NPC_ABS(0), D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => X_Logic0_port, D(25) => 
                           X_Logic0_port, D(24) => X_Logic0_port, D(23) => 
                           X_Logic0_port, D(22) => X_Logic0_port, D(21) => 
                           X_Logic0_port, D(20) => X_Logic0_port, D(19) => 
                           X_Logic0_port, D(18) => X_Logic0_port, D(17) => 
                           X_Logic0_port, D(16) => X_Logic0_port, D(15) => 
                           X_Logic0_port, D(14) => X_Logic0_port, D(13) => 
                           X_Logic0_port, D(12) => X_Logic0_port, D(11) => 
                           X_Logic0_port, D(10) => X_Logic0_port, D(9) => 
                           X_Logic0_port, D(8) => X_Logic0_port, D(7) => 
                           X_Logic0_port, D(6) => X_Logic0_port, D(5) => 
                           X_Logic0_port, D(4) => X_Logic0_port, D(3) => 
                           X_Logic0_port, D(2) => X_Logic0_port, D(1) => 
                           X_Logic0_port, D(0) => X_Logic0_port, S(1) => 
                           PC_SEL(1), S(0) => PC_SEL(0), Z(31) => PC_OUT(31), 
                           Z(30) => PC_OUT(30), Z(29) => PC_OUT(29), Z(28) => 
                           PC_OUT(28), Z(27) => PC_OUT(27), Z(26) => PC_OUT(26)
                           , Z(25) => PC_OUT(25), Z(24) => PC_OUT(24), Z(23) =>
                           PC_OUT(23), Z(22) => PC_OUT(22), Z(21) => PC_OUT(21)
                           , Z(20) => PC_OUT(20), Z(19) => PC_OUT(19), Z(18) =>
                           PC_OUT(18), Z(17) => PC_OUT(17), Z(16) => PC_OUT(16)
                           , Z(15) => PC_OUT(15), Z(14) => PC_OUT(14), Z(13) =>
                           PC_OUT(13), Z(12) => PC_OUT(12), Z(11) => PC_OUT(11)
                           , Z(10) => PC_OUT(10), Z(9) => PC_OUT(9), Z(8) => 
                           PC_OUT(8), Z(7) => PC_OUT(7), Z(6) => PC_OUT(6), 
                           Z(5) => PC_OUT(5), Z(4) => PC_OUT(4), Z(3) => 
                           PC_OUT(3), Z(2) => PC_OUT(2), Z(1) => PC_OUT(1), 
                           Z(0) => PC_OUT(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ff_0 is

   port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);

end ff_0;

architecture SYN_bhv of ff_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n3, CK => CLK, RN => RST, Q => Q, QN => n2);
   U2 : OAI21_X1 port map( B1 => n2, B2 => EN, A => n1, ZN => n3);
   U3 : NAND2_X1 port map( A1 => EN, A2 => D, ZN => n1);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute is

   port( CLK, RST, MUX_A_SEL : in std_logic;  MUX_B_SEL : in std_logic_vector 
         (1 downto 0);  ALU_OPC : in std_logic_vector (0 to 3);  ALU_OUTREG_EN 
         : in std_logic;  JUMP_TYPE : in std_logic_vector (1 downto 0);  PC_IN,
         A_IN, B_IN, IMM_IN : in std_logic_vector (31 downto 0);  ADD_WR_IN, 
         ADD_RS1_IN, ADD_RS2_IN, ADD_WR_MEM, ADD_WR_WB : in std_logic_vector (4
         downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;  OP_MEM, OP_WB : in 
         std_logic_vector (31 downto 0);  PC_SEL : out std_logic_vector (1 
         downto 0);  ZERO_FLAG : out std_logic;  NPC_ABS, NPC_REL, ALU_RES, 
         B_OUT : out std_logic_vector (31 downto 0);  ADD_WR_OUT : out 
         std_logic_vector (4 downto 0));

end Execute;

architecture SYN_struct of Execute is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component Execute_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component Execute_DW01_add_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component regn_N32_3
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_4
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N5_2
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N32_5
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_6
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component ALU_NBIT32
      port( OP1, OP2 : in std_logic_vector (31 downto 0);  ALU_OPC : in 
            std_logic_vector (0 to 3);  ALU_RES : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux41_NBIT32_3
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux21_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux41_NBIT32_4
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux41_NBIT32_0
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component FWD_Unit
      port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB : in 
            std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;
            FWDA, FWDB : out std_logic_vector (1 downto 0));
   end component;
   
   component regn_N2
      port( DIN : in std_logic_vector (1 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (1 downto 0));
   end component;
   
   component ff_1
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Branch_Cond_Unit_NBIT32
      port( RST : in std_logic;  A : in std_logic_vector (31 downto 0);  
            ALU_OPC : in std_logic_vector (0 to 3);  JUMP_TYPE : in 
            std_logic_vector (1 downto 0);  PC_SEL : out std_logic_vector (1 
            downto 0);  ZERO : out std_logic);
   end component;
   
   signal ZERO_FLAG_port, sig_RST, sig_NPC_ABS_31_port, sig_NPC_ABS_30_port, 
      sig_NPC_ABS_29_port, sig_NPC_ABS_28_port, sig_NPC_ABS_27_port, 
      sig_NPC_ABS_26_port, sig_NPC_ABS_25_port, sig_NPC_ABS_24_port, 
      sig_NPC_ABS_23_port, sig_NPC_ABS_22_port, sig_NPC_ABS_21_port, 
      sig_NPC_ABS_20_port, sig_NPC_ABS_19_port, sig_NPC_ABS_18_port, 
      sig_NPC_ABS_17_port, sig_NPC_ABS_16_port, sig_NPC_ABS_15_port, 
      sig_NPC_ABS_14_port, sig_NPC_ABS_13_port, sig_NPC_ABS_12_port, 
      sig_NPC_ABS_11_port, sig_NPC_ABS_10_port, sig_NPC_ABS_9_port, 
      sig_NPC_ABS_8_port, sig_NPC_ABS_7_port, sig_NPC_ABS_6_port, 
      sig_NPC_ABS_5_port, sig_NPC_ABS_4_port, sig_NPC_ABS_3_port, 
      sig_NPC_ABS_2_port, sig_NPC_ABS_1_port, sig_NPC_ABS_0_port, 
      sig_NPC_REL_31_port, sig_NPC_REL_30_port, sig_NPC_REL_29_port, 
      sig_NPC_REL_28_port, sig_NPC_REL_27_port, sig_NPC_REL_26_port, 
      sig_NPC_REL_25_port, sig_NPC_REL_24_port, sig_NPC_REL_23_port, 
      sig_NPC_REL_22_port, sig_NPC_REL_21_port, sig_NPC_REL_20_port, 
      sig_NPC_REL_19_port, sig_NPC_REL_18_port, sig_NPC_REL_17_port, 
      sig_NPC_REL_16_port, sig_NPC_REL_15_port, sig_NPC_REL_14_port, 
      sig_NPC_REL_13_port, sig_NPC_REL_12_port, sig_NPC_REL_11_port, 
      sig_NPC_REL_10_port, sig_NPC_REL_9_port, sig_NPC_REL_8_port, 
      sig_NPC_REL_7_port, sig_NPC_REL_6_port, sig_NPC_REL_5_port, 
      sig_NPC_REL_4_port, sig_NPC_REL_3_port, sig_NPC_REL_2_port, 
      sig_NPC_REL_1_port, sig_NPC_REL_0_port, sig_PC_SEL_1_port, 
      sig_PC_SEL_0_port, sig_ZERO_FLAG, FWDA_1_port, FWDA_0_port, FWDB_1_port, 
      FWDB_0_port, OP2_FW_31_port, OP2_FW_30_port, OP2_FW_29_port, 
      OP2_FW_28_port, OP2_FW_27_port, OP2_FW_26_port, OP2_FW_25_port, 
      OP2_FW_24_port, OP2_FW_23_port, OP2_FW_22_port, OP2_FW_21_port, 
      OP2_FW_20_port, OP2_FW_19_port, OP2_FW_18_port, OP2_FW_17_port, 
      OP2_FW_16_port, OP2_FW_15_port, OP2_FW_14_port, OP2_FW_13_port, 
      OP2_FW_12_port, OP2_FW_11_port, OP2_FW_10_port, OP2_FW_9_port, 
      OP2_FW_8_port, OP2_FW_7_port, OP2_FW_6_port, OP2_FW_5_port, OP2_FW_4_port
      , OP2_FW_3_port, OP2_FW_2_port, OP2_FW_1_port, OP2_FW_0_port, 
      sig_OP1_31_port, sig_OP1_30_port, sig_OP1_29_port, sig_OP1_28_port, 
      sig_OP1_27_port, sig_OP1_26_port, sig_OP1_25_port, sig_OP1_24_port, 
      sig_OP1_23_port, sig_OP1_22_port, sig_OP1_21_port, sig_OP1_20_port, 
      sig_OP1_19_port, sig_OP1_18_port, sig_OP1_17_port, sig_OP1_16_port, 
      sig_OP1_15_port, sig_OP1_14_port, sig_OP1_13_port, sig_OP1_12_port, 
      sig_OP1_11_port, sig_OP1_10_port, sig_OP1_9_port, sig_OP1_8_port, 
      sig_OP1_7_port, sig_OP1_6_port, sig_OP1_5_port, sig_OP1_4_port, 
      sig_OP1_3_port, sig_OP1_2_port, sig_OP1_1_port, sig_OP1_0_port, 
      sig_OP2_31_port, sig_OP2_30_port, sig_OP2_29_port, sig_OP2_28_port, 
      sig_OP2_27_port, sig_OP2_26_port, sig_OP2_25_port, sig_OP2_24_port, 
      sig_OP2_23_port, sig_OP2_22_port, sig_OP2_21_port, sig_OP2_20_port, 
      sig_OP2_19_port, sig_OP2_18_port, sig_OP2_17_port, sig_OP2_16_port, 
      sig_OP2_15_port, sig_OP2_14_port, sig_OP2_13_port, sig_OP2_12_port, 
      sig_OP2_11_port, sig_OP2_10_port, sig_OP2_9_port, sig_OP2_8_port, 
      sig_OP2_7_port, sig_OP2_6_port, sig_OP2_5_port, sig_OP2_4_port, 
      sig_OP2_3_port, sig_OP2_2_port, sig_OP2_1_port, sig_OP2_0_port, 
      sig_ALU_RES_31_port, sig_ALU_RES_30_port, sig_ALU_RES_29_port, 
      sig_ALU_RES_28_port, sig_ALU_RES_27_port, sig_ALU_RES_26_port, 
      sig_ALU_RES_25_port, sig_ALU_RES_24_port, sig_ALU_RES_23_port, 
      sig_ALU_RES_22_port, sig_ALU_RES_21_port, sig_ALU_RES_20_port, 
      sig_ALU_RES_19_port, sig_ALU_RES_18_port, sig_ALU_RES_17_port, 
      sig_ALU_RES_16_port, sig_ALU_RES_15_port, sig_ALU_RES_14_port, 
      sig_ALU_RES_13_port, sig_ALU_RES_12_port, sig_ALU_RES_11_port, 
      sig_ALU_RES_10_port, sig_ALU_RES_9_port, sig_ALU_RES_8_port, 
      sig_ALU_RES_7_port, sig_ALU_RES_6_port, sig_ALU_RES_5_port, 
      sig_ALU_RES_4_port, sig_ALU_RES_3_port, sig_ALU_RES_2_port, 
      sig_ALU_RES_1_port, sig_ALU_RES_0_port, N9, N8, N7, N6, N5, N4, N31, N30,
      N3, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N2, N19, N18, N17, 
      N16, N15, N14, N13, N12, N11, N10, N1, N0, n1_port, n2_port, n3_port, 
      n4_port, n5_port, n6_port, n7_port, n_1943, n_1944 : std_logic;

begin
   ZERO_FLAG <= ZERO_FLAG_port;
   
   n7_port <= '1';
   n6_port <= '0';
   Branch_Cond : Branch_Cond_Unit_NBIT32 port map( RST => sig_RST, A(31) => 
                           sig_NPC_ABS_31_port, A(30) => sig_NPC_ABS_30_port, 
                           A(29) => sig_NPC_ABS_29_port, A(28) => 
                           sig_NPC_ABS_28_port, A(27) => sig_NPC_ABS_27_port, 
                           A(26) => sig_NPC_ABS_26_port, A(25) => 
                           sig_NPC_ABS_25_port, A(24) => sig_NPC_ABS_24_port, 
                           A(23) => sig_NPC_ABS_23_port, A(22) => 
                           sig_NPC_ABS_22_port, A(21) => sig_NPC_ABS_21_port, 
                           A(20) => sig_NPC_ABS_20_port, A(19) => 
                           sig_NPC_ABS_19_port, A(18) => sig_NPC_ABS_18_port, 
                           A(17) => sig_NPC_ABS_17_port, A(16) => 
                           sig_NPC_ABS_16_port, A(15) => sig_NPC_ABS_15_port, 
                           A(14) => sig_NPC_ABS_14_port, A(13) => 
                           sig_NPC_ABS_13_port, A(12) => sig_NPC_ABS_12_port, 
                           A(11) => sig_NPC_ABS_11_port, A(10) => 
                           sig_NPC_ABS_10_port, A(9) => sig_NPC_ABS_9_port, 
                           A(8) => sig_NPC_ABS_8_port, A(7) => 
                           sig_NPC_ABS_7_port, A(6) => sig_NPC_ABS_6_port, A(5)
                           => sig_NPC_ABS_5_port, A(4) => sig_NPC_ABS_4_port, 
                           A(3) => sig_NPC_ABS_3_port, A(2) => 
                           sig_NPC_ABS_2_port, A(1) => sig_NPC_ABS_1_port, A(0)
                           => sig_NPC_ABS_0_port, ALU_OPC(0) => ALU_OPC(0), 
                           ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => ALU_OPC(2), 
                           ALU_OPC(3) => ALU_OPC(3), JUMP_TYPE(1) => 
                           JUMP_TYPE(1), JUMP_TYPE(0) => JUMP_TYPE(0), 
                           PC_SEL(1) => sig_PC_SEL_1_port, PC_SEL(0) => 
                           sig_PC_SEL_0_port, ZERO => sig_ZERO_FLAG);
   ff0 : ff_1 port map( D => sig_ZERO_FLAG, CLK => CLK, EN => n7_port, RST => 
                           RST, Q => ZERO_FLAG_port);
   reg0 : regn_N2 port map( DIN(1) => sig_PC_SEL_1_port, DIN(0) => 
                           sig_PC_SEL_0_port, CLK => CLK, EN => n7_port, RST =>
                           RST, DOUT(1) => PC_SEL(1), DOUT(0) => PC_SEL(0));
   FWD : FWD_Unit port map( RST => sig_RST, ADD_RS1(4) => ADD_RS1_IN(4), 
                           ADD_RS1(3) => ADD_RS1_IN(3), ADD_RS1(2) => 
                           ADD_RS1_IN(2), ADD_RS1(1) => ADD_RS1_IN(1), 
                           ADD_RS1(0) => ADD_RS1_IN(0), ADD_RS2(4) => 
                           ADD_RS2_IN(4), ADD_RS2(3) => ADD_RS2_IN(3), 
                           ADD_RS2(2) => ADD_RS2_IN(2), ADD_RS2(1) => 
                           ADD_RS2_IN(1), ADD_RS2(0) => ADD_RS2_IN(0), 
                           ADD_WR_MEM(4) => ADD_WR_MEM(4), ADD_WR_MEM(3) => 
                           ADD_WR_MEM(3), ADD_WR_MEM(2) => ADD_WR_MEM(2), 
                           ADD_WR_MEM(1) => ADD_WR_MEM(1), ADD_WR_MEM(0) => 
                           ADD_WR_MEM(0), ADD_WR_WB(4) => ADD_WR_WB(4), 
                           ADD_WR_WB(3) => ADD_WR_WB(3), ADD_WR_WB(2) => 
                           ADD_WR_WB(2), ADD_WR_WB(1) => ADD_WR_WB(1), 
                           ADD_WR_WB(0) => ADD_WR_WB(0), RF_WE_MEM => RF_WE_MEM
                           , RF_WE_WB => RF_WE_WB, FWDA(1) => FWDA_1_port, 
                           FWDA(0) => FWDA_0_port, FWDB(1) => FWDB_1_port, 
                           FWDB(0) => FWDB_0_port);
   FW1 : mux41_NBIT32_0 port map( A(31) => A_IN(31), A(30) => A_IN(30), A(29) 
                           => A_IN(29), A(28) => A_IN(28), A(27) => A_IN(27), 
                           A(26) => A_IN(26), A(25) => A_IN(25), A(24) => 
                           A_IN(24), A(23) => A_IN(23), A(22) => A_IN(22), 
                           A(21) => A_IN(21), A(20) => A_IN(20), A(19) => 
                           A_IN(19), A(18) => A_IN(18), A(17) => A_IN(17), 
                           A(16) => A_IN(16), A(15) => A_IN(15), A(14) => 
                           A_IN(14), A(13) => A_IN(13), A(12) => A_IN(12), 
                           A(11) => A_IN(11), A(10) => A_IN(10), A(9) => 
                           A_IN(9), A(8) => A_IN(8), A(7) => A_IN(7), A(6) => 
                           A_IN(6), A(5) => A_IN(5), A(4) => A_IN(4), A(3) => 
                           A_IN(3), A(2) => A_IN(2), A(1) => A_IN(1), A(0) => 
                           A_IN(0), B(31) => OP_WB(31), B(30) => OP_WB(30), 
                           B(29) => OP_WB(29), B(28) => OP_WB(28), B(27) => 
                           OP_WB(27), B(26) => OP_WB(26), B(25) => OP_WB(25), 
                           B(24) => OP_WB(24), B(23) => OP_WB(23), B(22) => 
                           OP_WB(22), B(21) => OP_WB(21), B(20) => OP_WB(20), 
                           B(19) => OP_WB(19), B(18) => OP_WB(18), B(17) => 
                           OP_WB(17), B(16) => OP_WB(16), B(15) => OP_WB(15), 
                           B(14) => OP_WB(14), B(13) => OP_WB(13), B(12) => 
                           OP_WB(12), B(11) => OP_WB(11), B(10) => OP_WB(10), 
                           B(9) => OP_WB(9), B(8) => OP_WB(8), B(7) => OP_WB(7)
                           , B(6) => OP_WB(6), B(5) => OP_WB(5), B(4) => 
                           OP_WB(4), B(3) => OP_WB(3), B(2) => OP_WB(2), B(1) 
                           => OP_WB(1), B(0) => OP_WB(0), C(31) => OP_MEM(31), 
                           C(30) => OP_MEM(30), C(29) => OP_MEM(29), C(28) => 
                           OP_MEM(28), C(27) => OP_MEM(27), C(26) => OP_MEM(26)
                           , C(25) => OP_MEM(25), C(24) => OP_MEM(24), C(23) =>
                           OP_MEM(23), C(22) => OP_MEM(22), C(21) => OP_MEM(21)
                           , C(20) => OP_MEM(20), C(19) => OP_MEM(19), C(18) =>
                           OP_MEM(18), C(17) => OP_MEM(17), C(16) => OP_MEM(16)
                           , C(15) => OP_MEM(15), C(14) => OP_MEM(14), C(13) =>
                           OP_MEM(13), C(12) => OP_MEM(12), C(11) => OP_MEM(11)
                           , C(10) => OP_MEM(10), C(9) => OP_MEM(9), C(8) => 
                           OP_MEM(8), C(7) => OP_MEM(7), C(6) => OP_MEM(6), 
                           C(5) => OP_MEM(5), C(4) => OP_MEM(4), C(3) => 
                           OP_MEM(3), C(2) => OP_MEM(2), C(1) => OP_MEM(1), 
                           C(0) => OP_MEM(0), D(31) => n6_port, D(30) => 
                           n6_port, D(29) => n6_port, D(28) => n6_port, D(27) 
                           => n6_port, D(26) => n6_port, D(25) => n6_port, 
                           D(24) => n6_port, D(23) => n6_port, D(22) => n6_port
                           , D(21) => n6_port, D(20) => n6_port, D(19) => 
                           n6_port, D(18) => n6_port, D(17) => n6_port, D(16) 
                           => n6_port, D(15) => n6_port, D(14) => n6_port, 
                           D(13) => n6_port, D(12) => n6_port, D(11) => n6_port
                           , D(10) => n6_port, D(9) => n6_port, D(8) => n6_port
                           , D(7) => n6_port, D(6) => n6_port, D(5) => n6_port,
                           D(4) => n6_port, D(3) => n6_port, D(2) => n6_port, 
                           D(1) => n6_port, D(0) => n6_port, S(1) => 
                           FWDA_1_port, S(0) => FWDA_0_port, Z(31) => 
                           sig_NPC_ABS_31_port, Z(30) => sig_NPC_ABS_30_port, 
                           Z(29) => sig_NPC_ABS_29_port, Z(28) => 
                           sig_NPC_ABS_28_port, Z(27) => sig_NPC_ABS_27_port, 
                           Z(26) => sig_NPC_ABS_26_port, Z(25) => 
                           sig_NPC_ABS_25_port, Z(24) => sig_NPC_ABS_24_port, 
                           Z(23) => sig_NPC_ABS_23_port, Z(22) => 
                           sig_NPC_ABS_22_port, Z(21) => sig_NPC_ABS_21_port, 
                           Z(20) => sig_NPC_ABS_20_port, Z(19) => 
                           sig_NPC_ABS_19_port, Z(18) => sig_NPC_ABS_18_port, 
                           Z(17) => sig_NPC_ABS_17_port, Z(16) => 
                           sig_NPC_ABS_16_port, Z(15) => sig_NPC_ABS_15_port, 
                           Z(14) => sig_NPC_ABS_14_port, Z(13) => 
                           sig_NPC_ABS_13_port, Z(12) => sig_NPC_ABS_12_port, 
                           Z(11) => sig_NPC_ABS_11_port, Z(10) => 
                           sig_NPC_ABS_10_port, Z(9) => sig_NPC_ABS_9_port, 
                           Z(8) => sig_NPC_ABS_8_port, Z(7) => 
                           sig_NPC_ABS_7_port, Z(6) => sig_NPC_ABS_6_port, Z(5)
                           => sig_NPC_ABS_5_port, Z(4) => sig_NPC_ABS_4_port, 
                           Z(3) => sig_NPC_ABS_3_port, Z(2) => 
                           sig_NPC_ABS_2_port, Z(1) => sig_NPC_ABS_1_port, Z(0)
                           => sig_NPC_ABS_0_port);
   FW2 : mux41_NBIT32_4 port map( A(31) => B_IN(31), A(30) => B_IN(30), A(29) 
                           => B_IN(29), A(28) => B_IN(28), A(27) => B_IN(27), 
                           A(26) => B_IN(26), A(25) => B_IN(25), A(24) => 
                           B_IN(24), A(23) => B_IN(23), A(22) => B_IN(22), 
                           A(21) => B_IN(21), A(20) => B_IN(20), A(19) => 
                           B_IN(19), A(18) => B_IN(18), A(17) => B_IN(17), 
                           A(16) => B_IN(16), A(15) => B_IN(15), A(14) => 
                           B_IN(14), A(13) => B_IN(13), A(12) => B_IN(12), 
                           A(11) => B_IN(11), A(10) => B_IN(10), A(9) => 
                           B_IN(9), A(8) => B_IN(8), A(7) => B_IN(7), A(6) => 
                           B_IN(6), A(5) => B_IN(5), A(4) => B_IN(4), A(3) => 
                           B_IN(3), A(2) => B_IN(2), A(1) => B_IN(1), A(0) => 
                           B_IN(0), B(31) => OP_WB(31), B(30) => OP_WB(30), 
                           B(29) => OP_WB(29), B(28) => OP_WB(28), B(27) => 
                           OP_WB(27), B(26) => OP_WB(26), B(25) => OP_WB(25), 
                           B(24) => OP_WB(24), B(23) => OP_WB(23), B(22) => 
                           OP_WB(22), B(21) => OP_WB(21), B(20) => OP_WB(20), 
                           B(19) => OP_WB(19), B(18) => OP_WB(18), B(17) => 
                           OP_WB(17), B(16) => OP_WB(16), B(15) => OP_WB(15), 
                           B(14) => OP_WB(14), B(13) => OP_WB(13), B(12) => 
                           OP_WB(12), B(11) => OP_WB(11), B(10) => OP_WB(10), 
                           B(9) => OP_WB(9), B(8) => OP_WB(8), B(7) => OP_WB(7)
                           , B(6) => OP_WB(6), B(5) => OP_WB(5), B(4) => 
                           OP_WB(4), B(3) => OP_WB(3), B(2) => OP_WB(2), B(1) 
                           => OP_WB(1), B(0) => OP_WB(0), C(31) => OP_MEM(31), 
                           C(30) => OP_MEM(30), C(29) => OP_MEM(29), C(28) => 
                           OP_MEM(28), C(27) => OP_MEM(27), C(26) => OP_MEM(26)
                           , C(25) => OP_MEM(25), C(24) => OP_MEM(24), C(23) =>
                           OP_MEM(23), C(22) => OP_MEM(22), C(21) => OP_MEM(21)
                           , C(20) => OP_MEM(20), C(19) => OP_MEM(19), C(18) =>
                           OP_MEM(18), C(17) => OP_MEM(17), C(16) => OP_MEM(16)
                           , C(15) => OP_MEM(15), C(14) => OP_MEM(14), C(13) =>
                           OP_MEM(13), C(12) => OP_MEM(12), C(11) => OP_MEM(11)
                           , C(10) => OP_MEM(10), C(9) => OP_MEM(9), C(8) => 
                           OP_MEM(8), C(7) => OP_MEM(7), C(6) => OP_MEM(6), 
                           C(5) => OP_MEM(5), C(4) => OP_MEM(4), C(3) => 
                           OP_MEM(3), C(2) => OP_MEM(2), C(1) => OP_MEM(1), 
                           C(0) => OP_MEM(0), D(31) => n6_port, D(30) => 
                           n6_port, D(29) => n6_port, D(28) => n6_port, D(27) 
                           => n6_port, D(26) => n6_port, D(25) => n6_port, 
                           D(24) => n6_port, D(23) => n6_port, D(22) => n6_port
                           , D(21) => n6_port, D(20) => n6_port, D(19) => 
                           n6_port, D(18) => n6_port, D(17) => n6_port, D(16) 
                           => n6_port, D(15) => n6_port, D(14) => n6_port, 
                           D(13) => n6_port, D(12) => n6_port, D(11) => n6_port
                           , D(10) => n6_port, D(9) => n6_port, D(8) => n6_port
                           , D(7) => n6_port, D(6) => n6_port, D(5) => n6_port,
                           D(4) => n6_port, D(3) => n6_port, D(2) => n6_port, 
                           D(1) => n6_port, D(0) => n6_port, S(1) => 
                           FWDB_1_port, S(0) => FWDB_0_port, Z(31) => 
                           OP2_FW_31_port, Z(30) => OP2_FW_30_port, Z(29) => 
                           OP2_FW_29_port, Z(28) => OP2_FW_28_port, Z(27) => 
                           OP2_FW_27_port, Z(26) => OP2_FW_26_port, Z(25) => 
                           OP2_FW_25_port, Z(24) => OP2_FW_24_port, Z(23) => 
                           OP2_FW_23_port, Z(22) => OP2_FW_22_port, Z(21) => 
                           OP2_FW_21_port, Z(20) => OP2_FW_20_port, Z(19) => 
                           OP2_FW_19_port, Z(18) => OP2_FW_18_port, Z(17) => 
                           OP2_FW_17_port, Z(16) => OP2_FW_16_port, Z(15) => 
                           OP2_FW_15_port, Z(14) => OP2_FW_14_port, Z(13) => 
                           OP2_FW_13_port, Z(12) => OP2_FW_12_port, Z(11) => 
                           OP2_FW_11_port, Z(10) => OP2_FW_10_port, Z(9) => 
                           OP2_FW_9_port, Z(8) => OP2_FW_8_port, Z(7) => 
                           OP2_FW_7_port, Z(6) => OP2_FW_6_port, Z(5) => 
                           OP2_FW_5_port, Z(4) => OP2_FW_4_port, Z(3) => 
                           OP2_FW_3_port, Z(2) => OP2_FW_2_port, Z(1) => 
                           OP2_FW_1_port, Z(0) => OP2_FW_0_port);
   muxA : mux21_NBIT32_3 port map( A(31) => sig_NPC_ABS_31_port, A(30) => 
                           sig_NPC_ABS_30_port, A(29) => sig_NPC_ABS_29_port, 
                           A(28) => sig_NPC_ABS_28_port, A(27) => 
                           sig_NPC_ABS_27_port, A(26) => sig_NPC_ABS_26_port, 
                           A(25) => sig_NPC_ABS_25_port, A(24) => 
                           sig_NPC_ABS_24_port, A(23) => sig_NPC_ABS_23_port, 
                           A(22) => sig_NPC_ABS_22_port, A(21) => 
                           sig_NPC_ABS_21_port, A(20) => sig_NPC_ABS_20_port, 
                           A(19) => sig_NPC_ABS_19_port, A(18) => 
                           sig_NPC_ABS_18_port, A(17) => sig_NPC_ABS_17_port, 
                           A(16) => sig_NPC_ABS_16_port, A(15) => 
                           sig_NPC_ABS_15_port, A(14) => sig_NPC_ABS_14_port, 
                           A(13) => sig_NPC_ABS_13_port, A(12) => 
                           sig_NPC_ABS_12_port, A(11) => sig_NPC_ABS_11_port, 
                           A(10) => sig_NPC_ABS_10_port, A(9) => 
                           sig_NPC_ABS_9_port, A(8) => sig_NPC_ABS_8_port, A(7)
                           => sig_NPC_ABS_7_port, A(6) => sig_NPC_ABS_6_port, 
                           A(5) => sig_NPC_ABS_5_port, A(4) => 
                           sig_NPC_ABS_4_port, A(3) => sig_NPC_ABS_3_port, A(2)
                           => sig_NPC_ABS_2_port, A(1) => sig_NPC_ABS_1_port, 
                           A(0) => sig_NPC_ABS_0_port, B(31) => PC_IN(31), 
                           B(30) => PC_IN(30), B(29) => PC_IN(29), B(28) => 
                           PC_IN(28), B(27) => PC_IN(27), B(26) => PC_IN(26), 
                           B(25) => PC_IN(25), B(24) => PC_IN(24), B(23) => 
                           PC_IN(23), B(22) => PC_IN(22), B(21) => PC_IN(21), 
                           B(20) => PC_IN(20), B(19) => PC_IN(19), B(18) => 
                           PC_IN(18), B(17) => PC_IN(17), B(16) => PC_IN(16), 
                           B(15) => PC_IN(15), B(14) => PC_IN(14), B(13) => 
                           PC_IN(13), B(12) => PC_IN(12), B(11) => PC_IN(11), 
                           B(10) => PC_IN(10), B(9) => PC_IN(9), B(8) => 
                           PC_IN(8), B(7) => PC_IN(7), B(6) => PC_IN(6), B(5) 
                           => PC_IN(5), B(4) => PC_IN(4), B(3) => PC_IN(3), 
                           B(2) => PC_IN(2), B(1) => PC_IN(1), B(0) => PC_IN(0)
                           , S => MUX_A_SEL, Z(31) => sig_OP1_31_port, Z(30) =>
                           sig_OP1_30_port, Z(29) => sig_OP1_29_port, Z(28) => 
                           sig_OP1_28_port, Z(27) => sig_OP1_27_port, Z(26) => 
                           sig_OP1_26_port, Z(25) => sig_OP1_25_port, Z(24) => 
                           sig_OP1_24_port, Z(23) => sig_OP1_23_port, Z(22) => 
                           sig_OP1_22_port, Z(21) => sig_OP1_21_port, Z(20) => 
                           sig_OP1_20_port, Z(19) => sig_OP1_19_port, Z(18) => 
                           sig_OP1_18_port, Z(17) => sig_OP1_17_port, Z(16) => 
                           sig_OP1_16_port, Z(15) => sig_OP1_15_port, Z(14) => 
                           sig_OP1_14_port, Z(13) => sig_OP1_13_port, Z(12) => 
                           sig_OP1_12_port, Z(11) => sig_OP1_11_port, Z(10) => 
                           sig_OP1_10_port, Z(9) => sig_OP1_9_port, Z(8) => 
                           sig_OP1_8_port, Z(7) => sig_OP1_7_port, Z(6) => 
                           sig_OP1_6_port, Z(5) => sig_OP1_5_port, Z(4) => 
                           sig_OP1_4_port, Z(3) => sig_OP1_3_port, Z(2) => 
                           sig_OP1_2_port, Z(1) => sig_OP1_1_port, Z(0) => 
                           sig_OP1_0_port);
   muxB : mux41_NBIT32_3 port map( A(31) => OP2_FW_31_port, A(30) => 
                           OP2_FW_30_port, A(29) => OP2_FW_29_port, A(28) => 
                           OP2_FW_28_port, A(27) => OP2_FW_27_port, A(26) => 
                           OP2_FW_26_port, A(25) => OP2_FW_25_port, A(24) => 
                           OP2_FW_24_port, A(23) => OP2_FW_23_port, A(22) => 
                           OP2_FW_22_port, A(21) => OP2_FW_21_port, A(20) => 
                           OP2_FW_20_port, A(19) => OP2_FW_19_port, A(18) => 
                           OP2_FW_18_port, A(17) => OP2_FW_17_port, A(16) => 
                           OP2_FW_16_port, A(15) => OP2_FW_15_port, A(14) => 
                           OP2_FW_14_port, A(13) => OP2_FW_13_port, A(12) => 
                           OP2_FW_12_port, A(11) => OP2_FW_11_port, A(10) => 
                           OP2_FW_10_port, A(9) => OP2_FW_9_port, A(8) => 
                           OP2_FW_8_port, A(7) => OP2_FW_7_port, A(6) => 
                           OP2_FW_6_port, A(5) => OP2_FW_5_port, A(4) => 
                           OP2_FW_4_port, A(3) => OP2_FW_3_port, A(2) => 
                           OP2_FW_2_port, A(1) => OP2_FW_1_port, A(0) => 
                           OP2_FW_0_port, B(31) => IMM_IN(31), B(30) => 
                           IMM_IN(30), B(29) => IMM_IN(29), B(28) => IMM_IN(28)
                           , B(27) => IMM_IN(27), B(26) => IMM_IN(26), B(25) =>
                           IMM_IN(25), B(24) => IMM_IN(24), B(23) => IMM_IN(23)
                           , B(22) => IMM_IN(22), B(21) => IMM_IN(21), B(20) =>
                           IMM_IN(20), B(19) => IMM_IN(19), B(18) => IMM_IN(18)
                           , B(17) => IMM_IN(17), B(16) => IMM_IN(16), B(15) =>
                           IMM_IN(15), B(14) => IMM_IN(14), B(13) => IMM_IN(13)
                           , B(12) => IMM_IN(12), B(11) => IMM_IN(11), B(10) =>
                           IMM_IN(10), B(9) => IMM_IN(9), B(8) => IMM_IN(8), 
                           B(7) => IMM_IN(7), B(6) => IMM_IN(6), B(5) => 
                           IMM_IN(5), B(4) => IMM_IN(4), B(3) => IMM_IN(3), 
                           B(2) => IMM_IN(2), B(1) => IMM_IN(1), B(0) => 
                           IMM_IN(0), C(31) => n6_port, C(30) => n6_port, C(29)
                           => n6_port, C(28) => n6_port, C(27) => n6_port, 
                           C(26) => n6_port, C(25) => n6_port, C(24) => n6_port
                           , C(23) => n6_port, C(22) => n6_port, C(21) => 
                           n6_port, C(20) => n6_port, C(19) => n6_port, C(18) 
                           => n6_port, C(17) => n6_port, C(16) => n6_port, 
                           C(15) => n6_port, C(14) => n6_port, C(13) => n6_port
                           , C(12) => n6_port, C(11) => n6_port, C(10) => 
                           n6_port, C(9) => n6_port, C(8) => n6_port, C(7) => 
                           n6_port, C(6) => n6_port, C(5) => n6_port, C(4) => 
                           n6_port, C(3) => n6_port, C(2) => n7_port, C(1) => 
                           n6_port, C(0) => n6_port, D(31) => n6_port, D(30) =>
                           n6_port, D(29) => n6_port, D(28) => n6_port, D(27) 
                           => n6_port, D(26) => n6_port, D(25) => n6_port, 
                           D(24) => n6_port, D(23) => n6_port, D(22) => n6_port
                           , D(21) => n6_port, D(20) => n6_port, D(19) => 
                           n6_port, D(18) => n6_port, D(17) => n6_port, D(16) 
                           => n6_port, D(15) => n6_port, D(14) => n6_port, 
                           D(13) => n6_port, D(12) => n6_port, D(11) => n6_port
                           , D(10) => n6_port, D(9) => n6_port, D(8) => n6_port
                           , D(7) => n6_port, D(6) => n6_port, D(5) => n6_port,
                           D(4) => n6_port, D(3) => n6_port, D(2) => n6_port, 
                           D(1) => n6_port, D(0) => n6_port, S(1) => 
                           MUX_B_SEL(1), S(0) => MUX_B_SEL(0), Z(31) => 
                           sig_OP2_31_port, Z(30) => sig_OP2_30_port, Z(29) => 
                           sig_OP2_29_port, Z(28) => sig_OP2_28_port, Z(27) => 
                           sig_OP2_27_port, Z(26) => sig_OP2_26_port, Z(25) => 
                           sig_OP2_25_port, Z(24) => sig_OP2_24_port, Z(23) => 
                           sig_OP2_23_port, Z(22) => sig_OP2_22_port, Z(21) => 
                           sig_OP2_21_port, Z(20) => sig_OP2_20_port, Z(19) => 
                           sig_OP2_19_port, Z(18) => sig_OP2_18_port, Z(17) => 
                           sig_OP2_17_port, Z(16) => sig_OP2_16_port, Z(15) => 
                           sig_OP2_15_port, Z(14) => sig_OP2_14_port, Z(13) => 
                           sig_OP2_13_port, Z(12) => sig_OP2_12_port, Z(11) => 
                           sig_OP2_11_port, Z(10) => sig_OP2_10_port, Z(9) => 
                           sig_OP2_9_port, Z(8) => sig_OP2_8_port, Z(7) => 
                           sig_OP2_7_port, Z(6) => sig_OP2_6_port, Z(5) => 
                           sig_OP2_5_port, Z(4) => sig_OP2_4_port, Z(3) => 
                           sig_OP2_3_port, Z(2) => sig_OP2_2_port, Z(1) => 
                           sig_OP2_1_port, Z(0) => sig_OP2_0_port);
   alu0 : ALU_NBIT32 port map( OP1(31) => sig_OP1_31_port, OP1(30) => 
                           sig_OP1_30_port, OP1(29) => sig_OP1_29_port, OP1(28)
                           => sig_OP1_28_port, OP1(27) => sig_OP1_27_port, 
                           OP1(26) => sig_OP1_26_port, OP1(25) => 
                           sig_OP1_25_port, OP1(24) => sig_OP1_24_port, OP1(23)
                           => sig_OP1_23_port, OP1(22) => sig_OP1_22_port, 
                           OP1(21) => sig_OP1_21_port, OP1(20) => 
                           sig_OP1_20_port, OP1(19) => sig_OP1_19_port, OP1(18)
                           => sig_OP1_18_port, OP1(17) => sig_OP1_17_port, 
                           OP1(16) => sig_OP1_16_port, OP1(15) => 
                           sig_OP1_15_port, OP1(14) => sig_OP1_14_port, OP1(13)
                           => sig_OP1_13_port, OP1(12) => sig_OP1_12_port, 
                           OP1(11) => sig_OP1_11_port, OP1(10) => 
                           sig_OP1_10_port, OP1(9) => sig_OP1_9_port, OP1(8) =>
                           sig_OP1_8_port, OP1(7) => sig_OP1_7_port, OP1(6) => 
                           sig_OP1_6_port, OP1(5) => sig_OP1_5_port, OP1(4) => 
                           sig_OP1_4_port, OP1(3) => sig_OP1_3_port, OP1(2) => 
                           sig_OP1_2_port, OP1(1) => sig_OP1_1_port, OP1(0) => 
                           sig_OP1_0_port, OP2(31) => sig_OP2_31_port, OP2(30) 
                           => sig_OP2_30_port, OP2(29) => sig_OP2_29_port, 
                           OP2(28) => sig_OP2_28_port, OP2(27) => 
                           sig_OP2_27_port, OP2(26) => sig_OP2_26_port, OP2(25)
                           => sig_OP2_25_port, OP2(24) => sig_OP2_24_port, 
                           OP2(23) => sig_OP2_23_port, OP2(22) => 
                           sig_OP2_22_port, OP2(21) => sig_OP2_21_port, OP2(20)
                           => sig_OP2_20_port, OP2(19) => sig_OP2_19_port, 
                           OP2(18) => sig_OP2_18_port, OP2(17) => 
                           sig_OP2_17_port, OP2(16) => sig_OP2_16_port, OP2(15)
                           => sig_OP2_15_port, OP2(14) => sig_OP2_14_port, 
                           OP2(13) => sig_OP2_13_port, OP2(12) => 
                           sig_OP2_12_port, OP2(11) => sig_OP2_11_port, OP2(10)
                           => sig_OP2_10_port, OP2(9) => sig_OP2_9_port, OP2(8)
                           => sig_OP2_8_port, OP2(7) => sig_OP2_7_port, OP2(6) 
                           => sig_OP2_6_port, OP2(5) => sig_OP2_5_port, OP2(4) 
                           => sig_OP2_4_port, OP2(3) => sig_OP2_3_port, OP2(2) 
                           => sig_OP2_2_port, OP2(1) => sig_OP2_1_port, OP2(0) 
                           => sig_OP2_0_port, ALU_OPC(0) => ALU_OPC(0), 
                           ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => ALU_OPC(2), 
                           ALU_OPC(3) => ALU_OPC(3), ALU_RES(31) => 
                           sig_ALU_RES_31_port, ALU_RES(30) => 
                           sig_ALU_RES_30_port, ALU_RES(29) => 
                           sig_ALU_RES_29_port, ALU_RES(28) => 
                           sig_ALU_RES_28_port, ALU_RES(27) => 
                           sig_ALU_RES_27_port, ALU_RES(26) => 
                           sig_ALU_RES_26_port, ALU_RES(25) => 
                           sig_ALU_RES_25_port, ALU_RES(24) => 
                           sig_ALU_RES_24_port, ALU_RES(23) => 
                           sig_ALU_RES_23_port, ALU_RES(22) => 
                           sig_ALU_RES_22_port, ALU_RES(21) => 
                           sig_ALU_RES_21_port, ALU_RES(20) => 
                           sig_ALU_RES_20_port, ALU_RES(19) => 
                           sig_ALU_RES_19_port, ALU_RES(18) => 
                           sig_ALU_RES_18_port, ALU_RES(17) => 
                           sig_ALU_RES_17_port, ALU_RES(16) => 
                           sig_ALU_RES_16_port, ALU_RES(15) => 
                           sig_ALU_RES_15_port, ALU_RES(14) => 
                           sig_ALU_RES_14_port, ALU_RES(13) => 
                           sig_ALU_RES_13_port, ALU_RES(12) => 
                           sig_ALU_RES_12_port, ALU_RES(11) => 
                           sig_ALU_RES_11_port, ALU_RES(10) => 
                           sig_ALU_RES_10_port, ALU_RES(9) => 
                           sig_ALU_RES_9_port, ALU_RES(8) => sig_ALU_RES_8_port
                           , ALU_RES(7) => sig_ALU_RES_7_port, ALU_RES(6) => 
                           sig_ALU_RES_6_port, ALU_RES(5) => sig_ALU_RES_5_port
                           , ALU_RES(4) => sig_ALU_RES_4_port, ALU_RES(3) => 
                           sig_ALU_RES_3_port, ALU_RES(2) => sig_ALU_RES_2_port
                           , ALU_RES(1) => sig_ALU_RES_1_port, ALU_RES(0) => 
                           sig_ALU_RES_0_port);
   alureg : regn_N32_6 port map( DIN(31) => sig_ALU_RES_31_port, DIN(30) => 
                           sig_ALU_RES_30_port, DIN(29) => sig_ALU_RES_29_port,
                           DIN(28) => sig_ALU_RES_28_port, DIN(27) => 
                           sig_ALU_RES_27_port, DIN(26) => sig_ALU_RES_26_port,
                           DIN(25) => sig_ALU_RES_25_port, DIN(24) => 
                           sig_ALU_RES_24_port, DIN(23) => sig_ALU_RES_23_port,
                           DIN(22) => sig_ALU_RES_22_port, DIN(21) => 
                           sig_ALU_RES_21_port, DIN(20) => sig_ALU_RES_20_port,
                           DIN(19) => sig_ALU_RES_19_port, DIN(18) => 
                           sig_ALU_RES_18_port, DIN(17) => sig_ALU_RES_17_port,
                           DIN(16) => sig_ALU_RES_16_port, DIN(15) => 
                           sig_ALU_RES_15_port, DIN(14) => sig_ALU_RES_14_port,
                           DIN(13) => sig_ALU_RES_13_port, DIN(12) => 
                           sig_ALU_RES_12_port, DIN(11) => sig_ALU_RES_11_port,
                           DIN(10) => sig_ALU_RES_10_port, DIN(9) => 
                           sig_ALU_RES_9_port, DIN(8) => sig_ALU_RES_8_port, 
                           DIN(7) => sig_ALU_RES_7_port, DIN(6) => 
                           sig_ALU_RES_6_port, DIN(5) => sig_ALU_RES_5_port, 
                           DIN(4) => sig_ALU_RES_4_port, DIN(3) => 
                           sig_ALU_RES_3_port, DIN(2) => sig_ALU_RES_2_port, 
                           DIN(1) => sig_ALU_RES_1_port, DIN(0) => 
                           sig_ALU_RES_0_port, CLK => CLK, EN => ALU_OUTREG_EN,
                           RST => RST, DOUT(31) => ALU_RES(31), DOUT(30) => 
                           ALU_RES(30), DOUT(29) => ALU_RES(29), DOUT(28) => 
                           ALU_RES(28), DOUT(27) => ALU_RES(27), DOUT(26) => 
                           ALU_RES(26), DOUT(25) => ALU_RES(25), DOUT(24) => 
                           ALU_RES(24), DOUT(23) => ALU_RES(23), DOUT(22) => 
                           ALU_RES(22), DOUT(21) => ALU_RES(21), DOUT(20) => 
                           ALU_RES(20), DOUT(19) => ALU_RES(19), DOUT(18) => 
                           ALU_RES(18), DOUT(17) => ALU_RES(17), DOUT(16) => 
                           ALU_RES(16), DOUT(15) => ALU_RES(15), DOUT(14) => 
                           ALU_RES(14), DOUT(13) => ALU_RES(13), DOUT(12) => 
                           ALU_RES(12), DOUT(11) => ALU_RES(11), DOUT(10) => 
                           ALU_RES(10), DOUT(9) => ALU_RES(9), DOUT(8) => 
                           ALU_RES(8), DOUT(7) => ALU_RES(7), DOUT(6) => 
                           ALU_RES(6), DOUT(5) => ALU_RES(5), DOUT(4) => 
                           ALU_RES(4), DOUT(3) => ALU_RES(3), DOUT(2) => 
                           ALU_RES(2), DOUT(1) => ALU_RES(1), DOUT(0) => 
                           ALU_RES(0));
   B_reg : regn_N32_5 port map( DIN(31) => OP2_FW_31_port, DIN(30) => 
                           OP2_FW_30_port, DIN(29) => OP2_FW_29_port, DIN(28) 
                           => OP2_FW_28_port, DIN(27) => OP2_FW_27_port, 
                           DIN(26) => OP2_FW_26_port, DIN(25) => OP2_FW_25_port
                           , DIN(24) => OP2_FW_24_port, DIN(23) => 
                           OP2_FW_23_port, DIN(22) => OP2_FW_22_port, DIN(21) 
                           => OP2_FW_21_port, DIN(20) => OP2_FW_20_port, 
                           DIN(19) => OP2_FW_19_port, DIN(18) => OP2_FW_18_port
                           , DIN(17) => OP2_FW_17_port, DIN(16) => 
                           OP2_FW_16_port, DIN(15) => OP2_FW_15_port, DIN(14) 
                           => OP2_FW_14_port, DIN(13) => OP2_FW_13_port, 
                           DIN(12) => OP2_FW_12_port, DIN(11) => OP2_FW_11_port
                           , DIN(10) => OP2_FW_10_port, DIN(9) => OP2_FW_9_port
                           , DIN(8) => OP2_FW_8_port, DIN(7) => OP2_FW_7_port, 
                           DIN(6) => OP2_FW_6_port, DIN(5) => OP2_FW_5_port, 
                           DIN(4) => OP2_FW_4_port, DIN(3) => OP2_FW_3_port, 
                           DIN(2) => OP2_FW_2_port, DIN(1) => OP2_FW_1_port, 
                           DIN(0) => OP2_FW_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => B_OUT(31), 
                           DOUT(30) => B_OUT(30), DOUT(29) => B_OUT(29), 
                           DOUT(28) => B_OUT(28), DOUT(27) => B_OUT(27), 
                           DOUT(26) => B_OUT(26), DOUT(25) => B_OUT(25), 
                           DOUT(24) => B_OUT(24), DOUT(23) => B_OUT(23), 
                           DOUT(22) => B_OUT(22), DOUT(21) => B_OUT(21), 
                           DOUT(20) => B_OUT(20), DOUT(19) => B_OUT(19), 
                           DOUT(18) => B_OUT(18), DOUT(17) => B_OUT(17), 
                           DOUT(16) => B_OUT(16), DOUT(15) => B_OUT(15), 
                           DOUT(14) => B_OUT(14), DOUT(13) => B_OUT(13), 
                           DOUT(12) => B_OUT(12), DOUT(11) => B_OUT(11), 
                           DOUT(10) => B_OUT(10), DOUT(9) => B_OUT(9), DOUT(8) 
                           => B_OUT(8), DOUT(7) => B_OUT(7), DOUT(6) => 
                           B_OUT(6), DOUT(5) => B_OUT(5), DOUT(4) => B_OUT(4), 
                           DOUT(3) => B_OUT(3), DOUT(2) => B_OUT(2), DOUT(1) =>
                           B_OUT(1), DOUT(0) => B_OUT(0));
   ADD_WR_reg : regn_N5_2 port map( DIN(4) => ADD_WR_IN(4), DIN(3) => 
                           ADD_WR_IN(3), DIN(2) => ADD_WR_IN(2), DIN(1) => 
                           ADD_WR_IN(1), DIN(0) => ADD_WR_IN(0), CLK => CLK, EN
                           => ALU_OUTREG_EN, RST => RST, DOUT(4) => 
                           ADD_WR_OUT(4), DOUT(3) => ADD_WR_OUT(3), DOUT(2) => 
                           ADD_WR_OUT(2), DOUT(1) => ADD_WR_OUT(1), DOUT(0) => 
                           ADD_WR_OUT(0));
   NPC_ABS_reg : regn_N32_4 port map( DIN(31) => sig_NPC_ABS_31_port, DIN(30) 
                           => sig_NPC_ABS_30_port, DIN(29) => 
                           sig_NPC_ABS_29_port, DIN(28) => sig_NPC_ABS_28_port,
                           DIN(27) => sig_NPC_ABS_27_port, DIN(26) => 
                           sig_NPC_ABS_26_port, DIN(25) => sig_NPC_ABS_25_port,
                           DIN(24) => sig_NPC_ABS_24_port, DIN(23) => 
                           sig_NPC_ABS_23_port, DIN(22) => sig_NPC_ABS_22_port,
                           DIN(21) => sig_NPC_ABS_21_port, DIN(20) => 
                           sig_NPC_ABS_20_port, DIN(19) => sig_NPC_ABS_19_port,
                           DIN(18) => sig_NPC_ABS_18_port, DIN(17) => 
                           sig_NPC_ABS_17_port, DIN(16) => sig_NPC_ABS_16_port,
                           DIN(15) => sig_NPC_ABS_15_port, DIN(14) => 
                           sig_NPC_ABS_14_port, DIN(13) => sig_NPC_ABS_13_port,
                           DIN(12) => sig_NPC_ABS_12_port, DIN(11) => 
                           sig_NPC_ABS_11_port, DIN(10) => sig_NPC_ABS_10_port,
                           DIN(9) => sig_NPC_ABS_9_port, DIN(8) => 
                           sig_NPC_ABS_8_port, DIN(7) => sig_NPC_ABS_7_port, 
                           DIN(6) => sig_NPC_ABS_6_port, DIN(5) => 
                           sig_NPC_ABS_5_port, DIN(4) => sig_NPC_ABS_4_port, 
                           DIN(3) => sig_NPC_ABS_3_port, DIN(2) => 
                           sig_NPC_ABS_2_port, DIN(1) => sig_NPC_ABS_1_port, 
                           DIN(0) => sig_NPC_ABS_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => NPC_ABS(31), 
                           DOUT(30) => NPC_ABS(30), DOUT(29) => NPC_ABS(29), 
                           DOUT(28) => NPC_ABS(28), DOUT(27) => NPC_ABS(27), 
                           DOUT(26) => NPC_ABS(26), DOUT(25) => NPC_ABS(25), 
                           DOUT(24) => NPC_ABS(24), DOUT(23) => NPC_ABS(23), 
                           DOUT(22) => NPC_ABS(22), DOUT(21) => NPC_ABS(21), 
                           DOUT(20) => NPC_ABS(20), DOUT(19) => NPC_ABS(19), 
                           DOUT(18) => NPC_ABS(18), DOUT(17) => NPC_ABS(17), 
                           DOUT(16) => NPC_ABS(16), DOUT(15) => NPC_ABS(15), 
                           DOUT(14) => NPC_ABS(14), DOUT(13) => NPC_ABS(13), 
                           DOUT(12) => NPC_ABS(12), DOUT(11) => NPC_ABS(11), 
                           DOUT(10) => NPC_ABS(10), DOUT(9) => NPC_ABS(9), 
                           DOUT(8) => NPC_ABS(8), DOUT(7) => NPC_ABS(7), 
                           DOUT(6) => NPC_ABS(6), DOUT(5) => NPC_ABS(5), 
                           DOUT(4) => NPC_ABS(4), DOUT(3) => NPC_ABS(3), 
                           DOUT(2) => NPC_ABS(2), DOUT(1) => NPC_ABS(1), 
                           DOUT(0) => NPC_ABS(0));
   NPC_REL_reg : regn_N32_3 port map( DIN(31) => sig_NPC_REL_31_port, DIN(30) 
                           => sig_NPC_REL_30_port, DIN(29) => 
                           sig_NPC_REL_29_port, DIN(28) => sig_NPC_REL_28_port,
                           DIN(27) => sig_NPC_REL_27_port, DIN(26) => 
                           sig_NPC_REL_26_port, DIN(25) => sig_NPC_REL_25_port,
                           DIN(24) => sig_NPC_REL_24_port, DIN(23) => 
                           sig_NPC_REL_23_port, DIN(22) => sig_NPC_REL_22_port,
                           DIN(21) => sig_NPC_REL_21_port, DIN(20) => 
                           sig_NPC_REL_20_port, DIN(19) => sig_NPC_REL_19_port,
                           DIN(18) => sig_NPC_REL_18_port, DIN(17) => 
                           sig_NPC_REL_17_port, DIN(16) => sig_NPC_REL_16_port,
                           DIN(15) => sig_NPC_REL_15_port, DIN(14) => 
                           sig_NPC_REL_14_port, DIN(13) => sig_NPC_REL_13_port,
                           DIN(12) => sig_NPC_REL_12_port, DIN(11) => 
                           sig_NPC_REL_11_port, DIN(10) => sig_NPC_REL_10_port,
                           DIN(9) => sig_NPC_REL_9_port, DIN(8) => 
                           sig_NPC_REL_8_port, DIN(7) => sig_NPC_REL_7_port, 
                           DIN(6) => sig_NPC_REL_6_port, DIN(5) => 
                           sig_NPC_REL_5_port, DIN(4) => sig_NPC_REL_4_port, 
                           DIN(3) => sig_NPC_REL_3_port, DIN(2) => 
                           sig_NPC_REL_2_port, DIN(1) => sig_NPC_REL_1_port, 
                           DIN(0) => sig_NPC_REL_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => NPC_REL(31), 
                           DOUT(30) => NPC_REL(30), DOUT(29) => NPC_REL(29), 
                           DOUT(28) => NPC_REL(28), DOUT(27) => NPC_REL(27), 
                           DOUT(26) => NPC_REL(26), DOUT(25) => NPC_REL(25), 
                           DOUT(24) => NPC_REL(24), DOUT(23) => NPC_REL(23), 
                           DOUT(22) => NPC_REL(22), DOUT(21) => NPC_REL(21), 
                           DOUT(20) => NPC_REL(20), DOUT(19) => NPC_REL(19), 
                           DOUT(18) => NPC_REL(18), DOUT(17) => NPC_REL(17), 
                           DOUT(16) => NPC_REL(16), DOUT(15) => NPC_REL(15), 
                           DOUT(14) => NPC_REL(14), DOUT(13) => NPC_REL(13), 
                           DOUT(12) => NPC_REL(12), DOUT(11) => NPC_REL(11), 
                           DOUT(10) => NPC_REL(10), DOUT(9) => NPC_REL(9), 
                           DOUT(8) => NPC_REL(8), DOUT(7) => NPC_REL(7), 
                           DOUT(6) => NPC_REL(6), DOUT(5) => NPC_REL(5), 
                           DOUT(4) => NPC_REL(4), DOUT(3) => NPC_REL(3), 
                           DOUT(2) => NPC_REL(2), DOUT(1) => NPC_REL(1), 
                           DOUT(0) => NPC_REL(0));
   add_1_root_add_0_root_add_118_2 : Execute_DW01_add_1 port map( A(31) => 
                           n2_port, A(30) => n2_port, A(29) => n2_port, A(28) 
                           => n2_port, A(27) => n2_port, A(26) => n2_port, 
                           A(25) => n2_port, A(24) => n2_port, A(23) => n2_port
                           , A(22) => n2_port, A(21) => n2_port, A(20) => 
                           n2_port, A(19) => n2_port, A(18) => n2_port, A(17) 
                           => n2_port, A(16) => n2_port, A(15) => n2_port, 
                           A(14) => n2_port, A(13) => n2_port, A(12) => n2_port
                           , A(11) => n2_port, A(10) => n2_port, A(9) => 
                           n2_port, A(8) => n2_port, A(7) => n2_port, A(6) => 
                           n2_port, A(5) => n2_port, A(4) => n2_port, A(3) => 
                           n2_port, A(2) => n3_port, A(1) => n2_port, A(0) => 
                           n2_port, B(31) => IMM_IN(31), B(30) => IMM_IN(30), 
                           B(29) => IMM_IN(29), B(28) => IMM_IN(28), B(27) => 
                           IMM_IN(27), B(26) => IMM_IN(26), B(25) => IMM_IN(25)
                           , B(24) => IMM_IN(24), B(23) => IMM_IN(23), B(22) =>
                           IMM_IN(22), B(21) => IMM_IN(21), B(20) => IMM_IN(20)
                           , B(19) => IMM_IN(19), B(18) => IMM_IN(18), B(17) =>
                           IMM_IN(17), B(16) => IMM_IN(16), B(15) => IMM_IN(15)
                           , B(14) => IMM_IN(14), B(13) => IMM_IN(13), B(12) =>
                           IMM_IN(12), B(11) => IMM_IN(11), B(10) => IMM_IN(10)
                           , B(9) => IMM_IN(9), B(8) => IMM_IN(8), B(7) => 
                           IMM_IN(7), B(6) => IMM_IN(6), B(5) => IMM_IN(5), 
                           B(4) => IMM_IN(4), B(3) => IMM_IN(3), B(2) => 
                           IMM_IN(2), B(1) => IMM_IN(1), B(0) => IMM_IN(0), CI 
                           => n4_port, SUM(31) => N31, SUM(30) => N30, SUM(29) 
                           => N29, SUM(28) => N28, SUM(27) => N27, SUM(26) => 
                           N26, SUM(25) => N25, SUM(24) => N24, SUM(23) => N23,
                           SUM(22) => N22, SUM(21) => N21, SUM(20) => N20, 
                           SUM(19) => N19, SUM(18) => N18, SUM(17) => N17, 
                           SUM(16) => N16, SUM(15) => N15, SUM(14) => N14, 
                           SUM(13) => N13, SUM(12) => N12, SUM(11) => N11, 
                           SUM(10) => N10, SUM(9) => N9, SUM(8) => N8, SUM(7) 
                           => N7, SUM(6) => N6, SUM(5) => N5, SUM(4) => N4, 
                           SUM(3) => N3, SUM(2) => N2, SUM(1) => N1, SUM(0) => 
                           N0, CO => n_1943);
   add_0_root_add_0_root_add_118_2 : Execute_DW01_add_0 port map( A(31) => 
                           PC_IN(31), A(30) => PC_IN(30), A(29) => PC_IN(29), 
                           A(28) => PC_IN(28), A(27) => PC_IN(27), A(26) => 
                           PC_IN(26), A(25) => PC_IN(25), A(24) => PC_IN(24), 
                           A(23) => PC_IN(23), A(22) => PC_IN(22), A(21) => 
                           PC_IN(21), A(20) => PC_IN(20), A(19) => PC_IN(19), 
                           A(18) => PC_IN(18), A(17) => PC_IN(17), A(16) => 
                           PC_IN(16), A(15) => PC_IN(15), A(14) => PC_IN(14), 
                           A(13) => PC_IN(13), A(12) => PC_IN(12), A(11) => 
                           PC_IN(11), A(10) => PC_IN(10), A(9) => PC_IN(9), 
                           A(8) => PC_IN(8), A(7) => PC_IN(7), A(6) => PC_IN(6)
                           , A(5) => PC_IN(5), A(4) => PC_IN(4), A(3) => 
                           PC_IN(3), A(2) => PC_IN(2), A(1) => PC_IN(1), A(0) 
                           => PC_IN(0), B(31) => N31, B(30) => N30, B(29) => 
                           N29, B(28) => N28, B(27) => N27, B(26) => N26, B(25)
                           => N25, B(24) => N24, B(23) => N23, B(22) => N22, 
                           B(21) => N21, B(20) => N20, B(19) => N19, B(18) => 
                           N18, B(17) => N17, B(16) => N16, B(15) => N15, B(14)
                           => N14, B(13) => N13, B(12) => N12, B(11) => N11, 
                           B(10) => N10, B(9) => N9, B(8) => N8, B(7) => N7, 
                           B(6) => N6, B(5) => N5, B(4) => N4, B(3) => N3, B(2)
                           => N2, B(1) => N1, B(0) => N0, CI => n5_port, 
                           SUM(31) => sig_NPC_REL_31_port, SUM(30) => 
                           sig_NPC_REL_30_port, SUM(29) => sig_NPC_REL_29_port,
                           SUM(28) => sig_NPC_REL_28_port, SUM(27) => 
                           sig_NPC_REL_27_port, SUM(26) => sig_NPC_REL_26_port,
                           SUM(25) => sig_NPC_REL_25_port, SUM(24) => 
                           sig_NPC_REL_24_port, SUM(23) => sig_NPC_REL_23_port,
                           SUM(22) => sig_NPC_REL_22_port, SUM(21) => 
                           sig_NPC_REL_21_port, SUM(20) => sig_NPC_REL_20_port,
                           SUM(19) => sig_NPC_REL_19_port, SUM(18) => 
                           sig_NPC_REL_18_port, SUM(17) => sig_NPC_REL_17_port,
                           SUM(16) => sig_NPC_REL_16_port, SUM(15) => 
                           sig_NPC_REL_15_port, SUM(14) => sig_NPC_REL_14_port,
                           SUM(13) => sig_NPC_REL_13_port, SUM(12) => 
                           sig_NPC_REL_12_port, SUM(11) => sig_NPC_REL_11_port,
                           SUM(10) => sig_NPC_REL_10_port, SUM(9) => 
                           sig_NPC_REL_9_port, SUM(8) => sig_NPC_REL_8_port, 
                           SUM(7) => sig_NPC_REL_7_port, SUM(6) => 
                           sig_NPC_REL_6_port, SUM(5) => sig_NPC_REL_5_port, 
                           SUM(4) => sig_NPC_REL_4_port, SUM(3) => 
                           sig_NPC_REL_3_port, SUM(2) => sig_NPC_REL_2_port, 
                           SUM(1) => sig_NPC_REL_1_port, SUM(0) => 
                           sig_NPC_REL_0_port, CO => n_1944);
   U3 : NOR2_X1 port map( A1 => ZERO_FLAG_port, A2 => n1_port, ZN => sig_RST);
   U4 : INV_X1 port map( A => RST, ZN => n1_port);
   n2_port <= '0';
   n3_port <= '1';
   n4_port <= '0';
   n5_port <= '0';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Decode is

   port( CLK, RST, REG_LATCH_EN, RD1, RD2, RF_WE, ZERO_FLAG : in std_logic;  
         PC_IN, INS_IN : in std_logic_vector (31 downto 0);  ADD_WR : in 
         std_logic_vector (4 downto 0);  DATA_WR_IN : in std_logic_vector (31 
         downto 0);  PC_OUT, A_OUT, B_OUT, IMM_OUT : out std_logic_vector (31 
         downto 0);  ADD_RS1_HDU, ADD_RS2_HDU, ADD_WR_OUT, ADD_RS1_OUT, 
         ADD_RS2_OUT : out std_logic_vector (4 downto 0));

end Decode;

architecture SYN_struct of Decode is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component register_file_NBIT_ADD5_NBIT_DATA32
      port( CLK, RST, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RS1, 
            ADD_RS2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component regn_N5_3
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N5_4
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N5_0
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N32_7
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_8
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component instruction_decomposition
      port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype :
            in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : out std_logic_vector (4 
            downto 0);  IMM : out std_logic_vector (31 downto 0));
   end component;
   
   component instruction_type
      port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype :
            out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic1_port, ADD_RS1_HDU_4_port, ADD_RS1_HDU_3_port, 
      ADD_RS1_HDU_2_port, ADD_RS1_HDU_1_port, ADD_RS1_HDU_0_port, 
      ADD_RS2_HDU_4_port, ADD_RS2_HDU_3_port, ADD_RS2_HDU_2_port, 
      ADD_RS2_HDU_1_port, ADD_RS2_HDU_0_port, sig_RST, sig_Rtype, sig_Itype, 
      sig_Jtype, sig_ADD_WR_4_port, sig_ADD_WR_3_port, sig_ADD_WR_2_port, 
      sig_ADD_WR_1_port, sig_ADD_WR_0_port, sig_IMM_31_port, sig_IMM_30_port, 
      sig_IMM_29_port, sig_IMM_28_port, sig_IMM_27_port, sig_IMM_26_port, 
      sig_IMM_25_port, sig_IMM_24_port, sig_IMM_23_port, sig_IMM_22_port, 
      sig_IMM_21_port, sig_IMM_20_port, sig_IMM_19_port, sig_IMM_18_port, 
      sig_IMM_17_port, sig_IMM_16_port, sig_IMM_15_port, sig_IMM_14_port, 
      sig_IMM_13_port, sig_IMM_12_port, sig_IMM_11_port, sig_IMM_10_port, 
      sig_IMM_9_port, sig_IMM_8_port, sig_IMM_7_port, sig_IMM_6_port, 
      sig_IMM_5_port, sig_IMM_4_port, sig_IMM_3_port, sig_IMM_2_port, 
      sig_IMM_1_port, sig_IMM_0_port, n1 : std_logic;

begin
   ADD_RS1_HDU <= ( ADD_RS1_HDU_4_port, ADD_RS1_HDU_3_port, ADD_RS1_HDU_2_port,
      ADD_RS1_HDU_1_port, ADD_RS1_HDU_0_port );
   ADD_RS2_HDU <= ( ADD_RS2_HDU_4_port, ADD_RS2_HDU_3_port, ADD_RS2_HDU_2_port,
      ADD_RS2_HDU_1_port, ADD_RS2_HDU_0_port );
   
   X_Logic1_port <= '1';
   U2 : NOR2_X2 port map( A1 => ZERO_FLAG, A2 => n1, ZN => sig_RST);
   ins_type : instruction_type port map( INST_IN(31) => INS_IN(31), INST_IN(30)
                           => INS_IN(30), INST_IN(29) => INS_IN(29), 
                           INST_IN(28) => INS_IN(28), INST_IN(27) => INS_IN(27)
                           , INST_IN(26) => INS_IN(26), INST_IN(25) => 
                           INS_IN(25), INST_IN(24) => INS_IN(24), INST_IN(23) 
                           => INS_IN(23), INST_IN(22) => INS_IN(22), 
                           INST_IN(21) => INS_IN(21), INST_IN(20) => INS_IN(20)
                           , INST_IN(19) => INS_IN(19), INST_IN(18) => 
                           INS_IN(18), INST_IN(17) => INS_IN(17), INST_IN(16) 
                           => INS_IN(16), INST_IN(15) => INS_IN(15), 
                           INST_IN(14) => INS_IN(14), INST_IN(13) => INS_IN(13)
                           , INST_IN(12) => INS_IN(12), INST_IN(11) => 
                           INS_IN(11), INST_IN(10) => INS_IN(10), INST_IN(9) =>
                           INS_IN(9), INST_IN(8) => INS_IN(8), INST_IN(7) => 
                           INS_IN(7), INST_IN(6) => INS_IN(6), INST_IN(5) => 
                           INS_IN(5), INST_IN(4) => INS_IN(4), INST_IN(3) => 
                           INS_IN(3), INST_IN(2) => INS_IN(2), INST_IN(1) => 
                           INS_IN(1), INST_IN(0) => INS_IN(0), Rtype => 
                           sig_Rtype, Itype => sig_Itype, Jtype => sig_Jtype);
   ins_dec : instruction_decomposition port map( INST_IN(31) => INS_IN(31), 
                           INST_IN(30) => INS_IN(30), INST_IN(29) => INS_IN(29)
                           , INST_IN(28) => INS_IN(28), INST_IN(27) => 
                           INS_IN(27), INST_IN(26) => INS_IN(26), INST_IN(25) 
                           => INS_IN(25), INST_IN(24) => INS_IN(24), 
                           INST_IN(23) => INS_IN(23), INST_IN(22) => INS_IN(22)
                           , INST_IN(21) => INS_IN(21), INST_IN(20) => 
                           INS_IN(20), INST_IN(19) => INS_IN(19), INST_IN(18) 
                           => INS_IN(18), INST_IN(17) => INS_IN(17), 
                           INST_IN(16) => INS_IN(16), INST_IN(15) => INS_IN(15)
                           , INST_IN(14) => INS_IN(14), INST_IN(13) => 
                           INS_IN(13), INST_IN(12) => INS_IN(12), INST_IN(11) 
                           => INS_IN(11), INST_IN(10) => INS_IN(10), INST_IN(9)
                           => INS_IN(9), INST_IN(8) => INS_IN(8), INST_IN(7) =>
                           INS_IN(7), INST_IN(6) => INS_IN(6), INST_IN(5) => 
                           INS_IN(5), INST_IN(4) => INS_IN(4), INST_IN(3) => 
                           INS_IN(3), INST_IN(2) => INS_IN(2), INST_IN(1) => 
                           INS_IN(1), INST_IN(0) => INS_IN(0), Rtype => 
                           sig_Rtype, Itype => sig_Itype, Jtype => sig_Jtype, 
                           ADD_RS1(4) => ADD_RS1_HDU_4_port, ADD_RS1(3) => 
                           ADD_RS1_HDU_3_port, ADD_RS1(2) => ADD_RS1_HDU_2_port
                           , ADD_RS1(1) => ADD_RS1_HDU_1_port, ADD_RS1(0) => 
                           ADD_RS1_HDU_0_port, ADD_RS2(4) => ADD_RS2_HDU_4_port
                           , ADD_RS2(3) => ADD_RS2_HDU_3_port, ADD_RS2(2) => 
                           ADD_RS2_HDU_2_port, ADD_RS2(1) => ADD_RS2_HDU_1_port
                           , ADD_RS2(0) => ADD_RS2_HDU_0_port, ADD_WR(4) => 
                           sig_ADD_WR_4_port, ADD_WR(3) => sig_ADD_WR_3_port, 
                           ADD_WR(2) => sig_ADD_WR_2_port, ADD_WR(1) => 
                           sig_ADD_WR_1_port, ADD_WR(0) => sig_ADD_WR_0_port, 
                           IMM(31) => sig_IMM_31_port, IMM(30) => 
                           sig_IMM_30_port, IMM(29) => sig_IMM_29_port, IMM(28)
                           => sig_IMM_28_port, IMM(27) => sig_IMM_27_port, 
                           IMM(26) => sig_IMM_26_port, IMM(25) => 
                           sig_IMM_25_port, IMM(24) => sig_IMM_24_port, IMM(23)
                           => sig_IMM_23_port, IMM(22) => sig_IMM_22_port, 
                           IMM(21) => sig_IMM_21_port, IMM(20) => 
                           sig_IMM_20_port, IMM(19) => sig_IMM_19_port, IMM(18)
                           => sig_IMM_18_port, IMM(17) => sig_IMM_17_port, 
                           IMM(16) => sig_IMM_16_port, IMM(15) => 
                           sig_IMM_15_port, IMM(14) => sig_IMM_14_port, IMM(13)
                           => sig_IMM_13_port, IMM(12) => sig_IMM_12_port, 
                           IMM(11) => sig_IMM_11_port, IMM(10) => 
                           sig_IMM_10_port, IMM(9) => sig_IMM_9_port, IMM(8) =>
                           sig_IMM_8_port, IMM(7) => sig_IMM_7_port, IMM(6) => 
                           sig_IMM_6_port, IMM(5) => sig_IMM_5_port, IMM(4) => 
                           sig_IMM_4_port, IMM(3) => sig_IMM_3_port, IMM(2) => 
                           sig_IMM_2_port, IMM(1) => sig_IMM_1_port, IMM(0) => 
                           sig_IMM_0_port);
   regPC : regn_N32_8 port map( DIN(31) => PC_IN(31), DIN(30) => PC_IN(30), 
                           DIN(29) => PC_IN(29), DIN(28) => PC_IN(28), DIN(27) 
                           => PC_IN(27), DIN(26) => PC_IN(26), DIN(25) => 
                           PC_IN(25), DIN(24) => PC_IN(24), DIN(23) => 
                           PC_IN(23), DIN(22) => PC_IN(22), DIN(21) => 
                           PC_IN(21), DIN(20) => PC_IN(20), DIN(19) => 
                           PC_IN(19), DIN(18) => PC_IN(18), DIN(17) => 
                           PC_IN(17), DIN(16) => PC_IN(16), DIN(15) => 
                           PC_IN(15), DIN(14) => PC_IN(14), DIN(13) => 
                           PC_IN(13), DIN(12) => PC_IN(12), DIN(11) => 
                           PC_IN(11), DIN(10) => PC_IN(10), DIN(9) => PC_IN(9),
                           DIN(8) => PC_IN(8), DIN(7) => PC_IN(7), DIN(6) => 
                           PC_IN(6), DIN(5) => PC_IN(5), DIN(4) => PC_IN(4), 
                           DIN(3) => PC_IN(3), DIN(2) => PC_IN(2), DIN(1) => 
                           PC_IN(1), DIN(0) => PC_IN(0), CLK => CLK, EN => 
                           X_Logic1_port, RST => sig_RST, DOUT(31) => 
                           PC_OUT(31), DOUT(30) => PC_OUT(30), DOUT(29) => 
                           PC_OUT(29), DOUT(28) => PC_OUT(28), DOUT(27) => 
                           PC_OUT(27), DOUT(26) => PC_OUT(26), DOUT(25) => 
                           PC_OUT(25), DOUT(24) => PC_OUT(24), DOUT(23) => 
                           PC_OUT(23), DOUT(22) => PC_OUT(22), DOUT(21) => 
                           PC_OUT(21), DOUT(20) => PC_OUT(20), DOUT(19) => 
                           PC_OUT(19), DOUT(18) => PC_OUT(18), DOUT(17) => 
                           PC_OUT(17), DOUT(16) => PC_OUT(16), DOUT(15) => 
                           PC_OUT(15), DOUT(14) => PC_OUT(14), DOUT(13) => 
                           PC_OUT(13), DOUT(12) => PC_OUT(12), DOUT(11) => 
                           PC_OUT(11), DOUT(10) => PC_OUT(10), DOUT(9) => 
                           PC_OUT(9), DOUT(8) => PC_OUT(8), DOUT(7) => 
                           PC_OUT(7), DOUT(6) => PC_OUT(6), DOUT(5) => 
                           PC_OUT(5), DOUT(4) => PC_OUT(4), DOUT(3) => 
                           PC_OUT(3), DOUT(2) => PC_OUT(2), DOUT(1) => 
                           PC_OUT(1), DOUT(0) => PC_OUT(0));
   regIMM : regn_N32_7 port map( DIN(31) => sig_IMM_31_port, DIN(30) => 
                           sig_IMM_30_port, DIN(29) => sig_IMM_29_port, DIN(28)
                           => sig_IMM_28_port, DIN(27) => sig_IMM_27_port, 
                           DIN(26) => sig_IMM_26_port, DIN(25) => 
                           sig_IMM_25_port, DIN(24) => sig_IMM_24_port, DIN(23)
                           => sig_IMM_23_port, DIN(22) => sig_IMM_22_port, 
                           DIN(21) => sig_IMM_21_port, DIN(20) => 
                           sig_IMM_20_port, DIN(19) => sig_IMM_19_port, DIN(18)
                           => sig_IMM_18_port, DIN(17) => sig_IMM_17_port, 
                           DIN(16) => sig_IMM_16_port, DIN(15) => 
                           sig_IMM_15_port, DIN(14) => sig_IMM_14_port, DIN(13)
                           => sig_IMM_13_port, DIN(12) => sig_IMM_12_port, 
                           DIN(11) => sig_IMM_11_port, DIN(10) => 
                           sig_IMM_10_port, DIN(9) => sig_IMM_9_port, DIN(8) =>
                           sig_IMM_8_port, DIN(7) => sig_IMM_7_port, DIN(6) => 
                           sig_IMM_6_port, DIN(5) => sig_IMM_5_port, DIN(4) => 
                           sig_IMM_4_port, DIN(3) => sig_IMM_3_port, DIN(2) => 
                           sig_IMM_2_port, DIN(1) => sig_IMM_1_port, DIN(0) => 
                           sig_IMM_0_port, CLK => CLK, EN => REG_LATCH_EN, RST 
                           => sig_RST, DOUT(31) => IMM_OUT(31), DOUT(30) => 
                           IMM_OUT(30), DOUT(29) => IMM_OUT(29), DOUT(28) => 
                           IMM_OUT(28), DOUT(27) => IMM_OUT(27), DOUT(26) => 
                           IMM_OUT(26), DOUT(25) => IMM_OUT(25), DOUT(24) => 
                           IMM_OUT(24), DOUT(23) => IMM_OUT(23), DOUT(22) => 
                           IMM_OUT(22), DOUT(21) => IMM_OUT(21), DOUT(20) => 
                           IMM_OUT(20), DOUT(19) => IMM_OUT(19), DOUT(18) => 
                           IMM_OUT(18), DOUT(17) => IMM_OUT(17), DOUT(16) => 
                           IMM_OUT(16), DOUT(15) => IMM_OUT(15), DOUT(14) => 
                           IMM_OUT(14), DOUT(13) => IMM_OUT(13), DOUT(12) => 
                           IMM_OUT(12), DOUT(11) => IMM_OUT(11), DOUT(10) => 
                           IMM_OUT(10), DOUT(9) => IMM_OUT(9), DOUT(8) => 
                           IMM_OUT(8), DOUT(7) => IMM_OUT(7), DOUT(6) => 
                           IMM_OUT(6), DOUT(5) => IMM_OUT(5), DOUT(4) => 
                           IMM_OUT(4), DOUT(3) => IMM_OUT(3), DOUT(2) => 
                           IMM_OUT(2), DOUT(1) => IMM_OUT(1), DOUT(0) => 
                           IMM_OUT(0));
   regWR : regn_N5_0 port map( DIN(4) => sig_ADD_WR_4_port, DIN(3) => 
                           sig_ADD_WR_3_port, DIN(2) => sig_ADD_WR_2_port, 
                           DIN(1) => sig_ADD_WR_1_port, DIN(0) => 
                           sig_ADD_WR_0_port, CLK => CLK, EN => REG_LATCH_EN, 
                           RST => sig_RST, DOUT(4) => ADD_WR_OUT(4), DOUT(3) =>
                           ADD_WR_OUT(3), DOUT(2) => ADD_WR_OUT(2), DOUT(1) => 
                           ADD_WR_OUT(1), DOUT(0) => ADD_WR_OUT(0));
   regRS1 : regn_N5_4 port map( DIN(4) => ADD_RS1_HDU_4_port, DIN(3) => 
                           ADD_RS1_HDU_3_port, DIN(2) => ADD_RS1_HDU_2_port, 
                           DIN(1) => ADD_RS1_HDU_1_port, DIN(0) => 
                           ADD_RS1_HDU_0_port, CLK => CLK, EN => REG_LATCH_EN, 
                           RST => sig_RST, DOUT(4) => ADD_RS1_OUT(4), DOUT(3) 
                           => ADD_RS1_OUT(3), DOUT(2) => ADD_RS1_OUT(2), 
                           DOUT(1) => ADD_RS1_OUT(1), DOUT(0) => ADD_RS1_OUT(0)
                           );
   regRS2 : regn_N5_3 port map( DIN(4) => ADD_RS2_HDU_4_port, DIN(3) => 
                           ADD_RS2_HDU_3_port, DIN(2) => ADD_RS2_HDU_2_port, 
                           DIN(1) => ADD_RS2_HDU_1_port, DIN(0) => 
                           ADD_RS2_HDU_0_port, CLK => CLK, EN => REG_LATCH_EN, 
                           RST => sig_RST, DOUT(4) => ADD_RS2_OUT(4), DOUT(3) 
                           => ADD_RS2_OUT(3), DOUT(2) => ADD_RS2_OUT(2), 
                           DOUT(1) => ADD_RS2_OUT(1), DOUT(0) => ADD_RS2_OUT(0)
                           );
   rf : register_file_NBIT_ADD5_NBIT_DATA32 port map( CLK => CLK, RST => RST, 
                           ENABLE => REG_LATCH_EN, RD1 => RD1, RD2 => RD2, WR 
                           => RF_WE, ADD_WR(4) => ADD_WR(4), ADD_WR(3) => 
                           ADD_WR(3), ADD_WR(2) => ADD_WR(2), ADD_WR(1) => 
                           ADD_WR(1), ADD_WR(0) => ADD_WR(0), ADD_RS1(4) => 
                           ADD_RS1_HDU_4_port, ADD_RS1(3) => ADD_RS1_HDU_3_port
                           , ADD_RS1(2) => ADD_RS1_HDU_2_port, ADD_RS1(1) => 
                           ADD_RS1_HDU_1_port, ADD_RS1(0) => ADD_RS1_HDU_0_port
                           , ADD_RS2(4) => ADD_RS2_HDU_4_port, ADD_RS2(3) => 
                           ADD_RS2_HDU_3_port, ADD_RS2(2) => ADD_RS2_HDU_2_port
                           , ADD_RS2(1) => ADD_RS2_HDU_1_port, ADD_RS2(0) => 
                           ADD_RS2_HDU_0_port, DATAIN(31) => DATA_WR_IN(31), 
                           DATAIN(30) => DATA_WR_IN(30), DATAIN(29) => 
                           DATA_WR_IN(29), DATAIN(28) => DATA_WR_IN(28), 
                           DATAIN(27) => DATA_WR_IN(27), DATAIN(26) => 
                           DATA_WR_IN(26), DATAIN(25) => DATA_WR_IN(25), 
                           DATAIN(24) => DATA_WR_IN(24), DATAIN(23) => 
                           DATA_WR_IN(23), DATAIN(22) => DATA_WR_IN(22), 
                           DATAIN(21) => DATA_WR_IN(21), DATAIN(20) => 
                           DATA_WR_IN(20), DATAIN(19) => DATA_WR_IN(19), 
                           DATAIN(18) => DATA_WR_IN(18), DATAIN(17) => 
                           DATA_WR_IN(17), DATAIN(16) => DATA_WR_IN(16), 
                           DATAIN(15) => DATA_WR_IN(15), DATAIN(14) => 
                           DATA_WR_IN(14), DATAIN(13) => DATA_WR_IN(13), 
                           DATAIN(12) => DATA_WR_IN(12), DATAIN(11) => 
                           DATA_WR_IN(11), DATAIN(10) => DATA_WR_IN(10), 
                           DATAIN(9) => DATA_WR_IN(9), DATAIN(8) => 
                           DATA_WR_IN(8), DATAIN(7) => DATA_WR_IN(7), DATAIN(6)
                           => DATA_WR_IN(6), DATAIN(5) => DATA_WR_IN(5), 
                           DATAIN(4) => DATA_WR_IN(4), DATAIN(3) => 
                           DATA_WR_IN(3), DATAIN(2) => DATA_WR_IN(2), DATAIN(1)
                           => DATA_WR_IN(1), DATAIN(0) => DATA_WR_IN(0), 
                           OUT1(31) => A_OUT(31), OUT1(30) => A_OUT(30), 
                           OUT1(29) => A_OUT(29), OUT1(28) => A_OUT(28), 
                           OUT1(27) => A_OUT(27), OUT1(26) => A_OUT(26), 
                           OUT1(25) => A_OUT(25), OUT1(24) => A_OUT(24), 
                           OUT1(23) => A_OUT(23), OUT1(22) => A_OUT(22), 
                           OUT1(21) => A_OUT(21), OUT1(20) => A_OUT(20), 
                           OUT1(19) => A_OUT(19), OUT1(18) => A_OUT(18), 
                           OUT1(17) => A_OUT(17), OUT1(16) => A_OUT(16), 
                           OUT1(15) => A_OUT(15), OUT1(14) => A_OUT(14), 
                           OUT1(13) => A_OUT(13), OUT1(12) => A_OUT(12), 
                           OUT1(11) => A_OUT(11), OUT1(10) => A_OUT(10), 
                           OUT1(9) => A_OUT(9), OUT1(8) => A_OUT(8), OUT1(7) =>
                           A_OUT(7), OUT1(6) => A_OUT(6), OUT1(5) => A_OUT(5), 
                           OUT1(4) => A_OUT(4), OUT1(3) => A_OUT(3), OUT1(2) =>
                           A_OUT(2), OUT1(1) => A_OUT(1), OUT1(0) => A_OUT(0), 
                           OUT2(31) => B_OUT(31), OUT2(30) => B_OUT(30), 
                           OUT2(29) => B_OUT(29), OUT2(28) => B_OUT(28), 
                           OUT2(27) => B_OUT(27), OUT2(26) => B_OUT(26), 
                           OUT2(25) => B_OUT(25), OUT2(24) => B_OUT(24), 
                           OUT2(23) => B_OUT(23), OUT2(22) => B_OUT(22), 
                           OUT2(21) => B_OUT(21), OUT2(20) => B_OUT(20), 
                           OUT2(19) => B_OUT(19), OUT2(18) => B_OUT(18), 
                           OUT2(17) => B_OUT(17), OUT2(16) => B_OUT(16), 
                           OUT2(15) => B_OUT(15), OUT2(14) => B_OUT(14), 
                           OUT2(13) => B_OUT(13), OUT2(12) => B_OUT(12), 
                           OUT2(11) => B_OUT(11), OUT2(10) => B_OUT(10), 
                           OUT2(9) => B_OUT(9), OUT2(8) => B_OUT(8), OUT2(7) =>
                           B_OUT(7), OUT2(6) => B_OUT(6), OUT2(5) => B_OUT(5), 
                           OUT2(4) => B_OUT(4), OUT2(3) => B_OUT(3), OUT2(2) =>
                           B_OUT(2), OUT2(1) => B_OUT(1), OUT2(0) => B_OUT(0));
   U3 : INV_X1 port map( A => RST, ZN => n1);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Fetch is

   port( CLK, RST, ZERO_FLAG : in std_logic;  PC_EXT, INS_IN : in 
         std_logic_vector (31 downto 0);  Bubble_in : in std_logic;  HDU_INS_IN
         , HDU_PC_IN, HDU_NPC_IN : in std_logic_vector (31 downto 0);  PC_OUT, 
         ADDR_OUT, NPC_OUT, INS_OUT : out std_logic_vector (31 downto 0));

end Fetch;

architecture SYN_struct of Fetch is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component Fetch_DW01_add_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component regn_N32_9
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_10
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_0
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, ADDR_OUT_31_port, ADDR_OUT_30_port, n19, 
      ADDR_OUT_28_port, ADDR_OUT_27_port, ADDR_OUT_26_port, ADDR_OUT_25_port, 
      ADDR_OUT_24_port, n20, ADDR_OUT_22_port, ADDR_OUT_21_port, 
      ADDR_OUT_20_port, ADDR_OUT_19_port, ADDR_OUT_18_port, n21, n22, 
      ADDR_OUT_15_port, n23, ADDR_OUT_13_port, n24, ADDR_OUT_11_port, 
      ADDR_OUT_10_port, n25, n26, n27, n28, n29, n30, n31, n32, ADDR_OUT_1_port
      , ADDR_OUT_0_port, sig_RST, sig_NPC_31_port, sig_NPC_30_port, 
      sig_NPC_29_port, sig_NPC_28_port, sig_NPC_27_port, sig_NPC_26_port, 
      sig_NPC_25_port, sig_NPC_24_port, sig_NPC_23_port, sig_NPC_22_port, 
      sig_NPC_21_port, sig_NPC_20_port, sig_NPC_19_port, sig_NPC_18_port, 
      sig_NPC_17_port, sig_NPC_16_port, sig_NPC_15_port, sig_NPC_14_port, 
      sig_NPC_13_port, sig_NPC_12_port, sig_NPC_11_port, sig_NPC_10_port, 
      sig_NPC_9_port, sig_NPC_8_port, sig_NPC_7_port, sig_NPC_6_port, 
      sig_NPC_5_port, sig_NPC_4_port, sig_NPC_3_port, sig_NPC_2_port, 
      sig_NPC_1_port, sig_NPC_0_port, PC_MUX_OUT_31_port, PC_MUX_OUT_30_port, 
      PC_MUX_OUT_29_port, PC_MUX_OUT_28_port, PC_MUX_OUT_27_port, 
      PC_MUX_OUT_26_port, PC_MUX_OUT_25_port, PC_MUX_OUT_24_port, 
      PC_MUX_OUT_23_port, PC_MUX_OUT_22_port, PC_MUX_OUT_21_port, 
      PC_MUX_OUT_20_port, PC_MUX_OUT_19_port, PC_MUX_OUT_18_port, 
      PC_MUX_OUT_17_port, PC_MUX_OUT_16_port, PC_MUX_OUT_15_port, 
      PC_MUX_OUT_14_port, PC_MUX_OUT_13_port, PC_MUX_OUT_12_port, 
      PC_MUX_OUT_11_port, PC_MUX_OUT_10_port, PC_MUX_OUT_9_port, 
      PC_MUX_OUT_8_port, PC_MUX_OUT_7_port, PC_MUX_OUT_6_port, 
      PC_MUX_OUT_5_port, PC_MUX_OUT_4_port, PC_MUX_OUT_3_port, 
      PC_MUX_OUT_2_port, PC_MUX_OUT_1_port, PC_MUX_OUT_0_port, sig_INS_31_port,
      sig_INS_30_port, sig_INS_29_port, sig_INS_28_port, sig_INS_27_port, 
      sig_INS_26_port, sig_INS_25_port, sig_INS_24_port, sig_INS_23_port, 
      sig_INS_22_port, sig_INS_21_port, sig_INS_20_port, sig_INS_19_port, 
      sig_INS_18_port, sig_INS_17_port, sig_INS_16_port, sig_INS_15_port, 
      sig_INS_14_port, sig_INS_13_port, sig_INS_12_port, sig_INS_11_port, 
      sig_INS_10_port, sig_INS_9_port, sig_INS_8_port, sig_INS_7_port, 
      sig_INS_6_port, sig_INS_5_port, sig_INS_4_port, sig_INS_3_port, 
      sig_INS_2_port, sig_INS_1_port, sig_INS_0_port, n1, n2, n3, 
      ADDR_OUT_8_port, ADDR_OUT_29_port, ADDR_OUT_7_port, ADDR_OUT_2_port, 
      ADDR_OUT_23_port, ADDR_OUT_12_port, ADDR_OUT_6_port, ADDR_OUT_3_port, 
      ADDR_OUT_17_port, ADDR_OUT_16_port, ADDR_OUT_5_port, ADDR_OUT_14_port, 
      ADDR_OUT_4_port, ADDR_OUT_9_port, n18, n_1945 : std_logic;

begin
   ADDR_OUT <= ( ADDR_OUT_31_port, ADDR_OUT_30_port, ADDR_OUT_29_port, 
      ADDR_OUT_28_port, ADDR_OUT_27_port, ADDR_OUT_26_port, ADDR_OUT_25_port, 
      ADDR_OUT_24_port, ADDR_OUT_23_port, ADDR_OUT_22_port, ADDR_OUT_21_port, 
      ADDR_OUT_20_port, ADDR_OUT_19_port, ADDR_OUT_18_port, ADDR_OUT_17_port, 
      ADDR_OUT_16_port, ADDR_OUT_15_port, ADDR_OUT_14_port, ADDR_OUT_13_port, 
      ADDR_OUT_12_port, ADDR_OUT_11_port, ADDR_OUT_10_port, ADDR_OUT_9_port, 
      ADDR_OUT_8_port, ADDR_OUT_7_port, ADDR_OUT_6_port, ADDR_OUT_5_port, 
      ADDR_OUT_4_port, ADDR_OUT_3_port, ADDR_OUT_2_port, ADDR_OUT_1_port, 
      ADDR_OUT_0_port );
   
   X_Logic1_port <= '1';
   n1 <= '0';
   n2 <= '1';
   n3 <= '0';
   NPC_or_NPC_HDU : mux21_NBIT32_0 port map( A(31) => PC_EXT(31), A(30) => 
                           PC_EXT(30), A(29) => PC_EXT(29), A(28) => PC_EXT(28)
                           , A(27) => PC_EXT(27), A(26) => PC_EXT(26), A(25) =>
                           PC_EXT(25), A(24) => PC_EXT(24), A(23) => PC_EXT(23)
                           , A(22) => PC_EXT(22), A(21) => PC_EXT(21), A(20) =>
                           PC_EXT(20), A(19) => PC_EXT(19), A(18) => PC_EXT(18)
                           , A(17) => PC_EXT(17), A(16) => PC_EXT(16), A(15) =>
                           PC_EXT(15), A(14) => PC_EXT(14), A(13) => PC_EXT(13)
                           , A(12) => PC_EXT(12), A(11) => PC_EXT(11), A(10) =>
                           PC_EXT(10), A(9) => PC_EXT(9), A(8) => PC_EXT(8), 
                           A(7) => PC_EXT(7), A(6) => PC_EXT(6), A(5) => 
                           PC_EXT(5), A(4) => PC_EXT(4), A(3) => PC_EXT(3), 
                           A(2) => PC_EXT(2), A(1) => PC_EXT(1), A(0) => 
                           PC_EXT(0), B(31) => HDU_NPC_IN(31), B(30) => 
                           HDU_NPC_IN(30), B(29) => HDU_NPC_IN(29), B(28) => 
                           HDU_NPC_IN(28), B(27) => HDU_NPC_IN(27), B(26) => 
                           HDU_NPC_IN(26), B(25) => HDU_NPC_IN(25), B(24) => 
                           HDU_NPC_IN(24), B(23) => HDU_NPC_IN(23), B(22) => 
                           HDU_NPC_IN(22), B(21) => HDU_NPC_IN(21), B(20) => 
                           HDU_NPC_IN(20), B(19) => HDU_NPC_IN(19), B(18) => 
                           HDU_NPC_IN(18), B(17) => HDU_NPC_IN(17), B(16) => 
                           HDU_NPC_IN(16), B(15) => HDU_NPC_IN(15), B(14) => 
                           HDU_NPC_IN(14), B(13) => HDU_NPC_IN(13), B(12) => 
                           HDU_NPC_IN(12), B(11) => HDU_NPC_IN(11), B(10) => 
                           HDU_NPC_IN(10), B(9) => HDU_NPC_IN(9), B(8) => 
                           HDU_NPC_IN(8), B(7) => HDU_NPC_IN(7), B(6) => 
                           HDU_NPC_IN(6), B(5) => HDU_NPC_IN(5), B(4) => 
                           HDU_NPC_IN(4), B(3) => HDU_NPC_IN(3), B(2) => 
                           HDU_NPC_IN(2), B(1) => HDU_NPC_IN(1), B(0) => 
                           HDU_NPC_IN(0), S => Bubble_in, Z(31) => 
                           sig_NPC_31_port, Z(30) => sig_NPC_30_port, Z(29) => 
                           sig_NPC_29_port, Z(28) => sig_NPC_28_port, Z(27) => 
                           sig_NPC_27_port, Z(26) => sig_NPC_26_port, Z(25) => 
                           sig_NPC_25_port, Z(24) => sig_NPC_24_port, Z(23) => 
                           sig_NPC_23_port, Z(22) => sig_NPC_22_port, Z(21) => 
                           sig_NPC_21_port, Z(20) => sig_NPC_20_port, Z(19) => 
                           sig_NPC_19_port, Z(18) => sig_NPC_18_port, Z(17) => 
                           sig_NPC_17_port, Z(16) => sig_NPC_16_port, Z(15) => 
                           sig_NPC_15_port, Z(14) => sig_NPC_14_port, Z(13) => 
                           sig_NPC_13_port, Z(12) => sig_NPC_12_port, Z(11) => 
                           sig_NPC_11_port, Z(10) => sig_NPC_10_port, Z(9) => 
                           sig_NPC_9_port, Z(8) => sig_NPC_8_port, Z(7) => 
                           sig_NPC_7_port, Z(6) => sig_NPC_6_port, Z(5) => 
                           sig_NPC_5_port, Z(4) => sig_NPC_4_port, Z(3) => 
                           sig_NPC_3_port, Z(2) => sig_NPC_2_port, Z(1) => 
                           sig_NPC_1_port, Z(0) => sig_NPC_0_port);
   PC_or_PC_HDU : mux21_NBIT32_5 port map( A(31) => ADDR_OUT_31_port, A(30) => 
                           ADDR_OUT_30_port, A(29) => ADDR_OUT_29_port, A(28) 
                           => ADDR_OUT_28_port, A(27) => ADDR_OUT_27_port, 
                           A(26) => ADDR_OUT_26_port, A(25) => ADDR_OUT_25_port
                           , A(24) => ADDR_OUT_24_port, A(23) => 
                           ADDR_OUT_23_port, A(22) => ADDR_OUT_22_port, A(21) 
                           => ADDR_OUT_21_port, A(20) => ADDR_OUT_20_port, 
                           A(19) => ADDR_OUT_19_port, A(18) => ADDR_OUT_18_port
                           , A(17) => ADDR_OUT_17_port, A(16) => 
                           ADDR_OUT_16_port, A(15) => ADDR_OUT_15_port, A(14) 
                           => ADDR_OUT_14_port, A(13) => ADDR_OUT_13_port, 
                           A(12) => ADDR_OUT_12_port, A(11) => ADDR_OUT_11_port
                           , A(10) => ADDR_OUT_10_port, A(9) => ADDR_OUT_9_port
                           , A(8) => ADDR_OUT_8_port, A(7) => ADDR_OUT_7_port, 
                           A(6) => ADDR_OUT_6_port, A(5) => ADDR_OUT_5_port, 
                           A(4) => ADDR_OUT_4_port, A(3) => ADDR_OUT_3_port, 
                           A(2) => ADDR_OUT_2_port, A(1) => ADDR_OUT_1_port, 
                           A(0) => ADDR_OUT_0_port, B(31) => HDU_PC_IN(31), 
                           B(30) => HDU_PC_IN(30), B(29) => HDU_PC_IN(29), 
                           B(28) => HDU_PC_IN(28), B(27) => HDU_PC_IN(27), 
                           B(26) => HDU_PC_IN(26), B(25) => HDU_PC_IN(25), 
                           B(24) => HDU_PC_IN(24), B(23) => HDU_PC_IN(23), 
                           B(22) => HDU_PC_IN(22), B(21) => HDU_PC_IN(21), 
                           B(20) => HDU_PC_IN(20), B(19) => HDU_PC_IN(19), 
                           B(18) => HDU_PC_IN(18), B(17) => HDU_PC_IN(17), 
                           B(16) => HDU_PC_IN(16), B(15) => HDU_PC_IN(15), 
                           B(14) => HDU_PC_IN(14), B(13) => HDU_PC_IN(13), 
                           B(12) => HDU_PC_IN(12), B(11) => HDU_PC_IN(11), 
                           B(10) => HDU_PC_IN(10), B(9) => HDU_PC_IN(9), B(8) 
                           => HDU_PC_IN(8), B(7) => HDU_PC_IN(7), B(6) => 
                           HDU_PC_IN(6), B(5) => HDU_PC_IN(5), B(4) => 
                           HDU_PC_IN(4), B(3) => HDU_PC_IN(3), B(2) => 
                           HDU_PC_IN(2), B(1) => HDU_PC_IN(1), B(0) => 
                           HDU_PC_IN(0), S => Bubble_in, Z(31) => 
                           PC_MUX_OUT_31_port, Z(30) => PC_MUX_OUT_30_port, 
                           Z(29) => PC_MUX_OUT_29_port, Z(28) => 
                           PC_MUX_OUT_28_port, Z(27) => PC_MUX_OUT_27_port, 
                           Z(26) => PC_MUX_OUT_26_port, Z(25) => 
                           PC_MUX_OUT_25_port, Z(24) => PC_MUX_OUT_24_port, 
                           Z(23) => PC_MUX_OUT_23_port, Z(22) => 
                           PC_MUX_OUT_22_port, Z(21) => PC_MUX_OUT_21_port, 
                           Z(20) => PC_MUX_OUT_20_port, Z(19) => 
                           PC_MUX_OUT_19_port, Z(18) => PC_MUX_OUT_18_port, 
                           Z(17) => PC_MUX_OUT_17_port, Z(16) => 
                           PC_MUX_OUT_16_port, Z(15) => PC_MUX_OUT_15_port, 
                           Z(14) => PC_MUX_OUT_14_port, Z(13) => 
                           PC_MUX_OUT_13_port, Z(12) => PC_MUX_OUT_12_port, 
                           Z(11) => PC_MUX_OUT_11_port, Z(10) => 
                           PC_MUX_OUT_10_port, Z(9) => PC_MUX_OUT_9_port, Z(8) 
                           => PC_MUX_OUT_8_port, Z(7) => PC_MUX_OUT_7_port, 
                           Z(6) => PC_MUX_OUT_6_port, Z(5) => PC_MUX_OUT_5_port
                           , Z(4) => PC_MUX_OUT_4_port, Z(3) => 
                           PC_MUX_OUT_3_port, Z(2) => PC_MUX_OUT_2_port, Z(1) 
                           => PC_MUX_OUT_1_port, Z(0) => PC_MUX_OUT_0_port);
   INS_or_HDU_INS : mux21_NBIT32_4 port map( A(31) => INS_IN(31), A(30) => 
                           INS_IN(30), A(29) => INS_IN(29), A(28) => INS_IN(28)
                           , A(27) => INS_IN(27), A(26) => INS_IN(26), A(25) =>
                           INS_IN(25), A(24) => INS_IN(24), A(23) => INS_IN(23)
                           , A(22) => INS_IN(22), A(21) => INS_IN(21), A(20) =>
                           INS_IN(20), A(19) => INS_IN(19), A(18) => INS_IN(18)
                           , A(17) => INS_IN(17), A(16) => INS_IN(16), A(15) =>
                           INS_IN(15), A(14) => INS_IN(14), A(13) => INS_IN(13)
                           , A(12) => INS_IN(12), A(11) => INS_IN(11), A(10) =>
                           INS_IN(10), A(9) => INS_IN(9), A(8) => INS_IN(8), 
                           A(7) => INS_IN(7), A(6) => INS_IN(6), A(5) => 
                           INS_IN(5), A(4) => INS_IN(4), A(3) => INS_IN(3), 
                           A(2) => INS_IN(2), A(1) => INS_IN(1), A(0) => 
                           INS_IN(0), B(31) => HDU_INS_IN(31), B(30) => 
                           HDU_INS_IN(30), B(29) => HDU_INS_IN(29), B(28) => 
                           HDU_INS_IN(28), B(27) => HDU_INS_IN(27), B(26) => 
                           HDU_INS_IN(26), B(25) => HDU_INS_IN(25), B(24) => 
                           HDU_INS_IN(24), B(23) => HDU_INS_IN(23), B(22) => 
                           HDU_INS_IN(22), B(21) => HDU_INS_IN(21), B(20) => 
                           HDU_INS_IN(20), B(19) => HDU_INS_IN(19), B(18) => 
                           HDU_INS_IN(18), B(17) => HDU_INS_IN(17), B(16) => 
                           HDU_INS_IN(16), B(15) => HDU_INS_IN(15), B(14) => 
                           HDU_INS_IN(14), B(13) => HDU_INS_IN(13), B(12) => 
                           HDU_INS_IN(12), B(11) => HDU_INS_IN(11), B(10) => 
                           HDU_INS_IN(10), B(9) => HDU_INS_IN(9), B(8) => 
                           HDU_INS_IN(8), B(7) => HDU_INS_IN(7), B(6) => 
                           HDU_INS_IN(6), B(5) => HDU_INS_IN(5), B(4) => 
                           HDU_INS_IN(4), B(3) => HDU_INS_IN(3), B(2) => 
                           HDU_INS_IN(2), B(1) => HDU_INS_IN(1), B(0) => 
                           HDU_INS_IN(0), S => Bubble_in, Z(31) => 
                           sig_INS_31_port, Z(30) => sig_INS_30_port, Z(29) => 
                           sig_INS_29_port, Z(28) => sig_INS_28_port, Z(27) => 
                           sig_INS_27_port, Z(26) => sig_INS_26_port, Z(25) => 
                           sig_INS_25_port, Z(24) => sig_INS_24_port, Z(23) => 
                           sig_INS_23_port, Z(22) => sig_INS_22_port, Z(21) => 
                           sig_INS_21_port, Z(20) => sig_INS_20_port, Z(19) => 
                           sig_INS_19_port, Z(18) => sig_INS_18_port, Z(17) => 
                           sig_INS_17_port, Z(16) => sig_INS_16_port, Z(15) => 
                           sig_INS_15_port, Z(14) => sig_INS_14_port, Z(13) => 
                           sig_INS_13_port, Z(12) => sig_INS_12_port, Z(11) => 
                           sig_INS_11_port, Z(10) => sig_INS_10_port, Z(9) => 
                           sig_INS_9_port, Z(8) => sig_INS_8_port, Z(7) => 
                           sig_INS_7_port, Z(6) => sig_INS_6_port, Z(5) => 
                           sig_INS_5_port, Z(4) => sig_INS_4_port, Z(3) => 
                           sig_INS_3_port, Z(2) => sig_INS_2_port, Z(1) => 
                           sig_INS_1_port, Z(0) => sig_INS_0_port);
   PC : regn_N32_0 port map( DIN(31) => sig_NPC_31_port, DIN(30) => 
                           sig_NPC_30_port, DIN(29) => sig_NPC_29_port, DIN(28)
                           => sig_NPC_28_port, DIN(27) => sig_NPC_27_port, 
                           DIN(26) => sig_NPC_26_port, DIN(25) => 
                           sig_NPC_25_port, DIN(24) => sig_NPC_24_port, DIN(23)
                           => sig_NPC_23_port, DIN(22) => sig_NPC_22_port, 
                           DIN(21) => sig_NPC_21_port, DIN(20) => 
                           sig_NPC_20_port, DIN(19) => sig_NPC_19_port, DIN(18)
                           => sig_NPC_18_port, DIN(17) => sig_NPC_17_port, 
                           DIN(16) => sig_NPC_16_port, DIN(15) => 
                           sig_NPC_15_port, DIN(14) => sig_NPC_14_port, DIN(13)
                           => sig_NPC_13_port, DIN(12) => sig_NPC_12_port, 
                           DIN(11) => sig_NPC_11_port, DIN(10) => 
                           sig_NPC_10_port, DIN(9) => sig_NPC_9_port, DIN(8) =>
                           sig_NPC_8_port, DIN(7) => sig_NPC_7_port, DIN(6) => 
                           sig_NPC_6_port, DIN(5) => sig_NPC_5_port, DIN(4) => 
                           sig_NPC_4_port, DIN(3) => sig_NPC_3_port, DIN(2) => 
                           sig_NPC_2_port, DIN(1) => sig_NPC_1_port, DIN(0) => 
                           sig_NPC_0_port, CLK => CLK, EN => X_Logic1_port, RST
                           => RST, DOUT(31) => ADDR_OUT_31_port, DOUT(30) => 
                           ADDR_OUT_30_port, DOUT(29) => n19, DOUT(28) => 
                           ADDR_OUT_28_port, DOUT(27) => ADDR_OUT_27_port, 
                           DOUT(26) => ADDR_OUT_26_port, DOUT(25) => 
                           ADDR_OUT_25_port, DOUT(24) => ADDR_OUT_24_port, 
                           DOUT(23) => n20, DOUT(22) => ADDR_OUT_22_port, 
                           DOUT(21) => ADDR_OUT_21_port, DOUT(20) => 
                           ADDR_OUT_20_port, DOUT(19) => ADDR_OUT_19_port, 
                           DOUT(18) => ADDR_OUT_18_port, DOUT(17) => n21, 
                           DOUT(16) => n22, DOUT(15) => ADDR_OUT_15_port, 
                           DOUT(14) => n23, DOUT(13) => ADDR_OUT_13_port, 
                           DOUT(12) => n24, DOUT(11) => ADDR_OUT_11_port, 
                           DOUT(10) => ADDR_OUT_10_port, DOUT(9) => n25, 
                           DOUT(8) => n26, DOUT(7) => n27, DOUT(6) => n28, 
                           DOUT(5) => n29, DOUT(4) => n30, DOUT(3) => n31, 
                           DOUT(2) => n32, DOUT(1) => ADDR_OUT_1_port, DOUT(0) 
                           => ADDR_OUT_0_port);
   PC_reg : regn_N32_10 port map( DIN(31) => PC_MUX_OUT_31_port, DIN(30) => 
                           PC_MUX_OUT_30_port, DIN(29) => PC_MUX_OUT_29_port, 
                           DIN(28) => PC_MUX_OUT_28_port, DIN(27) => 
                           PC_MUX_OUT_27_port, DIN(26) => PC_MUX_OUT_26_port, 
                           DIN(25) => PC_MUX_OUT_25_port, DIN(24) => 
                           PC_MUX_OUT_24_port, DIN(23) => PC_MUX_OUT_23_port, 
                           DIN(22) => PC_MUX_OUT_22_port, DIN(21) => 
                           PC_MUX_OUT_21_port, DIN(20) => PC_MUX_OUT_20_port, 
                           DIN(19) => PC_MUX_OUT_19_port, DIN(18) => 
                           PC_MUX_OUT_18_port, DIN(17) => PC_MUX_OUT_17_port, 
                           DIN(16) => PC_MUX_OUT_16_port, DIN(15) => 
                           PC_MUX_OUT_15_port, DIN(14) => PC_MUX_OUT_14_port, 
                           DIN(13) => PC_MUX_OUT_13_port, DIN(12) => 
                           PC_MUX_OUT_12_port, DIN(11) => PC_MUX_OUT_11_port, 
                           DIN(10) => PC_MUX_OUT_10_port, DIN(9) => 
                           PC_MUX_OUT_9_port, DIN(8) => PC_MUX_OUT_8_port, 
                           DIN(7) => PC_MUX_OUT_7_port, DIN(6) => 
                           PC_MUX_OUT_6_port, DIN(5) => PC_MUX_OUT_5_port, 
                           DIN(4) => PC_MUX_OUT_4_port, DIN(3) => 
                           PC_MUX_OUT_3_port, DIN(2) => PC_MUX_OUT_2_port, 
                           DIN(1) => PC_MUX_OUT_1_port, DIN(0) => 
                           PC_MUX_OUT_0_port, CLK => CLK, EN => X_Logic1_port, 
                           RST => sig_RST, DOUT(31) => PC_OUT(31), DOUT(30) => 
                           PC_OUT(30), DOUT(29) => PC_OUT(29), DOUT(28) => 
                           PC_OUT(28), DOUT(27) => PC_OUT(27), DOUT(26) => 
                           PC_OUT(26), DOUT(25) => PC_OUT(25), DOUT(24) => 
                           PC_OUT(24), DOUT(23) => PC_OUT(23), DOUT(22) => 
                           PC_OUT(22), DOUT(21) => PC_OUT(21), DOUT(20) => 
                           PC_OUT(20), DOUT(19) => PC_OUT(19), DOUT(18) => 
                           PC_OUT(18), DOUT(17) => PC_OUT(17), DOUT(16) => 
                           PC_OUT(16), DOUT(15) => PC_OUT(15), DOUT(14) => 
                           PC_OUT(14), DOUT(13) => PC_OUT(13), DOUT(12) => 
                           PC_OUT(12), DOUT(11) => PC_OUT(11), DOUT(10) => 
                           PC_OUT(10), DOUT(9) => PC_OUT(9), DOUT(8) => 
                           PC_OUT(8), DOUT(7) => PC_OUT(7), DOUT(6) => 
                           PC_OUT(6), DOUT(5) => PC_OUT(5), DOUT(4) => 
                           PC_OUT(4), DOUT(3) => PC_OUT(3), DOUT(2) => 
                           PC_OUT(2), DOUT(1) => PC_OUT(1), DOUT(0) => 
                           PC_OUT(0));
   IR : regn_N32_9 port map( DIN(31) => sig_INS_31_port, DIN(30) => 
                           sig_INS_30_port, DIN(29) => sig_INS_29_port, DIN(28)
                           => sig_INS_28_port, DIN(27) => sig_INS_27_port, 
                           DIN(26) => sig_INS_26_port, DIN(25) => 
                           sig_INS_25_port, DIN(24) => sig_INS_24_port, DIN(23)
                           => sig_INS_23_port, DIN(22) => sig_INS_22_port, 
                           DIN(21) => sig_INS_21_port, DIN(20) => 
                           sig_INS_20_port, DIN(19) => sig_INS_19_port, DIN(18)
                           => sig_INS_18_port, DIN(17) => sig_INS_17_port, 
                           DIN(16) => sig_INS_16_port, DIN(15) => 
                           sig_INS_15_port, DIN(14) => sig_INS_14_port, DIN(13)
                           => sig_INS_13_port, DIN(12) => sig_INS_12_port, 
                           DIN(11) => sig_INS_11_port, DIN(10) => 
                           sig_INS_10_port, DIN(9) => sig_INS_9_port, DIN(8) =>
                           sig_INS_8_port, DIN(7) => sig_INS_7_port, DIN(6) => 
                           sig_INS_6_port, DIN(5) => sig_INS_5_port, DIN(4) => 
                           sig_INS_4_port, DIN(3) => sig_INS_3_port, DIN(2) => 
                           sig_INS_2_port, DIN(1) => sig_INS_1_port, DIN(0) => 
                           sig_INS_0_port, CLK => CLK, EN => X_Logic1_port, RST
                           => sig_RST, DOUT(31) => INS_OUT(31), DOUT(30) => 
                           INS_OUT(30), DOUT(29) => INS_OUT(29), DOUT(28) => 
                           INS_OUT(28), DOUT(27) => INS_OUT(27), DOUT(26) => 
                           INS_OUT(26), DOUT(25) => INS_OUT(25), DOUT(24) => 
                           INS_OUT(24), DOUT(23) => INS_OUT(23), DOUT(22) => 
                           INS_OUT(22), DOUT(21) => INS_OUT(21), DOUT(20) => 
                           INS_OUT(20), DOUT(19) => INS_OUT(19), DOUT(18) => 
                           INS_OUT(18), DOUT(17) => INS_OUT(17), DOUT(16) => 
                           INS_OUT(16), DOUT(15) => INS_OUT(15), DOUT(14) => 
                           INS_OUT(14), DOUT(13) => INS_OUT(13), DOUT(12) => 
                           INS_OUT(12), DOUT(11) => INS_OUT(11), DOUT(10) => 
                           INS_OUT(10), DOUT(9) => INS_OUT(9), DOUT(8) => 
                           INS_OUT(8), DOUT(7) => INS_OUT(7), DOUT(6) => 
                           INS_OUT(6), DOUT(5) => INS_OUT(5), DOUT(4) => 
                           INS_OUT(4), DOUT(3) => INS_OUT(3), DOUT(2) => 
                           INS_OUT(2), DOUT(1) => INS_OUT(1), DOUT(0) => 
                           INS_OUT(0));
   add_54 : Fetch_DW01_add_1 port map( A(31) => ADDR_OUT_31_port, A(30) => 
                           ADDR_OUT_30_port, A(29) => n19, A(28) => 
                           ADDR_OUT_28_port, A(27) => ADDR_OUT_27_port, A(26) 
                           => ADDR_OUT_26_port, A(25) => ADDR_OUT_25_port, 
                           A(24) => ADDR_OUT_24_port, A(23) => n20, A(22) => 
                           ADDR_OUT_22_port, A(21) => ADDR_OUT_21_port, A(20) 
                           => ADDR_OUT_20_port, A(19) => ADDR_OUT_19_port, 
                           A(18) => ADDR_OUT_18_port, A(17) => n21, A(16) => 
                           n22, A(15) => ADDR_OUT_15_port, A(14) => n23, A(13) 
                           => ADDR_OUT_13_port, A(12) => n24, A(11) => 
                           ADDR_OUT_11_port, A(10) => ADDR_OUT_10_port, A(9) =>
                           n25, A(8) => n26, A(7) => n27, A(6) => n28, A(5) => 
                           n29, A(4) => n30, A(3) => n31, A(2) => n32, A(1) => 
                           ADDR_OUT_1_port, A(0) => ADDR_OUT_0_port, B(31) => 
                           n1, B(30) => n1, B(29) => n1, B(28) => n1, B(27) => 
                           n1, B(26) => n1, B(25) => n1, B(24) => n1, B(23) => 
                           n1, B(22) => n1, B(21) => n1, B(20) => n1, B(19) => 
                           n1, B(18) => n1, B(17) => n1, B(16) => n1, B(15) => 
                           n1, B(14) => n1, B(13) => n1, B(12) => n1, B(11) => 
                           n1, B(10) => n1, B(9) => n1, B(8) => n1, B(7) => n1,
                           B(6) => n1, B(5) => n1, B(4) => n1, B(3) => n1, B(2)
                           => n2, B(1) => n1, B(0) => n1, CI => n3, SUM(31) => 
                           NPC_OUT(31), SUM(30) => NPC_OUT(30), SUM(29) => 
                           NPC_OUT(29), SUM(28) => NPC_OUT(28), SUM(27) => 
                           NPC_OUT(27), SUM(26) => NPC_OUT(26), SUM(25) => 
                           NPC_OUT(25), SUM(24) => NPC_OUT(24), SUM(23) => 
                           NPC_OUT(23), SUM(22) => NPC_OUT(22), SUM(21) => 
                           NPC_OUT(21), SUM(20) => NPC_OUT(20), SUM(19) => 
                           NPC_OUT(19), SUM(18) => NPC_OUT(18), SUM(17) => 
                           NPC_OUT(17), SUM(16) => NPC_OUT(16), SUM(15) => 
                           NPC_OUT(15), SUM(14) => NPC_OUT(14), SUM(13) => 
                           NPC_OUT(13), SUM(12) => NPC_OUT(12), SUM(11) => 
                           NPC_OUT(11), SUM(10) => NPC_OUT(10), SUM(9) => 
                           NPC_OUT(9), SUM(8) => NPC_OUT(8), SUM(7) => 
                           NPC_OUT(7), SUM(6) => NPC_OUT(6), SUM(5) => 
                           NPC_OUT(5), SUM(4) => NPC_OUT(4), SUM(3) => 
                           NPC_OUT(3), SUM(2) => NPC_OUT(2), SUM(1) => 
                           NPC_OUT(1), SUM(0) => NPC_OUT(0), CO => n_1945);
   U6 : CLKBUF_X1 port map( A => n26, Z => ADDR_OUT_8_port);
   U7 : CLKBUF_X1 port map( A => n19, Z => ADDR_OUT_29_port);
   U8 : CLKBUF_X1 port map( A => n27, Z => ADDR_OUT_7_port);
   U9 : CLKBUF_X1 port map( A => n32, Z => ADDR_OUT_2_port);
   U10 : CLKBUF_X1 port map( A => n20, Z => ADDR_OUT_23_port);
   U11 : CLKBUF_X1 port map( A => n24, Z => ADDR_OUT_12_port);
   U12 : CLKBUF_X1 port map( A => n28, Z => ADDR_OUT_6_port);
   U13 : CLKBUF_X1 port map( A => n31, Z => ADDR_OUT_3_port);
   U14 : CLKBUF_X1 port map( A => n21, Z => ADDR_OUT_17_port);
   U15 : CLKBUF_X1 port map( A => n22, Z => ADDR_OUT_16_port);
   U16 : NOR2_X1 port map( A1 => ZERO_FLAG, A2 => n18, ZN => sig_RST);
   U17 : CLKBUF_X1 port map( A => n29, Z => ADDR_OUT_5_port);
   U18 : CLKBUF_X1 port map( A => n23, Z => ADDR_OUT_14_port);
   U19 : CLKBUF_X1 port map( A => n30, Z => ADDR_OUT_4_port);
   U20 : CLKBUF_X1 port map( A => n25, Z => ADDR_OUT_9_port);
   U21 : INV_X1 port map( A => RST, ZN => n18);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity hardwired_cu_NBIT32 is

   port( REG_LATCH_EN, RD1, RD2, MUX_A_SEL : out std_logic;  MUX_B_SEL : out 
         std_logic_vector (1 downto 0);  ALU_OPC : out std_logic_vector (0 to 
         3);  ALU_OUTREG_EN, DRAM_R_IN : out std_logic;  JUMP_TYPE : out 
         std_logic_vector (1 downto 0);  MEM_EN_IN, DRAM_W_IN, RF_WE, 
         DRAM_EN_IN, WB_MUX_SEL : out std_logic;  INS_IN : in std_logic_vector 
         (31 downto 0);  Bubble, Clk, Rst : in std_logic);

end hardwired_cu_NBIT32;

architecture SYN_bhv of hardwired_cu_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal AluOP_E_3_port, AluOP_E_2_port, AluOP_E_1_port, AluOP_E_0_port, N24, 
      N25, N26, N27, n19, n20, n21, n22, n23, n24_port, n25_port, n26_port, 
      n27_port, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40
      , n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, 
      n55, n56, n58, n59, n60, n61, n62, n63, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n_1946, n_1947, n_1948, 
      n_1949, n_1950, n_1951, n_1952, n_1953 : std_logic;

begin
   
   AluOP_E_reg_3_inst : DFFR_X1 port map( D => N27, CK => Clk, RN => Rst, Q => 
                           AluOP_E_3_port, QN => n_1946);
   AluOP_E_reg_2_inst : DFFR_X1 port map( D => N26, CK => Clk, RN => Rst, Q => 
                           AluOP_E_2_port, QN => n_1947);
   AluOP_E_reg_1_inst : DFFR_X1 port map( D => N25, CK => Clk, RN => Rst, Q => 
                           AluOP_E_1_port, QN => n_1948);
   AluOP_E_reg_0_inst : DFFR_X1 port map( D => N24, CK => Clk, RN => Rst, Q => 
                           AluOP_E_0_port, QN => n_1949);
   WB_MUX_SEL <= '0';
   DRAM_EN_IN <= '0';
   RF_WE <= '0';
   DRAM_W_IN <= '0';
   MEM_EN_IN <= '0';
   JUMP_TYPE(0) <= '0';
   JUMP_TYPE(1) <= '0';
   DRAM_R_IN <= '0';
   ALU_OUTREG_EN <= '0';
   MUX_B_SEL(0) <= '0';
   MUX_B_SEL(1) <= '0';
   MUX_A_SEL <= '0';
   RD2 <= '0';
   RD1 <= '0';
   REG_LATCH_EN <= '0';
   U74 : XOR2_X1 port map( A => n2, B => INS_IN(1), Z => n33);
   U75 : NAND3_X1 port map( A1 => n16, A2 => n13, A3 => INS_IN(30), ZN => n37);
   U76 : OAI33_X1 port map( A1 => n26_port, A2 => n13, A3 => n17, B1 => n46, B2
                           => INS_IN(30), B3 => INS_IN(28), ZN => n43);
   U77 : OAI33_X1 port map( A1 => n24_port, A2 => n25_port, A3 => n17, B1 => n3
                           , B2 => n8, B3 => n34, ZN => n50);
   U78 : OAI33_X1 port map( A1 => n12, A2 => n56, A3 => n11, B1 => n27_port, B2
                           => INS_IN(30), B3 => n25_port, ZN => n55);
   U79 : NAND3_X1 port map( A1 => n51, A2 => n7, A3 => INS_IN(5), ZN => n35);
   U80 : OAI33_X1 port map( A1 => n58, A2 => n13, A3 => n17, B1 => n59, B2 => 
                           n39, B3 => n6, ZN => n48);
   U81 : NAND3_X1 port map( A1 => INS_IN(3), A2 => n51, A3 => INS_IN(5), ZN => 
                           n39);
   U82 : NAND3_X1 port map( A1 => n15, A2 => n18, A3 => INS_IN(28), ZN => 
                           n24_port);
   U83 : NAND3_X1 port map( A1 => n10, A2 => n13, A3 => n63, ZN => n34);
   U84 : NAND3_X1 port map( A1 => n16, A2 => n17, A3 => INS_IN(28), ZN => n36);
   ALU_OPC_reg_3_inst : DFFR_X1 port map( D => AluOP_E_3_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(0), QN => n_1950);
   ALU_OPC_reg_2_inst : DFFR_X1 port map( D => AluOP_E_2_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(1), QN => n_1951);
   ALU_OPC_reg_1_inst : DFFR_X1 port map( D => AluOP_E_1_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(2), QN => n_1952);
   ALU_OPC_reg_0_inst : DFFR_X1 port map( D => AluOP_E_0_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(3), QN => n_1953);
   U18 : INV_X1 port map( A => n25_port, ZN => n10);
   U19 : NAND2_X1 port map( A1 => n12, A2 => n11, ZN => n25_port);
   U20 : AOI21_X1 port map( B1 => n40, B2 => n41, A => Bubble, ZN => N25);
   U21 : AOI211_X1 port map( C1 => n14, C2 => n10, A => n38, B => n48, ZN => 
                           n40);
   U22 : AOI221_X1 port map( B1 => n42, B2 => n5, C1 => n16, C2 => n43, A => 
                           n44, ZN => n41);
   U23 : INV_X1 port map( A => n47, ZN => n5);
   U24 : AOI21_X1 port map( B1 => n28, B2 => n29, A => Bubble, ZN => N26);
   U25 : AOI21_X1 port map( B1 => n20, B2 => n6, A => n38, ZN => n28);
   U26 : NOR3_X1 port map( A1 => n30, A2 => n31, A3 => n32, ZN => n29);
   U27 : AOI21_X1 port map( B1 => n36, B2 => n37, A => n26_port, ZN => n30);
   U28 : INV_X1 port map( A => n36, ZN => n14);
   U29 : INV_X1 port map( A => n27_port, ZN => n16);
   U30 : OR2_X1 port map( A1 => n49, A2 => n50, ZN => n38);
   U31 : INV_X1 port map( A => n52, ZN => n3);
   U32 : INV_X1 port map( A => n51, ZN => n8);
   U33 : NAND2_X1 port map( A1 => n16, A2 => n10, ZN => n58);
   U34 : OR3_X1 port map( A1 => INS_IN(0), A2 => INS_IN(1), A3 => n34, ZN => 
                           n59);
   U35 : NOR4_X1 port map( A1 => INS_IN(6), A2 => INS_IN(4), A3 => INS_IN(10), 
                           A4 => n62, ZN => n51);
   U36 : OR3_X1 port map( A1 => INS_IN(9), A2 => INS_IN(8), A3 => INS_IN(7), ZN
                           => n62);
   U37 : NAND2_X1 port map( A1 => INS_IN(27), A2 => n11, ZN => n46);
   U38 : NOR3_X1 port map( A1 => INS_IN(29), A2 => INS_IN(31), A3 => INS_IN(30)
                           , ZN => n63);
   U39 : NOR4_X1 port map( A1 => n2, A2 => n39, A3 => n34, A4 => INS_IN(1), ZN 
                           => n20);
   U40 : NOR4_X1 port map( A1 => n6, A2 => INS_IN(0), A3 => INS_IN(3), A4 => 
                           INS_IN(5), ZN => n52);
   U41 : NOR4_X1 port map( A1 => n33, A2 => n34, A3 => n6, A4 => n35, ZN => n32
                           );
   U42 : NOR4_X1 port map( A1 => INS_IN(1), A2 => n4, A3 => n34, A4 => n6, ZN 
                           => n44);
   U43 : INV_X1 port map( A => n45, ZN => n4);
   U44 : OAI21_X1 port map( B1 => n35, B2 => INS_IN(0), A => n39, ZN => n45);
   U45 : NOR3_X1 port map( A1 => n34, A2 => INS_IN(0), A3 => n35, ZN => n42);
   U46 : INV_X1 port map( A => INS_IN(3), ZN => n7);
   U47 : NOR3_X1 port map( A1 => n36, A2 => INS_IN(26), A3 => n12, ZN => n31);
   U48 : INV_X1 port map( A => INS_IN(2), ZN => n6);
   U49 : INV_X1 port map( A => INS_IN(30), ZN => n17);
   U50 : AOI22_X1 port map( A1 => n15, A2 => n18, B1 => INS_IN(31), B2 => n17, 
                           ZN => n56);
   U51 : NAND2_X1 port map( A1 => INS_IN(26), A2 => n12, ZN => n26_port);
   U52 : INV_X1 port map( A => INS_IN(27), ZN => n12);
   U53 : AOI21_X1 port map( B1 => n53, B2 => n54, A => Bubble, ZN => N24);
   U54 : AOI211_X1 port map( C1 => n14, C2 => n10, A => n49, B => n23, ZN => 
                           n53);
   U55 : AOI221_X1 port map( B1 => n42, B2 => n47, C1 => n55, C2 => n13, A => 
                           n31, ZN => n54);
   U56 : INV_X1 port map( A => INS_IN(28), ZN => n13);
   U57 : NAND2_X1 port map( A1 => INS_IN(29), A2 => n18, ZN => n27_port);
   U58 : OR2_X1 port map( A1 => n48, A2 => n1, ZN => n23);
   U59 : NOR3_X1 port map( A1 => n26_port, A2 => INS_IN(30), A3 => n24_port, ZN
                           => n1);
   U60 : NAND2_X1 port map( A1 => INS_IN(1), A2 => n6, ZN => n47);
   U61 : INV_X1 port map( A => INS_IN(31), ZN => n18);
   U62 : INV_X1 port map( A => INS_IN(26), ZN => n11);
   U63 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => n49);
   U64 : OR4_X1 port map( A1 => n12, A2 => n24_port, A3 => n17, A4 => 
                           INS_IN(26), ZN => n61);
   U65 : NAND4_X1 port map( A1 => INS_IN(1), A2 => n52, A3 => n9, A4 => n51, ZN
                           => n60);
   U66 : INV_X1 port map( A => n34, ZN => n9);
   U67 : NOR2_X1 port map( A1 => Bubble, A2 => n19, ZN => N27);
   U68 : NOR4_X1 port map( A1 => n20, A2 => n21, A3 => n22, A4 => n23, ZN => 
                           n19);
   U69 : NOR3_X1 port map( A1 => n26_port, A2 => n27_port, A3 => n17, ZN => n21
                           );
   U70 : NOR3_X1 port map( A1 => n24_port, A2 => INS_IN(30), A3 => n25_port, ZN
                           => n22);
   U71 : INV_X1 port map( A => INS_IN(0), ZN => n2);
   U72 : INV_X1 port map( A => INS_IN(29), ZN => n15);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Datapath is

   port( CLK, RST : in std_logic;  INS_IN, DATA_IN : in std_logic_vector (31 
         downto 0);  REG_LATCH_EN, RD1, RD2, MUX_A_SEL : in std_logic;  
         MUX_B_SEL : in std_logic_vector (1 downto 0);  ALU_OPC : in 
         std_logic_vector (0 to 3);  ALU_OUTREG_EN : in std_logic;  JUMP_TYPE :
         in std_logic_vector (1 downto 0);  DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, 
         RF_WE, DRAM_EN_IN, WB_MUX_SEL : in std_logic;  INS_OUT, IRAM_ADDR_OUT,
         DRAM_ADDR_OUT, DATA_OUT : out std_logic_vector (31 downto 0);  
         DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble_out : out std_logic);

end Datapath;

architecture SYN_struct of Datapath is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HazardDetection
      port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : in std_logic_vector
            (4 downto 0);  DRAM_R : in std_logic;  INS_IN, PC_IN : in 
            std_logic_vector (31 downto 0);  Bubble : out std_logic;  
            HDU_INS_OUT, HDU_PC_OUT, HDU_NPC_OUT : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Writeback
      port( WB_MUX_SEL : in std_logic;  DATA_IN, ALU_RES_IN : in 
            std_logic_vector (31 downto 0);  ADD_WR_IN : in std_logic_vector (4
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0);  
            ADD_WR_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component ff_2
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Memory
      port( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, DRAM_EN_IN : in 
            std_logic;  PC_SEL : in std_logic_vector (1 downto 0);  NPC_IN, 
            NPC_ABS, NPC_REL, ALU_RES_IN, B_IN : in std_logic_vector (31 downto
            0);  ADD_WR_IN : in std_logic_vector (4 downto 0);  DRAM_DATA_IN : 
            in std_logic_vector (31 downto 0);  PC_OUT : out std_logic_vector 
            (31 downto 0);  DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT : out std_logic
            ;  DRAM_ADDR_OUT, DRAM_DATA_OUT, DATA_OUT, ALU_RES_OUT, OP_MEM : 
            out std_logic_vector (31 downto 0);  ADD_WR_MEM, ADD_WR_OUT : out 
            std_logic_vector (4 downto 0));
   end component;
   
   component ff_0
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Execute
      port( CLK, RST, MUX_A_SEL : in std_logic;  MUX_B_SEL : in 
            std_logic_vector (1 downto 0);  ALU_OPC : in std_logic_vector (0 to
            3);  ALU_OUTREG_EN : in std_logic;  JUMP_TYPE : in std_logic_vector
            (1 downto 0);  PC_IN, A_IN, B_IN, IMM_IN : in std_logic_vector (31 
            downto 0);  ADD_WR_IN, ADD_RS1_IN, ADD_RS2_IN, ADD_WR_MEM, 
            ADD_WR_WB : in std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB 
            : in std_logic;  OP_MEM, OP_WB : in std_logic_vector (31 downto 0);
            PC_SEL : out std_logic_vector (1 downto 0);  ZERO_FLAG : out 
            std_logic;  NPC_ABS, NPC_REL, ALU_RES, B_OUT : out std_logic_vector
            (31 downto 0);  ADD_WR_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component Decode
      port( CLK, RST, REG_LATCH_EN, RD1, RD2, RF_WE, ZERO_FLAG : in std_logic; 
            PC_IN, INS_IN : in std_logic_vector (31 downto 0);  ADD_WR : in 
            std_logic_vector (4 downto 0);  DATA_WR_IN : in std_logic_vector 
            (31 downto 0);  PC_OUT, A_OUT, B_OUT, IMM_OUT : out 
            std_logic_vector (31 downto 0);  ADD_RS1_HDU, ADD_RS2_HDU, 
            ADD_WR_OUT, ADD_RS1_OUT, ADD_RS2_OUT : out std_logic_vector (4 
            downto 0));
   end component;
   
   component Fetch
      port( CLK, RST, ZERO_FLAG : in std_logic;  PC_EXT, INS_IN : in 
            std_logic_vector (31 downto 0);  Bubble_in : in std_logic;  
            HDU_INS_IN, HDU_PC_IN, HDU_NPC_IN : in std_logic_vector (31 downto 
            0);  PC_OUT, ADDR_OUT, NPC_OUT, INS_OUT : out std_logic_vector (31 
            downto 0));
   end component;
   
   signal X_Logic1_port, INS_OUT_31_port, INS_OUT_30_port, INS_OUT_29_port, 
      INS_OUT_28_port, INS_OUT_27_port, INS_OUT_26_port, INS_OUT_25_port, 
      INS_OUT_24_port, INS_OUT_23_port, INS_OUT_22_port, INS_OUT_21_port, 
      INS_OUT_20_port, INS_OUT_19_port, INS_OUT_18_port, INS_OUT_17_port, 
      INS_OUT_16_port, INS_OUT_15_port, INS_OUT_14_port, INS_OUT_13_port, 
      INS_OUT_12_port, INS_OUT_11_port, INS_OUT_10_port, INS_OUT_9_port, 
      INS_OUT_8_port, INS_OUT_7_port, INS_OUT_6_port, INS_OUT_5_port, 
      INS_OUT_4_port, INS_OUT_3_port, INS_OUT_2_port, INS_OUT_1_port, 
      INS_OUT_0_port, n2, ZERO_FLAG_EX, PC_MEM_OUT_31_port, PC_MEM_OUT_30_port,
      PC_MEM_OUT_29_port, PC_MEM_OUT_28_port, PC_MEM_OUT_27_port, 
      PC_MEM_OUT_26_port, PC_MEM_OUT_25_port, PC_MEM_OUT_24_port, 
      PC_MEM_OUT_23_port, PC_MEM_OUT_22_port, PC_MEM_OUT_21_port, 
      PC_MEM_OUT_20_port, PC_MEM_OUT_19_port, PC_MEM_OUT_18_port, 
      PC_MEM_OUT_17_port, PC_MEM_OUT_16_port, PC_MEM_OUT_15_port, 
      PC_MEM_OUT_14_port, PC_MEM_OUT_13_port, PC_MEM_OUT_12_port, 
      PC_MEM_OUT_11_port, PC_MEM_OUT_10_port, PC_MEM_OUT_9_port, 
      PC_MEM_OUT_8_port, PC_MEM_OUT_7_port, PC_MEM_OUT_6_port, 
      PC_MEM_OUT_5_port, PC_MEM_OUT_4_port, PC_MEM_OUT_3_port, 
      PC_MEM_OUT_2_port, PC_MEM_OUT_1_port, PC_MEM_OUT_0_port, 
      sig_HDU_INS_OUT_31_port, sig_HDU_INS_OUT_30_port, sig_HDU_INS_OUT_29_port
      , sig_HDU_INS_OUT_28_port, sig_HDU_INS_OUT_27_port, 
      sig_HDU_INS_OUT_26_port, sig_HDU_INS_OUT_25_port, sig_HDU_INS_OUT_24_port
      , sig_HDU_INS_OUT_23_port, sig_HDU_INS_OUT_22_port, 
      sig_HDU_INS_OUT_21_port, sig_HDU_INS_OUT_20_port, sig_HDU_INS_OUT_19_port
      , sig_HDU_INS_OUT_18_port, sig_HDU_INS_OUT_17_port, 
      sig_HDU_INS_OUT_16_port, sig_HDU_INS_OUT_15_port, sig_HDU_INS_OUT_14_port
      , sig_HDU_INS_OUT_13_port, sig_HDU_INS_OUT_12_port, 
      sig_HDU_INS_OUT_11_port, sig_HDU_INS_OUT_10_port, sig_HDU_INS_OUT_9_port,
      sig_HDU_INS_OUT_8_port, sig_HDU_INS_OUT_7_port, sig_HDU_INS_OUT_6_port, 
      sig_HDU_INS_OUT_5_port, sig_HDU_INS_OUT_4_port, sig_HDU_INS_OUT_3_port, 
      sig_HDU_INS_OUT_2_port, sig_HDU_INS_OUT_1_port, sig_HDU_INS_OUT_0_port, 
      sig_HDU_PC_OUT_31_port, sig_HDU_PC_OUT_30_port, sig_HDU_PC_OUT_29_port, 
      sig_HDU_PC_OUT_28_port, sig_HDU_PC_OUT_27_port, sig_HDU_PC_OUT_26_port, 
      sig_HDU_PC_OUT_25_port, sig_HDU_PC_OUT_24_port, sig_HDU_PC_OUT_23_port, 
      sig_HDU_PC_OUT_22_port, sig_HDU_PC_OUT_21_port, sig_HDU_PC_OUT_20_port, 
      sig_HDU_PC_OUT_19_port, sig_HDU_PC_OUT_18_port, sig_HDU_PC_OUT_17_port, 
      sig_HDU_PC_OUT_16_port, sig_HDU_PC_OUT_15_port, sig_HDU_PC_OUT_14_port, 
      sig_HDU_PC_OUT_13_port, sig_HDU_PC_OUT_12_port, sig_HDU_PC_OUT_11_port, 
      sig_HDU_PC_OUT_10_port, sig_HDU_PC_OUT_9_port, sig_HDU_PC_OUT_8_port, 
      sig_HDU_PC_OUT_7_port, sig_HDU_PC_OUT_6_port, sig_HDU_PC_OUT_5_port, 
      sig_HDU_PC_OUT_4_port, sig_HDU_PC_OUT_3_port, sig_HDU_PC_OUT_2_port, 
      sig_HDU_PC_OUT_1_port, sig_HDU_PC_OUT_0_port, sig_HDU_NPC_OUT_31_port, 
      sig_HDU_NPC_OUT_30_port, sig_HDU_NPC_OUT_29_port, sig_HDU_NPC_OUT_28_port
      , sig_HDU_NPC_OUT_27_port, sig_HDU_NPC_OUT_26_port, 
      sig_HDU_NPC_OUT_25_port, sig_HDU_NPC_OUT_24_port, sig_HDU_NPC_OUT_23_port
      , sig_HDU_NPC_OUT_22_port, sig_HDU_NPC_OUT_21_port, 
      sig_HDU_NPC_OUT_20_port, sig_HDU_NPC_OUT_19_port, sig_HDU_NPC_OUT_18_port
      , sig_HDU_NPC_OUT_17_port, sig_HDU_NPC_OUT_16_port, 
      sig_HDU_NPC_OUT_15_port, sig_HDU_NPC_OUT_14_port, sig_HDU_NPC_OUT_13_port
      , sig_HDU_NPC_OUT_12_port, sig_HDU_NPC_OUT_11_port, 
      sig_HDU_NPC_OUT_10_port, sig_HDU_NPC_OUT_9_port, sig_HDU_NPC_OUT_8_port, 
      sig_HDU_NPC_OUT_7_port, sig_HDU_NPC_OUT_6_port, sig_HDU_NPC_OUT_5_port, 
      sig_HDU_NPC_OUT_4_port, sig_HDU_NPC_OUT_3_port, sig_HDU_NPC_OUT_2_port, 
      sig_HDU_NPC_OUT_1_port, sig_HDU_NPC_OUT_0_port, PC_FETCH_OUT_31_port, 
      PC_FETCH_OUT_30_port, PC_FETCH_OUT_29_port, PC_FETCH_OUT_28_port, 
      PC_FETCH_OUT_27_port, PC_FETCH_OUT_26_port, PC_FETCH_OUT_25_port, 
      PC_FETCH_OUT_24_port, PC_FETCH_OUT_23_port, PC_FETCH_OUT_22_port, 
      PC_FETCH_OUT_21_port, PC_FETCH_OUT_20_port, PC_FETCH_OUT_19_port, 
      PC_FETCH_OUT_18_port, PC_FETCH_OUT_17_port, PC_FETCH_OUT_16_port, 
      PC_FETCH_OUT_15_port, PC_FETCH_OUT_14_port, PC_FETCH_OUT_13_port, 
      PC_FETCH_OUT_12_port, PC_FETCH_OUT_11_port, PC_FETCH_OUT_10_port, 
      PC_FETCH_OUT_9_port, PC_FETCH_OUT_8_port, PC_FETCH_OUT_7_port, 
      PC_FETCH_OUT_6_port, PC_FETCH_OUT_5_port, PC_FETCH_OUT_4_port, 
      PC_FETCH_OUT_3_port, PC_FETCH_OUT_2_port, PC_FETCH_OUT_1_port, 
      PC_FETCH_OUT_0_port, NPC_FETCH_OUT_31_port, NPC_FETCH_OUT_30_port, 
      NPC_FETCH_OUT_29_port, NPC_FETCH_OUT_28_port, NPC_FETCH_OUT_27_port, 
      NPC_FETCH_OUT_26_port, NPC_FETCH_OUT_25_port, NPC_FETCH_OUT_24_port, 
      NPC_FETCH_OUT_23_port, NPC_FETCH_OUT_22_port, NPC_FETCH_OUT_21_port, 
      NPC_FETCH_OUT_20_port, NPC_FETCH_OUT_19_port, NPC_FETCH_OUT_18_port, 
      NPC_FETCH_OUT_17_port, NPC_FETCH_OUT_16_port, NPC_FETCH_OUT_15_port, 
      NPC_FETCH_OUT_14_port, NPC_FETCH_OUT_13_port, NPC_FETCH_OUT_12_port, 
      NPC_FETCH_OUT_11_port, NPC_FETCH_OUT_10_port, NPC_FETCH_OUT_9_port, 
      NPC_FETCH_OUT_8_port, NPC_FETCH_OUT_7_port, NPC_FETCH_OUT_6_port, 
      NPC_FETCH_OUT_5_port, NPC_FETCH_OUT_4_port, NPC_FETCH_OUT_3_port, 
      NPC_FETCH_OUT_2_port, NPC_FETCH_OUT_1_port, NPC_FETCH_OUT_0_port, 
      RF_WE_WB, ADD_WR_WB_4_port, ADD_WR_WB_3_port, ADD_WR_WB_2_port, 
      ADD_WR_WB_1_port, ADD_WR_WB_0_port, OP_WB_31_port, OP_WB_30_port, 
      OP_WB_29_port, OP_WB_28_port, OP_WB_27_port, OP_WB_26_port, OP_WB_25_port
      , OP_WB_24_port, OP_WB_23_port, OP_WB_22_port, OP_WB_21_port, 
      OP_WB_20_port, OP_WB_19_port, OP_WB_18_port, OP_WB_17_port, OP_WB_16_port
      , OP_WB_15_port, OP_WB_14_port, OP_WB_13_port, OP_WB_12_port, 
      OP_WB_11_port, OP_WB_10_port, OP_WB_9_port, OP_WB_8_port, OP_WB_7_port, 
      OP_WB_6_port, OP_WB_5_port, OP_WB_4_port, OP_WB_3_port, OP_WB_2_port, 
      OP_WB_1_port, OP_WB_0_port, PC_DECODE_OUT_31_port, PC_DECODE_OUT_30_port,
      PC_DECODE_OUT_29_port, PC_DECODE_OUT_28_port, PC_DECODE_OUT_27_port, 
      PC_DECODE_OUT_26_port, PC_DECODE_OUT_25_port, PC_DECODE_OUT_24_port, 
      PC_DECODE_OUT_23_port, PC_DECODE_OUT_22_port, PC_DECODE_OUT_21_port, 
      PC_DECODE_OUT_20_port, PC_DECODE_OUT_19_port, PC_DECODE_OUT_18_port, 
      PC_DECODE_OUT_17_port, PC_DECODE_OUT_16_port, PC_DECODE_OUT_15_port, 
      PC_DECODE_OUT_14_port, PC_DECODE_OUT_13_port, PC_DECODE_OUT_12_port, 
      PC_DECODE_OUT_11_port, PC_DECODE_OUT_10_port, PC_DECODE_OUT_9_port, 
      PC_DECODE_OUT_8_port, PC_DECODE_OUT_7_port, PC_DECODE_OUT_6_port, 
      PC_DECODE_OUT_5_port, PC_DECODE_OUT_4_port, PC_DECODE_OUT_3_port, 
      PC_DECODE_OUT_2_port, PC_DECODE_OUT_1_port, PC_DECODE_OUT_0_port, 
      A_DECODE_OUT_31_port, A_DECODE_OUT_30_port, A_DECODE_OUT_29_port, 
      A_DECODE_OUT_28_port, A_DECODE_OUT_27_port, A_DECODE_OUT_26_port, 
      A_DECODE_OUT_25_port, A_DECODE_OUT_24_port, A_DECODE_OUT_23_port, 
      A_DECODE_OUT_22_port, A_DECODE_OUT_21_port, A_DECODE_OUT_20_port, 
      A_DECODE_OUT_19_port, A_DECODE_OUT_18_port, A_DECODE_OUT_17_port, 
      A_DECODE_OUT_16_port, A_DECODE_OUT_15_port, A_DECODE_OUT_14_port, 
      A_DECODE_OUT_13_port, A_DECODE_OUT_12_port, A_DECODE_OUT_11_port, 
      A_DECODE_OUT_10_port, A_DECODE_OUT_9_port, A_DECODE_OUT_8_port, 
      A_DECODE_OUT_7_port, A_DECODE_OUT_6_port, A_DECODE_OUT_5_port, 
      A_DECODE_OUT_4_port, A_DECODE_OUT_3_port, A_DECODE_OUT_2_port, 
      A_DECODE_OUT_1_port, A_DECODE_OUT_0_port, B_DECODE_OUT_31_port, 
      B_DECODE_OUT_30_port, B_DECODE_OUT_29_port, B_DECODE_OUT_28_port, 
      B_DECODE_OUT_27_port, B_DECODE_OUT_26_port, B_DECODE_OUT_25_port, 
      B_DECODE_OUT_24_port, B_DECODE_OUT_23_port, B_DECODE_OUT_22_port, 
      B_DECODE_OUT_21_port, B_DECODE_OUT_20_port, B_DECODE_OUT_19_port, 
      B_DECODE_OUT_18_port, B_DECODE_OUT_17_port, B_DECODE_OUT_16_port, 
      B_DECODE_OUT_15_port, B_DECODE_OUT_14_port, B_DECODE_OUT_13_port, 
      B_DECODE_OUT_12_port, B_DECODE_OUT_11_port, B_DECODE_OUT_10_port, 
      B_DECODE_OUT_9_port, B_DECODE_OUT_8_port, B_DECODE_OUT_7_port, 
      B_DECODE_OUT_6_port, B_DECODE_OUT_5_port, B_DECODE_OUT_4_port, 
      B_DECODE_OUT_3_port, B_DECODE_OUT_2_port, B_DECODE_OUT_1_port, 
      B_DECODE_OUT_0_port, IMM_DECODE_OUT_31_port, IMM_DECODE_OUT_30_port, 
      IMM_DECODE_OUT_29_port, IMM_DECODE_OUT_28_port, IMM_DECODE_OUT_27_port, 
      IMM_DECODE_OUT_26_port, IMM_DECODE_OUT_25_port, IMM_DECODE_OUT_24_port, 
      IMM_DECODE_OUT_23_port, IMM_DECODE_OUT_22_port, IMM_DECODE_OUT_21_port, 
      IMM_DECODE_OUT_20_port, IMM_DECODE_OUT_19_port, IMM_DECODE_OUT_18_port, 
      IMM_DECODE_OUT_17_port, IMM_DECODE_OUT_16_port, IMM_DECODE_OUT_15_port, 
      IMM_DECODE_OUT_14_port, IMM_DECODE_OUT_13_port, IMM_DECODE_OUT_12_port, 
      IMM_DECODE_OUT_11_port, IMM_DECODE_OUT_10_port, IMM_DECODE_OUT_9_port, 
      IMM_DECODE_OUT_8_port, IMM_DECODE_OUT_7_port, IMM_DECODE_OUT_6_port, 
      IMM_DECODE_OUT_5_port, IMM_DECODE_OUT_4_port, IMM_DECODE_OUT_3_port, 
      IMM_DECODE_OUT_2_port, IMM_DECODE_OUT_1_port, IMM_DECODE_OUT_0_port, 
      ADD_RS1_HDU_4_port, ADD_RS1_HDU_3_port, ADD_RS1_HDU_2_port, 
      ADD_RS1_HDU_1_port, ADD_RS1_HDU_0_port, ADD_RS2_HDU_4_port, 
      ADD_RS2_HDU_3_port, ADD_RS2_HDU_2_port, ADD_RS2_HDU_1_port, 
      ADD_RS2_HDU_0_port, ADD_WR_DECODE_OUT_4_port, ADD_WR_DECODE_OUT_3_port, 
      ADD_WR_DECODE_OUT_2_port, ADD_WR_DECODE_OUT_1_port, 
      ADD_WR_DECODE_OUT_0_port, ADD_RS1_DECODE_OUT_4_port, 
      ADD_RS1_DECODE_OUT_3_port, ADD_RS1_DECODE_OUT_2_port, 
      ADD_RS1_DECODE_OUT_1_port, ADD_RS1_DECODE_OUT_0_port, 
      ADD_RS2_DECODE_OUT_4_port, ADD_RS2_DECODE_OUT_3_port, 
      ADD_RS2_DECODE_OUT_2_port, ADD_RS2_DECODE_OUT_1_port, 
      ADD_RS2_DECODE_OUT_0_port, ADD_WR_MEM_4_port, ADD_WR_MEM_3_port, 
      ADD_WR_MEM_2_port, ADD_WR_MEM_1_port, ADD_WR_MEM_0_port, OP_MEM_31_port, 
      OP_MEM_30_port, OP_MEM_29_port, OP_MEM_28_port, OP_MEM_27_port, 
      OP_MEM_26_port, OP_MEM_25_port, OP_MEM_24_port, OP_MEM_23_port, 
      OP_MEM_22_port, OP_MEM_21_port, OP_MEM_20_port, OP_MEM_19_port, 
      OP_MEM_18_port, OP_MEM_17_port, OP_MEM_16_port, OP_MEM_15_port, 
      OP_MEM_14_port, OP_MEM_13_port, OP_MEM_12_port, OP_MEM_11_port, 
      OP_MEM_10_port, OP_MEM_9_port, OP_MEM_8_port, OP_MEM_7_port, 
      OP_MEM_6_port, OP_MEM_5_port, OP_MEM_4_port, OP_MEM_3_port, OP_MEM_2_port
      , OP_MEM_1_port, OP_MEM_0_port, PC_SEL_EX_1_port, PC_SEL_EX_0_port, 
      NPC_ABS_EX_31_port, NPC_ABS_EX_30_port, NPC_ABS_EX_29_port, 
      NPC_ABS_EX_28_port, NPC_ABS_EX_27_port, NPC_ABS_EX_26_port, 
      NPC_ABS_EX_25_port, NPC_ABS_EX_24_port, NPC_ABS_EX_23_port, 
      NPC_ABS_EX_22_port, NPC_ABS_EX_21_port, NPC_ABS_EX_20_port, 
      NPC_ABS_EX_19_port, NPC_ABS_EX_18_port, NPC_ABS_EX_17_port, 
      NPC_ABS_EX_16_port, NPC_ABS_EX_15_port, NPC_ABS_EX_14_port, 
      NPC_ABS_EX_13_port, NPC_ABS_EX_12_port, NPC_ABS_EX_11_port, 
      NPC_ABS_EX_10_port, NPC_ABS_EX_9_port, NPC_ABS_EX_8_port, 
      NPC_ABS_EX_7_port, NPC_ABS_EX_6_port, NPC_ABS_EX_5_port, 
      NPC_ABS_EX_4_port, NPC_ABS_EX_3_port, NPC_ABS_EX_2_port, 
      NPC_ABS_EX_1_port, NPC_ABS_EX_0_port, NPC_REL_EX_31_port, 
      NPC_REL_EX_30_port, NPC_REL_EX_29_port, NPC_REL_EX_28_port, 
      NPC_REL_EX_27_port, NPC_REL_EX_26_port, NPC_REL_EX_25_port, 
      NPC_REL_EX_24_port, NPC_REL_EX_23_port, NPC_REL_EX_22_port, 
      NPC_REL_EX_21_port, NPC_REL_EX_20_port, NPC_REL_EX_19_port, 
      NPC_REL_EX_18_port, NPC_REL_EX_17_port, NPC_REL_EX_16_port, 
      NPC_REL_EX_15_port, NPC_REL_EX_14_port, NPC_REL_EX_13_port, 
      NPC_REL_EX_12_port, NPC_REL_EX_11_port, NPC_REL_EX_10_port, 
      NPC_REL_EX_9_port, NPC_REL_EX_8_port, NPC_REL_EX_7_port, 
      NPC_REL_EX_6_port, NPC_REL_EX_5_port, NPC_REL_EX_4_port, 
      NPC_REL_EX_3_port, NPC_REL_EX_2_port, NPC_REL_EX_1_port, 
      NPC_REL_EX_0_port, ALU_RES_EX_31_port, ALU_RES_EX_30_port, 
      ALU_RES_EX_29_port, ALU_RES_EX_28_port, ALU_RES_EX_27_port, 
      ALU_RES_EX_26_port, ALU_RES_EX_25_port, ALU_RES_EX_24_port, 
      ALU_RES_EX_23_port, ALU_RES_EX_22_port, ALU_RES_EX_21_port, 
      ALU_RES_EX_20_port, ALU_RES_EX_19_port, ALU_RES_EX_18_port, 
      ALU_RES_EX_17_port, ALU_RES_EX_16_port, ALU_RES_EX_15_port, 
      ALU_RES_EX_14_port, ALU_RES_EX_13_port, ALU_RES_EX_12_port, 
      ALU_RES_EX_11_port, ALU_RES_EX_10_port, ALU_RES_EX_9_port, 
      ALU_RES_EX_8_port, ALU_RES_EX_7_port, ALU_RES_EX_6_port, 
      ALU_RES_EX_5_port, ALU_RES_EX_4_port, ALU_RES_EX_3_port, 
      ALU_RES_EX_2_port, ALU_RES_EX_1_port, ALU_RES_EX_0_port, B_EX_OUT_31_port
      , B_EX_OUT_30_port, B_EX_OUT_29_port, B_EX_OUT_28_port, B_EX_OUT_27_port,
      B_EX_OUT_26_port, B_EX_OUT_25_port, B_EX_OUT_24_port, B_EX_OUT_23_port, 
      B_EX_OUT_22_port, B_EX_OUT_21_port, B_EX_OUT_20_port, B_EX_OUT_19_port, 
      B_EX_OUT_18_port, B_EX_OUT_17_port, B_EX_OUT_16_port, B_EX_OUT_15_port, 
      B_EX_OUT_14_port, B_EX_OUT_13_port, B_EX_OUT_12_port, B_EX_OUT_11_port, 
      B_EX_OUT_10_port, B_EX_OUT_9_port, B_EX_OUT_8_port, B_EX_OUT_7_port, 
      B_EX_OUT_6_port, B_EX_OUT_5_port, B_EX_OUT_4_port, B_EX_OUT_3_port, 
      B_EX_OUT_2_port, B_EX_OUT_1_port, B_EX_OUT_0_port, ADD_WR_EX_OUT_4_port, 
      ADD_WR_EX_OUT_3_port, ADD_WR_EX_OUT_2_port, ADD_WR_EX_OUT_1_port, 
      ADD_WR_EX_OUT_0_port, DRAM_R_MEM, DATA_MEM_OUT_31_port, 
      DATA_MEM_OUT_30_port, DATA_MEM_OUT_29_port, DATA_MEM_OUT_28_port, 
      DATA_MEM_OUT_27_port, DATA_MEM_OUT_26_port, DATA_MEM_OUT_25_port, 
      DATA_MEM_OUT_24_port, DATA_MEM_OUT_23_port, DATA_MEM_OUT_22_port, 
      DATA_MEM_OUT_21_port, DATA_MEM_OUT_20_port, DATA_MEM_OUT_19_port, 
      DATA_MEM_OUT_18_port, DATA_MEM_OUT_17_port, DATA_MEM_OUT_16_port, 
      DATA_MEM_OUT_15_port, DATA_MEM_OUT_14_port, DATA_MEM_OUT_13_port, 
      DATA_MEM_OUT_12_port, DATA_MEM_OUT_11_port, DATA_MEM_OUT_10_port, 
      DATA_MEM_OUT_9_port, DATA_MEM_OUT_8_port, DATA_MEM_OUT_7_port, 
      DATA_MEM_OUT_6_port, DATA_MEM_OUT_5_port, DATA_MEM_OUT_4_port, 
      DATA_MEM_OUT_3_port, DATA_MEM_OUT_2_port, DATA_MEM_OUT_1_port, 
      DATA_MEM_OUT_0_port, ALU_RES_MEM_31_port, ALU_RES_MEM_30_port, 
      ALU_RES_MEM_29_port, ALU_RES_MEM_28_port, ALU_RES_MEM_27_port, 
      ALU_RES_MEM_26_port, ALU_RES_MEM_25_port, ALU_RES_MEM_24_port, 
      ALU_RES_MEM_23_port, ALU_RES_MEM_22_port, ALU_RES_MEM_21_port, 
      ALU_RES_MEM_20_port, ALU_RES_MEM_19_port, ALU_RES_MEM_18_port, 
      ALU_RES_MEM_17_port, ALU_RES_MEM_16_port, ALU_RES_MEM_15_port, 
      ALU_RES_MEM_14_port, ALU_RES_MEM_13_port, ALU_RES_MEM_12_port, 
      ALU_RES_MEM_11_port, ALU_RES_MEM_10_port, ALU_RES_MEM_9_port, 
      ALU_RES_MEM_8_port, ALU_RES_MEM_7_port, ALU_RES_MEM_6_port, 
      ALU_RES_MEM_5_port, ALU_RES_MEM_4_port, ALU_RES_MEM_3_port, 
      ALU_RES_MEM_2_port, ALU_RES_MEM_1_port, ALU_RES_MEM_0_port, 
      ADD_WR_MEM_OUT_4_port, ADD_WR_MEM_OUT_3_port, ADD_WR_MEM_OUT_2_port, 
      ADD_WR_MEM_OUT_1_port, ADD_WR_MEM_OUT_0_port, Bubble_out_port : std_logic
      ;

begin
   INS_OUT <= ( INS_OUT_31_port, INS_OUT_30_port, INS_OUT_29_port, 
      INS_OUT_28_port, INS_OUT_27_port, INS_OUT_26_port, INS_OUT_25_port, 
      INS_OUT_24_port, INS_OUT_23_port, INS_OUT_22_port, INS_OUT_21_port, 
      INS_OUT_20_port, INS_OUT_19_port, INS_OUT_18_port, INS_OUT_17_port, 
      INS_OUT_16_port, INS_OUT_15_port, INS_OUT_14_port, INS_OUT_13_port, 
      INS_OUT_12_port, INS_OUT_11_port, INS_OUT_10_port, INS_OUT_9_port, 
      INS_OUT_8_port, INS_OUT_7_port, INS_OUT_6_port, INS_OUT_5_port, 
      INS_OUT_4_port, INS_OUT_3_port, INS_OUT_2_port, INS_OUT_1_port, 
      INS_OUT_0_port );
   Bubble_out <= Bubble_out_port;
   
   X_Logic1_port <= '1';
   FetchStage : Fetch port map( CLK => CLK, RST => RST, ZERO_FLAG => 
                           ZERO_FLAG_EX, PC_EXT(31) => PC_MEM_OUT_31_port, 
                           PC_EXT(30) => PC_MEM_OUT_30_port, PC_EXT(29) => 
                           PC_MEM_OUT_29_port, PC_EXT(28) => PC_MEM_OUT_28_port
                           , PC_EXT(27) => PC_MEM_OUT_27_port, PC_EXT(26) => 
                           PC_MEM_OUT_26_port, PC_EXT(25) => PC_MEM_OUT_25_port
                           , PC_EXT(24) => PC_MEM_OUT_24_port, PC_EXT(23) => 
                           PC_MEM_OUT_23_port, PC_EXT(22) => PC_MEM_OUT_22_port
                           , PC_EXT(21) => PC_MEM_OUT_21_port, PC_EXT(20) => 
                           PC_MEM_OUT_20_port, PC_EXT(19) => PC_MEM_OUT_19_port
                           , PC_EXT(18) => PC_MEM_OUT_18_port, PC_EXT(17) => 
                           PC_MEM_OUT_17_port, PC_EXT(16) => PC_MEM_OUT_16_port
                           , PC_EXT(15) => PC_MEM_OUT_15_port, PC_EXT(14) => 
                           PC_MEM_OUT_14_port, PC_EXT(13) => PC_MEM_OUT_13_port
                           , PC_EXT(12) => PC_MEM_OUT_12_port, PC_EXT(11) => 
                           PC_MEM_OUT_11_port, PC_EXT(10) => PC_MEM_OUT_10_port
                           , PC_EXT(9) => PC_MEM_OUT_9_port, PC_EXT(8) => 
                           PC_MEM_OUT_8_port, PC_EXT(7) => PC_MEM_OUT_7_port, 
                           PC_EXT(6) => PC_MEM_OUT_6_port, PC_EXT(5) => 
                           PC_MEM_OUT_5_port, PC_EXT(4) => PC_MEM_OUT_4_port, 
                           PC_EXT(3) => PC_MEM_OUT_3_port, PC_EXT(2) => 
                           PC_MEM_OUT_2_port, PC_EXT(1) => PC_MEM_OUT_1_port, 
                           PC_EXT(0) => PC_MEM_OUT_0_port, INS_IN(31) => 
                           INS_IN(31), INS_IN(30) => INS_IN(30), INS_IN(29) => 
                           INS_IN(29), INS_IN(28) => INS_IN(28), INS_IN(27) => 
                           INS_IN(27), INS_IN(26) => INS_IN(26), INS_IN(25) => 
                           INS_IN(25), INS_IN(24) => INS_IN(24), INS_IN(23) => 
                           INS_IN(23), INS_IN(22) => INS_IN(22), INS_IN(21) => 
                           INS_IN(21), INS_IN(20) => INS_IN(20), INS_IN(19) => 
                           INS_IN(19), INS_IN(18) => INS_IN(18), INS_IN(17) => 
                           INS_IN(17), INS_IN(16) => INS_IN(16), INS_IN(15) => 
                           INS_IN(15), INS_IN(14) => INS_IN(14), INS_IN(13) => 
                           INS_IN(13), INS_IN(12) => INS_IN(12), INS_IN(11) => 
                           INS_IN(11), INS_IN(10) => INS_IN(10), INS_IN(9) => 
                           INS_IN(9), INS_IN(8) => INS_IN(8), INS_IN(7) => 
                           INS_IN(7), INS_IN(6) => INS_IN(6), INS_IN(5) => 
                           INS_IN(5), INS_IN(4) => INS_IN(4), INS_IN(3) => 
                           INS_IN(3), INS_IN(2) => INS_IN(2), INS_IN(1) => 
                           INS_IN(1), INS_IN(0) => INS_IN(0), Bubble_in => 
                           Bubble_out_port, HDU_INS_IN(31) => 
                           sig_HDU_INS_OUT_31_port, HDU_INS_IN(30) => 
                           sig_HDU_INS_OUT_30_port, HDU_INS_IN(29) => 
                           sig_HDU_INS_OUT_29_port, HDU_INS_IN(28) => 
                           sig_HDU_INS_OUT_28_port, HDU_INS_IN(27) => 
                           sig_HDU_INS_OUT_27_port, HDU_INS_IN(26) => 
                           sig_HDU_INS_OUT_26_port, HDU_INS_IN(25) => 
                           sig_HDU_INS_OUT_25_port, HDU_INS_IN(24) => 
                           sig_HDU_INS_OUT_24_port, HDU_INS_IN(23) => 
                           sig_HDU_INS_OUT_23_port, HDU_INS_IN(22) => 
                           sig_HDU_INS_OUT_22_port, HDU_INS_IN(21) => 
                           sig_HDU_INS_OUT_21_port, HDU_INS_IN(20) => 
                           sig_HDU_INS_OUT_20_port, HDU_INS_IN(19) => 
                           sig_HDU_INS_OUT_19_port, HDU_INS_IN(18) => 
                           sig_HDU_INS_OUT_18_port, HDU_INS_IN(17) => 
                           sig_HDU_INS_OUT_17_port, HDU_INS_IN(16) => 
                           sig_HDU_INS_OUT_16_port, HDU_INS_IN(15) => 
                           sig_HDU_INS_OUT_15_port, HDU_INS_IN(14) => 
                           sig_HDU_INS_OUT_14_port, HDU_INS_IN(13) => 
                           sig_HDU_INS_OUT_13_port, HDU_INS_IN(12) => 
                           sig_HDU_INS_OUT_12_port, HDU_INS_IN(11) => 
                           sig_HDU_INS_OUT_11_port, HDU_INS_IN(10) => 
                           sig_HDU_INS_OUT_10_port, HDU_INS_IN(9) => 
                           sig_HDU_INS_OUT_9_port, HDU_INS_IN(8) => 
                           sig_HDU_INS_OUT_8_port, HDU_INS_IN(7) => 
                           sig_HDU_INS_OUT_7_port, HDU_INS_IN(6) => 
                           sig_HDU_INS_OUT_6_port, HDU_INS_IN(5) => 
                           sig_HDU_INS_OUT_5_port, HDU_INS_IN(4) => 
                           sig_HDU_INS_OUT_4_port, HDU_INS_IN(3) => 
                           sig_HDU_INS_OUT_3_port, HDU_INS_IN(2) => 
                           sig_HDU_INS_OUT_2_port, HDU_INS_IN(1) => 
                           sig_HDU_INS_OUT_1_port, HDU_INS_IN(0) => 
                           sig_HDU_INS_OUT_0_port, HDU_PC_IN(31) => 
                           sig_HDU_PC_OUT_31_port, HDU_PC_IN(30) => 
                           sig_HDU_PC_OUT_30_port, HDU_PC_IN(29) => 
                           sig_HDU_PC_OUT_29_port, HDU_PC_IN(28) => 
                           sig_HDU_PC_OUT_28_port, HDU_PC_IN(27) => 
                           sig_HDU_PC_OUT_27_port, HDU_PC_IN(26) => 
                           sig_HDU_PC_OUT_26_port, HDU_PC_IN(25) => 
                           sig_HDU_PC_OUT_25_port, HDU_PC_IN(24) => 
                           sig_HDU_PC_OUT_24_port, HDU_PC_IN(23) => 
                           sig_HDU_PC_OUT_23_port, HDU_PC_IN(22) => 
                           sig_HDU_PC_OUT_22_port, HDU_PC_IN(21) => 
                           sig_HDU_PC_OUT_21_port, HDU_PC_IN(20) => 
                           sig_HDU_PC_OUT_20_port, HDU_PC_IN(19) => 
                           sig_HDU_PC_OUT_19_port, HDU_PC_IN(18) => 
                           sig_HDU_PC_OUT_18_port, HDU_PC_IN(17) => 
                           sig_HDU_PC_OUT_17_port, HDU_PC_IN(16) => 
                           sig_HDU_PC_OUT_16_port, HDU_PC_IN(15) => 
                           sig_HDU_PC_OUT_15_port, HDU_PC_IN(14) => 
                           sig_HDU_PC_OUT_14_port, HDU_PC_IN(13) => 
                           sig_HDU_PC_OUT_13_port, HDU_PC_IN(12) => 
                           sig_HDU_PC_OUT_12_port, HDU_PC_IN(11) => 
                           sig_HDU_PC_OUT_11_port, HDU_PC_IN(10) => 
                           sig_HDU_PC_OUT_10_port, HDU_PC_IN(9) => 
                           sig_HDU_PC_OUT_9_port, HDU_PC_IN(8) => 
                           sig_HDU_PC_OUT_8_port, HDU_PC_IN(7) => 
                           sig_HDU_PC_OUT_7_port, HDU_PC_IN(6) => 
                           sig_HDU_PC_OUT_6_port, HDU_PC_IN(5) => 
                           sig_HDU_PC_OUT_5_port, HDU_PC_IN(4) => 
                           sig_HDU_PC_OUT_4_port, HDU_PC_IN(3) => 
                           sig_HDU_PC_OUT_3_port, HDU_PC_IN(2) => 
                           sig_HDU_PC_OUT_2_port, HDU_PC_IN(1) => 
                           sig_HDU_PC_OUT_1_port, HDU_PC_IN(0) => 
                           sig_HDU_PC_OUT_0_port, HDU_NPC_IN(31) => 
                           sig_HDU_NPC_OUT_31_port, HDU_NPC_IN(30) => 
                           sig_HDU_NPC_OUT_30_port, HDU_NPC_IN(29) => 
                           sig_HDU_NPC_OUT_29_port, HDU_NPC_IN(28) => 
                           sig_HDU_NPC_OUT_28_port, HDU_NPC_IN(27) => 
                           sig_HDU_NPC_OUT_27_port, HDU_NPC_IN(26) => 
                           sig_HDU_NPC_OUT_26_port, HDU_NPC_IN(25) => 
                           sig_HDU_NPC_OUT_25_port, HDU_NPC_IN(24) => 
                           sig_HDU_NPC_OUT_24_port, HDU_NPC_IN(23) => 
                           sig_HDU_NPC_OUT_23_port, HDU_NPC_IN(22) => 
                           sig_HDU_NPC_OUT_22_port, HDU_NPC_IN(21) => 
                           sig_HDU_NPC_OUT_21_port, HDU_NPC_IN(20) => 
                           sig_HDU_NPC_OUT_20_port, HDU_NPC_IN(19) => 
                           sig_HDU_NPC_OUT_19_port, HDU_NPC_IN(18) => 
                           sig_HDU_NPC_OUT_18_port, HDU_NPC_IN(17) => 
                           sig_HDU_NPC_OUT_17_port, HDU_NPC_IN(16) => 
                           sig_HDU_NPC_OUT_16_port, HDU_NPC_IN(15) => 
                           sig_HDU_NPC_OUT_15_port, HDU_NPC_IN(14) => 
                           sig_HDU_NPC_OUT_14_port, HDU_NPC_IN(13) => 
                           sig_HDU_NPC_OUT_13_port, HDU_NPC_IN(12) => 
                           sig_HDU_NPC_OUT_12_port, HDU_NPC_IN(11) => 
                           sig_HDU_NPC_OUT_11_port, HDU_NPC_IN(10) => 
                           sig_HDU_NPC_OUT_10_port, HDU_NPC_IN(9) => 
                           sig_HDU_NPC_OUT_9_port, HDU_NPC_IN(8) => 
                           sig_HDU_NPC_OUT_8_port, HDU_NPC_IN(7) => 
                           sig_HDU_NPC_OUT_7_port, HDU_NPC_IN(6) => 
                           sig_HDU_NPC_OUT_6_port, HDU_NPC_IN(5) => 
                           sig_HDU_NPC_OUT_5_port, HDU_NPC_IN(4) => 
                           sig_HDU_NPC_OUT_4_port, HDU_NPC_IN(3) => 
                           sig_HDU_NPC_OUT_3_port, HDU_NPC_IN(2) => 
                           sig_HDU_NPC_OUT_2_port, HDU_NPC_IN(1) => 
                           sig_HDU_NPC_OUT_1_port, HDU_NPC_IN(0) => 
                           sig_HDU_NPC_OUT_0_port, PC_OUT(31) => 
                           PC_FETCH_OUT_31_port, PC_OUT(30) => 
                           PC_FETCH_OUT_30_port, PC_OUT(29) => 
                           PC_FETCH_OUT_29_port, PC_OUT(28) => 
                           PC_FETCH_OUT_28_port, PC_OUT(27) => 
                           PC_FETCH_OUT_27_port, PC_OUT(26) => 
                           PC_FETCH_OUT_26_port, PC_OUT(25) => 
                           PC_FETCH_OUT_25_port, PC_OUT(24) => 
                           PC_FETCH_OUT_24_port, PC_OUT(23) => 
                           PC_FETCH_OUT_23_port, PC_OUT(22) => 
                           PC_FETCH_OUT_22_port, PC_OUT(21) => 
                           PC_FETCH_OUT_21_port, PC_OUT(20) => 
                           PC_FETCH_OUT_20_port, PC_OUT(19) => 
                           PC_FETCH_OUT_19_port, PC_OUT(18) => 
                           PC_FETCH_OUT_18_port, PC_OUT(17) => 
                           PC_FETCH_OUT_17_port, PC_OUT(16) => 
                           PC_FETCH_OUT_16_port, PC_OUT(15) => 
                           PC_FETCH_OUT_15_port, PC_OUT(14) => 
                           PC_FETCH_OUT_14_port, PC_OUT(13) => 
                           PC_FETCH_OUT_13_port, PC_OUT(12) => 
                           PC_FETCH_OUT_12_port, PC_OUT(11) => 
                           PC_FETCH_OUT_11_port, PC_OUT(10) => 
                           PC_FETCH_OUT_10_port, PC_OUT(9) => 
                           PC_FETCH_OUT_9_port, PC_OUT(8) => 
                           PC_FETCH_OUT_8_port, PC_OUT(7) => 
                           PC_FETCH_OUT_7_port, PC_OUT(6) => 
                           PC_FETCH_OUT_6_port, PC_OUT(5) => 
                           PC_FETCH_OUT_5_port, PC_OUT(4) => 
                           PC_FETCH_OUT_4_port, PC_OUT(3) => 
                           PC_FETCH_OUT_3_port, PC_OUT(2) => 
                           PC_FETCH_OUT_2_port, PC_OUT(1) => 
                           PC_FETCH_OUT_1_port, PC_OUT(0) => 
                           PC_FETCH_OUT_0_port, ADDR_OUT(31) => 
                           IRAM_ADDR_OUT(31), ADDR_OUT(30) => IRAM_ADDR_OUT(30)
                           , ADDR_OUT(29) => IRAM_ADDR_OUT(29), ADDR_OUT(28) =>
                           IRAM_ADDR_OUT(28), ADDR_OUT(27) => IRAM_ADDR_OUT(27)
                           , ADDR_OUT(26) => IRAM_ADDR_OUT(26), ADDR_OUT(25) =>
                           IRAM_ADDR_OUT(25), ADDR_OUT(24) => IRAM_ADDR_OUT(24)
                           , ADDR_OUT(23) => IRAM_ADDR_OUT(23), ADDR_OUT(22) =>
                           IRAM_ADDR_OUT(22), ADDR_OUT(21) => IRAM_ADDR_OUT(21)
                           , ADDR_OUT(20) => IRAM_ADDR_OUT(20), ADDR_OUT(19) =>
                           IRAM_ADDR_OUT(19), ADDR_OUT(18) => IRAM_ADDR_OUT(18)
                           , ADDR_OUT(17) => IRAM_ADDR_OUT(17), ADDR_OUT(16) =>
                           IRAM_ADDR_OUT(16), ADDR_OUT(15) => IRAM_ADDR_OUT(15)
                           , ADDR_OUT(14) => IRAM_ADDR_OUT(14), ADDR_OUT(13) =>
                           IRAM_ADDR_OUT(13), ADDR_OUT(12) => IRAM_ADDR_OUT(12)
                           , ADDR_OUT(11) => IRAM_ADDR_OUT(11), ADDR_OUT(10) =>
                           IRAM_ADDR_OUT(10), ADDR_OUT(9) => IRAM_ADDR_OUT(9), 
                           ADDR_OUT(8) => IRAM_ADDR_OUT(8), ADDR_OUT(7) => 
                           IRAM_ADDR_OUT(7), ADDR_OUT(6) => IRAM_ADDR_OUT(6), 
                           ADDR_OUT(5) => IRAM_ADDR_OUT(5), ADDR_OUT(4) => 
                           IRAM_ADDR_OUT(4), ADDR_OUT(3) => IRAM_ADDR_OUT(3), 
                           ADDR_OUT(2) => IRAM_ADDR_OUT(2), ADDR_OUT(1) => 
                           IRAM_ADDR_OUT(1), ADDR_OUT(0) => IRAM_ADDR_OUT(0), 
                           NPC_OUT(31) => NPC_FETCH_OUT_31_port, NPC_OUT(30) =>
                           NPC_FETCH_OUT_30_port, NPC_OUT(29) => 
                           NPC_FETCH_OUT_29_port, NPC_OUT(28) => 
                           NPC_FETCH_OUT_28_port, NPC_OUT(27) => 
                           NPC_FETCH_OUT_27_port, NPC_OUT(26) => 
                           NPC_FETCH_OUT_26_port, NPC_OUT(25) => 
                           NPC_FETCH_OUT_25_port, NPC_OUT(24) => 
                           NPC_FETCH_OUT_24_port, NPC_OUT(23) => 
                           NPC_FETCH_OUT_23_port, NPC_OUT(22) => 
                           NPC_FETCH_OUT_22_port, NPC_OUT(21) => 
                           NPC_FETCH_OUT_21_port, NPC_OUT(20) => 
                           NPC_FETCH_OUT_20_port, NPC_OUT(19) => 
                           NPC_FETCH_OUT_19_port, NPC_OUT(18) => 
                           NPC_FETCH_OUT_18_port, NPC_OUT(17) => 
                           NPC_FETCH_OUT_17_port, NPC_OUT(16) => 
                           NPC_FETCH_OUT_16_port, NPC_OUT(15) => 
                           NPC_FETCH_OUT_15_port, NPC_OUT(14) => 
                           NPC_FETCH_OUT_14_port, NPC_OUT(13) => 
                           NPC_FETCH_OUT_13_port, NPC_OUT(12) => 
                           NPC_FETCH_OUT_12_port, NPC_OUT(11) => 
                           NPC_FETCH_OUT_11_port, NPC_OUT(10) => 
                           NPC_FETCH_OUT_10_port, NPC_OUT(9) => 
                           NPC_FETCH_OUT_9_port, NPC_OUT(8) => 
                           NPC_FETCH_OUT_8_port, NPC_OUT(7) => 
                           NPC_FETCH_OUT_7_port, NPC_OUT(6) => 
                           NPC_FETCH_OUT_6_port, NPC_OUT(5) => 
                           NPC_FETCH_OUT_5_port, NPC_OUT(4) => 
                           NPC_FETCH_OUT_4_port, NPC_OUT(3) => 
                           NPC_FETCH_OUT_3_port, NPC_OUT(2) => 
                           NPC_FETCH_OUT_2_port, NPC_OUT(1) => 
                           NPC_FETCH_OUT_1_port, NPC_OUT(0) => 
                           NPC_FETCH_OUT_0_port, INS_OUT(31) => INS_OUT_31_port
                           , INS_OUT(30) => INS_OUT_30_port, INS_OUT(29) => 
                           INS_OUT_29_port, INS_OUT(28) => INS_OUT_28_port, 
                           INS_OUT(27) => INS_OUT_27_port, INS_OUT(26) => 
                           INS_OUT_26_port, INS_OUT(25) => INS_OUT_25_port, 
                           INS_OUT(24) => INS_OUT_24_port, INS_OUT(23) => 
                           INS_OUT_23_port, INS_OUT(22) => INS_OUT_22_port, 
                           INS_OUT(21) => INS_OUT_21_port, INS_OUT(20) => 
                           INS_OUT_20_port, INS_OUT(19) => INS_OUT_19_port, 
                           INS_OUT(18) => INS_OUT_18_port, INS_OUT(17) => 
                           INS_OUT_17_port, INS_OUT(16) => INS_OUT_16_port, 
                           INS_OUT(15) => INS_OUT_15_port, INS_OUT(14) => 
                           INS_OUT_14_port, INS_OUT(13) => INS_OUT_13_port, 
                           INS_OUT(12) => INS_OUT_12_port, INS_OUT(11) => 
                           INS_OUT_11_port, INS_OUT(10) => INS_OUT_10_port, 
                           INS_OUT(9) => INS_OUT_9_port, INS_OUT(8) => 
                           INS_OUT_8_port, INS_OUT(7) => INS_OUT_7_port, 
                           INS_OUT(6) => INS_OUT_6_port, INS_OUT(5) => 
                           INS_OUT_5_port, INS_OUT(4) => INS_OUT_4_port, 
                           INS_OUT(3) => INS_OUT_3_port, INS_OUT(2) => 
                           INS_OUT_2_port, INS_OUT(1) => INS_OUT_1_port, 
                           INS_OUT(0) => INS_OUT_0_port);
   DecodeStage : Decode port map( CLK => CLK, RST => RST, REG_LATCH_EN => 
                           REG_LATCH_EN, RD1 => RD1, RD2 => RD2, RF_WE => 
                           RF_WE_WB, ZERO_FLAG => ZERO_FLAG_EX, PC_IN(31) => 
                           PC_FETCH_OUT_31_port, PC_IN(30) => 
                           PC_FETCH_OUT_30_port, PC_IN(29) => 
                           PC_FETCH_OUT_29_port, PC_IN(28) => 
                           PC_FETCH_OUT_28_port, PC_IN(27) => 
                           PC_FETCH_OUT_27_port, PC_IN(26) => 
                           PC_FETCH_OUT_26_port, PC_IN(25) => 
                           PC_FETCH_OUT_25_port, PC_IN(24) => 
                           PC_FETCH_OUT_24_port, PC_IN(23) => 
                           PC_FETCH_OUT_23_port, PC_IN(22) => 
                           PC_FETCH_OUT_22_port, PC_IN(21) => 
                           PC_FETCH_OUT_21_port, PC_IN(20) => 
                           PC_FETCH_OUT_20_port, PC_IN(19) => 
                           PC_FETCH_OUT_19_port, PC_IN(18) => 
                           PC_FETCH_OUT_18_port, PC_IN(17) => 
                           PC_FETCH_OUT_17_port, PC_IN(16) => 
                           PC_FETCH_OUT_16_port, PC_IN(15) => 
                           PC_FETCH_OUT_15_port, PC_IN(14) => 
                           PC_FETCH_OUT_14_port, PC_IN(13) => 
                           PC_FETCH_OUT_13_port, PC_IN(12) => 
                           PC_FETCH_OUT_12_port, PC_IN(11) => 
                           PC_FETCH_OUT_11_port, PC_IN(10) => 
                           PC_FETCH_OUT_10_port, PC_IN(9) => 
                           PC_FETCH_OUT_9_port, PC_IN(8) => PC_FETCH_OUT_8_port
                           , PC_IN(7) => PC_FETCH_OUT_7_port, PC_IN(6) => 
                           PC_FETCH_OUT_6_port, PC_IN(5) => PC_FETCH_OUT_5_port
                           , PC_IN(4) => PC_FETCH_OUT_4_port, PC_IN(3) => 
                           PC_FETCH_OUT_3_port, PC_IN(2) => PC_FETCH_OUT_2_port
                           , PC_IN(1) => PC_FETCH_OUT_1_port, PC_IN(0) => 
                           PC_FETCH_OUT_0_port, INS_IN(31) => INS_OUT_31_port, 
                           INS_IN(30) => INS_OUT_30_port, INS_IN(29) => 
                           INS_OUT_29_port, INS_IN(28) => INS_OUT_28_port, 
                           INS_IN(27) => INS_OUT_27_port, INS_IN(26) => 
                           INS_OUT_26_port, INS_IN(25) => INS_OUT_25_port, 
                           INS_IN(24) => INS_OUT_24_port, INS_IN(23) => 
                           INS_OUT_23_port, INS_IN(22) => INS_OUT_22_port, 
                           INS_IN(21) => INS_OUT_21_port, INS_IN(20) => 
                           INS_OUT_20_port, INS_IN(19) => INS_OUT_19_port, 
                           INS_IN(18) => INS_OUT_18_port, INS_IN(17) => 
                           INS_OUT_17_port, INS_IN(16) => INS_OUT_16_port, 
                           INS_IN(15) => INS_OUT_15_port, INS_IN(14) => 
                           INS_OUT_14_port, INS_IN(13) => INS_OUT_13_port, 
                           INS_IN(12) => INS_OUT_12_port, INS_IN(11) => 
                           INS_OUT_11_port, INS_IN(10) => INS_OUT_10_port, 
                           INS_IN(9) => INS_OUT_9_port, INS_IN(8) => 
                           INS_OUT_8_port, INS_IN(7) => INS_OUT_7_port, 
                           INS_IN(6) => INS_OUT_6_port, INS_IN(5) => 
                           INS_OUT_5_port, INS_IN(4) => INS_OUT_4_port, 
                           INS_IN(3) => INS_OUT_3_port, INS_IN(2) => 
                           INS_OUT_2_port, INS_IN(1) => INS_OUT_1_port, 
                           INS_IN(0) => INS_OUT_0_port, ADD_WR(4) => 
                           ADD_WR_WB_4_port, ADD_WR(3) => ADD_WR_WB_3_port, 
                           ADD_WR(2) => ADD_WR_WB_2_port, ADD_WR(1) => 
                           ADD_WR_WB_1_port, ADD_WR(0) => ADD_WR_WB_0_port, 
                           DATA_WR_IN(31) => OP_WB_31_port, DATA_WR_IN(30) => 
                           OP_WB_30_port, DATA_WR_IN(29) => OP_WB_29_port, 
                           DATA_WR_IN(28) => OP_WB_28_port, DATA_WR_IN(27) => 
                           OP_WB_27_port, DATA_WR_IN(26) => OP_WB_26_port, 
                           DATA_WR_IN(25) => OP_WB_25_port, DATA_WR_IN(24) => 
                           OP_WB_24_port, DATA_WR_IN(23) => OP_WB_23_port, 
                           DATA_WR_IN(22) => OP_WB_22_port, DATA_WR_IN(21) => 
                           OP_WB_21_port, DATA_WR_IN(20) => OP_WB_20_port, 
                           DATA_WR_IN(19) => OP_WB_19_port, DATA_WR_IN(18) => 
                           OP_WB_18_port, DATA_WR_IN(17) => OP_WB_17_port, 
                           DATA_WR_IN(16) => OP_WB_16_port, DATA_WR_IN(15) => 
                           OP_WB_15_port, DATA_WR_IN(14) => OP_WB_14_port, 
                           DATA_WR_IN(13) => OP_WB_13_port, DATA_WR_IN(12) => 
                           OP_WB_12_port, DATA_WR_IN(11) => OP_WB_11_port, 
                           DATA_WR_IN(10) => OP_WB_10_port, DATA_WR_IN(9) => 
                           OP_WB_9_port, DATA_WR_IN(8) => OP_WB_8_port, 
                           DATA_WR_IN(7) => OP_WB_7_port, DATA_WR_IN(6) => 
                           OP_WB_6_port, DATA_WR_IN(5) => OP_WB_5_port, 
                           DATA_WR_IN(4) => OP_WB_4_port, DATA_WR_IN(3) => 
                           OP_WB_3_port, DATA_WR_IN(2) => OP_WB_2_port, 
                           DATA_WR_IN(1) => OP_WB_1_port, DATA_WR_IN(0) => 
                           OP_WB_0_port, PC_OUT(31) => PC_DECODE_OUT_31_port, 
                           PC_OUT(30) => PC_DECODE_OUT_30_port, PC_OUT(29) => 
                           PC_DECODE_OUT_29_port, PC_OUT(28) => 
                           PC_DECODE_OUT_28_port, PC_OUT(27) => 
                           PC_DECODE_OUT_27_port, PC_OUT(26) => 
                           PC_DECODE_OUT_26_port, PC_OUT(25) => 
                           PC_DECODE_OUT_25_port, PC_OUT(24) => 
                           PC_DECODE_OUT_24_port, PC_OUT(23) => 
                           PC_DECODE_OUT_23_port, PC_OUT(22) => 
                           PC_DECODE_OUT_22_port, PC_OUT(21) => 
                           PC_DECODE_OUT_21_port, PC_OUT(20) => 
                           PC_DECODE_OUT_20_port, PC_OUT(19) => 
                           PC_DECODE_OUT_19_port, PC_OUT(18) => 
                           PC_DECODE_OUT_18_port, PC_OUT(17) => 
                           PC_DECODE_OUT_17_port, PC_OUT(16) => 
                           PC_DECODE_OUT_16_port, PC_OUT(15) => 
                           PC_DECODE_OUT_15_port, PC_OUT(14) => 
                           PC_DECODE_OUT_14_port, PC_OUT(13) => 
                           PC_DECODE_OUT_13_port, PC_OUT(12) => 
                           PC_DECODE_OUT_12_port, PC_OUT(11) => 
                           PC_DECODE_OUT_11_port, PC_OUT(10) => 
                           PC_DECODE_OUT_10_port, PC_OUT(9) => 
                           PC_DECODE_OUT_9_port, PC_OUT(8) => 
                           PC_DECODE_OUT_8_port, PC_OUT(7) => 
                           PC_DECODE_OUT_7_port, PC_OUT(6) => 
                           PC_DECODE_OUT_6_port, PC_OUT(5) => 
                           PC_DECODE_OUT_5_port, PC_OUT(4) => 
                           PC_DECODE_OUT_4_port, PC_OUT(3) => 
                           PC_DECODE_OUT_3_port, PC_OUT(2) => 
                           PC_DECODE_OUT_2_port, PC_OUT(1) => 
                           PC_DECODE_OUT_1_port, PC_OUT(0) => 
                           PC_DECODE_OUT_0_port, A_OUT(31) => 
                           A_DECODE_OUT_31_port, A_OUT(30) => 
                           A_DECODE_OUT_30_port, A_OUT(29) => 
                           A_DECODE_OUT_29_port, A_OUT(28) => 
                           A_DECODE_OUT_28_port, A_OUT(27) => 
                           A_DECODE_OUT_27_port, A_OUT(26) => 
                           A_DECODE_OUT_26_port, A_OUT(25) => 
                           A_DECODE_OUT_25_port, A_OUT(24) => 
                           A_DECODE_OUT_24_port, A_OUT(23) => 
                           A_DECODE_OUT_23_port, A_OUT(22) => 
                           A_DECODE_OUT_22_port, A_OUT(21) => 
                           A_DECODE_OUT_21_port, A_OUT(20) => 
                           A_DECODE_OUT_20_port, A_OUT(19) => 
                           A_DECODE_OUT_19_port, A_OUT(18) => 
                           A_DECODE_OUT_18_port, A_OUT(17) => 
                           A_DECODE_OUT_17_port, A_OUT(16) => 
                           A_DECODE_OUT_16_port, A_OUT(15) => 
                           A_DECODE_OUT_15_port, A_OUT(14) => 
                           A_DECODE_OUT_14_port, A_OUT(13) => 
                           A_DECODE_OUT_13_port, A_OUT(12) => 
                           A_DECODE_OUT_12_port, A_OUT(11) => 
                           A_DECODE_OUT_11_port, A_OUT(10) => 
                           A_DECODE_OUT_10_port, A_OUT(9) => 
                           A_DECODE_OUT_9_port, A_OUT(8) => A_DECODE_OUT_8_port
                           , A_OUT(7) => A_DECODE_OUT_7_port, A_OUT(6) => 
                           A_DECODE_OUT_6_port, A_OUT(5) => A_DECODE_OUT_5_port
                           , A_OUT(4) => A_DECODE_OUT_4_port, A_OUT(3) => 
                           A_DECODE_OUT_3_port, A_OUT(2) => A_DECODE_OUT_2_port
                           , A_OUT(1) => A_DECODE_OUT_1_port, A_OUT(0) => 
                           A_DECODE_OUT_0_port, B_OUT(31) => 
                           B_DECODE_OUT_31_port, B_OUT(30) => 
                           B_DECODE_OUT_30_port, B_OUT(29) => 
                           B_DECODE_OUT_29_port, B_OUT(28) => 
                           B_DECODE_OUT_28_port, B_OUT(27) => 
                           B_DECODE_OUT_27_port, B_OUT(26) => 
                           B_DECODE_OUT_26_port, B_OUT(25) => 
                           B_DECODE_OUT_25_port, B_OUT(24) => 
                           B_DECODE_OUT_24_port, B_OUT(23) => 
                           B_DECODE_OUT_23_port, B_OUT(22) => 
                           B_DECODE_OUT_22_port, B_OUT(21) => 
                           B_DECODE_OUT_21_port, B_OUT(20) => 
                           B_DECODE_OUT_20_port, B_OUT(19) => 
                           B_DECODE_OUT_19_port, B_OUT(18) => 
                           B_DECODE_OUT_18_port, B_OUT(17) => 
                           B_DECODE_OUT_17_port, B_OUT(16) => 
                           B_DECODE_OUT_16_port, B_OUT(15) => 
                           B_DECODE_OUT_15_port, B_OUT(14) => 
                           B_DECODE_OUT_14_port, B_OUT(13) => 
                           B_DECODE_OUT_13_port, B_OUT(12) => 
                           B_DECODE_OUT_12_port, B_OUT(11) => 
                           B_DECODE_OUT_11_port, B_OUT(10) => 
                           B_DECODE_OUT_10_port, B_OUT(9) => 
                           B_DECODE_OUT_9_port, B_OUT(8) => B_DECODE_OUT_8_port
                           , B_OUT(7) => B_DECODE_OUT_7_port, B_OUT(6) => 
                           B_DECODE_OUT_6_port, B_OUT(5) => B_DECODE_OUT_5_port
                           , B_OUT(4) => B_DECODE_OUT_4_port, B_OUT(3) => 
                           B_DECODE_OUT_3_port, B_OUT(2) => B_DECODE_OUT_2_port
                           , B_OUT(1) => B_DECODE_OUT_1_port, B_OUT(0) => 
                           B_DECODE_OUT_0_port, IMM_OUT(31) => 
                           IMM_DECODE_OUT_31_port, IMM_OUT(30) => 
                           IMM_DECODE_OUT_30_port, IMM_OUT(29) => 
                           IMM_DECODE_OUT_29_port, IMM_OUT(28) => 
                           IMM_DECODE_OUT_28_port, IMM_OUT(27) => 
                           IMM_DECODE_OUT_27_port, IMM_OUT(26) => 
                           IMM_DECODE_OUT_26_port, IMM_OUT(25) => 
                           IMM_DECODE_OUT_25_port, IMM_OUT(24) => 
                           IMM_DECODE_OUT_24_port, IMM_OUT(23) => 
                           IMM_DECODE_OUT_23_port, IMM_OUT(22) => 
                           IMM_DECODE_OUT_22_port, IMM_OUT(21) => 
                           IMM_DECODE_OUT_21_port, IMM_OUT(20) => 
                           IMM_DECODE_OUT_20_port, IMM_OUT(19) => 
                           IMM_DECODE_OUT_19_port, IMM_OUT(18) => 
                           IMM_DECODE_OUT_18_port, IMM_OUT(17) => 
                           IMM_DECODE_OUT_17_port, IMM_OUT(16) => 
                           IMM_DECODE_OUT_16_port, IMM_OUT(15) => 
                           IMM_DECODE_OUT_15_port, IMM_OUT(14) => 
                           IMM_DECODE_OUT_14_port, IMM_OUT(13) => 
                           IMM_DECODE_OUT_13_port, IMM_OUT(12) => 
                           IMM_DECODE_OUT_12_port, IMM_OUT(11) => 
                           IMM_DECODE_OUT_11_port, IMM_OUT(10) => 
                           IMM_DECODE_OUT_10_port, IMM_OUT(9) => 
                           IMM_DECODE_OUT_9_port, IMM_OUT(8) => 
                           IMM_DECODE_OUT_8_port, IMM_OUT(7) => 
                           IMM_DECODE_OUT_7_port, IMM_OUT(6) => 
                           IMM_DECODE_OUT_6_port, IMM_OUT(5) => 
                           IMM_DECODE_OUT_5_port, IMM_OUT(4) => 
                           IMM_DECODE_OUT_4_port, IMM_OUT(3) => 
                           IMM_DECODE_OUT_3_port, IMM_OUT(2) => 
                           IMM_DECODE_OUT_2_port, IMM_OUT(1) => 
                           IMM_DECODE_OUT_1_port, IMM_OUT(0) => 
                           IMM_DECODE_OUT_0_port, ADD_RS1_HDU(4) => 
                           ADD_RS1_HDU_4_port, ADD_RS1_HDU(3) => 
                           ADD_RS1_HDU_3_port, ADD_RS1_HDU(2) => 
                           ADD_RS1_HDU_2_port, ADD_RS1_HDU(1) => 
                           ADD_RS1_HDU_1_port, ADD_RS1_HDU(0) => 
                           ADD_RS1_HDU_0_port, ADD_RS2_HDU(4) => 
                           ADD_RS2_HDU_4_port, ADD_RS2_HDU(3) => 
                           ADD_RS2_HDU_3_port, ADD_RS2_HDU(2) => 
                           ADD_RS2_HDU_2_port, ADD_RS2_HDU(1) => 
                           ADD_RS2_HDU_1_port, ADD_RS2_HDU(0) => 
                           ADD_RS2_HDU_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_DECODE_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_DECODE_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_DECODE_OUT_0_port, ADD_RS1_OUT(4) => 
                           ADD_RS1_DECODE_OUT_4_port, ADD_RS1_OUT(3) => 
                           ADD_RS1_DECODE_OUT_3_port, ADD_RS1_OUT(2) => 
                           ADD_RS1_DECODE_OUT_2_port, ADD_RS1_OUT(1) => 
                           ADD_RS1_DECODE_OUT_1_port, ADD_RS1_OUT(0) => 
                           ADD_RS1_DECODE_OUT_0_port, ADD_RS2_OUT(4) => 
                           ADD_RS2_DECODE_OUT_4_port, ADD_RS2_OUT(3) => 
                           ADD_RS2_DECODE_OUT_3_port, ADD_RS2_OUT(2) => 
                           ADD_RS2_DECODE_OUT_2_port, ADD_RS2_OUT(1) => 
                           ADD_RS2_DECODE_OUT_1_port, ADD_RS2_OUT(0) => 
                           ADD_RS2_DECODE_OUT_0_port);
   ExecuteStage : Execute port map( CLK => CLK, RST => RST, MUX_A_SEL => 
                           MUX_A_SEL, MUX_B_SEL(1) => MUX_B_SEL(1), 
                           MUX_B_SEL(0) => MUX_B_SEL(0), ALU_OPC(0) => 
                           ALU_OPC(0), ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => 
                           ALU_OPC(2), ALU_OPC(3) => ALU_OPC(3), ALU_OUTREG_EN 
                           => ALU_OUTREG_EN, JUMP_TYPE(1) => JUMP_TYPE(1), 
                           JUMP_TYPE(0) => JUMP_TYPE(0), PC_IN(31) => 
                           PC_DECODE_OUT_31_port, PC_IN(30) => 
                           PC_DECODE_OUT_30_port, PC_IN(29) => 
                           PC_DECODE_OUT_29_port, PC_IN(28) => 
                           PC_DECODE_OUT_28_port, PC_IN(27) => 
                           PC_DECODE_OUT_27_port, PC_IN(26) => 
                           PC_DECODE_OUT_26_port, PC_IN(25) => 
                           PC_DECODE_OUT_25_port, PC_IN(24) => 
                           PC_DECODE_OUT_24_port, PC_IN(23) => 
                           PC_DECODE_OUT_23_port, PC_IN(22) => 
                           PC_DECODE_OUT_22_port, PC_IN(21) => 
                           PC_DECODE_OUT_21_port, PC_IN(20) => 
                           PC_DECODE_OUT_20_port, PC_IN(19) => 
                           PC_DECODE_OUT_19_port, PC_IN(18) => 
                           PC_DECODE_OUT_18_port, PC_IN(17) => 
                           PC_DECODE_OUT_17_port, PC_IN(16) => 
                           PC_DECODE_OUT_16_port, PC_IN(15) => 
                           PC_DECODE_OUT_15_port, PC_IN(14) => 
                           PC_DECODE_OUT_14_port, PC_IN(13) => 
                           PC_DECODE_OUT_13_port, PC_IN(12) => 
                           PC_DECODE_OUT_12_port, PC_IN(11) => 
                           PC_DECODE_OUT_11_port, PC_IN(10) => 
                           PC_DECODE_OUT_10_port, PC_IN(9) => 
                           PC_DECODE_OUT_9_port, PC_IN(8) => 
                           PC_DECODE_OUT_8_port, PC_IN(7) => 
                           PC_DECODE_OUT_7_port, PC_IN(6) => 
                           PC_DECODE_OUT_6_port, PC_IN(5) => 
                           PC_DECODE_OUT_5_port, PC_IN(4) => 
                           PC_DECODE_OUT_4_port, PC_IN(3) => 
                           PC_DECODE_OUT_3_port, PC_IN(2) => 
                           PC_DECODE_OUT_2_port, PC_IN(1) => 
                           PC_DECODE_OUT_1_port, PC_IN(0) => 
                           PC_DECODE_OUT_0_port, A_IN(31) => 
                           A_DECODE_OUT_31_port, A_IN(30) => 
                           A_DECODE_OUT_30_port, A_IN(29) => 
                           A_DECODE_OUT_29_port, A_IN(28) => 
                           A_DECODE_OUT_28_port, A_IN(27) => 
                           A_DECODE_OUT_27_port, A_IN(26) => 
                           A_DECODE_OUT_26_port, A_IN(25) => 
                           A_DECODE_OUT_25_port, A_IN(24) => 
                           A_DECODE_OUT_24_port, A_IN(23) => 
                           A_DECODE_OUT_23_port, A_IN(22) => 
                           A_DECODE_OUT_22_port, A_IN(21) => 
                           A_DECODE_OUT_21_port, A_IN(20) => 
                           A_DECODE_OUT_20_port, A_IN(19) => 
                           A_DECODE_OUT_19_port, A_IN(18) => 
                           A_DECODE_OUT_18_port, A_IN(17) => 
                           A_DECODE_OUT_17_port, A_IN(16) => 
                           A_DECODE_OUT_16_port, A_IN(15) => 
                           A_DECODE_OUT_15_port, A_IN(14) => 
                           A_DECODE_OUT_14_port, A_IN(13) => 
                           A_DECODE_OUT_13_port, A_IN(12) => 
                           A_DECODE_OUT_12_port, A_IN(11) => 
                           A_DECODE_OUT_11_port, A_IN(10) => 
                           A_DECODE_OUT_10_port, A_IN(9) => A_DECODE_OUT_9_port
                           , A_IN(8) => A_DECODE_OUT_8_port, A_IN(7) => 
                           A_DECODE_OUT_7_port, A_IN(6) => A_DECODE_OUT_6_port,
                           A_IN(5) => A_DECODE_OUT_5_port, A_IN(4) => 
                           A_DECODE_OUT_4_port, A_IN(3) => A_DECODE_OUT_3_port,
                           A_IN(2) => A_DECODE_OUT_2_port, A_IN(1) => 
                           A_DECODE_OUT_1_port, A_IN(0) => A_DECODE_OUT_0_port,
                           B_IN(31) => B_DECODE_OUT_31_port, B_IN(30) => 
                           B_DECODE_OUT_30_port, B_IN(29) => 
                           B_DECODE_OUT_29_port, B_IN(28) => 
                           B_DECODE_OUT_28_port, B_IN(27) => 
                           B_DECODE_OUT_27_port, B_IN(26) => 
                           B_DECODE_OUT_26_port, B_IN(25) => 
                           B_DECODE_OUT_25_port, B_IN(24) => 
                           B_DECODE_OUT_24_port, B_IN(23) => 
                           B_DECODE_OUT_23_port, B_IN(22) => 
                           B_DECODE_OUT_22_port, B_IN(21) => 
                           B_DECODE_OUT_21_port, B_IN(20) => 
                           B_DECODE_OUT_20_port, B_IN(19) => 
                           B_DECODE_OUT_19_port, B_IN(18) => 
                           B_DECODE_OUT_18_port, B_IN(17) => 
                           B_DECODE_OUT_17_port, B_IN(16) => 
                           B_DECODE_OUT_16_port, B_IN(15) => 
                           B_DECODE_OUT_15_port, B_IN(14) => 
                           B_DECODE_OUT_14_port, B_IN(13) => 
                           B_DECODE_OUT_13_port, B_IN(12) => 
                           B_DECODE_OUT_12_port, B_IN(11) => 
                           B_DECODE_OUT_11_port, B_IN(10) => 
                           B_DECODE_OUT_10_port, B_IN(9) => B_DECODE_OUT_9_port
                           , B_IN(8) => B_DECODE_OUT_8_port, B_IN(7) => 
                           B_DECODE_OUT_7_port, B_IN(6) => B_DECODE_OUT_6_port,
                           B_IN(5) => B_DECODE_OUT_5_port, B_IN(4) => 
                           B_DECODE_OUT_4_port, B_IN(3) => B_DECODE_OUT_3_port,
                           B_IN(2) => B_DECODE_OUT_2_port, B_IN(1) => 
                           B_DECODE_OUT_1_port, B_IN(0) => B_DECODE_OUT_0_port,
                           IMM_IN(31) => IMM_DECODE_OUT_31_port, IMM_IN(30) => 
                           IMM_DECODE_OUT_30_port, IMM_IN(29) => 
                           IMM_DECODE_OUT_29_port, IMM_IN(28) => 
                           IMM_DECODE_OUT_28_port, IMM_IN(27) => 
                           IMM_DECODE_OUT_27_port, IMM_IN(26) => 
                           IMM_DECODE_OUT_26_port, IMM_IN(25) => 
                           IMM_DECODE_OUT_25_port, IMM_IN(24) => 
                           IMM_DECODE_OUT_24_port, IMM_IN(23) => 
                           IMM_DECODE_OUT_23_port, IMM_IN(22) => 
                           IMM_DECODE_OUT_22_port, IMM_IN(21) => 
                           IMM_DECODE_OUT_21_port, IMM_IN(20) => 
                           IMM_DECODE_OUT_20_port, IMM_IN(19) => 
                           IMM_DECODE_OUT_19_port, IMM_IN(18) => 
                           IMM_DECODE_OUT_18_port, IMM_IN(17) => 
                           IMM_DECODE_OUT_17_port, IMM_IN(16) => 
                           IMM_DECODE_OUT_16_port, IMM_IN(15) => 
                           IMM_DECODE_OUT_15_port, IMM_IN(14) => 
                           IMM_DECODE_OUT_14_port, IMM_IN(13) => 
                           IMM_DECODE_OUT_13_port, IMM_IN(12) => 
                           IMM_DECODE_OUT_12_port, IMM_IN(11) => 
                           IMM_DECODE_OUT_11_port, IMM_IN(10) => 
                           IMM_DECODE_OUT_10_port, IMM_IN(9) => 
                           IMM_DECODE_OUT_9_port, IMM_IN(8) => 
                           IMM_DECODE_OUT_8_port, IMM_IN(7) => 
                           IMM_DECODE_OUT_7_port, IMM_IN(6) => 
                           IMM_DECODE_OUT_6_port, IMM_IN(5) => 
                           IMM_DECODE_OUT_5_port, IMM_IN(4) => 
                           IMM_DECODE_OUT_4_port, IMM_IN(3) => 
                           IMM_DECODE_OUT_3_port, IMM_IN(2) => 
                           IMM_DECODE_OUT_2_port, IMM_IN(1) => 
                           IMM_DECODE_OUT_1_port, IMM_IN(0) => 
                           IMM_DECODE_OUT_0_port, ADD_WR_IN(4) => 
                           ADD_WR_DECODE_OUT_4_port, ADD_WR_IN(3) => 
                           ADD_WR_DECODE_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_DECODE_OUT_0_port, ADD_RS1_IN(4) => 
                           ADD_RS1_DECODE_OUT_4_port, ADD_RS1_IN(3) => 
                           ADD_RS1_DECODE_OUT_3_port, ADD_RS1_IN(2) => 
                           ADD_RS1_DECODE_OUT_2_port, ADD_RS1_IN(1) => 
                           ADD_RS1_DECODE_OUT_1_port, ADD_RS1_IN(0) => 
                           ADD_RS1_DECODE_OUT_0_port, ADD_RS2_IN(4) => 
                           ADD_RS2_DECODE_OUT_4_port, ADD_RS2_IN(3) => 
                           ADD_RS2_DECODE_OUT_3_port, ADD_RS2_IN(2) => 
                           ADD_RS2_DECODE_OUT_2_port, ADD_RS2_IN(1) => 
                           ADD_RS2_DECODE_OUT_1_port, ADD_RS2_IN(0) => 
                           ADD_RS2_DECODE_OUT_0_port, ADD_WR_MEM(4) => 
                           ADD_WR_MEM_4_port, ADD_WR_MEM(3) => 
                           ADD_WR_MEM_3_port, ADD_WR_MEM(2) => 
                           ADD_WR_MEM_2_port, ADD_WR_MEM(1) => 
                           ADD_WR_MEM_1_port, ADD_WR_MEM(0) => 
                           ADD_WR_MEM_0_port, ADD_WR_WB(4) => ADD_WR_WB_4_port,
                           ADD_WR_WB(3) => ADD_WR_WB_3_port, ADD_WR_WB(2) => 
                           ADD_WR_WB_2_port, ADD_WR_WB(1) => ADD_WR_WB_1_port, 
                           ADD_WR_WB(0) => ADD_WR_WB_0_port, RF_WE_MEM => RF_WE
                           , RF_WE_WB => RF_WE_WB, OP_MEM(31) => OP_MEM_31_port
                           , OP_MEM(30) => OP_MEM_30_port, OP_MEM(29) => 
                           OP_MEM_29_port, OP_MEM(28) => OP_MEM_28_port, 
                           OP_MEM(27) => OP_MEM_27_port, OP_MEM(26) => 
                           OP_MEM_26_port, OP_MEM(25) => OP_MEM_25_port, 
                           OP_MEM(24) => OP_MEM_24_port, OP_MEM(23) => 
                           OP_MEM_23_port, OP_MEM(22) => OP_MEM_22_port, 
                           OP_MEM(21) => OP_MEM_21_port, OP_MEM(20) => 
                           OP_MEM_20_port, OP_MEM(19) => OP_MEM_19_port, 
                           OP_MEM(18) => OP_MEM_18_port, OP_MEM(17) => 
                           OP_MEM_17_port, OP_MEM(16) => OP_MEM_16_port, 
                           OP_MEM(15) => OP_MEM_15_port, OP_MEM(14) => 
                           OP_MEM_14_port, OP_MEM(13) => OP_MEM_13_port, 
                           OP_MEM(12) => OP_MEM_12_port, OP_MEM(11) => 
                           OP_MEM_11_port, OP_MEM(10) => OP_MEM_10_port, 
                           OP_MEM(9) => OP_MEM_9_port, OP_MEM(8) => 
                           OP_MEM_8_port, OP_MEM(7) => OP_MEM_7_port, OP_MEM(6)
                           => OP_MEM_6_port, OP_MEM(5) => OP_MEM_5_port, 
                           OP_MEM(4) => OP_MEM_4_port, OP_MEM(3) => 
                           OP_MEM_3_port, OP_MEM(2) => OP_MEM_2_port, OP_MEM(1)
                           => OP_MEM_1_port, OP_MEM(0) => OP_MEM_0_port, 
                           OP_WB(31) => OP_WB_31_port, OP_WB(30) => 
                           OP_WB_30_port, OP_WB(29) => OP_WB_29_port, OP_WB(28)
                           => OP_WB_28_port, OP_WB(27) => OP_WB_27_port, 
                           OP_WB(26) => OP_WB_26_port, OP_WB(25) => 
                           OP_WB_25_port, OP_WB(24) => OP_WB_24_port, OP_WB(23)
                           => OP_WB_23_port, OP_WB(22) => OP_WB_22_port, 
                           OP_WB(21) => OP_WB_21_port, OP_WB(20) => 
                           OP_WB_20_port, OP_WB(19) => OP_WB_19_port, OP_WB(18)
                           => OP_WB_18_port, OP_WB(17) => OP_WB_17_port, 
                           OP_WB(16) => OP_WB_16_port, OP_WB(15) => 
                           OP_WB_15_port, OP_WB(14) => OP_WB_14_port, OP_WB(13)
                           => OP_WB_13_port, OP_WB(12) => OP_WB_12_port, 
                           OP_WB(11) => OP_WB_11_port, OP_WB(10) => 
                           OP_WB_10_port, OP_WB(9) => OP_WB_9_port, OP_WB(8) =>
                           OP_WB_8_port, OP_WB(7) => OP_WB_7_port, OP_WB(6) => 
                           OP_WB_6_port, OP_WB(5) => OP_WB_5_port, OP_WB(4) => 
                           OP_WB_4_port, OP_WB(3) => OP_WB_3_port, OP_WB(2) => 
                           OP_WB_2_port, OP_WB(1) => OP_WB_1_port, OP_WB(0) => 
                           OP_WB_0_port, PC_SEL(1) => PC_SEL_EX_1_port, 
                           PC_SEL(0) => PC_SEL_EX_0_port, ZERO_FLAG => 
                           ZERO_FLAG_EX, NPC_ABS(31) => NPC_ABS_EX_31_port, 
                           NPC_ABS(30) => NPC_ABS_EX_30_port, NPC_ABS(29) => 
                           NPC_ABS_EX_29_port, NPC_ABS(28) => 
                           NPC_ABS_EX_28_port, NPC_ABS(27) => 
                           NPC_ABS_EX_27_port, NPC_ABS(26) => 
                           NPC_ABS_EX_26_port, NPC_ABS(25) => 
                           NPC_ABS_EX_25_port, NPC_ABS(24) => 
                           NPC_ABS_EX_24_port, NPC_ABS(23) => 
                           NPC_ABS_EX_23_port, NPC_ABS(22) => 
                           NPC_ABS_EX_22_port, NPC_ABS(21) => 
                           NPC_ABS_EX_21_port, NPC_ABS(20) => 
                           NPC_ABS_EX_20_port, NPC_ABS(19) => 
                           NPC_ABS_EX_19_port, NPC_ABS(18) => 
                           NPC_ABS_EX_18_port, NPC_ABS(17) => 
                           NPC_ABS_EX_17_port, NPC_ABS(16) => 
                           NPC_ABS_EX_16_port, NPC_ABS(15) => 
                           NPC_ABS_EX_15_port, NPC_ABS(14) => 
                           NPC_ABS_EX_14_port, NPC_ABS(13) => 
                           NPC_ABS_EX_13_port, NPC_ABS(12) => 
                           NPC_ABS_EX_12_port, NPC_ABS(11) => 
                           NPC_ABS_EX_11_port, NPC_ABS(10) => 
                           NPC_ABS_EX_10_port, NPC_ABS(9) => NPC_ABS_EX_9_port,
                           NPC_ABS(8) => NPC_ABS_EX_8_port, NPC_ABS(7) => 
                           NPC_ABS_EX_7_port, NPC_ABS(6) => NPC_ABS_EX_6_port, 
                           NPC_ABS(5) => NPC_ABS_EX_5_port, NPC_ABS(4) => 
                           NPC_ABS_EX_4_port, NPC_ABS(3) => NPC_ABS_EX_3_port, 
                           NPC_ABS(2) => NPC_ABS_EX_2_port, NPC_ABS(1) => 
                           NPC_ABS_EX_1_port, NPC_ABS(0) => NPC_ABS_EX_0_port, 
                           NPC_REL(31) => NPC_REL_EX_31_port, NPC_REL(30) => 
                           NPC_REL_EX_30_port, NPC_REL(29) => 
                           NPC_REL_EX_29_port, NPC_REL(28) => 
                           NPC_REL_EX_28_port, NPC_REL(27) => 
                           NPC_REL_EX_27_port, NPC_REL(26) => 
                           NPC_REL_EX_26_port, NPC_REL(25) => 
                           NPC_REL_EX_25_port, NPC_REL(24) => 
                           NPC_REL_EX_24_port, NPC_REL(23) => 
                           NPC_REL_EX_23_port, NPC_REL(22) => 
                           NPC_REL_EX_22_port, NPC_REL(21) => 
                           NPC_REL_EX_21_port, NPC_REL(20) => 
                           NPC_REL_EX_20_port, NPC_REL(19) => 
                           NPC_REL_EX_19_port, NPC_REL(18) => 
                           NPC_REL_EX_18_port, NPC_REL(17) => 
                           NPC_REL_EX_17_port, NPC_REL(16) => 
                           NPC_REL_EX_16_port, NPC_REL(15) => 
                           NPC_REL_EX_15_port, NPC_REL(14) => 
                           NPC_REL_EX_14_port, NPC_REL(13) => 
                           NPC_REL_EX_13_port, NPC_REL(12) => 
                           NPC_REL_EX_12_port, NPC_REL(11) => 
                           NPC_REL_EX_11_port, NPC_REL(10) => 
                           NPC_REL_EX_10_port, NPC_REL(9) => NPC_REL_EX_9_port,
                           NPC_REL(8) => NPC_REL_EX_8_port, NPC_REL(7) => 
                           NPC_REL_EX_7_port, NPC_REL(6) => NPC_REL_EX_6_port, 
                           NPC_REL(5) => NPC_REL_EX_5_port, NPC_REL(4) => 
                           NPC_REL_EX_4_port, NPC_REL(3) => NPC_REL_EX_3_port, 
                           NPC_REL(2) => NPC_REL_EX_2_port, NPC_REL(1) => 
                           NPC_REL_EX_1_port, NPC_REL(0) => NPC_REL_EX_0_port, 
                           ALU_RES(31) => ALU_RES_EX_31_port, ALU_RES(30) => 
                           ALU_RES_EX_30_port, ALU_RES(29) => 
                           ALU_RES_EX_29_port, ALU_RES(28) => 
                           ALU_RES_EX_28_port, ALU_RES(27) => 
                           ALU_RES_EX_27_port, ALU_RES(26) => 
                           ALU_RES_EX_26_port, ALU_RES(25) => 
                           ALU_RES_EX_25_port, ALU_RES(24) => 
                           ALU_RES_EX_24_port, ALU_RES(23) => 
                           ALU_RES_EX_23_port, ALU_RES(22) => 
                           ALU_RES_EX_22_port, ALU_RES(21) => 
                           ALU_RES_EX_21_port, ALU_RES(20) => 
                           ALU_RES_EX_20_port, ALU_RES(19) => 
                           ALU_RES_EX_19_port, ALU_RES(18) => 
                           ALU_RES_EX_18_port, ALU_RES(17) => 
                           ALU_RES_EX_17_port, ALU_RES(16) => 
                           ALU_RES_EX_16_port, ALU_RES(15) => 
                           ALU_RES_EX_15_port, ALU_RES(14) => 
                           ALU_RES_EX_14_port, ALU_RES(13) => 
                           ALU_RES_EX_13_port, ALU_RES(12) => 
                           ALU_RES_EX_12_port, ALU_RES(11) => 
                           ALU_RES_EX_11_port, ALU_RES(10) => 
                           ALU_RES_EX_10_port, ALU_RES(9) => ALU_RES_EX_9_port,
                           ALU_RES(8) => ALU_RES_EX_8_port, ALU_RES(7) => 
                           ALU_RES_EX_7_port, ALU_RES(6) => ALU_RES_EX_6_port, 
                           ALU_RES(5) => ALU_RES_EX_5_port, ALU_RES(4) => 
                           ALU_RES_EX_4_port, ALU_RES(3) => ALU_RES_EX_3_port, 
                           ALU_RES(2) => ALU_RES_EX_2_port, ALU_RES(1) => 
                           ALU_RES_EX_1_port, ALU_RES(0) => ALU_RES_EX_0_port, 
                           B_OUT(31) => B_EX_OUT_31_port, B_OUT(30) => 
                           B_EX_OUT_30_port, B_OUT(29) => B_EX_OUT_29_port, 
                           B_OUT(28) => B_EX_OUT_28_port, B_OUT(27) => 
                           B_EX_OUT_27_port, B_OUT(26) => B_EX_OUT_26_port, 
                           B_OUT(25) => B_EX_OUT_25_port, B_OUT(24) => 
                           B_EX_OUT_24_port, B_OUT(23) => B_EX_OUT_23_port, 
                           B_OUT(22) => B_EX_OUT_22_port, B_OUT(21) => 
                           B_EX_OUT_21_port, B_OUT(20) => B_EX_OUT_20_port, 
                           B_OUT(19) => B_EX_OUT_19_port, B_OUT(18) => 
                           B_EX_OUT_18_port, B_OUT(17) => B_EX_OUT_17_port, 
                           B_OUT(16) => B_EX_OUT_16_port, B_OUT(15) => 
                           B_EX_OUT_15_port, B_OUT(14) => B_EX_OUT_14_port, 
                           B_OUT(13) => B_EX_OUT_13_port, B_OUT(12) => 
                           B_EX_OUT_12_port, B_OUT(11) => B_EX_OUT_11_port, 
                           B_OUT(10) => B_EX_OUT_10_port, B_OUT(9) => 
                           B_EX_OUT_9_port, B_OUT(8) => B_EX_OUT_8_port, 
                           B_OUT(7) => B_EX_OUT_7_port, B_OUT(6) => 
                           B_EX_OUT_6_port, B_OUT(5) => B_EX_OUT_5_port, 
                           B_OUT(4) => B_EX_OUT_4_port, B_OUT(3) => 
                           B_EX_OUT_3_port, B_OUT(2) => B_EX_OUT_2_port, 
                           B_OUT(1) => B_EX_OUT_1_port, B_OUT(0) => 
                           B_EX_OUT_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_EX_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_EX_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_EX_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_EX_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_EX_OUT_0_port);
   DRAM_R_ff : ff_0 port map( D => DRAM_R_IN, CLK => CLK, EN => X_Logic1_port, 
                           RST => RST, Q => DRAM_R_MEM);
   MemoryStage : Memory port map( CLK => CLK, RST => RST, MEM_EN_IN => 
                           MEM_EN_IN, DRAM_R_IN => DRAM_R_MEM, DRAM_W_IN => 
                           DRAM_W_IN, DRAM_EN_IN => DRAM_EN_IN, PC_SEL(1) => 
                           PC_SEL_EX_1_port, PC_SEL(0) => PC_SEL_EX_0_port, 
                           NPC_IN(31) => NPC_FETCH_OUT_31_port, NPC_IN(30) => 
                           NPC_FETCH_OUT_30_port, NPC_IN(29) => 
                           NPC_FETCH_OUT_29_port, NPC_IN(28) => 
                           NPC_FETCH_OUT_28_port, NPC_IN(27) => 
                           NPC_FETCH_OUT_27_port, NPC_IN(26) => 
                           NPC_FETCH_OUT_26_port, NPC_IN(25) => 
                           NPC_FETCH_OUT_25_port, NPC_IN(24) => 
                           NPC_FETCH_OUT_24_port, NPC_IN(23) => 
                           NPC_FETCH_OUT_23_port, NPC_IN(22) => 
                           NPC_FETCH_OUT_22_port, NPC_IN(21) => 
                           NPC_FETCH_OUT_21_port, NPC_IN(20) => 
                           NPC_FETCH_OUT_20_port, NPC_IN(19) => 
                           NPC_FETCH_OUT_19_port, NPC_IN(18) => 
                           NPC_FETCH_OUT_18_port, NPC_IN(17) => 
                           NPC_FETCH_OUT_17_port, NPC_IN(16) => 
                           NPC_FETCH_OUT_16_port, NPC_IN(15) => 
                           NPC_FETCH_OUT_15_port, NPC_IN(14) => 
                           NPC_FETCH_OUT_14_port, NPC_IN(13) => 
                           NPC_FETCH_OUT_13_port, NPC_IN(12) => 
                           NPC_FETCH_OUT_12_port, NPC_IN(11) => 
                           NPC_FETCH_OUT_11_port, NPC_IN(10) => 
                           NPC_FETCH_OUT_10_port, NPC_IN(9) => 
                           NPC_FETCH_OUT_9_port, NPC_IN(8) => 
                           NPC_FETCH_OUT_8_port, NPC_IN(7) => 
                           NPC_FETCH_OUT_7_port, NPC_IN(6) => 
                           NPC_FETCH_OUT_6_port, NPC_IN(5) => 
                           NPC_FETCH_OUT_5_port, NPC_IN(4) => 
                           NPC_FETCH_OUT_4_port, NPC_IN(3) => 
                           NPC_FETCH_OUT_3_port, NPC_IN(2) => 
                           NPC_FETCH_OUT_2_port, NPC_IN(1) => 
                           NPC_FETCH_OUT_1_port, NPC_IN(0) => 
                           NPC_FETCH_OUT_0_port, NPC_ABS(31) => 
                           NPC_ABS_EX_31_port, NPC_ABS(30) => 
                           NPC_ABS_EX_30_port, NPC_ABS(29) => 
                           NPC_ABS_EX_29_port, NPC_ABS(28) => 
                           NPC_ABS_EX_28_port, NPC_ABS(27) => 
                           NPC_ABS_EX_27_port, NPC_ABS(26) => 
                           NPC_ABS_EX_26_port, NPC_ABS(25) => 
                           NPC_ABS_EX_25_port, NPC_ABS(24) => 
                           NPC_ABS_EX_24_port, NPC_ABS(23) => 
                           NPC_ABS_EX_23_port, NPC_ABS(22) => 
                           NPC_ABS_EX_22_port, NPC_ABS(21) => 
                           NPC_ABS_EX_21_port, NPC_ABS(20) => 
                           NPC_ABS_EX_20_port, NPC_ABS(19) => 
                           NPC_ABS_EX_19_port, NPC_ABS(18) => 
                           NPC_ABS_EX_18_port, NPC_ABS(17) => 
                           NPC_ABS_EX_17_port, NPC_ABS(16) => 
                           NPC_ABS_EX_16_port, NPC_ABS(15) => 
                           NPC_ABS_EX_15_port, NPC_ABS(14) => 
                           NPC_ABS_EX_14_port, NPC_ABS(13) => 
                           NPC_ABS_EX_13_port, NPC_ABS(12) => 
                           NPC_ABS_EX_12_port, NPC_ABS(11) => 
                           NPC_ABS_EX_11_port, NPC_ABS(10) => 
                           NPC_ABS_EX_10_port, NPC_ABS(9) => NPC_ABS_EX_9_port,
                           NPC_ABS(8) => NPC_ABS_EX_8_port, NPC_ABS(7) => 
                           NPC_ABS_EX_7_port, NPC_ABS(6) => NPC_ABS_EX_6_port, 
                           NPC_ABS(5) => NPC_ABS_EX_5_port, NPC_ABS(4) => 
                           NPC_ABS_EX_4_port, NPC_ABS(3) => NPC_ABS_EX_3_port, 
                           NPC_ABS(2) => NPC_ABS_EX_2_port, NPC_ABS(1) => 
                           NPC_ABS_EX_1_port, NPC_ABS(0) => NPC_ABS_EX_0_port, 
                           NPC_REL(31) => NPC_REL_EX_31_port, NPC_REL(30) => 
                           NPC_REL_EX_30_port, NPC_REL(29) => 
                           NPC_REL_EX_29_port, NPC_REL(28) => 
                           NPC_REL_EX_28_port, NPC_REL(27) => 
                           NPC_REL_EX_27_port, NPC_REL(26) => 
                           NPC_REL_EX_26_port, NPC_REL(25) => 
                           NPC_REL_EX_25_port, NPC_REL(24) => 
                           NPC_REL_EX_24_port, NPC_REL(23) => 
                           NPC_REL_EX_23_port, NPC_REL(22) => 
                           NPC_REL_EX_22_port, NPC_REL(21) => 
                           NPC_REL_EX_21_port, NPC_REL(20) => 
                           NPC_REL_EX_20_port, NPC_REL(19) => 
                           NPC_REL_EX_19_port, NPC_REL(18) => 
                           NPC_REL_EX_18_port, NPC_REL(17) => 
                           NPC_REL_EX_17_port, NPC_REL(16) => 
                           NPC_REL_EX_16_port, NPC_REL(15) => 
                           NPC_REL_EX_15_port, NPC_REL(14) => 
                           NPC_REL_EX_14_port, NPC_REL(13) => 
                           NPC_REL_EX_13_port, NPC_REL(12) => 
                           NPC_REL_EX_12_port, NPC_REL(11) => 
                           NPC_REL_EX_11_port, NPC_REL(10) => 
                           NPC_REL_EX_10_port, NPC_REL(9) => NPC_REL_EX_9_port,
                           NPC_REL(8) => NPC_REL_EX_8_port, NPC_REL(7) => 
                           NPC_REL_EX_7_port, NPC_REL(6) => NPC_REL_EX_6_port, 
                           NPC_REL(5) => NPC_REL_EX_5_port, NPC_REL(4) => 
                           NPC_REL_EX_4_port, NPC_REL(3) => NPC_REL_EX_3_port, 
                           NPC_REL(2) => NPC_REL_EX_2_port, NPC_REL(1) => 
                           NPC_REL_EX_1_port, NPC_REL(0) => NPC_REL_EX_0_port, 
                           ALU_RES_IN(31) => ALU_RES_EX_31_port, ALU_RES_IN(30)
                           => ALU_RES_EX_30_port, ALU_RES_IN(29) => 
                           ALU_RES_EX_29_port, ALU_RES_IN(28) => 
                           ALU_RES_EX_28_port, ALU_RES_IN(27) => 
                           ALU_RES_EX_27_port, ALU_RES_IN(26) => 
                           ALU_RES_EX_26_port, ALU_RES_IN(25) => 
                           ALU_RES_EX_25_port, ALU_RES_IN(24) => 
                           ALU_RES_EX_24_port, ALU_RES_IN(23) => 
                           ALU_RES_EX_23_port, ALU_RES_IN(22) => 
                           ALU_RES_EX_22_port, ALU_RES_IN(21) => 
                           ALU_RES_EX_21_port, ALU_RES_IN(20) => 
                           ALU_RES_EX_20_port, ALU_RES_IN(19) => 
                           ALU_RES_EX_19_port, ALU_RES_IN(18) => 
                           ALU_RES_EX_18_port, ALU_RES_IN(17) => 
                           ALU_RES_EX_17_port, ALU_RES_IN(16) => 
                           ALU_RES_EX_16_port, ALU_RES_IN(15) => 
                           ALU_RES_EX_15_port, ALU_RES_IN(14) => 
                           ALU_RES_EX_14_port, ALU_RES_IN(13) => 
                           ALU_RES_EX_13_port, ALU_RES_IN(12) => 
                           ALU_RES_EX_12_port, ALU_RES_IN(11) => 
                           ALU_RES_EX_11_port, ALU_RES_IN(10) => 
                           ALU_RES_EX_10_port, ALU_RES_IN(9) => 
                           ALU_RES_EX_9_port, ALU_RES_IN(8) => 
                           ALU_RES_EX_8_port, ALU_RES_IN(7) => 
                           ALU_RES_EX_7_port, ALU_RES_IN(6) => 
                           ALU_RES_EX_6_port, ALU_RES_IN(5) => 
                           ALU_RES_EX_5_port, ALU_RES_IN(4) => 
                           ALU_RES_EX_4_port, ALU_RES_IN(3) => 
                           ALU_RES_EX_3_port, ALU_RES_IN(2) => 
                           ALU_RES_EX_2_port, ALU_RES_IN(1) => 
                           ALU_RES_EX_1_port, ALU_RES_IN(0) => 
                           ALU_RES_EX_0_port, B_IN(31) => B_EX_OUT_31_port, 
                           B_IN(30) => B_EX_OUT_30_port, B_IN(29) => 
                           B_EX_OUT_29_port, B_IN(28) => B_EX_OUT_28_port, 
                           B_IN(27) => B_EX_OUT_27_port, B_IN(26) => 
                           B_EX_OUT_26_port, B_IN(25) => B_EX_OUT_25_port, 
                           B_IN(24) => B_EX_OUT_24_port, B_IN(23) => 
                           B_EX_OUT_23_port, B_IN(22) => B_EX_OUT_22_port, 
                           B_IN(21) => B_EX_OUT_21_port, B_IN(20) => 
                           B_EX_OUT_20_port, B_IN(19) => B_EX_OUT_19_port, 
                           B_IN(18) => B_EX_OUT_18_port, B_IN(17) => 
                           B_EX_OUT_17_port, B_IN(16) => B_EX_OUT_16_port, 
                           B_IN(15) => B_EX_OUT_15_port, B_IN(14) => 
                           B_EX_OUT_14_port, B_IN(13) => B_EX_OUT_13_port, 
                           B_IN(12) => B_EX_OUT_12_port, B_IN(11) => 
                           B_EX_OUT_11_port, B_IN(10) => B_EX_OUT_10_port, 
                           B_IN(9) => B_EX_OUT_9_port, B_IN(8) => 
                           B_EX_OUT_8_port, B_IN(7) => B_EX_OUT_7_port, B_IN(6)
                           => B_EX_OUT_6_port, B_IN(5) => B_EX_OUT_5_port, 
                           B_IN(4) => B_EX_OUT_4_port, B_IN(3) => 
                           B_EX_OUT_3_port, B_IN(2) => B_EX_OUT_2_port, B_IN(1)
                           => B_EX_OUT_1_port, B_IN(0) => B_EX_OUT_0_port, 
                           ADD_WR_IN(4) => ADD_WR_EX_OUT_4_port, ADD_WR_IN(3) 
                           => ADD_WR_EX_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_EX_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_EX_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_EX_OUT_0_port, DRAM_DATA_IN(31) => 
                           DATA_IN(31), DRAM_DATA_IN(30) => DATA_IN(30), 
                           DRAM_DATA_IN(29) => DATA_IN(29), DRAM_DATA_IN(28) =>
                           DATA_IN(28), DRAM_DATA_IN(27) => DATA_IN(27), 
                           DRAM_DATA_IN(26) => DATA_IN(26), DRAM_DATA_IN(25) =>
                           DATA_IN(25), DRAM_DATA_IN(24) => DATA_IN(24), 
                           DRAM_DATA_IN(23) => DATA_IN(23), DRAM_DATA_IN(22) =>
                           DATA_IN(22), DRAM_DATA_IN(21) => DATA_IN(21), 
                           DRAM_DATA_IN(20) => DATA_IN(20), DRAM_DATA_IN(19) =>
                           DATA_IN(19), DRAM_DATA_IN(18) => DATA_IN(18), 
                           DRAM_DATA_IN(17) => DATA_IN(17), DRAM_DATA_IN(16) =>
                           DATA_IN(16), DRAM_DATA_IN(15) => DATA_IN(15), 
                           DRAM_DATA_IN(14) => DATA_IN(14), DRAM_DATA_IN(13) =>
                           DATA_IN(13), DRAM_DATA_IN(12) => DATA_IN(12), 
                           DRAM_DATA_IN(11) => DATA_IN(11), DRAM_DATA_IN(10) =>
                           DATA_IN(10), DRAM_DATA_IN(9) => DATA_IN(9), 
                           DRAM_DATA_IN(8) => DATA_IN(8), DRAM_DATA_IN(7) => 
                           DATA_IN(7), DRAM_DATA_IN(6) => DATA_IN(6), 
                           DRAM_DATA_IN(5) => DATA_IN(5), DRAM_DATA_IN(4) => 
                           DATA_IN(4), DRAM_DATA_IN(3) => DATA_IN(3), 
                           DRAM_DATA_IN(2) => DATA_IN(2), DRAM_DATA_IN(1) => 
                           DATA_IN(1), DRAM_DATA_IN(0) => DATA_IN(0), 
                           PC_OUT(31) => PC_MEM_OUT_31_port, PC_OUT(30) => 
                           PC_MEM_OUT_30_port, PC_OUT(29) => PC_MEM_OUT_29_port
                           , PC_OUT(28) => PC_MEM_OUT_28_port, PC_OUT(27) => 
                           PC_MEM_OUT_27_port, PC_OUT(26) => PC_MEM_OUT_26_port
                           , PC_OUT(25) => PC_MEM_OUT_25_port, PC_OUT(24) => 
                           PC_MEM_OUT_24_port, PC_OUT(23) => PC_MEM_OUT_23_port
                           , PC_OUT(22) => PC_MEM_OUT_22_port, PC_OUT(21) => 
                           PC_MEM_OUT_21_port, PC_OUT(20) => PC_MEM_OUT_20_port
                           , PC_OUT(19) => PC_MEM_OUT_19_port, PC_OUT(18) => 
                           PC_MEM_OUT_18_port, PC_OUT(17) => PC_MEM_OUT_17_port
                           , PC_OUT(16) => PC_MEM_OUT_16_port, PC_OUT(15) => 
                           PC_MEM_OUT_15_port, PC_OUT(14) => PC_MEM_OUT_14_port
                           , PC_OUT(13) => PC_MEM_OUT_13_port, PC_OUT(12) => 
                           PC_MEM_OUT_12_port, PC_OUT(11) => PC_MEM_OUT_11_port
                           , PC_OUT(10) => PC_MEM_OUT_10_port, PC_OUT(9) => 
                           PC_MEM_OUT_9_port, PC_OUT(8) => PC_MEM_OUT_8_port, 
                           PC_OUT(7) => PC_MEM_OUT_7_port, PC_OUT(6) => 
                           PC_MEM_OUT_6_port, PC_OUT(5) => PC_MEM_OUT_5_port, 
                           PC_OUT(4) => PC_MEM_OUT_4_port, PC_OUT(3) => 
                           PC_MEM_OUT_3_port, PC_OUT(2) => PC_MEM_OUT_2_port, 
                           PC_OUT(1) => PC_MEM_OUT_1_port, PC_OUT(0) => 
                           PC_MEM_OUT_0_port, DRAM_EN_OUT => DRAM_EN_OUT, 
                           DRAM_R_OUT => DRAM_R_OUT, DRAM_W_OUT => DRAM_W_OUT, 
                           DRAM_ADDR_OUT(31) => DRAM_ADDR_OUT(31), 
                           DRAM_ADDR_OUT(30) => DRAM_ADDR_OUT(30), 
                           DRAM_ADDR_OUT(29) => DRAM_ADDR_OUT(29), 
                           DRAM_ADDR_OUT(28) => DRAM_ADDR_OUT(28), 
                           DRAM_ADDR_OUT(27) => DRAM_ADDR_OUT(27), 
                           DRAM_ADDR_OUT(26) => DRAM_ADDR_OUT(26), 
                           DRAM_ADDR_OUT(25) => DRAM_ADDR_OUT(25), 
                           DRAM_ADDR_OUT(24) => DRAM_ADDR_OUT(24), 
                           DRAM_ADDR_OUT(23) => DRAM_ADDR_OUT(23), 
                           DRAM_ADDR_OUT(22) => DRAM_ADDR_OUT(22), 
                           DRAM_ADDR_OUT(21) => DRAM_ADDR_OUT(21), 
                           DRAM_ADDR_OUT(20) => DRAM_ADDR_OUT(20), 
                           DRAM_ADDR_OUT(19) => DRAM_ADDR_OUT(19), 
                           DRAM_ADDR_OUT(18) => DRAM_ADDR_OUT(18), 
                           DRAM_ADDR_OUT(17) => DRAM_ADDR_OUT(17), 
                           DRAM_ADDR_OUT(16) => DRAM_ADDR_OUT(16), 
                           DRAM_ADDR_OUT(15) => DRAM_ADDR_OUT(15), 
                           DRAM_ADDR_OUT(14) => DRAM_ADDR_OUT(14), 
                           DRAM_ADDR_OUT(13) => DRAM_ADDR_OUT(13), 
                           DRAM_ADDR_OUT(12) => DRAM_ADDR_OUT(12), 
                           DRAM_ADDR_OUT(11) => DRAM_ADDR_OUT(11), 
                           DRAM_ADDR_OUT(10) => DRAM_ADDR_OUT(10), 
                           DRAM_ADDR_OUT(9) => DRAM_ADDR_OUT(9), 
                           DRAM_ADDR_OUT(8) => DRAM_ADDR_OUT(8), 
                           DRAM_ADDR_OUT(7) => DRAM_ADDR_OUT(7), 
                           DRAM_ADDR_OUT(6) => DRAM_ADDR_OUT(6), 
                           DRAM_ADDR_OUT(5) => DRAM_ADDR_OUT(5), 
                           DRAM_ADDR_OUT(4) => DRAM_ADDR_OUT(4), 
                           DRAM_ADDR_OUT(3) => DRAM_ADDR_OUT(3), 
                           DRAM_ADDR_OUT(2) => DRAM_ADDR_OUT(2), 
                           DRAM_ADDR_OUT(1) => DRAM_ADDR_OUT(1), 
                           DRAM_ADDR_OUT(0) => DRAM_ADDR_OUT(0), 
                           DRAM_DATA_OUT(31) => DATA_OUT(31), DRAM_DATA_OUT(30)
                           => DATA_OUT(30), DRAM_DATA_OUT(29) => DATA_OUT(29), 
                           DRAM_DATA_OUT(28) => DATA_OUT(28), DRAM_DATA_OUT(27)
                           => DATA_OUT(27), DRAM_DATA_OUT(26) => DATA_OUT(26), 
                           DRAM_DATA_OUT(25) => DATA_OUT(25), DRAM_DATA_OUT(24)
                           => DATA_OUT(24), DRAM_DATA_OUT(23) => DATA_OUT(23), 
                           DRAM_DATA_OUT(22) => DATA_OUT(22), DRAM_DATA_OUT(21)
                           => DATA_OUT(21), DRAM_DATA_OUT(20) => DATA_OUT(20), 
                           DRAM_DATA_OUT(19) => DATA_OUT(19), DRAM_DATA_OUT(18)
                           => DATA_OUT(18), DRAM_DATA_OUT(17) => DATA_OUT(17), 
                           DRAM_DATA_OUT(16) => DATA_OUT(16), DRAM_DATA_OUT(15)
                           => DATA_OUT(15), DRAM_DATA_OUT(14) => DATA_OUT(14), 
                           DRAM_DATA_OUT(13) => DATA_OUT(13), DRAM_DATA_OUT(12)
                           => DATA_OUT(12), DRAM_DATA_OUT(11) => DATA_OUT(11), 
                           DRAM_DATA_OUT(10) => DATA_OUT(10), DRAM_DATA_OUT(9) 
                           => DATA_OUT(9), DRAM_DATA_OUT(8) => DATA_OUT(8), 
                           DRAM_DATA_OUT(7) => DATA_OUT(7), DRAM_DATA_OUT(6) =>
                           DATA_OUT(6), DRAM_DATA_OUT(5) => DATA_OUT(5), 
                           DRAM_DATA_OUT(4) => DATA_OUT(4), DRAM_DATA_OUT(3) =>
                           DATA_OUT(3), DRAM_DATA_OUT(2) => DATA_OUT(2), 
                           DRAM_DATA_OUT(1) => DATA_OUT(1), DRAM_DATA_OUT(0) =>
                           DATA_OUT(0), DATA_OUT(31) => DATA_MEM_OUT_31_port, 
                           DATA_OUT(30) => DATA_MEM_OUT_30_port, DATA_OUT(29) 
                           => DATA_MEM_OUT_29_port, DATA_OUT(28) => 
                           DATA_MEM_OUT_28_port, DATA_OUT(27) => 
                           DATA_MEM_OUT_27_port, DATA_OUT(26) => 
                           DATA_MEM_OUT_26_port, DATA_OUT(25) => 
                           DATA_MEM_OUT_25_port, DATA_OUT(24) => 
                           DATA_MEM_OUT_24_port, DATA_OUT(23) => 
                           DATA_MEM_OUT_23_port, DATA_OUT(22) => 
                           DATA_MEM_OUT_22_port, DATA_OUT(21) => 
                           DATA_MEM_OUT_21_port, DATA_OUT(20) => 
                           DATA_MEM_OUT_20_port, DATA_OUT(19) => 
                           DATA_MEM_OUT_19_port, DATA_OUT(18) => 
                           DATA_MEM_OUT_18_port, DATA_OUT(17) => 
                           DATA_MEM_OUT_17_port, DATA_OUT(16) => 
                           DATA_MEM_OUT_16_port, DATA_OUT(15) => 
                           DATA_MEM_OUT_15_port, DATA_OUT(14) => 
                           DATA_MEM_OUT_14_port, DATA_OUT(13) => 
                           DATA_MEM_OUT_13_port, DATA_OUT(12) => 
                           DATA_MEM_OUT_12_port, DATA_OUT(11) => 
                           DATA_MEM_OUT_11_port, DATA_OUT(10) => 
                           DATA_MEM_OUT_10_port, DATA_OUT(9) => 
                           DATA_MEM_OUT_9_port, DATA_OUT(8) => 
                           DATA_MEM_OUT_8_port, DATA_OUT(7) => 
                           DATA_MEM_OUT_7_port, DATA_OUT(6) => 
                           DATA_MEM_OUT_6_port, DATA_OUT(5) => 
                           DATA_MEM_OUT_5_port, DATA_OUT(4) => 
                           DATA_MEM_OUT_4_port, DATA_OUT(3) => 
                           DATA_MEM_OUT_3_port, DATA_OUT(2) => 
                           DATA_MEM_OUT_2_port, DATA_OUT(1) => 
                           DATA_MEM_OUT_1_port, DATA_OUT(0) => 
                           DATA_MEM_OUT_0_port, ALU_RES_OUT(31) => 
                           ALU_RES_MEM_31_port, ALU_RES_OUT(30) => 
                           ALU_RES_MEM_30_port, ALU_RES_OUT(29) => 
                           ALU_RES_MEM_29_port, ALU_RES_OUT(28) => 
                           ALU_RES_MEM_28_port, ALU_RES_OUT(27) => 
                           ALU_RES_MEM_27_port, ALU_RES_OUT(26) => 
                           ALU_RES_MEM_26_port, ALU_RES_OUT(25) => 
                           ALU_RES_MEM_25_port, ALU_RES_OUT(24) => 
                           ALU_RES_MEM_24_port, ALU_RES_OUT(23) => 
                           ALU_RES_MEM_23_port, ALU_RES_OUT(22) => 
                           ALU_RES_MEM_22_port, ALU_RES_OUT(21) => 
                           ALU_RES_MEM_21_port, ALU_RES_OUT(20) => 
                           ALU_RES_MEM_20_port, ALU_RES_OUT(19) => 
                           ALU_RES_MEM_19_port, ALU_RES_OUT(18) => 
                           ALU_RES_MEM_18_port, ALU_RES_OUT(17) => 
                           ALU_RES_MEM_17_port, ALU_RES_OUT(16) => 
                           ALU_RES_MEM_16_port, ALU_RES_OUT(15) => 
                           ALU_RES_MEM_15_port, ALU_RES_OUT(14) => 
                           ALU_RES_MEM_14_port, ALU_RES_OUT(13) => 
                           ALU_RES_MEM_13_port, ALU_RES_OUT(12) => 
                           ALU_RES_MEM_12_port, ALU_RES_OUT(11) => 
                           ALU_RES_MEM_11_port, ALU_RES_OUT(10) => 
                           ALU_RES_MEM_10_port, ALU_RES_OUT(9) => 
                           ALU_RES_MEM_9_port, ALU_RES_OUT(8) => 
                           ALU_RES_MEM_8_port, ALU_RES_OUT(7) => 
                           ALU_RES_MEM_7_port, ALU_RES_OUT(6) => 
                           ALU_RES_MEM_6_port, ALU_RES_OUT(5) => 
                           ALU_RES_MEM_5_port, ALU_RES_OUT(4) => 
                           ALU_RES_MEM_4_port, ALU_RES_OUT(3) => 
                           ALU_RES_MEM_3_port, ALU_RES_OUT(2) => 
                           ALU_RES_MEM_2_port, ALU_RES_OUT(1) => 
                           ALU_RES_MEM_1_port, ALU_RES_OUT(0) => 
                           ALU_RES_MEM_0_port, OP_MEM(31) => OP_MEM_31_port, 
                           OP_MEM(30) => OP_MEM_30_port, OP_MEM(29) => 
                           OP_MEM_29_port, OP_MEM(28) => OP_MEM_28_port, 
                           OP_MEM(27) => OP_MEM_27_port, OP_MEM(26) => 
                           OP_MEM_26_port, OP_MEM(25) => OP_MEM_25_port, 
                           OP_MEM(24) => OP_MEM_24_port, OP_MEM(23) => 
                           OP_MEM_23_port, OP_MEM(22) => OP_MEM_22_port, 
                           OP_MEM(21) => OP_MEM_21_port, OP_MEM(20) => 
                           OP_MEM_20_port, OP_MEM(19) => OP_MEM_19_port, 
                           OP_MEM(18) => OP_MEM_18_port, OP_MEM(17) => 
                           OP_MEM_17_port, OP_MEM(16) => OP_MEM_16_port, 
                           OP_MEM(15) => OP_MEM_15_port, OP_MEM(14) => 
                           OP_MEM_14_port, OP_MEM(13) => OP_MEM_13_port, 
                           OP_MEM(12) => OP_MEM_12_port, OP_MEM(11) => 
                           OP_MEM_11_port, OP_MEM(10) => OP_MEM_10_port, 
                           OP_MEM(9) => OP_MEM_9_port, OP_MEM(8) => 
                           OP_MEM_8_port, OP_MEM(7) => OP_MEM_7_port, OP_MEM(6)
                           => OP_MEM_6_port, OP_MEM(5) => OP_MEM_5_port, 
                           OP_MEM(4) => OP_MEM_4_port, OP_MEM(3) => 
                           OP_MEM_3_port, OP_MEM(2) => OP_MEM_2_port, OP_MEM(1)
                           => OP_MEM_1_port, OP_MEM(0) => OP_MEM_0_port, 
                           ADD_WR_MEM(4) => ADD_WR_MEM_4_port, ADD_WR_MEM(3) =>
                           ADD_WR_MEM_3_port, ADD_WR_MEM(2) => 
                           ADD_WR_MEM_2_port, ADD_WR_MEM(1) => 
                           ADD_WR_MEM_1_port, ADD_WR_MEM(0) => 
                           ADD_WR_MEM_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_MEM_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_MEM_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_MEM_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_MEM_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_MEM_OUT_0_port);
   RF_WE_ff : ff_2 port map( D => RF_WE, CLK => CLK, EN => X_Logic1_port, RST 
                           => RST, Q => RF_WE_WB);
   WritebackStage : Writeback port map( WB_MUX_SEL => WB_MUX_SEL, DATA_IN(31) 
                           => DATA_MEM_OUT_31_port, DATA_IN(30) => 
                           DATA_MEM_OUT_30_port, DATA_IN(29) => 
                           DATA_MEM_OUT_29_port, DATA_IN(28) => 
                           DATA_MEM_OUT_28_port, DATA_IN(27) => 
                           DATA_MEM_OUT_27_port, DATA_IN(26) => 
                           DATA_MEM_OUT_26_port, DATA_IN(25) => 
                           DATA_MEM_OUT_25_port, DATA_IN(24) => 
                           DATA_MEM_OUT_24_port, DATA_IN(23) => 
                           DATA_MEM_OUT_23_port, DATA_IN(22) => 
                           DATA_MEM_OUT_22_port, DATA_IN(21) => 
                           DATA_MEM_OUT_21_port, DATA_IN(20) => 
                           DATA_MEM_OUT_20_port, DATA_IN(19) => 
                           DATA_MEM_OUT_19_port, DATA_IN(18) => 
                           DATA_MEM_OUT_18_port, DATA_IN(17) => 
                           DATA_MEM_OUT_17_port, DATA_IN(16) => 
                           DATA_MEM_OUT_16_port, DATA_IN(15) => 
                           DATA_MEM_OUT_15_port, DATA_IN(14) => 
                           DATA_MEM_OUT_14_port, DATA_IN(13) => 
                           DATA_MEM_OUT_13_port, DATA_IN(12) => 
                           DATA_MEM_OUT_12_port, DATA_IN(11) => 
                           DATA_MEM_OUT_11_port, DATA_IN(10) => 
                           DATA_MEM_OUT_10_port, DATA_IN(9) => 
                           DATA_MEM_OUT_9_port, DATA_IN(8) => 
                           DATA_MEM_OUT_8_port, DATA_IN(7) => 
                           DATA_MEM_OUT_7_port, DATA_IN(6) => 
                           DATA_MEM_OUT_6_port, DATA_IN(5) => 
                           DATA_MEM_OUT_5_port, DATA_IN(4) => 
                           DATA_MEM_OUT_4_port, DATA_IN(3) => 
                           DATA_MEM_OUT_3_port, DATA_IN(2) => 
                           DATA_MEM_OUT_2_port, DATA_IN(1) => 
                           DATA_MEM_OUT_1_port, DATA_IN(0) => 
                           DATA_MEM_OUT_0_port, ALU_RES_IN(31) => 
                           ALU_RES_MEM_31_port, ALU_RES_IN(30) => 
                           ALU_RES_MEM_30_port, ALU_RES_IN(29) => 
                           ALU_RES_MEM_29_port, ALU_RES_IN(28) => 
                           ALU_RES_MEM_28_port, ALU_RES_IN(27) => 
                           ALU_RES_MEM_27_port, ALU_RES_IN(26) => 
                           ALU_RES_MEM_26_port, ALU_RES_IN(25) => 
                           ALU_RES_MEM_25_port, ALU_RES_IN(24) => 
                           ALU_RES_MEM_24_port, ALU_RES_IN(23) => 
                           ALU_RES_MEM_23_port, ALU_RES_IN(22) => 
                           ALU_RES_MEM_22_port, ALU_RES_IN(21) => 
                           ALU_RES_MEM_21_port, ALU_RES_IN(20) => 
                           ALU_RES_MEM_20_port, ALU_RES_IN(19) => 
                           ALU_RES_MEM_19_port, ALU_RES_IN(18) => 
                           ALU_RES_MEM_18_port, ALU_RES_IN(17) => 
                           ALU_RES_MEM_17_port, ALU_RES_IN(16) => 
                           ALU_RES_MEM_16_port, ALU_RES_IN(15) => 
                           ALU_RES_MEM_15_port, ALU_RES_IN(14) => 
                           ALU_RES_MEM_14_port, ALU_RES_IN(13) => 
                           ALU_RES_MEM_13_port, ALU_RES_IN(12) => 
                           ALU_RES_MEM_12_port, ALU_RES_IN(11) => 
                           ALU_RES_MEM_11_port, ALU_RES_IN(10) => 
                           ALU_RES_MEM_10_port, ALU_RES_IN(9) => 
                           ALU_RES_MEM_9_port, ALU_RES_IN(8) => 
                           ALU_RES_MEM_8_port, ALU_RES_IN(7) => 
                           ALU_RES_MEM_7_port, ALU_RES_IN(6) => 
                           ALU_RES_MEM_6_port, ALU_RES_IN(5) => 
                           ALU_RES_MEM_5_port, ALU_RES_IN(4) => 
                           ALU_RES_MEM_4_port, ALU_RES_IN(3) => 
                           ALU_RES_MEM_3_port, ALU_RES_IN(2) => 
                           ALU_RES_MEM_2_port, ALU_RES_IN(1) => 
                           ALU_RES_MEM_1_port, ALU_RES_IN(0) => 
                           ALU_RES_MEM_0_port, ADD_WR_IN(4) => 
                           ADD_WR_MEM_OUT_4_port, ADD_WR_IN(3) => 
                           ADD_WR_MEM_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_MEM_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_MEM_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_MEM_OUT_0_port, DATA_OUT(31) => OP_WB_31_port
                           , DATA_OUT(30) => OP_WB_30_port, DATA_OUT(29) => 
                           OP_WB_29_port, DATA_OUT(28) => OP_WB_28_port, 
                           DATA_OUT(27) => OP_WB_27_port, DATA_OUT(26) => 
                           OP_WB_26_port, DATA_OUT(25) => OP_WB_25_port, 
                           DATA_OUT(24) => OP_WB_24_port, DATA_OUT(23) => 
                           OP_WB_23_port, DATA_OUT(22) => OP_WB_22_port, 
                           DATA_OUT(21) => OP_WB_21_port, DATA_OUT(20) => 
                           OP_WB_20_port, DATA_OUT(19) => OP_WB_19_port, 
                           DATA_OUT(18) => OP_WB_18_port, DATA_OUT(17) => 
                           OP_WB_17_port, DATA_OUT(16) => OP_WB_16_port, 
                           DATA_OUT(15) => OP_WB_15_port, DATA_OUT(14) => 
                           OP_WB_14_port, DATA_OUT(13) => OP_WB_13_port, 
                           DATA_OUT(12) => OP_WB_12_port, DATA_OUT(11) => 
                           OP_WB_11_port, DATA_OUT(10) => OP_WB_10_port, 
                           DATA_OUT(9) => OP_WB_9_port, DATA_OUT(8) => 
                           OP_WB_8_port, DATA_OUT(7) => OP_WB_7_port, 
                           DATA_OUT(6) => OP_WB_6_port, DATA_OUT(5) => 
                           OP_WB_5_port, DATA_OUT(4) => OP_WB_4_port, 
                           DATA_OUT(3) => OP_WB_3_port, DATA_OUT(2) => 
                           OP_WB_2_port, DATA_OUT(1) => OP_WB_1_port, 
                           DATA_OUT(0) => OP_WB_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_WB_4_port, ADD_WR_OUT(3) => ADD_WR_WB_3_port,
                           ADD_WR_OUT(2) => ADD_WR_WB_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_WB_1_port, ADD_WR_OUT(0) => ADD_WR_WB_0_port)
                           ;
   HDU : HazardDetection port map( RST => RST, ADD_RS1(4) => ADD_RS1_HDU_4_port
                           , ADD_RS1(3) => ADD_RS1_HDU_3_port, ADD_RS1(2) => 
                           ADD_RS1_HDU_2_port, ADD_RS1(1) => ADD_RS1_HDU_1_port
                           , ADD_RS1(0) => ADD_RS1_HDU_0_port, ADD_RS2(4) => 
                           ADD_RS2_HDU_4_port, ADD_RS2(3) => ADD_RS2_HDU_3_port
                           , ADD_RS2(2) => ADD_RS2_HDU_2_port, ADD_RS2(1) => 
                           ADD_RS2_HDU_1_port, ADD_RS2(0) => ADD_RS2_HDU_0_port
                           , ADD_WR(4) => ADD_WR_DECODE_OUT_4_port, ADD_WR(3) 
                           => ADD_WR_DECODE_OUT_3_port, ADD_WR(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR(0) => 
                           ADD_WR_DECODE_OUT_0_port, DRAM_R => DRAM_R_IN, 
                           INS_IN(31) => INS_OUT_31_port, INS_IN(30) => 
                           INS_OUT_30_port, INS_IN(29) => INS_OUT_29_port, 
                           INS_IN(28) => INS_OUT_28_port, INS_IN(27) => 
                           INS_OUT_27_port, INS_IN(26) => INS_OUT_26_port, 
                           INS_IN(25) => INS_OUT_25_port, INS_IN(24) => 
                           INS_OUT_24_port, INS_IN(23) => INS_OUT_23_port, 
                           INS_IN(22) => INS_OUT_22_port, INS_IN(21) => 
                           INS_OUT_21_port, INS_IN(20) => INS_OUT_20_port, 
                           INS_IN(19) => INS_OUT_19_port, INS_IN(18) => 
                           INS_OUT_18_port, INS_IN(17) => INS_OUT_17_port, 
                           INS_IN(16) => INS_OUT_16_port, INS_IN(15) => 
                           INS_OUT_15_port, INS_IN(14) => INS_OUT_14_port, 
                           INS_IN(13) => INS_OUT_13_port, INS_IN(12) => 
                           INS_OUT_12_port, INS_IN(11) => INS_OUT_11_port, 
                           INS_IN(10) => INS_OUT_10_port, INS_IN(9) => 
                           INS_OUT_9_port, INS_IN(8) => INS_OUT_8_port, 
                           INS_IN(7) => INS_OUT_7_port, INS_IN(6) => 
                           INS_OUT_6_port, INS_IN(5) => INS_OUT_5_port, 
                           INS_IN(4) => INS_OUT_4_port, INS_IN(3) => 
                           INS_OUT_3_port, INS_IN(2) => INS_OUT_2_port, 
                           INS_IN(1) => INS_OUT_1_port, INS_IN(0) => 
                           INS_OUT_0_port, PC_IN(31) => PC_FETCH_OUT_31_port, 
                           PC_IN(30) => PC_FETCH_OUT_30_port, PC_IN(29) => 
                           PC_FETCH_OUT_29_port, PC_IN(28) => 
                           PC_FETCH_OUT_28_port, PC_IN(27) => 
                           PC_FETCH_OUT_27_port, PC_IN(26) => 
                           PC_FETCH_OUT_26_port, PC_IN(25) => 
                           PC_FETCH_OUT_25_port, PC_IN(24) => 
                           PC_FETCH_OUT_24_port, PC_IN(23) => 
                           PC_FETCH_OUT_23_port, PC_IN(22) => 
                           PC_FETCH_OUT_22_port, PC_IN(21) => 
                           PC_FETCH_OUT_21_port, PC_IN(20) => 
                           PC_FETCH_OUT_20_port, PC_IN(19) => 
                           PC_FETCH_OUT_19_port, PC_IN(18) => 
                           PC_FETCH_OUT_18_port, PC_IN(17) => 
                           PC_FETCH_OUT_17_port, PC_IN(16) => 
                           PC_FETCH_OUT_16_port, PC_IN(15) => 
                           PC_FETCH_OUT_15_port, PC_IN(14) => 
                           PC_FETCH_OUT_14_port, PC_IN(13) => 
                           PC_FETCH_OUT_13_port, PC_IN(12) => 
                           PC_FETCH_OUT_12_port, PC_IN(11) => 
                           PC_FETCH_OUT_11_port, PC_IN(10) => 
                           PC_FETCH_OUT_10_port, PC_IN(9) => 
                           PC_FETCH_OUT_9_port, PC_IN(8) => PC_FETCH_OUT_8_port
                           , PC_IN(7) => PC_FETCH_OUT_7_port, PC_IN(6) => 
                           PC_FETCH_OUT_6_port, PC_IN(5) => PC_FETCH_OUT_5_port
                           , PC_IN(4) => PC_FETCH_OUT_4_port, PC_IN(3) => 
                           PC_FETCH_OUT_3_port, PC_IN(2) => PC_FETCH_OUT_2_port
                           , PC_IN(1) => PC_FETCH_OUT_1_port, PC_IN(0) => 
                           PC_FETCH_OUT_0_port, Bubble => n2, HDU_INS_OUT(31) 
                           => sig_HDU_INS_OUT_31_port, HDU_INS_OUT(30) => 
                           sig_HDU_INS_OUT_30_port, HDU_INS_OUT(29) => 
                           sig_HDU_INS_OUT_29_port, HDU_INS_OUT(28) => 
                           sig_HDU_INS_OUT_28_port, HDU_INS_OUT(27) => 
                           sig_HDU_INS_OUT_27_port, HDU_INS_OUT(26) => 
                           sig_HDU_INS_OUT_26_port, HDU_INS_OUT(25) => 
                           sig_HDU_INS_OUT_25_port, HDU_INS_OUT(24) => 
                           sig_HDU_INS_OUT_24_port, HDU_INS_OUT(23) => 
                           sig_HDU_INS_OUT_23_port, HDU_INS_OUT(22) => 
                           sig_HDU_INS_OUT_22_port, HDU_INS_OUT(21) => 
                           sig_HDU_INS_OUT_21_port, HDU_INS_OUT(20) => 
                           sig_HDU_INS_OUT_20_port, HDU_INS_OUT(19) => 
                           sig_HDU_INS_OUT_19_port, HDU_INS_OUT(18) => 
                           sig_HDU_INS_OUT_18_port, HDU_INS_OUT(17) => 
                           sig_HDU_INS_OUT_17_port, HDU_INS_OUT(16) => 
                           sig_HDU_INS_OUT_16_port, HDU_INS_OUT(15) => 
                           sig_HDU_INS_OUT_15_port, HDU_INS_OUT(14) => 
                           sig_HDU_INS_OUT_14_port, HDU_INS_OUT(13) => 
                           sig_HDU_INS_OUT_13_port, HDU_INS_OUT(12) => 
                           sig_HDU_INS_OUT_12_port, HDU_INS_OUT(11) => 
                           sig_HDU_INS_OUT_11_port, HDU_INS_OUT(10) => 
                           sig_HDU_INS_OUT_10_port, HDU_INS_OUT(9) => 
                           sig_HDU_INS_OUT_9_port, HDU_INS_OUT(8) => 
                           sig_HDU_INS_OUT_8_port, HDU_INS_OUT(7) => 
                           sig_HDU_INS_OUT_7_port, HDU_INS_OUT(6) => 
                           sig_HDU_INS_OUT_6_port, HDU_INS_OUT(5) => 
                           sig_HDU_INS_OUT_5_port, HDU_INS_OUT(4) => 
                           sig_HDU_INS_OUT_4_port, HDU_INS_OUT(3) => 
                           sig_HDU_INS_OUT_3_port, HDU_INS_OUT(2) => 
                           sig_HDU_INS_OUT_2_port, HDU_INS_OUT(1) => 
                           sig_HDU_INS_OUT_1_port, HDU_INS_OUT(0) => 
                           sig_HDU_INS_OUT_0_port, HDU_PC_OUT(31) => 
                           sig_HDU_PC_OUT_31_port, HDU_PC_OUT(30) => 
                           sig_HDU_PC_OUT_30_port, HDU_PC_OUT(29) => 
                           sig_HDU_PC_OUT_29_port, HDU_PC_OUT(28) => 
                           sig_HDU_PC_OUT_28_port, HDU_PC_OUT(27) => 
                           sig_HDU_PC_OUT_27_port, HDU_PC_OUT(26) => 
                           sig_HDU_PC_OUT_26_port, HDU_PC_OUT(25) => 
                           sig_HDU_PC_OUT_25_port, HDU_PC_OUT(24) => 
                           sig_HDU_PC_OUT_24_port, HDU_PC_OUT(23) => 
                           sig_HDU_PC_OUT_23_port, HDU_PC_OUT(22) => 
                           sig_HDU_PC_OUT_22_port, HDU_PC_OUT(21) => 
                           sig_HDU_PC_OUT_21_port, HDU_PC_OUT(20) => 
                           sig_HDU_PC_OUT_20_port, HDU_PC_OUT(19) => 
                           sig_HDU_PC_OUT_19_port, HDU_PC_OUT(18) => 
                           sig_HDU_PC_OUT_18_port, HDU_PC_OUT(17) => 
                           sig_HDU_PC_OUT_17_port, HDU_PC_OUT(16) => 
                           sig_HDU_PC_OUT_16_port, HDU_PC_OUT(15) => 
                           sig_HDU_PC_OUT_15_port, HDU_PC_OUT(14) => 
                           sig_HDU_PC_OUT_14_port, HDU_PC_OUT(13) => 
                           sig_HDU_PC_OUT_13_port, HDU_PC_OUT(12) => 
                           sig_HDU_PC_OUT_12_port, HDU_PC_OUT(11) => 
                           sig_HDU_PC_OUT_11_port, HDU_PC_OUT(10) => 
                           sig_HDU_PC_OUT_10_port, HDU_PC_OUT(9) => 
                           sig_HDU_PC_OUT_9_port, HDU_PC_OUT(8) => 
                           sig_HDU_PC_OUT_8_port, HDU_PC_OUT(7) => 
                           sig_HDU_PC_OUT_7_port, HDU_PC_OUT(6) => 
                           sig_HDU_PC_OUT_6_port, HDU_PC_OUT(5) => 
                           sig_HDU_PC_OUT_5_port, HDU_PC_OUT(4) => 
                           sig_HDU_PC_OUT_4_port, HDU_PC_OUT(3) => 
                           sig_HDU_PC_OUT_3_port, HDU_PC_OUT(2) => 
                           sig_HDU_PC_OUT_2_port, HDU_PC_OUT(1) => 
                           sig_HDU_PC_OUT_1_port, HDU_PC_OUT(0) => 
                           sig_HDU_PC_OUT_0_port, HDU_NPC_OUT(31) => 
                           sig_HDU_NPC_OUT_31_port, HDU_NPC_OUT(30) => 
                           sig_HDU_NPC_OUT_30_port, HDU_NPC_OUT(29) => 
                           sig_HDU_NPC_OUT_29_port, HDU_NPC_OUT(28) => 
                           sig_HDU_NPC_OUT_28_port, HDU_NPC_OUT(27) => 
                           sig_HDU_NPC_OUT_27_port, HDU_NPC_OUT(26) => 
                           sig_HDU_NPC_OUT_26_port, HDU_NPC_OUT(25) => 
                           sig_HDU_NPC_OUT_25_port, HDU_NPC_OUT(24) => 
                           sig_HDU_NPC_OUT_24_port, HDU_NPC_OUT(23) => 
                           sig_HDU_NPC_OUT_23_port, HDU_NPC_OUT(22) => 
                           sig_HDU_NPC_OUT_22_port, HDU_NPC_OUT(21) => 
                           sig_HDU_NPC_OUT_21_port, HDU_NPC_OUT(20) => 
                           sig_HDU_NPC_OUT_20_port, HDU_NPC_OUT(19) => 
                           sig_HDU_NPC_OUT_19_port, HDU_NPC_OUT(18) => 
                           sig_HDU_NPC_OUT_18_port, HDU_NPC_OUT(17) => 
                           sig_HDU_NPC_OUT_17_port, HDU_NPC_OUT(16) => 
                           sig_HDU_NPC_OUT_16_port, HDU_NPC_OUT(15) => 
                           sig_HDU_NPC_OUT_15_port, HDU_NPC_OUT(14) => 
                           sig_HDU_NPC_OUT_14_port, HDU_NPC_OUT(13) => 
                           sig_HDU_NPC_OUT_13_port, HDU_NPC_OUT(12) => 
                           sig_HDU_NPC_OUT_12_port, HDU_NPC_OUT(11) => 
                           sig_HDU_NPC_OUT_11_port, HDU_NPC_OUT(10) => 
                           sig_HDU_NPC_OUT_10_port, HDU_NPC_OUT(9) => 
                           sig_HDU_NPC_OUT_9_port, HDU_NPC_OUT(8) => 
                           sig_HDU_NPC_OUT_8_port, HDU_NPC_OUT(7) => 
                           sig_HDU_NPC_OUT_7_port, HDU_NPC_OUT(6) => 
                           sig_HDU_NPC_OUT_6_port, HDU_NPC_OUT(5) => 
                           sig_HDU_NPC_OUT_5_port, HDU_NPC_OUT(4) => 
                           sig_HDU_NPC_OUT_4_port, HDU_NPC_OUT(3) => 
                           sig_HDU_NPC_OUT_3_port, HDU_NPC_OUT(2) => 
                           sig_HDU_NPC_OUT_2_port, HDU_NPC_OUT(1) => 
                           sig_HDU_NPC_OUT_1_port, HDU_NPC_OUT(0) => 
                           sig_HDU_NPC_OUT_0_port);
   U2 : BUF_X1 port map( A => n2, Z => Bubble_out_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( Clk, Rst : in std_logic);

end DLX;

architecture SYN_dlx_rtl of DLX is

   component DRAM
      port( En, Rst : in std_logic;  ADDR_IN, DATA_IN : in std_logic_vector (31
            downto 0);  DRAM_W, DRAM_R : in std_logic;  DATA_OUT : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component IRAM
      port( Rst : in std_logic;  Addr : in std_logic_vector (31 downto 0);  
            Iout : out std_logic_vector (31 downto 0));
   end component;
   
   component hardwired_cu_NBIT32
      port( REG_LATCH_EN, RD1, RD2, MUX_A_SEL : out std_logic;  MUX_B_SEL : out
            std_logic_vector (1 downto 0);  ALU_OPC : out std_logic_vector (0 
            to 3);  ALU_OUTREG_EN, DRAM_R_IN : out std_logic;  JUMP_TYPE : out 
            std_logic_vector (1 downto 0);  MEM_EN_IN, DRAM_W_IN, RF_WE, 
            DRAM_EN_IN, WB_MUX_SEL : out std_logic;  INS_IN : in 
            std_logic_vector (31 downto 0);  Bubble, Clk, Rst : in std_logic);
   end component;
   
   component Datapath
      port( CLK, RST : in std_logic;  INS_IN, DATA_IN : in std_logic_vector (31
            downto 0);  REG_LATCH_EN, RD1, RD2, MUX_A_SEL : in std_logic;  
            MUX_B_SEL : in std_logic_vector (1 downto 0);  ALU_OPC : in 
            std_logic_vector (0 to 3);  ALU_OUTREG_EN : in std_logic;  
            JUMP_TYPE : in std_logic_vector (1 downto 0);  DRAM_R_IN, MEM_EN_IN
            , DRAM_W_IN, RF_WE, DRAM_EN_IN, WB_MUX_SEL : in std_logic;  INS_OUT
            , IRAM_ADDR_OUT, DRAM_ADDR_OUT, DATA_OUT : out std_logic_vector (31
            downto 0);  DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble_out : out 
            std_logic);
   end component;
   
   signal INS_IN_31_port, INS_IN_30_port, INS_IN_29_port, INS_IN_28_port, 
      INS_IN_27_port, INS_IN_26_port, INS_IN_25_port, INS_IN_24_port, 
      INS_IN_23_port, INS_IN_22_port, INS_IN_21_port, INS_IN_20_port, 
      INS_IN_19_port, INS_IN_18_port, INS_IN_17_port, INS_IN_16_port, 
      INS_IN_15_port, INS_IN_14_port, INS_IN_13_port, INS_IN_12_port, 
      INS_IN_11_port, INS_IN_10_port, INS_IN_9_port, INS_IN_8_port, 
      INS_IN_7_port, INS_IN_6_port, INS_IN_5_port, INS_IN_4_port, INS_IN_3_port
      , INS_IN_2_port, INS_IN_1_port, INS_IN_0_port, DATA_IN_31_port, 
      DATA_IN_30_port, DATA_IN_29_port, DATA_IN_28_port, DATA_IN_27_port, 
      DATA_IN_26_port, DATA_IN_25_port, DATA_IN_24_port, DATA_IN_23_port, 
      DATA_IN_22_port, DATA_IN_21_port, DATA_IN_20_port, DATA_IN_19_port, 
      DATA_IN_18_port, DATA_IN_17_port, DATA_IN_16_port, DATA_IN_15_port, 
      DATA_IN_14_port, DATA_IN_13_port, DATA_IN_12_port, DATA_IN_11_port, 
      DATA_IN_10_port, DATA_IN_9_port, DATA_IN_8_port, DATA_IN_7_port, 
      DATA_IN_6_port, DATA_IN_5_port, DATA_IN_4_port, DATA_IN_3_port, 
      DATA_IN_2_port, DATA_IN_1_port, DATA_IN_0_port, REG_LATCH_EN, RD1, RD2, 
      MUX_A_SEL, MUX_B_SEL_1_port, MUX_B_SEL_0_port, ALU_OPC_3_port, 
      ALU_OPC_2_port, ALU_OPC_1_port, ALU_OPC_0_port, ALU_OUTREG_EN, 
      JUMP_TYPE_1_port, JUMP_TYPE_0_port, DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, 
      RF_WE, DRAM_EN_IN, WB_MUX_SEL, IRAM_ADDR_OUT_31_port, 
      IRAM_ADDR_OUT_30_port, IRAM_ADDR_OUT_29_port, IRAM_ADDR_OUT_28_port, 
      IRAM_ADDR_OUT_27_port, IRAM_ADDR_OUT_26_port, IRAM_ADDR_OUT_25_port, 
      IRAM_ADDR_OUT_24_port, IRAM_ADDR_OUT_23_port, IRAM_ADDR_OUT_22_port, 
      IRAM_ADDR_OUT_21_port, IRAM_ADDR_OUT_20_port, IRAM_ADDR_OUT_19_port, 
      IRAM_ADDR_OUT_18_port, IRAM_ADDR_OUT_17_port, IRAM_ADDR_OUT_16_port, 
      IRAM_ADDR_OUT_15_port, IRAM_ADDR_OUT_14_port, IRAM_ADDR_OUT_13_port, 
      IRAM_ADDR_OUT_12_port, IRAM_ADDR_OUT_11_port, IRAM_ADDR_OUT_10_port, 
      IRAM_ADDR_OUT_9_port, IRAM_ADDR_OUT_8_port, IRAM_ADDR_OUT_7_port, 
      IRAM_ADDR_OUT_6_port, IRAM_ADDR_OUT_5_port, IRAM_ADDR_OUT_4_port, 
      IRAM_ADDR_OUT_3_port, IRAM_ADDR_OUT_2_port, IRAM_ADDR_OUT_1_port, 
      IRAM_ADDR_OUT_0_port, DRAM_ADDR_OUT_31_port, DRAM_ADDR_OUT_30_port, 
      DRAM_ADDR_OUT_29_port, DRAM_ADDR_OUT_28_port, DRAM_ADDR_OUT_27_port, 
      DRAM_ADDR_OUT_26_port, DRAM_ADDR_OUT_25_port, DRAM_ADDR_OUT_24_port, 
      DRAM_ADDR_OUT_23_port, DRAM_ADDR_OUT_22_port, DRAM_ADDR_OUT_21_port, 
      DRAM_ADDR_OUT_20_port, DRAM_ADDR_OUT_19_port, DRAM_ADDR_OUT_18_port, 
      DRAM_ADDR_OUT_17_port, DRAM_ADDR_OUT_16_port, DRAM_ADDR_OUT_15_port, 
      DRAM_ADDR_OUT_14_port, DRAM_ADDR_OUT_13_port, DRAM_ADDR_OUT_12_port, 
      DRAM_ADDR_OUT_11_port, DRAM_ADDR_OUT_10_port, DRAM_ADDR_OUT_9_port, 
      DRAM_ADDR_OUT_8_port, DRAM_ADDR_OUT_7_port, DRAM_ADDR_OUT_6_port, 
      DRAM_ADDR_OUT_5_port, DRAM_ADDR_OUT_4_port, DRAM_ADDR_OUT_3_port, 
      DRAM_ADDR_OUT_2_port, DRAM_ADDR_OUT_1_port, DRAM_ADDR_OUT_0_port, 
      DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, DATA_OUT_28_port, 
      DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, DATA_OUT_24_port, 
      DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, DATA_OUT_20_port, 
      DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, DATA_OUT_16_port, 
      DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, DATA_OUT_12_port, 
      DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, DATA_OUT_8_port, 
      DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, DATA_OUT_4_port, 
      DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, DATA_OUT_0_port, 
      DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble, n_1954, n_1955, n_1956, 
      n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, 
      n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, 
      n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, 
      n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, 
      n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000 : 
      std_logic;

begin
   
   DP : Datapath port map( CLK => Clk, RST => Rst, INS_IN(31) => INS_IN_31_port
                           , INS_IN(30) => INS_IN_30_port, INS_IN(29) => 
                           INS_IN_29_port, INS_IN(28) => INS_IN_28_port, 
                           INS_IN(27) => INS_IN_27_port, INS_IN(26) => 
                           INS_IN_26_port, INS_IN(25) => INS_IN_25_port, 
                           INS_IN(24) => INS_IN_24_port, INS_IN(23) => 
                           INS_IN_23_port, INS_IN(22) => INS_IN_22_port, 
                           INS_IN(21) => INS_IN_21_port, INS_IN(20) => 
                           INS_IN_20_port, INS_IN(19) => INS_IN_19_port, 
                           INS_IN(18) => INS_IN_18_port, INS_IN(17) => 
                           INS_IN_17_port, INS_IN(16) => INS_IN_16_port, 
                           INS_IN(15) => INS_IN_15_port, INS_IN(14) => 
                           INS_IN_14_port, INS_IN(13) => INS_IN_13_port, 
                           INS_IN(12) => INS_IN_12_port, INS_IN(11) => 
                           INS_IN_11_port, INS_IN(10) => INS_IN_10_port, 
                           INS_IN(9) => INS_IN_9_port, INS_IN(8) => 
                           INS_IN_8_port, INS_IN(7) => INS_IN_7_port, INS_IN(6)
                           => INS_IN_6_port, INS_IN(5) => INS_IN_5_port, 
                           INS_IN(4) => INS_IN_4_port, INS_IN(3) => 
                           INS_IN_3_port, INS_IN(2) => INS_IN_2_port, INS_IN(1)
                           => INS_IN_1_port, INS_IN(0) => INS_IN_0_port, 
                           DATA_IN(31) => DATA_IN_31_port, DATA_IN(30) => 
                           DATA_IN_30_port, DATA_IN(29) => DATA_IN_29_port, 
                           DATA_IN(28) => DATA_IN_28_port, DATA_IN(27) => 
                           DATA_IN_27_port, DATA_IN(26) => DATA_IN_26_port, 
                           DATA_IN(25) => DATA_IN_25_port, DATA_IN(24) => 
                           DATA_IN_24_port, DATA_IN(23) => DATA_IN_23_port, 
                           DATA_IN(22) => DATA_IN_22_port, DATA_IN(21) => 
                           DATA_IN_21_port, DATA_IN(20) => DATA_IN_20_port, 
                           DATA_IN(19) => DATA_IN_19_port, DATA_IN(18) => 
                           DATA_IN_18_port, DATA_IN(17) => DATA_IN_17_port, 
                           DATA_IN(16) => DATA_IN_16_port, DATA_IN(15) => 
                           DATA_IN_15_port, DATA_IN(14) => DATA_IN_14_port, 
                           DATA_IN(13) => DATA_IN_13_port, DATA_IN(12) => 
                           DATA_IN_12_port, DATA_IN(11) => DATA_IN_11_port, 
                           DATA_IN(10) => DATA_IN_10_port, DATA_IN(9) => 
                           DATA_IN_9_port, DATA_IN(8) => DATA_IN_8_port, 
                           DATA_IN(7) => DATA_IN_7_port, DATA_IN(6) => 
                           DATA_IN_6_port, DATA_IN(5) => DATA_IN_5_port, 
                           DATA_IN(4) => DATA_IN_4_port, DATA_IN(3) => 
                           DATA_IN_3_port, DATA_IN(2) => DATA_IN_2_port, 
                           DATA_IN(1) => DATA_IN_1_port, DATA_IN(0) => 
                           DATA_IN_0_port, REG_LATCH_EN => REG_LATCH_EN, RD1 =>
                           RD1, RD2 => RD2, MUX_A_SEL => MUX_A_SEL, 
                           MUX_B_SEL(1) => MUX_B_SEL_1_port, MUX_B_SEL(0) => 
                           MUX_B_SEL_0_port, ALU_OPC(0) => ALU_OPC_3_port, 
                           ALU_OPC(1) => ALU_OPC_2_port, ALU_OPC(2) => 
                           ALU_OPC_1_port, ALU_OPC(3) => ALU_OPC_0_port, 
                           ALU_OUTREG_EN => ALU_OUTREG_EN, JUMP_TYPE(1) => 
                           JUMP_TYPE_1_port, JUMP_TYPE(0) => JUMP_TYPE_0_port, 
                           DRAM_R_IN => DRAM_R_IN, MEM_EN_IN => MEM_EN_IN, 
                           DRAM_W_IN => DRAM_W_IN, RF_WE => RF_WE, DRAM_EN_IN 
                           => DRAM_EN_IN, WB_MUX_SEL => WB_MUX_SEL, INS_OUT(31)
                           => n_1954, INS_OUT(30) => n_1955, INS_OUT(29) => 
                           n_1956, INS_OUT(28) => n_1957, INS_OUT(27) => n_1958
                           , INS_OUT(26) => n_1959, INS_OUT(25) => n_1960, 
                           INS_OUT(24) => n_1961, INS_OUT(23) => n_1962, 
                           INS_OUT(22) => n_1963, INS_OUT(21) => n_1964, 
                           INS_OUT(20) => n_1965, INS_OUT(19) => n_1966, 
                           INS_OUT(18) => n_1967, INS_OUT(17) => n_1968, 
                           INS_OUT(16) => n_1969, INS_OUT(15) => n_1970, 
                           INS_OUT(14) => n_1971, INS_OUT(13) => n_1972, 
                           INS_OUT(12) => n_1973, INS_OUT(11) => n_1974, 
                           INS_OUT(10) => n_1975, INS_OUT(9) => n_1976, 
                           INS_OUT(8) => n_1977, INS_OUT(7) => n_1978, 
                           INS_OUT(6) => n_1979, INS_OUT(5) => n_1980, 
                           INS_OUT(4) => n_1981, INS_OUT(3) => n_1982, 
                           INS_OUT(2) => n_1983, INS_OUT(1) => n_1984, 
                           INS_OUT(0) => n_1985, IRAM_ADDR_OUT(31) => 
                           IRAM_ADDR_OUT_31_port, IRAM_ADDR_OUT(30) => 
                           IRAM_ADDR_OUT_30_port, IRAM_ADDR_OUT(29) => 
                           IRAM_ADDR_OUT_29_port, IRAM_ADDR_OUT(28) => 
                           IRAM_ADDR_OUT_28_port, IRAM_ADDR_OUT(27) => 
                           IRAM_ADDR_OUT_27_port, IRAM_ADDR_OUT(26) => 
                           IRAM_ADDR_OUT_26_port, IRAM_ADDR_OUT(25) => 
                           IRAM_ADDR_OUT_25_port, IRAM_ADDR_OUT(24) => 
                           IRAM_ADDR_OUT_24_port, IRAM_ADDR_OUT(23) => 
                           IRAM_ADDR_OUT_23_port, IRAM_ADDR_OUT(22) => 
                           IRAM_ADDR_OUT_22_port, IRAM_ADDR_OUT(21) => 
                           IRAM_ADDR_OUT_21_port, IRAM_ADDR_OUT(20) => 
                           IRAM_ADDR_OUT_20_port, IRAM_ADDR_OUT(19) => 
                           IRAM_ADDR_OUT_19_port, IRAM_ADDR_OUT(18) => 
                           IRAM_ADDR_OUT_18_port, IRAM_ADDR_OUT(17) => 
                           IRAM_ADDR_OUT_17_port, IRAM_ADDR_OUT(16) => 
                           IRAM_ADDR_OUT_16_port, IRAM_ADDR_OUT(15) => 
                           IRAM_ADDR_OUT_15_port, IRAM_ADDR_OUT(14) => 
                           IRAM_ADDR_OUT_14_port, IRAM_ADDR_OUT(13) => 
                           IRAM_ADDR_OUT_13_port, IRAM_ADDR_OUT(12) => 
                           IRAM_ADDR_OUT_12_port, IRAM_ADDR_OUT(11) => 
                           IRAM_ADDR_OUT_11_port, IRAM_ADDR_OUT(10) => 
                           IRAM_ADDR_OUT_10_port, IRAM_ADDR_OUT(9) => 
                           IRAM_ADDR_OUT_9_port, IRAM_ADDR_OUT(8) => 
                           IRAM_ADDR_OUT_8_port, IRAM_ADDR_OUT(7) => 
                           IRAM_ADDR_OUT_7_port, IRAM_ADDR_OUT(6) => 
                           IRAM_ADDR_OUT_6_port, IRAM_ADDR_OUT(5) => 
                           IRAM_ADDR_OUT_5_port, IRAM_ADDR_OUT(4) => 
                           IRAM_ADDR_OUT_4_port, IRAM_ADDR_OUT(3) => 
                           IRAM_ADDR_OUT_3_port, IRAM_ADDR_OUT(2) => 
                           IRAM_ADDR_OUT_2_port, IRAM_ADDR_OUT(1) => 
                           IRAM_ADDR_OUT_1_port, IRAM_ADDR_OUT(0) => 
                           IRAM_ADDR_OUT_0_port, DRAM_ADDR_OUT(31) => 
                           DRAM_ADDR_OUT_31_port, DRAM_ADDR_OUT(30) => 
                           DRAM_ADDR_OUT_30_port, DRAM_ADDR_OUT(29) => 
                           DRAM_ADDR_OUT_29_port, DRAM_ADDR_OUT(28) => 
                           DRAM_ADDR_OUT_28_port, DRAM_ADDR_OUT(27) => 
                           DRAM_ADDR_OUT_27_port, DRAM_ADDR_OUT(26) => 
                           DRAM_ADDR_OUT_26_port, DRAM_ADDR_OUT(25) => 
                           DRAM_ADDR_OUT_25_port, DRAM_ADDR_OUT(24) => 
                           DRAM_ADDR_OUT_24_port, DRAM_ADDR_OUT(23) => 
                           DRAM_ADDR_OUT_23_port, DRAM_ADDR_OUT(22) => 
                           DRAM_ADDR_OUT_22_port, DRAM_ADDR_OUT(21) => 
                           DRAM_ADDR_OUT_21_port, DRAM_ADDR_OUT(20) => 
                           DRAM_ADDR_OUT_20_port, DRAM_ADDR_OUT(19) => 
                           DRAM_ADDR_OUT_19_port, DRAM_ADDR_OUT(18) => 
                           DRAM_ADDR_OUT_18_port, DRAM_ADDR_OUT(17) => 
                           DRAM_ADDR_OUT_17_port, DRAM_ADDR_OUT(16) => 
                           DRAM_ADDR_OUT_16_port, DRAM_ADDR_OUT(15) => 
                           DRAM_ADDR_OUT_15_port, DRAM_ADDR_OUT(14) => 
                           DRAM_ADDR_OUT_14_port, DRAM_ADDR_OUT(13) => 
                           DRAM_ADDR_OUT_13_port, DRAM_ADDR_OUT(12) => 
                           DRAM_ADDR_OUT_12_port, DRAM_ADDR_OUT(11) => 
                           DRAM_ADDR_OUT_11_port, DRAM_ADDR_OUT(10) => 
                           DRAM_ADDR_OUT_10_port, DRAM_ADDR_OUT(9) => 
                           DRAM_ADDR_OUT_9_port, DRAM_ADDR_OUT(8) => 
                           DRAM_ADDR_OUT_8_port, DRAM_ADDR_OUT(7) => 
                           DRAM_ADDR_OUT_7_port, DRAM_ADDR_OUT(6) => 
                           DRAM_ADDR_OUT_6_port, DRAM_ADDR_OUT(5) => 
                           DRAM_ADDR_OUT_5_port, DRAM_ADDR_OUT(4) => 
                           DRAM_ADDR_OUT_4_port, DRAM_ADDR_OUT(3) => 
                           DRAM_ADDR_OUT_3_port, DRAM_ADDR_OUT(2) => 
                           DRAM_ADDR_OUT_2_port, DRAM_ADDR_OUT(1) => 
                           DRAM_ADDR_OUT_1_port, DRAM_ADDR_OUT(0) => 
                           DRAM_ADDR_OUT_0_port, DATA_OUT(31) => 
                           DATA_OUT_31_port, DATA_OUT(30) => DATA_OUT_30_port, 
                           DATA_OUT(29) => DATA_OUT_29_port, DATA_OUT(28) => 
                           DATA_OUT_28_port, DATA_OUT(27) => DATA_OUT_27_port, 
                           DATA_OUT(26) => DATA_OUT_26_port, DATA_OUT(25) => 
                           DATA_OUT_25_port, DATA_OUT(24) => DATA_OUT_24_port, 
                           DATA_OUT(23) => DATA_OUT_23_port, DATA_OUT(22) => 
                           DATA_OUT_22_port, DATA_OUT(21) => DATA_OUT_21_port, 
                           DATA_OUT(20) => DATA_OUT_20_port, DATA_OUT(19) => 
                           DATA_OUT_19_port, DATA_OUT(18) => DATA_OUT_18_port, 
                           DATA_OUT(17) => DATA_OUT_17_port, DATA_OUT(16) => 
                           DATA_OUT_16_port, DATA_OUT(15) => DATA_OUT_15_port, 
                           DATA_OUT(14) => DATA_OUT_14_port, DATA_OUT(13) => 
                           DATA_OUT_13_port, DATA_OUT(12) => DATA_OUT_12_port, 
                           DATA_OUT(11) => DATA_OUT_11_port, DATA_OUT(10) => 
                           DATA_OUT_10_port, DATA_OUT(9) => DATA_OUT_9_port, 
                           DATA_OUT(8) => DATA_OUT_8_port, DATA_OUT(7) => 
                           DATA_OUT_7_port, DATA_OUT(6) => DATA_OUT_6_port, 
                           DATA_OUT(5) => DATA_OUT_5_port, DATA_OUT(4) => 
                           DATA_OUT_4_port, DATA_OUT(3) => DATA_OUT_3_port, 
                           DATA_OUT(2) => DATA_OUT_2_port, DATA_OUT(1) => 
                           DATA_OUT_1_port, DATA_OUT(0) => DATA_OUT_0_port, 
                           DRAM_EN_OUT => DRAM_EN_OUT, DRAM_R_OUT => DRAM_R_OUT
                           , DRAM_W_OUT => DRAM_W_OUT, Bubble_out => Bubble);
   CU : hardwired_cu_NBIT32 port map( REG_LATCH_EN => n_1986, RD1 => n_1987, 
                           RD2 => n_1988, MUX_A_SEL => n_1989, MUX_B_SEL(1) => 
                           n_1990, MUX_B_SEL(0) => n_1991, ALU_OPC(0) => 
                           ALU_OPC_3_port, ALU_OPC(1) => ALU_OPC_2_port, 
                           ALU_OPC(2) => ALU_OPC_1_port, ALU_OPC(3) => 
                           ALU_OPC_0_port, ALU_OUTREG_EN => n_1992, DRAM_R_IN 
                           => n_1993, JUMP_TYPE(1) => n_1994, JUMP_TYPE(0) => 
                           n_1995, MEM_EN_IN => n_1996, DRAM_W_IN => n_1997, 
                           RF_WE => n_1998, DRAM_EN_IN => n_1999, WB_MUX_SEL =>
                           n_2000, INS_IN(31) => INS_IN_31_port, INS_IN(30) => 
                           INS_IN_30_port, INS_IN(29) => INS_IN_29_port, 
                           INS_IN(28) => INS_IN_28_port, INS_IN(27) => 
                           INS_IN_27_port, INS_IN(26) => INS_IN_26_port, 
                           INS_IN(25) => INS_IN_25_port, INS_IN(24) => 
                           INS_IN_24_port, INS_IN(23) => INS_IN_23_port, 
                           INS_IN(22) => INS_IN_22_port, INS_IN(21) => 
                           INS_IN_21_port, INS_IN(20) => INS_IN_20_port, 
                           INS_IN(19) => INS_IN_19_port, INS_IN(18) => 
                           INS_IN_18_port, INS_IN(17) => INS_IN_17_port, 
                           INS_IN(16) => INS_IN_16_port, INS_IN(15) => 
                           INS_IN_15_port, INS_IN(14) => INS_IN_14_port, 
                           INS_IN(13) => INS_IN_13_port, INS_IN(12) => 
                           INS_IN_12_port, INS_IN(11) => INS_IN_11_port, 
                           INS_IN(10) => INS_IN_10_port, INS_IN(9) => 
                           INS_IN_9_port, INS_IN(8) => INS_IN_8_port, INS_IN(7)
                           => INS_IN_7_port, INS_IN(6) => INS_IN_6_port, 
                           INS_IN(5) => INS_IN_5_port, INS_IN(4) => 
                           INS_IN_4_port, INS_IN(3) => INS_IN_3_port, INS_IN(2)
                           => INS_IN_2_port, INS_IN(1) => INS_IN_1_port, 
                           INS_IN(0) => INS_IN_0_port, Bubble => Bubble, Clk =>
                           Clk, Rst => Rst);
   IRAM_I : IRAM port map( Rst => Rst, Addr(31) => IRAM_ADDR_OUT_31_port, 
                           Addr(30) => IRAM_ADDR_OUT_30_port, Addr(29) => 
                           IRAM_ADDR_OUT_29_port, Addr(28) => 
                           IRAM_ADDR_OUT_28_port, Addr(27) => 
                           IRAM_ADDR_OUT_27_port, Addr(26) => 
                           IRAM_ADDR_OUT_26_port, Addr(25) => 
                           IRAM_ADDR_OUT_25_port, Addr(24) => 
                           IRAM_ADDR_OUT_24_port, Addr(23) => 
                           IRAM_ADDR_OUT_23_port, Addr(22) => 
                           IRAM_ADDR_OUT_22_port, Addr(21) => 
                           IRAM_ADDR_OUT_21_port, Addr(20) => 
                           IRAM_ADDR_OUT_20_port, Addr(19) => 
                           IRAM_ADDR_OUT_19_port, Addr(18) => 
                           IRAM_ADDR_OUT_18_port, Addr(17) => 
                           IRAM_ADDR_OUT_17_port, Addr(16) => 
                           IRAM_ADDR_OUT_16_port, Addr(15) => 
                           IRAM_ADDR_OUT_15_port, Addr(14) => 
                           IRAM_ADDR_OUT_14_port, Addr(13) => 
                           IRAM_ADDR_OUT_13_port, Addr(12) => 
                           IRAM_ADDR_OUT_12_port, Addr(11) => 
                           IRAM_ADDR_OUT_11_port, Addr(10) => 
                           IRAM_ADDR_OUT_10_port, Addr(9) => 
                           IRAM_ADDR_OUT_9_port, Addr(8) => 
                           IRAM_ADDR_OUT_8_port, Addr(7) => 
                           IRAM_ADDR_OUT_7_port, Addr(6) => 
                           IRAM_ADDR_OUT_6_port, Addr(5) => 
                           IRAM_ADDR_OUT_5_port, Addr(4) => 
                           IRAM_ADDR_OUT_4_port, Addr(3) => 
                           IRAM_ADDR_OUT_3_port, Addr(2) => 
                           IRAM_ADDR_OUT_2_port, Addr(1) => 
                           IRAM_ADDR_OUT_1_port, Addr(0) => 
                           IRAM_ADDR_OUT_0_port, Iout(31) => INS_IN_31_port, 
                           Iout(30) => INS_IN_30_port, Iout(29) => 
                           INS_IN_29_port, Iout(28) => INS_IN_28_port, Iout(27)
                           => INS_IN_27_port, Iout(26) => INS_IN_26_port, 
                           Iout(25) => INS_IN_25_port, Iout(24) => 
                           INS_IN_24_port, Iout(23) => INS_IN_23_port, Iout(22)
                           => INS_IN_22_port, Iout(21) => INS_IN_21_port, 
                           Iout(20) => INS_IN_20_port, Iout(19) => 
                           INS_IN_19_port, Iout(18) => INS_IN_18_port, Iout(17)
                           => INS_IN_17_port, Iout(16) => INS_IN_16_port, 
                           Iout(15) => INS_IN_15_port, Iout(14) => 
                           INS_IN_14_port, Iout(13) => INS_IN_13_port, Iout(12)
                           => INS_IN_12_port, Iout(11) => INS_IN_11_port, 
                           Iout(10) => INS_IN_10_port, Iout(9) => INS_IN_9_port
                           , Iout(8) => INS_IN_8_port, Iout(7) => INS_IN_7_port
                           , Iout(6) => INS_IN_6_port, Iout(5) => INS_IN_5_port
                           , Iout(4) => INS_IN_4_port, Iout(3) => INS_IN_3_port
                           , Iout(2) => INS_IN_2_port, Iout(1) => INS_IN_1_port
                           , Iout(0) => INS_IN_0_port);
   DRAM_I : DRAM port map( En => DRAM_EN_OUT, Rst => Rst, ADDR_IN(31) => 
                           DRAM_ADDR_OUT_31_port, ADDR_IN(30) => 
                           DRAM_ADDR_OUT_30_port, ADDR_IN(29) => 
                           DRAM_ADDR_OUT_29_port, ADDR_IN(28) => 
                           DRAM_ADDR_OUT_28_port, ADDR_IN(27) => 
                           DRAM_ADDR_OUT_27_port, ADDR_IN(26) => 
                           DRAM_ADDR_OUT_26_port, ADDR_IN(25) => 
                           DRAM_ADDR_OUT_25_port, ADDR_IN(24) => 
                           DRAM_ADDR_OUT_24_port, ADDR_IN(23) => 
                           DRAM_ADDR_OUT_23_port, ADDR_IN(22) => 
                           DRAM_ADDR_OUT_22_port, ADDR_IN(21) => 
                           DRAM_ADDR_OUT_21_port, ADDR_IN(20) => 
                           DRAM_ADDR_OUT_20_port, ADDR_IN(19) => 
                           DRAM_ADDR_OUT_19_port, ADDR_IN(18) => 
                           DRAM_ADDR_OUT_18_port, ADDR_IN(17) => 
                           DRAM_ADDR_OUT_17_port, ADDR_IN(16) => 
                           DRAM_ADDR_OUT_16_port, ADDR_IN(15) => 
                           DRAM_ADDR_OUT_15_port, ADDR_IN(14) => 
                           DRAM_ADDR_OUT_14_port, ADDR_IN(13) => 
                           DRAM_ADDR_OUT_13_port, ADDR_IN(12) => 
                           DRAM_ADDR_OUT_12_port, ADDR_IN(11) => 
                           DRAM_ADDR_OUT_11_port, ADDR_IN(10) => 
                           DRAM_ADDR_OUT_10_port, ADDR_IN(9) => 
                           DRAM_ADDR_OUT_9_port, ADDR_IN(8) => 
                           DRAM_ADDR_OUT_8_port, ADDR_IN(7) => 
                           DRAM_ADDR_OUT_7_port, ADDR_IN(6) => 
                           DRAM_ADDR_OUT_6_port, ADDR_IN(5) => 
                           DRAM_ADDR_OUT_5_port, ADDR_IN(4) => 
                           DRAM_ADDR_OUT_4_port, ADDR_IN(3) => 
                           DRAM_ADDR_OUT_3_port, ADDR_IN(2) => 
                           DRAM_ADDR_OUT_2_port, ADDR_IN(1) => 
                           DRAM_ADDR_OUT_1_port, ADDR_IN(0) => 
                           DRAM_ADDR_OUT_0_port, DATA_IN(31) => 
                           DATA_OUT_31_port, DATA_IN(30) => DATA_OUT_30_port, 
                           DATA_IN(29) => DATA_OUT_29_port, DATA_IN(28) => 
                           DATA_OUT_28_port, DATA_IN(27) => DATA_OUT_27_port, 
                           DATA_IN(26) => DATA_OUT_26_port, DATA_IN(25) => 
                           DATA_OUT_25_port, DATA_IN(24) => DATA_OUT_24_port, 
                           DATA_IN(23) => DATA_OUT_23_port, DATA_IN(22) => 
                           DATA_OUT_22_port, DATA_IN(21) => DATA_OUT_21_port, 
                           DATA_IN(20) => DATA_OUT_20_port, DATA_IN(19) => 
                           DATA_OUT_19_port, DATA_IN(18) => DATA_OUT_18_port, 
                           DATA_IN(17) => DATA_OUT_17_port, DATA_IN(16) => 
                           DATA_OUT_16_port, DATA_IN(15) => DATA_OUT_15_port, 
                           DATA_IN(14) => DATA_OUT_14_port, DATA_IN(13) => 
                           DATA_OUT_13_port, DATA_IN(12) => DATA_OUT_12_port, 
                           DATA_IN(11) => DATA_OUT_11_port, DATA_IN(10) => 
                           DATA_OUT_10_port, DATA_IN(9) => DATA_OUT_9_port, 
                           DATA_IN(8) => DATA_OUT_8_port, DATA_IN(7) => 
                           DATA_OUT_7_port, DATA_IN(6) => DATA_OUT_6_port, 
                           DATA_IN(5) => DATA_OUT_5_port, DATA_IN(4) => 
                           DATA_OUT_4_port, DATA_IN(3) => DATA_OUT_3_port, 
                           DATA_IN(2) => DATA_OUT_2_port, DATA_IN(1) => 
                           DATA_OUT_1_port, DATA_IN(0) => DATA_OUT_0_port, 
                           DRAM_W => DRAM_W_OUT, DRAM_R => DRAM_R_OUT, 
                           DATA_OUT(31) => DATA_IN_31_port, DATA_OUT(30) => 
                           DATA_IN_30_port, DATA_OUT(29) => DATA_IN_29_port, 
                           DATA_OUT(28) => DATA_IN_28_port, DATA_OUT(27) => 
                           DATA_IN_27_port, DATA_OUT(26) => DATA_IN_26_port, 
                           DATA_OUT(25) => DATA_IN_25_port, DATA_OUT(24) => 
                           DATA_IN_24_port, DATA_OUT(23) => DATA_IN_23_port, 
                           DATA_OUT(22) => DATA_IN_22_port, DATA_OUT(21) => 
                           DATA_IN_21_port, DATA_OUT(20) => DATA_IN_20_port, 
                           DATA_OUT(19) => DATA_IN_19_port, DATA_OUT(18) => 
                           DATA_IN_18_port, DATA_OUT(17) => DATA_IN_17_port, 
                           DATA_OUT(16) => DATA_IN_16_port, DATA_OUT(15) => 
                           DATA_IN_15_port, DATA_OUT(14) => DATA_IN_14_port, 
                           DATA_OUT(13) => DATA_IN_13_port, DATA_OUT(12) => 
                           DATA_IN_12_port, DATA_OUT(11) => DATA_IN_11_port, 
                           DATA_OUT(10) => DATA_IN_10_port, DATA_OUT(9) => 
                           DATA_IN_9_port, DATA_OUT(8) => DATA_IN_8_port, 
                           DATA_OUT(7) => DATA_IN_7_port, DATA_OUT(6) => 
                           DATA_IN_6_port, DATA_OUT(5) => DATA_IN_5_port, 
                           DATA_OUT(4) => DATA_IN_4_port, DATA_OUT(3) => 
                           DATA_IN_3_port, DATA_OUT(2) => DATA_IN_2_port, 
                           DATA_OUT(1) => DATA_IN_1_port, DATA_OUT(0) => 
                           DATA_IN_0_port);
   WB_MUX_SEL <= '0';
   DRAM_EN_IN <= '0';
   RF_WE <= '0';
   DRAM_W_IN <= '0';
   MEM_EN_IN <= '0';
   JUMP_TYPE_0_port <= '0';
   JUMP_TYPE_1_port <= '0';
   DRAM_R_IN <= '0';
   ALU_OUTREG_EN <= '0';
   MUX_B_SEL_0_port <= '0';
   MUX_B_SEL_1_port <= '0';
   MUX_A_SEL <= '0';
   RD2 <= '0';
   RD1 <= '0';
   REG_LATCH_EN <= '0';

end SYN_dlx_rtl;
