
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type VHDLOUT_TYPE is range 0 to 5;
type aluOp is (NOP, ADDS, SUBS, ANDS, ORS, XORS, SLLS, SRLS, BEQZS, BNEZS, 
   SGES, SLES, NEQS);
attribute ENUM_ENCODING of aluOp : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010 1011 1100";
   
   -- Declarations for conversion functions.
   function integer_to_unsigned(arg, size : in INTEGER) return std_logic_vector
               ;
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 4 )) 
               return aluOp;
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX;

package body CONV_PACK_DLX is
   
   -- integer type to std_logic_vector function
   function integer_to_unsigned(arg, size : in INTEGER) return std_logic_vector
   is 
      variable result: std_logic_vector(size-1 downto 0);
      variable temp: INTEGER;
      -- synopsys built_in SYN_INTEGER_TO_UNSIGNED
   begin
      temp := arg;
      for i in 0 to size-1 loop
         if (temp mod 2) = 1 then
            result(i) := '1';
         else
            result(i) := '0';
         end if;
         temp := temp / 2;
      end loop;
      return result;
   end;
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 4 )) 
   return aluOp is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "0000" => return NOP;
         when "0001" => return ADDS;
         when "0010" => return SUBS;
         when "0011" => return ANDS;
         when "0100" => return ORS;
         when "0101" => return XORS;
         when "0110" => return SLLS;
         when "0111" => return SRLS;
         when "1000" => return BEQZS;
         when "1001" => return BNEZS;
         when "1010" => return SGES;
         when "1011" => return SLES;
         when "1100" => return NEQS;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "0000";
         when ADDS => return "0001";
         when SUBS => return "0010";
         when ANDS => return "0011";
         when ORS => return "0100";
         when XORS => return "0101";
         when SLLS => return "0110";
         when SRLS => return "0111";
         when BEQZS => return "1000";
         when BNEZS => return "1001";
         when SGES => return "1010";
         when SLES => return "1011";
         when NEQS => return "1100";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8;

architecture SYN_structural of SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   component carry_select_basic_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CSBI_1 : carry_select_basic_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) 
                           => A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), 
                           B(1) => B(1), B(0) => B(0), C_i => Ci(0), S(3) => 
                           S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CSBI_2 : carry_select_basic_N4_7 port map( A(3) => A(7), A(2) => A(6), A(1) 
                           => A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), 
                           B(1) => B(5), B(0) => B(4), C_i => Ci(1), S(3) => 
                           S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   CSBI_3 : carry_select_basic_N4_6 port map( A(3) => A(11), A(2) => A(10), 
                           A(1) => A(9), A(0) => A(8), B(3) => B(11), B(2) => 
                           B(10), B(1) => B(9), B(0) => B(8), C_i => Ci(2), 
                           S(3) => S(11), S(2) => S(10), S(1) => S(9), S(0) => 
                           S(8));
   CSBI_4 : carry_select_basic_N4_5 port map( A(3) => A(15), A(2) => A(14), 
                           A(1) => A(13), A(0) => A(12), B(3) => B(15), B(2) =>
                           B(14), B(1) => B(13), B(0) => B(12), C_i => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   CSBI_5 : carry_select_basic_N4_4 port map( A(3) => A(19), A(2) => A(18), 
                           A(1) => A(17), A(0) => A(16), B(3) => B(19), B(2) =>
                           B(18), B(1) => B(17), B(0) => B(16), C_i => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   CSBI_6 : carry_select_basic_N4_3 port map( A(3) => A(23), A(2) => A(22), 
                           A(1) => A(21), A(0) => A(20), B(3) => B(23), B(2) =>
                           B(22), B(1) => B(21), B(0) => B(20), C_i => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   CSBI_7 : carry_select_basic_N4_2 port map( A(3) => A(27), A(2) => A(26), 
                           A(1) => A(25), A(0) => A(24), B(3) => B(27), B(2) =>
                           B(26), B(1) => B(25), B(0) => B(24), C_i => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   CSBI_8 : carry_select_basic_N4_1 port map( A(3) => A(31), A(2) => A(30), 
                           A(1) => A(29), A(0) => A(28), B(3) => B(31), B(2) =>
                           B(30), B(1) => B(29), B(0) => B(28), C_i => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_generator_NBIT32_NBIT_PER_BLOCK4 is

   port( A, B : in std_logic_vector (32 downto 1);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end carry_generator_NBIT32_NBIT_PER_BLOCK4;

architecture SYN_struct of carry_generator_NBIT32_NBIT_PER_BLOCK4 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component PGblock_1
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_2
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_3
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_4
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_5
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_6
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_7
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_8
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_9
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_10
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_11
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_12
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_13
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_14
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_15
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_16
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_17
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_18
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_19
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_20
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_21
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_22
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_23
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_24
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_25
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_26
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_0
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component Gblock_1
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_2
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_3
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_4
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_5
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_6
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_7
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_8
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_0
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_net_1
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_2
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_3
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_4
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_5
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_6
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_7
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_8
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_9
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_10
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_11
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_12
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_13
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_14
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_15
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_16
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_17
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_18
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_19
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_20
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_21
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_22
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_23
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_24
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_25
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_26
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_27
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_28
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_29
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_30
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_0
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   signal Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port, G_1_1_port, n3, P_9_9_port, P_8_8_port, P_8_7_port,
      P_8_5_port, P_7_7_port, P_6_6_port, P_6_5_port, P_5_5_port, P_4_4_port, 
      P_4_3_port, P_3_3_port, P_32_32_port, P_32_31_port, P_32_29_port, 
      P_32_25_port, P_32_17_port, P_31_31_port, P_30_30_port, P_30_29_port, 
      P_2_2_port, P_29_29_port, P_28_28_port, P_28_27_port, P_28_25_port, 
      P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, P_25_25_port, 
      P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, P_23_23_port, 
      P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, P_20_19_port, 
      P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, P_17_17_port, 
      P_16_9_port, P_16_16_port, P_16_15_port, P_16_13_port, P_15_15_port, 
      P_14_14_port, P_14_13_port, P_13_13_port, P_12_9_port, P_12_12_port, 
      P_12_11_port, P_11_11_port, P_10_9_port, P_10_10_port, G_9_9_port, 
      G_8_8_port, G_8_7_port, G_8_5_port, G_7_7_port, G_6_6_port, G_6_5_port, 
      G_5_5_port, G_4_4_port, G_4_3_port, G_3_3_port, G_32_32_port, 
      G_32_31_port, G_32_29_port, G_32_25_port, G_32_17_port, G_31_31_port, 
      G_30_30_port, G_30_29_port, G_2_2_port, G_2_1_port, G_29_29_port, 
      G_28_28_port, G_28_27_port, G_28_25_port, G_28_17_port, G_27_27_port, 
      G_26_26_port, G_26_25_port, G_25_25_port, G_24_24_port, G_24_23_port, 
      G_24_21_port, G_24_17_port, G_23_23_port, G_22_22_port, G_22_21_port, 
      G_21_21_port, G_20_20_port, G_20_19_port, G_20_17_port, G_19_19_port, 
      G_18_18_port, G_18_17_port, G_17_17_port, G_16_9_port, G_16_16_port, 
      G_16_15_port, G_16_13_port, G_15_15_port, G_14_14_port, G_14_13_port, 
      G_13_13_port, G_12_9_port, G_12_12_port, G_12_11_port, G_11_11_port, 
      G_10_9_port, G_10_10_port, n4, n5 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port );
   
   PGnetblock_2 : PG_net_0 port map( a => A(2), b => B(2), p => P_2_2_port, g 
                           => G_2_2_port);
   PGnetblock_3 : PG_net_30 port map( a => A(3), b => B(3), p => P_3_3_port, g 
                           => G_3_3_port);
   PGnetblock_4 : PG_net_29 port map( a => A(4), b => B(4), p => P_4_4_port, g 
                           => G_4_4_port);
   PGnetblock_5 : PG_net_28 port map( a => A(5), b => B(5), p => P_5_5_port, g 
                           => G_5_5_port);
   PGnetblock_6 : PG_net_27 port map( a => A(6), b => B(6), p => P_6_6_port, g 
                           => G_6_6_port);
   PGnetblock_7 : PG_net_26 port map( a => A(7), b => B(7), p => P_7_7_port, g 
                           => G_7_7_port);
   PGnetblock_8 : PG_net_25 port map( a => A(8), b => B(8), p => P_8_8_port, g 
                           => G_8_8_port);
   PGnetblock_9 : PG_net_24 port map( a => A(9), b => B(9), p => P_9_9_port, g 
                           => G_9_9_port);
   PGnetblock_10 : PG_net_23 port map( a => A(10), b => B(10), p => 
                           P_10_10_port, g => G_10_10_port);
   PGnetblock_11 : PG_net_22 port map( a => A(11), b => B(11), p => 
                           P_11_11_port, g => G_11_11_port);
   PGnetblock_12 : PG_net_21 port map( a => A(12), b => B(12), p => 
                           P_12_12_port, g => G_12_12_port);
   PGnetblock_13 : PG_net_20 port map( a => A(13), b => B(13), p => 
                           P_13_13_port, g => G_13_13_port);
   PGnetblock_14 : PG_net_19 port map( a => A(14), b => B(14), p => 
                           P_14_14_port, g => G_14_14_port);
   PGnetblock_15 : PG_net_18 port map( a => A(15), b => B(15), p => 
                           P_15_15_port, g => G_15_15_port);
   PGnetblock_16 : PG_net_17 port map( a => A(16), b => B(16), p => 
                           P_16_16_port, g => G_16_16_port);
   PGnetblock_17 : PG_net_16 port map( a => A(17), b => B(17), p => 
                           P_17_17_port, g => G_17_17_port);
   PGnetblock_18 : PG_net_15 port map( a => A(18), b => B(18), p => 
                           P_18_18_port, g => G_18_18_port);
   PGnetblock_19 : PG_net_14 port map( a => A(19), b => B(19), p => 
                           P_19_19_port, g => G_19_19_port);
   PGnetblock_20 : PG_net_13 port map( a => A(20), b => B(20), p => 
                           P_20_20_port, g => G_20_20_port);
   PGnetblock_21 : PG_net_12 port map( a => A(21), b => B(21), p => 
                           P_21_21_port, g => G_21_21_port);
   PGnetblock_22 : PG_net_11 port map( a => A(22), b => B(22), p => 
                           P_22_22_port, g => G_22_22_port);
   PGnetblock_23 : PG_net_10 port map( a => A(23), b => B(23), p => 
                           P_23_23_port, g => G_23_23_port);
   PGnetblock_24 : PG_net_9 port map( a => A(24), b => B(24), p => P_24_24_port
                           , g => G_24_24_port);
   PGnetblock_25 : PG_net_8 port map( a => A(25), b => B(25), p => P_25_25_port
                           , g => G_25_25_port);
   PGnetblock_26 : PG_net_7 port map( a => A(26), b => B(26), p => P_26_26_port
                           , g => G_26_26_port);
   PGnetblock_27 : PG_net_6 port map( a => A(27), b => B(27), p => P_27_27_port
                           , g => G_27_27_port);
   PGnetblock_28 : PG_net_5 port map( a => A(28), b => B(28), p => P_28_28_port
                           , g => G_28_28_port);
   PGnetblock_29 : PG_net_4 port map( a => A(29), b => B(29), p => P_29_29_port
                           , g => G_29_29_port);
   PGnetblock_30 : PG_net_3 port map( a => A(30), b => B(30), p => P_30_30_port
                           , g => G_30_30_port);
   PGnetblock_31 : PG_net_2 port map( a => A(31), b => B(31), p => P_31_31_port
                           , g => G_31_31_port);
   PGnetblock_32 : PG_net_1 port map( a => A(32), b => B(32), p => P_32_32_port
                           , g => G_32_32_port);
   GB_low_1_2 : Gblock_0 port map( Pik => P_2_2_port, Gik => G_2_2_port, Gk_1j 
                           => G_1_1_port, Gij => G_2_1_port);
   GB_low_2_4 : Gblock_8 port map( Pik => P_4_3_port, Gik => G_4_3_port, Gk_1j 
                           => G_2_1_port, Gij => Co_0_port);
   GB_low_3_8 : Gblock_7 port map( Pik => P_8_5_port, Gik => G_8_5_port, Gk_1j 
                           => Co_0_port, Gij => Co_1_port);
   GB_high_4_16_0 : Gblock_6 port map( Pik => P_16_9_port, Gik => G_16_9_port, 
                           Gk_1j => Co_1_port, Gij => Co_3_port);
   GB_high_4_16_1 : Gblock_5 port map( Pik => P_12_9_port, Gik => G_12_9_port, 
                           Gk_1j => Co_1_port, Gij => Co_2_port);
   GB_high_5_32_0 : Gblock_4 port map( Pik => P_32_17_port, Gik => G_32_17_port
                           , Gk_1j => Co_3_port, Gij => Co_7_port);
   GB_high_5_32_1 : Gblock_3 port map( Pik => P_28_17_port, Gik => G_28_17_port
                           , Gk_1j => Co_3_port, Gij => Co_6_port);
   GB_high_5_32_2 : Gblock_2 port map( Pik => P_24_17_port, Gik => G_24_17_port
                           , Gk_1j => Co_3_port, Gij => Co_5_port);
   GB_high_5_32_3 : Gblock_1 port map( Pik => P_20_17_port, Gik => G_20_17_port
                           , Gk_1j => Co_3_port, Gij => Co_4_port);
   PGB_low_1_4 : PGblock_0 port map( Pik => P_4_4_port, Gik => G_4_4_port, 
                           Pk_1j => P_3_3_port, Gk_1j => G_3_3_port, Pij => 
                           P_4_3_port, Gij => G_4_3_port);
   PGB_low_1_6 : PGblock_26 port map( Pik => P_6_6_port, Gik => G_6_6_port, 
                           Pk_1j => P_5_5_port, Gk_1j => G_5_5_port, Pij => 
                           P_6_5_port, Gij => G_6_5_port);
   PGB_low_1_8 : PGblock_25 port map( Pik => P_8_8_port, Gik => G_8_8_port, 
                           Pk_1j => P_7_7_port, Gk_1j => G_7_7_port, Pij => 
                           P_8_7_port, Gij => G_8_7_port);
   PGB_low_1_10 : PGblock_24 port map( Pik => P_10_10_port, Gik => G_10_10_port
                           , Pk_1j => P_9_9_port, Gk_1j => G_9_9_port, Pij => 
                           P_10_9_port, Gij => G_10_9_port);
   PGB_low_1_12 : PGblock_23 port map( Pik => P_12_12_port, Gik => G_12_12_port
                           , Pk_1j => P_11_11_port, Gk_1j => G_11_11_port, Pij 
                           => P_12_11_port, Gij => G_12_11_port);
   PGB_low_1_14 : PGblock_22 port map( Pik => P_14_14_port, Gik => G_14_14_port
                           , Pk_1j => P_13_13_port, Gk_1j => G_13_13_port, Pij 
                           => P_14_13_port, Gij => G_14_13_port);
   PGB_low_1_16 : PGblock_21 port map( Pik => P_16_16_port, Gik => G_16_16_port
                           , Pk_1j => P_15_15_port, Gk_1j => G_15_15_port, Pij 
                           => P_16_15_port, Gij => G_16_15_port);
   PGB_low_1_18 : PGblock_20 port map( Pik => P_18_18_port, Gik => G_18_18_port
                           , Pk_1j => P_17_17_port, Gk_1j => G_17_17_port, Pij 
                           => P_18_17_port, Gij => G_18_17_port);
   PGB_low_1_20 : PGblock_19 port map( Pik => P_20_20_port, Gik => G_20_20_port
                           , Pk_1j => P_19_19_port, Gk_1j => G_19_19_port, Pij 
                           => P_20_19_port, Gij => G_20_19_port);
   PGB_low_1_22 : PGblock_18 port map( Pik => P_22_22_port, Gik => G_22_22_port
                           , Pk_1j => P_21_21_port, Gk_1j => G_21_21_port, Pij 
                           => P_22_21_port, Gij => G_22_21_port);
   PGB_low_1_24 : PGblock_17 port map( Pik => P_24_24_port, Gik => G_24_24_port
                           , Pk_1j => P_23_23_port, Gk_1j => G_23_23_port, Pij 
                           => P_24_23_port, Gij => G_24_23_port);
   PGB_low_1_26 : PGblock_16 port map( Pik => P_26_26_port, Gik => G_26_26_port
                           , Pk_1j => P_25_25_port, Gk_1j => G_25_25_port, Pij 
                           => P_26_25_port, Gij => G_26_25_port);
   PGB_low_1_28 : PGblock_15 port map( Pik => P_28_28_port, Gik => G_28_28_port
                           , Pk_1j => P_27_27_port, Gk_1j => G_27_27_port, Pij 
                           => P_28_27_port, Gij => G_28_27_port);
   PGB_low_1_30 : PGblock_14 port map( Pik => P_30_30_port, Gik => G_30_30_port
                           , Pk_1j => P_29_29_port, Gk_1j => G_29_29_port, Pij 
                           => P_30_29_port, Gij => G_30_29_port);
   PGB_low_1_32 : PGblock_13 port map( Pik => P_32_32_port, Gik => G_32_32_port
                           , Pk_1j => P_31_31_port, Gk_1j => G_31_31_port, Pij 
                           => P_32_31_port, Gij => G_32_31_port);
   PGB_low_2_8 : PGblock_12 port map( Pik => P_8_7_port, Gik => G_8_7_port, 
                           Pk_1j => P_6_5_port, Gk_1j => G_6_5_port, Pij => 
                           P_8_5_port, Gij => G_8_5_port);
   PGB_low_2_12 : PGblock_11 port map( Pik => P_12_11_port, Gik => G_12_11_port
                           , Pk_1j => P_10_9_port, Gk_1j => G_10_9_port, Pij =>
                           P_12_9_port, Gij => G_12_9_port);
   PGB_low_2_16 : PGblock_10 port map( Pik => P_16_15_port, Gik => G_16_15_port
                           , Pk_1j => P_14_13_port, Gk_1j => G_14_13_port, Pij 
                           => P_16_13_port, Gij => G_16_13_port);
   PGB_low_2_20 : PGblock_9 port map( Pik => P_20_19_port, Gik => G_20_19_port,
                           Pk_1j => P_18_17_port, Gk_1j => G_18_17_port, Pij =>
                           P_20_17_port, Gij => G_20_17_port);
   PGB_low_2_24 : PGblock_8 port map( Pik => P_24_23_port, Gik => G_24_23_port,
                           Pk_1j => P_22_21_port, Gk_1j => G_22_21_port, Pij =>
                           P_24_21_port, Gij => G_24_21_port);
   PGB_low_2_28 : PGblock_7 port map( Pik => P_28_27_port, Gik => G_28_27_port,
                           Pk_1j => P_26_25_port, Gk_1j => G_26_25_port, Pij =>
                           P_28_25_port, Gij => G_28_25_port);
   PGB_low_2_32 : PGblock_6 port map( Pik => P_32_31_port, Gik => G_32_31_port,
                           Pk_1j => P_30_29_port, Gk_1j => G_30_29_port, Pij =>
                           P_32_29_port, Gij => G_32_29_port);
   PGB_low_3_16 : PGblock_5 port map( Pik => P_16_13_port, Gik => G_16_13_port,
                           Pk_1j => P_12_9_port, Gk_1j => G_12_9_port, Pij => 
                           P_16_9_port, Gij => G_16_9_port);
   PGB_low_3_24 : PGblock_4 port map( Pik => P_24_21_port, Gik => G_24_21_port,
                           Pk_1j => P_20_17_port, Gk_1j => G_20_17_port, Pij =>
                           P_24_17_port, Gij => G_24_17_port);
   PGB_low_3_32 : PGblock_3 port map( Pik => P_32_29_port, Gik => G_32_29_port,
                           Pk_1j => P_28_25_port, Gk_1j => G_28_25_port, Pij =>
                           P_32_25_port, Gij => G_32_25_port);
   PGB_high_4_32_0 : PGblock_2 port map( Pik => P_32_25_port, Gik => 
                           G_32_25_port, Pk_1j => P_24_17_port, Gk_1j => 
                           G_24_17_port, Pij => P_32_17_port, Gij => 
                           G_32_17_port);
   PGB_high_4_32_1 : PGblock_1 port map( Pik => P_28_25_port, Gik => 
                           G_28_25_port, Pk_1j => P_24_17_port, Gk_1j => 
                           G_24_17_port, Pij => P_28_17_port, Gij => 
                           G_28_17_port);
   U1 : OAI21_X1 port map( B1 => n4, B2 => n5, A => n3, ZN => G_1_1_port);
   U2 : INV_X1 port map( A => A(1), ZN => n4);
   U3 : INV_X1 port map( A => B(1), ZN => n5);
   U4 : OAI21_X1 port map( B1 => A(1), B2 => B(1), A => Cin, ZN => n3);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity comparator_NBIT32_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end comparator_NBIT32_DW01_cmp6_0;

architecture SYN_rpl of comparator_NBIT32_DW01_cmp6_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal GT_port, GE_port, NE_port, n66, n67, n68, n69, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88
      , n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102
      , n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, LE_port, n206, n207, n208, n209, n210, n211, n212
      , n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
      n261, n262, n263, n264, n265, n266, n267 : std_logic;

begin
   GT <= GT_port;
   LE <= LE_port;
   GE <= GE_port;
   NE <= NE_port;
   
   U103 : XOR2_X1 port map( A => A(30), B => n208, Z => n70);
   U172 : NAND3_X1 port map( A1 => n197, A2 => n150, A3 => n147, ZN => n196);
   U176 : NAND3_X1 port map( A1 => n234, A2 => n199, A3 => n200, ZN => n197);
   U1 : INV_X1 port map( A => n142, ZN => n232);
   U2 : INV_X1 port map( A => n130, ZN => n228);
   U3 : INV_X1 port map( A => n118, ZN => n224);
   U4 : INV_X1 port map( A => n106, ZN => n220);
   U5 : INV_X1 port map( A => n94, ZN => n216);
   U6 : INV_X1 port map( A => n82, ZN => n212);
   U7 : NOR2_X1 port map( A1 => n193, A2 => n136, ZN => n135);
   U8 : NOR2_X1 port map( A1 => n187, A2 => n124, ZN => n123);
   U9 : NOR2_X1 port map( A1 => n181, A2 => n112, ZN => n111);
   U10 : NOR2_X1 port map( A1 => n175, A2 => n100, ZN => n99);
   U11 : NOR2_X1 port map( A1 => n169, A2 => n88, ZN => n87);
   U12 : NOR2_X1 port map( A1 => n163, A2 => n76, ZN => n75);
   U13 : OAI211_X1 port map( C1 => n161, C2 => n162, A => n78, B => n75, ZN => 
                           n160);
   U14 : NAND2_X1 port map( A1 => n210, A2 => n164, ZN => n162);
   U15 : AOI211_X1 port map( C1 => n165, C2 => n166, A => n82, B => n213, ZN =>
                           n161);
   U16 : INV_X1 port map( A => n79, ZN => n210);
   U17 : OAI211_X1 port map( C1 => n191, C2 => n192, A => n138, B => n135, ZN 
                           => n190);
   U18 : NAND2_X1 port map( A1 => n230, A2 => n194, ZN => n192);
   U19 : AOI211_X1 port map( C1 => n195, C2 => n196, A => n142, B => n233, ZN 
                           => n191);
   U20 : INV_X1 port map( A => n139, ZN => n230);
   U21 : OAI211_X1 port map( C1 => n185, C2 => n186, A => n126, B => n123, ZN 
                           => n184);
   U22 : NAND2_X1 port map( A1 => n226, A2 => n188, ZN => n186);
   U23 : AOI211_X1 port map( C1 => n189, C2 => n190, A => n130, B => n229, ZN 
                           => n185);
   U24 : INV_X1 port map( A => n127, ZN => n226);
   U25 : OAI211_X1 port map( C1 => n179, C2 => n180, A => n114, B => n111, ZN 
                           => n178);
   U26 : NAND2_X1 port map( A1 => n222, A2 => n182, ZN => n180);
   U27 : AOI211_X1 port map( C1 => n183, C2 => n184, A => n118, B => n225, ZN 
                           => n179);
   U28 : INV_X1 port map( A => n115, ZN => n222);
   U29 : OAI211_X1 port map( C1 => n173, C2 => n174, A => n102, B => n99, ZN =>
                           n172);
   U30 : NAND2_X1 port map( A1 => n218, A2 => n176, ZN => n174);
   U31 : AOI211_X1 port map( C1 => n177, C2 => n178, A => n106, B => n221, ZN 
                           => n173);
   U32 : INV_X1 port map( A => n103, ZN => n218);
   U33 : OAI211_X1 port map( C1 => n167, C2 => n168, A => n90, B => n87, ZN => 
                           n166);
   U34 : NAND2_X1 port map( A1 => n214, A2 => n170, ZN => n168);
   U35 : AOI211_X1 port map( C1 => n171, C2 => n172, A => n94, B => n217, ZN =>
                           n167);
   U36 : INV_X1 port map( A => n91, ZN => n214);
   U37 : AOI21_X1 port map( B1 => n143, B2 => n144, A => n145, ZN => n140);
   U38 : AOI21_X1 port map( B1 => n146, B2 => n147, A => n148, ZN => n143);
   U39 : AOI21_X1 port map( B1 => n149, B2 => n150, A => n151, ZN => n146);
   U40 : AOI21_X1 port map( B1 => n152, B2 => n153, A => n235, ZN => n149);
   U41 : AOI21_X1 port map( B1 => n131, B2 => n132, A => n133, ZN => n128);
   U42 : AOI21_X1 port map( B1 => n134, B2 => n135, A => n136, ZN => n131);
   U43 : AOI21_X1 port map( B1 => n137, B2 => n138, A => n139, ZN => n134);
   U44 : AOI21_X1 port map( B1 => n140, B2 => n232, A => n231, ZN => n137);
   U45 : AOI21_X1 port map( B1 => n119, B2 => n120, A => n121, ZN => n116);
   U46 : AOI21_X1 port map( B1 => n122, B2 => n123, A => n124, ZN => n119);
   U47 : AOI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n122);
   U48 : AOI21_X1 port map( B1 => n128, B2 => n228, A => n227, ZN => n125);
   U49 : AOI21_X1 port map( B1 => n107, B2 => n108, A => n109, ZN => n104);
   U50 : AOI21_X1 port map( B1 => n110, B2 => n111, A => n112, ZN => n107);
   U51 : AOI21_X1 port map( B1 => n113, B2 => n114, A => n115, ZN => n110);
   U52 : AOI21_X1 port map( B1 => n116, B2 => n224, A => n223, ZN => n113);
   U53 : AOI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n92);
   U54 : AOI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => n95);
   U55 : AOI21_X1 port map( B1 => n101, B2 => n102, A => n103, ZN => n98);
   U56 : AOI21_X1 port map( B1 => n104, B2 => n220, A => n219, ZN => n101);
   U57 : AOI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n80);
   U58 : AOI21_X1 port map( B1 => n86, B2 => n87, A => n88, ZN => n83);
   U59 : AOI21_X1 port map( B1 => n89, B2 => n90, A => n91, ZN => n86);
   U60 : AOI21_X1 port map( B1 => n92, B2 => n216, A => n215, ZN => n89);
   U61 : AOI21_X1 port map( B1 => n71, B2 => n72, A => n73, ZN => n69);
   U62 : AOI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => n71);
   U63 : AOI21_X1 port map( B1 => n77, B2 => n78, A => n79, ZN => n74);
   U64 : AOI21_X1 port map( B1 => n80, B2 => n212, A => n211, ZN => n77);
   U65 : NOR2_X1 port map( A1 => n198, A2 => n148, ZN => n147);
   U66 : NOR2_X1 port map( A1 => n198, A2 => n145, ZN => n195);
   U67 : NOR2_X1 port map( A1 => n193, A2 => n133, ZN => n189);
   U68 : NOR2_X1 port map( A1 => n187, A2 => n121, ZN => n183);
   U69 : NOR2_X1 port map( A1 => n181, A2 => n109, ZN => n177);
   U70 : NOR2_X1 port map( A1 => n175, A2 => n97, ZN => n171);
   U71 : NOR2_X1 port map( A1 => n169, A2 => n85, ZN => n165);
   U72 : NOR2_X1 port map( A1 => n163, A2 => n73, ZN => n159);
   U73 : NAND2_X1 port map( A1 => n194, A2 => n141, ZN => n142);
   U74 : NAND2_X1 port map( A1 => n188, A2 => n129, ZN => n130);
   U75 : NAND2_X1 port map( A1 => n182, A2 => n117, ZN => n118);
   U76 : NAND2_X1 port map( A1 => n176, A2 => n105, ZN => n106);
   U77 : NAND2_X1 port map( A1 => n170, A2 => n93, ZN => n94);
   U78 : NAND2_X1 port map( A1 => n164, A2 => n81, ZN => n82);
   U79 : AND2_X1 port map( A1 => n199, A2 => n154, ZN => n153);
   U80 : INV_X1 port map( A => GT_port, ZN => LE_port);
   U81 : INV_X1 port map( A => n108, ZN => n221);
   U82 : INV_X1 port map( A => n96, ZN => n217);
   U83 : INV_X1 port map( A => n84, ZN => n213);
   U84 : INV_X1 port map( A => n144, ZN => n233);
   U85 : INV_X1 port map( A => n132, ZN => n229);
   U86 : INV_X1 port map( A => n120, ZN => n225);
   U87 : INV_X1 port map( A => n141, ZN => n231);
   U88 : INV_X1 port map( A => n129, ZN => n227);
   U89 : INV_X1 port map( A => n117, ZN => n223);
   U90 : INV_X1 port map( A => n105, ZN => n219);
   U91 : INV_X1 port map( A => n93, ZN => n215);
   U92 : INV_X1 port map( A => n81, ZN => n211);
   U93 : INV_X1 port map( A => n154, ZN => n235);
   U94 : AOI21_X1 port map( B1 => n66, B2 => n207, A => n67, ZN => GE_port);
   U95 : INV_X1 port map( A => n68, ZN => n207);
   U96 : AOI22_X1 port map( A1 => B(30), A2 => n238, B1 => n69, B2 => n70, ZN 
                           => n68);
   U97 : INV_X1 port map( A => A(30), ZN => n238);
   U98 : OAI21_X1 port map( B1 => n67, B2 => n157, A => n66, ZN => GT_port);
   U99 : AOI22_X1 port map( A1 => A(30), A2 => n208, B1 => n158, B2 => n70, ZN 
                           => n157);
   U100 : AOI21_X1 port map( B1 => n159, B2 => n160, A => n209, ZN => n158);
   U101 : INV_X1 port map( A => n72, ZN => n209);
   U102 : INV_X1 port map( A => GE_port, ZN => LT);
   U104 : AOI22_X1 port map( A1 => n155, A2 => n237, B1 => A(1), B2 => n156, ZN
                           => n152);
   U105 : OR2_X1 port map( A1 => n156, A2 => A(1), ZN => n155);
   U106 : NAND2_X1 port map( A1 => B(0), A2 => n267, ZN => n156);
   U107 : NOR2_X1 port map( A1 => n267, A2 => B(0), ZN => n201);
   U108 : NOR2_X1 port map( A1 => n264, A2 => B(4), ZN => n198);
   U109 : NOR2_X1 port map( A1 => n260, A2 => B(8), ZN => n193);
   U110 : NOR2_X1 port map( A1 => n256, A2 => B(12), ZN => n187);
   U111 : NOR2_X1 port map( A1 => n252, A2 => B(16), ZN => n181);
   U112 : NOR2_X1 port map( A1 => n248, A2 => B(20), ZN => n175);
   U113 : NOR2_X1 port map( A1 => n244, A2 => B(24), ZN => n169);
   U114 : NOR2_X1 port map( A1 => n240, A2 => B(28), ZN => n163);
   U115 : NOR2_X1 port map( A1 => n263, A2 => B(5), ZN => n145);
   U116 : NOR2_X1 port map( A1 => n259, A2 => B(9), ZN => n133);
   U117 : NOR2_X1 port map( A1 => n255, A2 => B(13), ZN => n121);
   U118 : NOR2_X1 port map( A1 => n251, A2 => B(17), ZN => n109);
   U119 : NOR2_X1 port map( A1 => n247, A2 => B(21), ZN => n97);
   U120 : NOR2_X1 port map( A1 => n243, A2 => B(25), ZN => n85);
   U121 : NOR2_X1 port map( A1 => n239, A2 => B(29), ZN => n73);
   U122 : NOR2_X1 port map( A1 => n265, A2 => B(3), ZN => n151);
   U123 : NOR2_X1 port map( A1 => n261, A2 => B(7), ZN => n139);
   U124 : NOR2_X1 port map( A1 => n257, A2 => B(11), ZN => n127);
   U125 : NOR2_X1 port map( A1 => n253, A2 => B(15), ZN => n115);
   U126 : NOR2_X1 port map( A1 => n249, A2 => B(19), ZN => n103);
   U127 : NOR2_X1 port map( A1 => n245, A2 => B(23), ZN => n91);
   U128 : NOR2_X1 port map( A1 => n241, A2 => B(27), ZN => n79);
   U129 : NOR2_X1 port map( A1 => n206, A2 => A(31), ZN => n67);
   U130 : INV_X1 port map( A => NE_port, ZN => EQ);
   U131 : NAND2_X1 port map( A1 => LE_port, A2 => GE_port, ZN => NE_port);
   U132 : INV_X1 port map( A => n151, ZN => n234);
   U133 : OAI211_X1 port map( C1 => A(1), C2 => n201, A => n236, B => n153, ZN 
                           => n200);
   U134 : NAND2_X1 port map( A1 => B(7), A2 => n261, ZN => n138);
   U135 : NAND2_X1 port map( A1 => B(11), A2 => n257, ZN => n126);
   U136 : NAND2_X1 port map( A1 => B(15), A2 => n253, ZN => n114);
   U137 : NAND2_X1 port map( A1 => B(19), A2 => n249, ZN => n102);
   U138 : NAND2_X1 port map( A1 => B(23), A2 => n245, ZN => n90);
   U139 : NAND2_X1 port map( A1 => B(27), A2 => n241, ZN => n78);
   U140 : NAND2_X1 port map( A1 => B(5), A2 => n263, ZN => n144);
   U141 : NAND2_X1 port map( A1 => B(9), A2 => n259, ZN => n132);
   U142 : NAND2_X1 port map( A1 => B(13), A2 => n255, ZN => n120);
   U143 : NAND2_X1 port map( A1 => B(17), A2 => n251, ZN => n108);
   U144 : NAND2_X1 port map( A1 => B(21), A2 => n247, ZN => n96);
   U145 : NAND2_X1 port map( A1 => B(25), A2 => n243, ZN => n84);
   U146 : NAND2_X1 port map( A1 => B(29), A2 => n239, ZN => n72);
   U147 : NAND2_X1 port map( A1 => B(6), A2 => n262, ZN => n141);
   U148 : NAND2_X1 port map( A1 => B(10), A2 => n258, ZN => n129);
   U149 : NAND2_X1 port map( A1 => B(14), A2 => n254, ZN => n117);
   U150 : NAND2_X1 port map( A1 => B(18), A2 => n250, ZN => n105);
   U151 : NAND2_X1 port map( A1 => B(22), A2 => n246, ZN => n93);
   U152 : NAND2_X1 port map( A1 => B(26), A2 => n242, ZN => n81);
   U153 : NAND2_X1 port map( A1 => A(31), A2 => n206, ZN => n66);
   U154 : AND2_X1 port map( A1 => B(4), A2 => n264, ZN => n148);
   U155 : AND2_X1 port map( A1 => B(8), A2 => n260, ZN => n136);
   U156 : AND2_X1 port map( A1 => B(12), A2 => n256, ZN => n124);
   U157 : AND2_X1 port map( A1 => B(16), A2 => n252, ZN => n112);
   U158 : AND2_X1 port map( A1 => B(20), A2 => n248, ZN => n100);
   U159 : AND2_X1 port map( A1 => B(24), A2 => n244, ZN => n88);
   U160 : AND2_X1 port map( A1 => B(28), A2 => n240, ZN => n76);
   U161 : NAND2_X1 port map( A1 => B(3), A2 => n265, ZN => n150);
   U162 : NAND2_X1 port map( A1 => B(2), A2 => n266, ZN => n154);
   U163 : INV_X1 port map( A => A(0), ZN => n267);
   U164 : INV_X1 port map( A => A(3), ZN => n265);
   U165 : INV_X1 port map( A => A(5), ZN => n263);
   U166 : INV_X1 port map( A => A(7), ZN => n261);
   U167 : INV_X1 port map( A => A(9), ZN => n259);
   U168 : INV_X1 port map( A => A(11), ZN => n257);
   U169 : INV_X1 port map( A => A(13), ZN => n255);
   U170 : INV_X1 port map( A => A(15), ZN => n253);
   U171 : INV_X1 port map( A => A(17), ZN => n251);
   U173 : INV_X1 port map( A => A(19), ZN => n249);
   U174 : INV_X1 port map( A => A(21), ZN => n247);
   U175 : INV_X1 port map( A => A(23), ZN => n245);
   U177 : INV_X1 port map( A => A(25), ZN => n243);
   U178 : INV_X1 port map( A => A(29), ZN => n239);
   U179 : INV_X1 port map( A => A(27), ZN => n241);
   U180 : INV_X1 port map( A => B(31), ZN => n206);
   U181 : INV_X1 port map( A => B(1), ZN => n237);
   U182 : OR2_X1 port map( A1 => n262, A2 => B(6), ZN => n194);
   U183 : OR2_X1 port map( A1 => n258, A2 => B(10), ZN => n188);
   U184 : OR2_X1 port map( A1 => n254, A2 => B(14), ZN => n182);
   U185 : OR2_X1 port map( A1 => n250, A2 => B(18), ZN => n176);
   U186 : OR2_X1 port map( A1 => n246, A2 => B(22), ZN => n170);
   U187 : OR2_X1 port map( A1 => n242, A2 => B(26), ZN => n164);
   U188 : INV_X1 port map( A => B(30), ZN => n208);
   U189 : INV_X1 port map( A => A(2), ZN => n266);
   U190 : INV_X1 port map( A => A(6), ZN => n262);
   U191 : INV_X1 port map( A => A(10), ZN => n258);
   U192 : INV_X1 port map( A => A(14), ZN => n254);
   U193 : INV_X1 port map( A => A(18), ZN => n250);
   U194 : INV_X1 port map( A => A(22), ZN => n246);
   U195 : INV_X1 port map( A => A(26), ZN => n242);
   U196 : INV_X1 port map( A => A(4), ZN => n264);
   U197 : INV_X1 port map( A => A(8), ZN => n260);
   U198 : INV_X1 port map( A => A(12), ZN => n256);
   U199 : INV_X1 port map( A => A(16), ZN => n252);
   U200 : INV_X1 port map( A => A(20), ZN => n248);
   U201 : INV_X1 port map( A => A(24), ZN => n244);
   U202 : INV_X1 port map( A => A(28), ZN => n240);
   U203 : OR2_X1 port map( A1 => n266, A2 => B(2), ZN => n199);
   U204 : INV_X1 port map( A => n202, ZN => n236);
   U205 : AOI21_X1 port map( B1 => A(1), B2 => n201, A => n237, ZN => n202);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity P4Adder_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (31 downto 0);  Cout : out std_logic);

end P4Adder_NBIT32;

architecture SYN_struct of P4Adder_NBIT32 is

   component SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component carry_generator_NBIT32_NBIT_PER_BLOCK4
      port( A, B : in std_logic_vector (32 downto 1);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal Csum_7_port, Csum_6_port, Csum_5_port, Csum_4_port, Csum_3_port, 
      Csum_2_port, Csum_1_port : std_logic;

begin
   
   Carrygen0 : carry_generator_NBIT32_NBIT_PER_BLOCK4 port map( A(32) => A(31),
                           A(31) => A(30), A(30) => A(29), A(29) => A(28), 
                           A(28) => A(27), A(27) => A(26), A(26) => A(25), 
                           A(25) => A(24), A(24) => A(23), A(23) => A(22), 
                           A(22) => A(21), A(21) => A(20), A(20) => A(19), 
                           A(19) => A(18), A(18) => A(17), A(17) => A(16), 
                           A(16) => A(15), A(15) => A(14), A(14) => A(13), 
                           A(13) => A(12), A(12) => A(11), A(11) => A(10), 
                           A(10) => A(9), A(9) => A(8), A(8) => A(7), A(7) => 
                           A(6), A(6) => A(5), A(5) => A(4), A(4) => A(3), A(3)
                           => A(2), A(2) => A(1), A(1) => A(0), B(32) => B(31),
                           B(31) => B(30), B(30) => B(29), B(29) => B(28), 
                           B(28) => B(27), B(27) => B(26), B(26) => B(25), 
                           B(25) => B(24), B(24) => B(23), B(23) => B(22), 
                           B(22) => B(21), B(21) => B(20), B(20) => B(19), 
                           B(19) => B(18), B(18) => B(17), B(17) => B(16), 
                           B(16) => B(15), B(15) => B(14), B(14) => B(13), 
                           B(13) => B(12), B(12) => B(11), B(11) => B(10), 
                           B(10) => B(9), B(9) => B(8), B(8) => B(7), B(7) => 
                           B(6), B(6) => B(5), B(5) => B(4), B(4) => B(3), B(3)
                           => B(2), B(2) => B(1), B(1) => B(0), Cin => Cin, 
                           Co(7) => Cout, Co(6) => Csum_7_port, Co(5) => 
                           Csum_6_port, Co(4) => Csum_5_port, Co(3) => 
                           Csum_4_port, Co(2) => Csum_3_port, Co(1) => 
                           Csum_2_port, Co(0) => Csum_1_port);
   Sumgen0 : SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), Ci(7) => 
                           Csum_7_port, Ci(6) => Csum_6_port, Ci(5) => 
                           Csum_5_port, Ci(4) => Csum_4_port, Ci(3) => 
                           Csum_3_port, Ci(2) => Csum_2_port, Ci(1) => 
                           Csum_1_port, Ci(0) => Cin, S(31) => S(31), S(30) => 
                           S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           S(21), S(20) => S(20), S(19) => S(19), S(18) => 
                           S(18), S(17) => S(17), S(16) => S(16), S(15) => 
                           S(15), S(14) => S(14), S(13) => S(13), S(12) => 
                           S(12), S(11) => S(11), S(10) => S(10), S(9) => S(9),
                           S(8) => S(8), S(7) => S(7), S(6) => S(6), S(5) => 
                           S(5), S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1)
                           => S(1), S(0) => S(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity comparator_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  OPSel : in std_logic_vector
         (0 to 2);  RES : out std_logic_vector (31 downto 0));

end comparator_NBIT32;

architecture SYN_bhv of comparator_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component comparator_NBIT32_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   signal X_Logic0_port, N26, N27, N28, N29, N30, N31, n1, n6, n7, n8, n9, n11,
      n12, RES_0_port, n10, n13, n14 : std_logic;

begin
   RES <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, RES_0_port 
      );
   
   X_Logic0_port <= '0';
   n1 <= '0';
   r57 : comparator_NBIT32_DW01_cmp6_0 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), TC => n1, LT => N30, GT => N28, 
                           EQ => N26, LE => N31, GE => N29, NE => N27);
   U2 : AOI22_X1 port map( A1 => N30, A2 => n14, B1 => OPSel(2), B2 => N31, ZN 
                           => n9);
   U4 : AOI22_X1 port map( A1 => N26, A2 => n14, B1 => N27, B2 => OPSel(2), ZN 
                           => n12);
   U5 : AOI22_X1 port map( A1 => N28, A2 => n14, B1 => N29, B2 => OPSel(2), ZN 
                           => n11);
   U6 : INV_X1 port map( A => OPSel(0), ZN => n10);
   U7 : INV_X1 port map( A => OPSel(1), ZN => n13);
   U8 : INV_X1 port map( A => n6, ZN => RES_0_port);
   U9 : AOI21_X1 port map( B1 => n7, B2 => n10, A => n8, ZN => n6);
   U10 : NOR3_X1 port map( A1 => n10, A2 => OPSel(1), A3 => n9, ZN => n8);
   U11 : OAI22_X1 port map( A1 => n11, A2 => n13, B1 => OPSel(1), B2 => n12, ZN
                           => n7);
   U12 : INV_X1 port map( A => OPSel(2), ZN => n14);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HazardDetection_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end HazardDetection_DW01_sub_0;

architecture SYN_rpl of HazardDetection_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port,
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, carry_30_port, 
      carry_29_port, carry_28_port, carry_27_port, carry_26_port, carry_25_port
      , carry_24_port, carry_23_port, carry_22_port, carry_21_port, 
      carry_20_port, carry_19_port, carry_18_port, carry_17_port, carry_16_port
      , carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, n2, DIFF_2_port : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, A(1), A(0) );
   
   U1 : OR2_X1 port map( A1 => A(4), A2 => carry_4_port, ZN => carry_5_port);
   U2 : OR2_X1 port map( A1 => A(5), A2 => carry_5_port, ZN => carry_6_port);
   U3 : OR2_X1 port map( A1 => A(6), A2 => carry_6_port, ZN => carry_7_port);
   U4 : OR2_X1 port map( A1 => A(7), A2 => carry_7_port, ZN => carry_8_port);
   U5 : OR2_X1 port map( A1 => A(8), A2 => carry_8_port, ZN => carry_9_port);
   U6 : OR2_X1 port map( A1 => A(9), A2 => carry_9_port, ZN => carry_10_port);
   U7 : OR2_X1 port map( A1 => A(10), A2 => carry_10_port, ZN => carry_11_port)
                           ;
   U8 : OR2_X1 port map( A1 => A(11), A2 => carry_11_port, ZN => carry_12_port)
                           ;
   U9 : OR2_X1 port map( A1 => A(12), A2 => carry_12_port, ZN => carry_13_port)
                           ;
   U10 : OR2_X1 port map( A1 => A(13), A2 => carry_13_port, ZN => carry_14_port
                           );
   U11 : OR2_X1 port map( A1 => A(14), A2 => carry_14_port, ZN => carry_15_port
                           );
   U12 : OR2_X1 port map( A1 => A(15), A2 => carry_15_port, ZN => carry_16_port
                           );
   U13 : OR2_X1 port map( A1 => A(16), A2 => carry_16_port, ZN => carry_17_port
                           );
   U14 : OR2_X1 port map( A1 => A(17), A2 => carry_17_port, ZN => carry_18_port
                           );
   U15 : OR2_X1 port map( A1 => A(18), A2 => carry_18_port, ZN => carry_19_port
                           );
   U16 : OR2_X1 port map( A1 => A(19), A2 => carry_19_port, ZN => carry_20_port
                           );
   U17 : OR2_X1 port map( A1 => A(20), A2 => carry_20_port, ZN => carry_21_port
                           );
   U18 : OR2_X1 port map( A1 => A(21), A2 => carry_21_port, ZN => carry_22_port
                           );
   U19 : OR2_X1 port map( A1 => A(22), A2 => carry_22_port, ZN => carry_23_port
                           );
   U20 : OR2_X1 port map( A1 => A(23), A2 => carry_23_port, ZN => carry_24_port
                           );
   U21 : OR2_X1 port map( A1 => A(24), A2 => carry_24_port, ZN => carry_25_port
                           );
   U22 : OR2_X1 port map( A1 => A(25), A2 => carry_25_port, ZN => carry_26_port
                           );
   U23 : OR2_X1 port map( A1 => A(26), A2 => carry_26_port, ZN => carry_27_port
                           );
   U24 : OR2_X1 port map( A1 => A(27), A2 => carry_27_port, ZN => carry_28_port
                           );
   U25 : OR2_X1 port map( A1 => A(28), A2 => carry_28_port, ZN => carry_29_port
                           );
   U26 : OR2_X1 port map( A1 => A(29), A2 => carry_29_port, ZN => carry_30_port
                           );
   U27 : OR2_X1 port map( A1 => A(3), A2 => A(2), ZN => carry_4_port);
   U28 : XNOR2_X1 port map( A => A(4), B => carry_4_port, ZN => DIFF_4_port);
   U29 : XNOR2_X1 port map( A => A(5), B => carry_5_port, ZN => DIFF_5_port);
   U30 : XNOR2_X1 port map( A => A(6), B => carry_6_port, ZN => DIFF_6_port);
   U31 : XNOR2_X1 port map( A => A(7), B => carry_7_port, ZN => DIFF_7_port);
   U32 : XNOR2_X1 port map( A => A(8), B => carry_8_port, ZN => DIFF_8_port);
   U33 : XNOR2_X1 port map( A => A(9), B => carry_9_port, ZN => DIFF_9_port);
   U34 : XNOR2_X1 port map( A => A(10), B => carry_10_port, ZN => DIFF_10_port)
                           ;
   U35 : XNOR2_X1 port map( A => A(11), B => carry_11_port, ZN => DIFF_11_port)
                           ;
   U36 : XNOR2_X1 port map( A => A(12), B => carry_12_port, ZN => DIFF_12_port)
                           ;
   U37 : XNOR2_X1 port map( A => A(13), B => carry_13_port, ZN => DIFF_13_port)
                           ;
   U38 : XNOR2_X1 port map( A => A(14), B => carry_14_port, ZN => DIFF_14_port)
                           ;
   U39 : XNOR2_X1 port map( A => A(15), B => carry_15_port, ZN => DIFF_15_port)
                           ;
   U40 : XNOR2_X1 port map( A => A(16), B => carry_16_port, ZN => DIFF_16_port)
                           ;
   U41 : XNOR2_X1 port map( A => A(17), B => carry_17_port, ZN => DIFF_17_port)
                           ;
   U42 : XNOR2_X1 port map( A => A(18), B => carry_18_port, ZN => DIFF_18_port)
                           ;
   U43 : XNOR2_X1 port map( A => A(19), B => carry_19_port, ZN => DIFF_19_port)
                           ;
   U44 : XNOR2_X1 port map( A => A(20), B => carry_20_port, ZN => DIFF_20_port)
                           ;
   U45 : XNOR2_X1 port map( A => A(21), B => carry_21_port, ZN => DIFF_21_port)
                           ;
   U46 : XNOR2_X1 port map( A => A(22), B => carry_22_port, ZN => DIFF_22_port)
                           ;
   U47 : XNOR2_X1 port map( A => A(23), B => carry_23_port, ZN => DIFF_23_port)
                           ;
   U48 : XNOR2_X1 port map( A => A(24), B => carry_24_port, ZN => DIFF_24_port)
                           ;
   U49 : XNOR2_X1 port map( A => A(25), B => carry_25_port, ZN => DIFF_25_port)
                           ;
   U50 : XNOR2_X1 port map( A => A(26), B => carry_26_port, ZN => DIFF_26_port)
                           ;
   U51 : XNOR2_X1 port map( A => A(27), B => carry_27_port, ZN => DIFF_27_port)
                           ;
   U52 : XNOR2_X1 port map( A => A(28), B => carry_28_port, ZN => DIFF_28_port)
                           ;
   U53 : XNOR2_X1 port map( A => A(29), B => carry_29_port, ZN => DIFF_29_port)
                           ;
   U54 : XNOR2_X1 port map( A => A(30), B => carry_30_port, ZN => DIFF_30_port)
                           ;
   U55 : XOR2_X1 port map( A => A(31), B => n2, Z => DIFF_31_port);
   U56 : NOR2_X1 port map( A1 => A(30), A2 => carry_30_port, ZN => n2);
   U57 : XNOR2_X1 port map( A => A(3), B => A(2), ZN => DIFF_3_port);
   U58 : INV_X1 port map( A => A(2), ZN => DIFF_2_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Execute_DW01_add_0;

architecture SYN_rpl of Execute_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n2, n_1037 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1037, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n2, CO => carry_2_port, S
                           => SUM(1));
   U1 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U2 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n2);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute_DW01_add_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Execute_DW01_add_1;

architecture SYN_rpl of Execute_DW01_add_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_3_port, SUM_4_port, SUM_5_port, SUM_6_port, 
      SUM_7_port, SUM_8_port, SUM_9_port, SUM_10_port, SUM_11_port, SUM_12_port
      , SUM_13_port, SUM_14_port, SUM_15_port, SUM_16_port, SUM_17_port, 
      SUM_18_port, SUM_19_port, SUM_20_port, SUM_21_port, SUM_22_port, 
      SUM_23_port, SUM_24_port, SUM_25_port, SUM_26_port, SUM_27_port, 
      SUM_28_port, SUM_29_port, SUM_30_port, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n54, n55, n56, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, B(1), B(0) );
   
   U4 : XOR2_X1 port map( A => B(3), B => B(2), Z => SUM_3_port);
   U5 : XOR2_X1 port map( A => B(4), B => n30, Z => SUM_4_port);
   U6 : XOR2_X1 port map( A => B(5), B => n31, Z => SUM_5_port);
   U7 : XOR2_X1 port map( A => B(6), B => n32, Z => SUM_6_port);
   U8 : XOR2_X1 port map( A => B(7), B => n33, Z => SUM_7_port);
   U9 : XOR2_X1 port map( A => B(8), B => n34, Z => SUM_8_port);
   U10 : XOR2_X1 port map( A => B(9), B => n35, Z => SUM_9_port);
   U11 : XOR2_X1 port map( A => B(10), B => n36, Z => SUM_10_port);
   U12 : XOR2_X1 port map( A => B(11), B => n37, Z => SUM_11_port);
   U13 : XOR2_X1 port map( A => B(12), B => n38, Z => SUM_12_port);
   U14 : XOR2_X1 port map( A => B(13), B => n39, Z => SUM_13_port);
   U15 : XOR2_X1 port map( A => B(14), B => n40, Z => SUM_14_port);
   U16 : XOR2_X1 port map( A => B(15), B => n41, Z => SUM_15_port);
   U17 : XOR2_X1 port map( A => B(16), B => n42, Z => SUM_16_port);
   U18 : XOR2_X1 port map( A => B(17), B => n43, Z => SUM_17_port);
   U19 : XOR2_X1 port map( A => B(18), B => n44, Z => SUM_18_port);
   U20 : XOR2_X1 port map( A => B(19), B => n45, Z => SUM_19_port);
   U21 : XOR2_X1 port map( A => B(20), B => n46, Z => SUM_20_port);
   U22 : XOR2_X1 port map( A => B(21), B => n47, Z => SUM_21_port);
   U23 : XOR2_X1 port map( A => B(22), B => n48, Z => SUM_22_port);
   U24 : XOR2_X1 port map( A => B(23), B => n49, Z => SUM_23_port);
   U25 : XOR2_X1 port map( A => B(24), B => n50, Z => SUM_24_port);
   U26 : XOR2_X1 port map( A => B(25), B => n51, Z => SUM_25_port);
   U27 : XOR2_X1 port map( A => B(26), B => n52, Z => SUM_26_port);
   U28 : XOR2_X1 port map( A => B(27), B => n53, Z => SUM_27_port);
   U29 : XOR2_X1 port map( A => B(28), B => n54, Z => SUM_28_port);
   U30 : XOR2_X1 port map( A => B(29), B => n55, Z => SUM_29_port);
   U31 : XOR2_X1 port map( A => B(30), B => n56, Z => SUM_30_port);
   U1 : INV_X1 port map( A => B(2), ZN => SUM_2_port);
   U2 : AND2_X1 port map( A1 => B(29), A2 => n55, ZN => n56);
   U3 : AND2_X1 port map( A1 => B(4), A2 => n30, ZN => n31);
   U32 : AND2_X1 port map( A1 => B(5), A2 => n31, ZN => n32);
   U33 : AND2_X1 port map( A1 => B(6), A2 => n32, ZN => n33);
   U34 : AND2_X1 port map( A1 => B(7), A2 => n33, ZN => n34);
   U35 : AND2_X1 port map( A1 => B(8), A2 => n34, ZN => n35);
   U36 : AND2_X1 port map( A1 => B(9), A2 => n35, ZN => n36);
   U37 : AND2_X1 port map( A1 => B(10), A2 => n36, ZN => n37);
   U38 : AND2_X1 port map( A1 => B(11), A2 => n37, ZN => n38);
   U39 : AND2_X1 port map( A1 => B(12), A2 => n38, ZN => n39);
   U40 : AND2_X1 port map( A1 => B(13), A2 => n39, ZN => n40);
   U41 : AND2_X1 port map( A1 => B(14), A2 => n40, ZN => n41);
   U42 : AND2_X1 port map( A1 => B(15), A2 => n41, ZN => n42);
   U43 : AND2_X1 port map( A1 => B(16), A2 => n42, ZN => n43);
   U44 : AND2_X1 port map( A1 => B(17), A2 => n43, ZN => n44);
   U45 : AND2_X1 port map( A1 => B(18), A2 => n44, ZN => n45);
   U46 : AND2_X1 port map( A1 => B(19), A2 => n45, ZN => n46);
   U47 : AND2_X1 port map( A1 => B(20), A2 => n46, ZN => n47);
   U48 : AND2_X1 port map( A1 => B(21), A2 => n47, ZN => n48);
   U49 : AND2_X1 port map( A1 => B(22), A2 => n48, ZN => n49);
   U50 : AND2_X1 port map( A1 => B(23), A2 => n49, ZN => n50);
   U51 : AND2_X1 port map( A1 => B(24), A2 => n50, ZN => n51);
   U52 : AND2_X1 port map( A1 => B(25), A2 => n51, ZN => n52);
   U53 : AND2_X1 port map( A1 => B(26), A2 => n52, ZN => n53);
   U54 : AND2_X1 port map( A1 => B(27), A2 => n53, ZN => n54);
   U55 : AND2_X1 port map( A1 => B(28), A2 => n54, ZN => n55);
   U56 : AND2_X1 port map( A1 => B(3), A2 => B(2), ZN => n30);
   U57 : XNOR2_X1 port map( A => B(31), B => n57, ZN => SUM_31_port);
   U58 : NAND2_X1 port map( A1 => B(30), A2 => n56, ZN => n57);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_NBIT32 is

   port( OP1, OP2 : in std_logic_vector (31 downto 0);  ALU_OPC : in 
         std_logic_vector (0 to 3);  ALU_RES : out std_logic_vector (31 downto 
         0));

end ALU_NBIT32;

architecture SYN_struct of ALU_NBIT32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux21_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux41_NBIT32_1
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component P4Adder_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component shifter
      port( A, B : in std_logic_vector (31 downto 0);  LOGIC_ARITH, LEFT_RIGHT 
            : in std_logic;  RES : out std_logic_vector (31 downto 0));
   end component;
   
   component comparator_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  OPSel : in 
            std_logic_vector (0 to 2);  RES : out std_logic_vector (31 downto 
            0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal select_type_sig_1_port, select_type_sig_0_port, select_zero_sig, 
      ADD_SUB, A_ADD_31_port, A_ADD_30_port, A_ADD_29_port, A_ADD_28_port, 
      A_ADD_27_port, A_ADD_26_port, A_ADD_25_port, A_ADD_24_port, A_ADD_23_port
      , A_ADD_22_port, A_ADD_21_port, A_ADD_20_port, A_ADD_19_port, 
      A_ADD_18_port, A_ADD_17_port, A_ADD_16_port, A_ADD_15_port, A_ADD_14_port
      , A_ADD_13_port, A_ADD_12_port, A_ADD_11_port, A_ADD_10_port, 
      A_ADD_9_port, A_ADD_8_port, A_ADD_7_port, A_ADD_6_port, A_ADD_5_port, 
      A_ADD_4_port, A_ADD_3_port, A_ADD_2_port, A_ADD_1_port, A_ADD_0_port, 
      B_ADD_31_port, B_ADD_30_port, B_ADD_29_port, B_ADD_28_port, B_ADD_27_port
      , B_ADD_26_port, B_ADD_25_port, B_ADD_24_port, B_ADD_23_port, 
      B_ADD_22_port, B_ADD_21_port, B_ADD_20_port, B_ADD_19_port, B_ADD_18_port
      , B_ADD_17_port, B_ADD_16_port, B_ADD_15_port, B_ADD_14_port, 
      B_ADD_13_port, B_ADD_12_port, B_ADD_11_port, B_ADD_10_port, B_ADD_9_port,
      B_ADD_8_port, B_ADD_7_port, B_ADD_6_port, B_ADD_5_port, B_ADD_4_port, 
      B_ADD_3_port, B_ADD_2_port, B_ADD_1_port, B_ADD_0_port, LOGIC_RES_31_port
      , LOGIC_RES_30_port, LOGIC_RES_29_port, LOGIC_RES_28_port, 
      LOGIC_RES_27_port, LOGIC_RES_26_port, LOGIC_RES_25_port, 
      LOGIC_RES_24_port, LOGIC_RES_23_port, LOGIC_RES_22_port, 
      LOGIC_RES_21_port, LOGIC_RES_20_port, LOGIC_RES_19_port, 
      LOGIC_RES_18_port, LOGIC_RES_17_port, LOGIC_RES_16_port, 
      LOGIC_RES_15_port, LOGIC_RES_14_port, LOGIC_RES_13_port, 
      LOGIC_RES_12_port, LOGIC_RES_11_port, LOGIC_RES_10_port, LOGIC_RES_9_port
      , LOGIC_RES_8_port, LOGIC_RES_7_port, LOGIC_RES_6_port, LOGIC_RES_5_port,
      LOGIC_RES_4_port, LOGIC_RES_3_port, LOGIC_RES_2_port, LOGIC_RES_1_port, 
      LOGIC_RES_0_port, LEFT_RIGHT, A_SHF_31_port, A_SHF_30_port, A_SHF_29_port
      , A_SHF_28_port, A_SHF_27_port, A_SHF_26_port, A_SHF_25_port, 
      A_SHF_24_port, A_SHF_23_port, A_SHF_22_port, A_SHF_21_port, A_SHF_20_port
      , A_SHF_19_port, A_SHF_18_port, A_SHF_17_port, A_SHF_16_port, 
      A_SHF_15_port, A_SHF_14_port, A_SHF_13_port, A_SHF_12_port, A_SHF_11_port
      , A_SHF_10_port, A_SHF_9_port, A_SHF_8_port, A_SHF_7_port, A_SHF_6_port, 
      A_SHF_5_port, A_SHF_4_port, A_SHF_3_port, A_SHF_2_port, A_SHF_1_port, 
      A_SHF_0_port, B_SHF_31_port, B_SHF_30_port, B_SHF_29_port, B_SHF_28_port,
      B_SHF_27_port, B_SHF_26_port, B_SHF_25_port, B_SHF_24_port, B_SHF_23_port
      , B_SHF_22_port, B_SHF_21_port, B_SHF_20_port, B_SHF_19_port, 
      B_SHF_18_port, B_SHF_17_port, B_SHF_16_port, B_SHF_15_port, B_SHF_14_port
      , B_SHF_13_port, B_SHF_12_port, B_SHF_11_port, B_SHF_10_port, 
      B_SHF_9_port, B_SHF_8_port, B_SHF_7_port, B_SHF_6_port, B_SHF_5_port, 
      B_SHF_4_port, B_SHF_3_port, B_SHF_2_port, B_SHF_1_port, B_SHF_0_port, 
      OPSel_2_port, OPSel_1_port, OPSel_0_port, A_CMP_31_port, A_CMP_30_port, 
      A_CMP_29_port, A_CMP_28_port, A_CMP_27_port, A_CMP_26_port, A_CMP_25_port
      , A_CMP_24_port, A_CMP_23_port, A_CMP_22_port, A_CMP_21_port, 
      A_CMP_20_port, A_CMP_19_port, A_CMP_18_port, A_CMP_17_port, A_CMP_16_port
      , A_CMP_15_port, A_CMP_14_port, A_CMP_13_port, A_CMP_12_port, 
      A_CMP_11_port, A_CMP_10_port, A_CMP_9_port, A_CMP_8_port, A_CMP_7_port, 
      A_CMP_6_port, A_CMP_5_port, A_CMP_4_port, A_CMP_3_port, A_CMP_2_port, 
      A_CMP_1_port, A_CMP_0_port, B_CMP_31_port, B_CMP_30_port, B_CMP_29_port, 
      B_CMP_28_port, B_CMP_27_port, B_CMP_26_port, B_CMP_25_port, B_CMP_24_port
      , B_CMP_23_port, B_CMP_22_port, B_CMP_21_port, B_CMP_20_port, 
      B_CMP_19_port, B_CMP_18_port, B_CMP_17_port, B_CMP_16_port, B_CMP_15_port
      , B_CMP_14_port, B_CMP_13_port, B_CMP_12_port, B_CMP_11_port, 
      B_CMP_10_port, B_CMP_9_port, B_CMP_8_port, B_CMP_7_port, B_CMP_6_port, 
      B_CMP_5_port, B_CMP_4_port, B_CMP_3_port, B_CMP_2_port, B_CMP_1_port, 
      B_CMP_0_port, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185,
      N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, 
      N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, 
      N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, 
      N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, 
      N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, 
      COMP_RES_0_port, ADD_SUB_RES_31_port, ADD_SUB_RES_30_port, 
      ADD_SUB_RES_29_port, ADD_SUB_RES_28_port, ADD_SUB_RES_27_port, 
      ADD_SUB_RES_26_port, ADD_SUB_RES_25_port, ADD_SUB_RES_24_port, 
      ADD_SUB_RES_23_port, ADD_SUB_RES_22_port, ADD_SUB_RES_21_port, 
      ADD_SUB_RES_20_port, ADD_SUB_RES_19_port, ADD_SUB_RES_18_port, 
      ADD_SUB_RES_17_port, ADD_SUB_RES_16_port, ADD_SUB_RES_15_port, 
      ADD_SUB_RES_14_port, ADD_SUB_RES_13_port, ADD_SUB_RES_12_port, 
      ADD_SUB_RES_11_port, ADD_SUB_RES_10_port, ADD_SUB_RES_9_port, 
      ADD_SUB_RES_8_port, ADD_SUB_RES_7_port, ADD_SUB_RES_6_port, 
      ADD_SUB_RES_5_port, ADD_SUB_RES_4_port, ADD_SUB_RES_3_port, 
      ADD_SUB_RES_2_port, ADD_SUB_RES_1_port, ADD_SUB_RES_0_port, n149, n71, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, sig_intraMux_9_port
      , sig_intraMux_8_port, sig_intraMux_7_port, sig_intraMux_6_port, 
      sig_intraMux_5_port, sig_intraMux_4_port, sig_intraMux_3_port, 
      sig_intraMux_31_port, sig_intraMux_30_port, sig_intraMux_2_port, 
      sig_intraMux_29_port, sig_intraMux_28_port, sig_intraMux_27_port, 
      sig_intraMux_26_port, sig_intraMux_25_port, sig_intraMux_24_port, 
      sig_intraMux_23_port, sig_intraMux_22_port, sig_intraMux_21_port, 
      sig_intraMux_20_port, sig_intraMux_1_port, sig_intraMux_19_port, 
      sig_intraMux_18_port, sig_intraMux_17_port, sig_intraMux_16_port, 
      sig_intraMux_15_port, sig_intraMux_14_port, sig_intraMux_13_port, 
      sig_intraMux_12_port, sig_intraMux_11_port, sig_intraMux_10_port, 
      sig_intraMux_0_port, SHIFT_RES_9_port, SHIFT_RES_8_port, SHIFT_RES_7_port
      , SHIFT_RES_6_port, SHIFT_RES_5_port, SHIFT_RES_4_port, SHIFT_RES_3_port,
      SHIFT_RES_31_port, SHIFT_RES_30_port, SHIFT_RES_2_port, SHIFT_RES_29_port
      , SHIFT_RES_28_port, SHIFT_RES_27_port, SHIFT_RES_26_port, 
      SHIFT_RES_25_port, SHIFT_RES_24_port, SHIFT_RES_23_port, 
      SHIFT_RES_22_port, SHIFT_RES_21_port, SHIFT_RES_20_port, SHIFT_RES_1_port
      , SHIFT_RES_19_port, SHIFT_RES_18_port, SHIFT_RES_17_port, 
      SHIFT_RES_16_port, SHIFT_RES_15_port, SHIFT_RES_14_port, 
      SHIFT_RES_13_port, SHIFT_RES_12_port, SHIFT_RES_11_port, 
      SHIFT_RES_10_port, SHIFT_RES_0_port, n184_port, n185_port, n186_port, 
      n187_port, n188_port, n189_port, n190_port, n191_port, n192_port, 
      n193_port, n194_port, n195_port, n196_port, n197_port, n198_port, 
      n199_port, n200_port, n201_port, n202_port, n203_port, n204_port, 
      n205_port, n206_port, n207_port, n208_port, n209_port, n210_port, 
      n211_port, n212_port, n213_port, n214_port, n215_port, n216_port, 
      n217_port, n218_port, n219_port, n220_port, n221_port, n222_port, 
      n223_port, n224_port, n225_port, n226_port, n227_port, n228_port, 
      n229_port, n230_port, n231_port, n232_port, n233_port, n234_port, 
      n235_port, n236_port, n237_port, n238_port, n239_port, n240_port, 
      n241_port, n242_port, n243_port, n244_port, n245_port, n246, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
      n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, 
      n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, 
      n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, 
      n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, 
      n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, 
      n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, 
      n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, 
      n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, 
      n_1099, n_1100, n_1101, n_1102, n_1103 : std_logic;

begin
   
   B_CMP_reg_31_inst : DLH_X1 port map( G => n203_port, D => OP2(31), Q => 
                           B_CMP_31_port);
   B_CMP_reg_30_inst : DLH_X1 port map( G => n203_port, D => OP2(30), Q => 
                           B_CMP_30_port);
   B_CMP_reg_29_inst : DLH_X1 port map( G => n203_port, D => OP2(29), Q => 
                           B_CMP_29_port);
   B_CMP_reg_28_inst : DLH_X1 port map( G => n203_port, D => OP2(28), Q => 
                           B_CMP_28_port);
   B_CMP_reg_27_inst : DLH_X1 port map( G => n203_port, D => OP2(27), Q => 
                           B_CMP_27_port);
   B_CMP_reg_26_inst : DLH_X1 port map( G => n203_port, D => OP2(26), Q => 
                           B_CMP_26_port);
   B_CMP_reg_25_inst : DLH_X1 port map( G => n203_port, D => OP2(25), Q => 
                           B_CMP_25_port);
   B_CMP_reg_24_inst : DLH_X1 port map( G => n203_port, D => OP2(24), Q => 
                           B_CMP_24_port);
   B_CMP_reg_23_inst : DLH_X1 port map( G => n203_port, D => OP2(23), Q => 
                           B_CMP_23_port);
   B_CMP_reg_22_inst : DLH_X1 port map( G => n203_port, D => OP2(22), Q => 
                           B_CMP_22_port);
   B_CMP_reg_21_inst : DLH_X1 port map( G => n203_port, D => OP2(21), Q => 
                           B_CMP_21_port);
   B_CMP_reg_20_inst : DLH_X1 port map( G => n203_port, D => OP2(20), Q => 
                           B_CMP_20_port);
   B_CMP_reg_19_inst : DLH_X1 port map( G => n203_port, D => OP2(19), Q => 
                           B_CMP_19_port);
   B_CMP_reg_18_inst : DLH_X1 port map( G => n207_port, D => OP2(18), Q => 
                           B_CMP_18_port);
   B_CMP_reg_17_inst : DLH_X1 port map( G => n207_port, D => OP2(17), Q => 
                           B_CMP_17_port);
   B_CMP_reg_16_inst : DLH_X1 port map( G => n207_port, D => OP2(16), Q => 
                           B_CMP_16_port);
   B_CMP_reg_15_inst : DLH_X1 port map( G => n207_port, D => OP2(15), Q => 
                           B_CMP_15_port);
   B_CMP_reg_14_inst : DLH_X1 port map( G => n207_port, D => OP2(14), Q => 
                           B_CMP_14_port);
   B_CMP_reg_13_inst : DLH_X1 port map( G => n206_port, D => OP2(13), Q => 
                           B_CMP_13_port);
   B_CMP_reg_12_inst : DLH_X1 port map( G => n206_port, D => OP2(12), Q => 
                           B_CMP_12_port);
   B_CMP_reg_11_inst : DLH_X1 port map( G => n206_port, D => OP2(11), Q => 
                           B_CMP_11_port);
   B_CMP_reg_10_inst : DLH_X1 port map( G => n206_port, D => OP2(10), Q => 
                           B_CMP_10_port);
   B_CMP_reg_9_inst : DLH_X1 port map( G => n206_port, D => OP2(9), Q => 
                           B_CMP_9_port);
   B_CMP_reg_8_inst : DLH_X1 port map( G => n206_port, D => OP2(8), Q => 
                           B_CMP_8_port);
   B_CMP_reg_7_inst : DLH_X1 port map( G => n206_port, D => OP2(7), Q => 
                           B_CMP_7_port);
   B_CMP_reg_6_inst : DLH_X1 port map( G => n206_port, D => OP2(6), Q => 
                           B_CMP_6_port);
   B_CMP_reg_5_inst : DLH_X1 port map( G => n206_port, D => OP2(5), Q => 
                           B_CMP_5_port);
   B_CMP_reg_4_inst : DLH_X1 port map( G => n206_port, D => OP2(4), Q => 
                           B_CMP_4_port);
   B_CMP_reg_3_inst : DLH_X1 port map( G => n206_port, D => OP2(3), Q => 
                           B_CMP_3_port);
   B_CMP_reg_2_inst : DLH_X1 port map( G => n205_port, D => OP2(2), Q => 
                           B_CMP_2_port);
   B_CMP_reg_1_inst : DLH_X1 port map( G => n205_port, D => OP2(1), Q => 
                           B_CMP_1_port);
   B_CMP_reg_0_inst : DLH_X1 port map( G => n205_port, D => OP2(0), Q => 
                           B_CMP_0_port);
   select_zero_sig_reg : DLH_X1 port map( G => N176, D => N177, Q => 
                           select_zero_sig);
   ADD_SUB_reg : DLH_X1 port map( G => n215_port, D => n184_port, Q => ADD_SUB)
                           ;
   A_ADD_reg_31_inst : DLH_X1 port map( G => n215_port, D => OP1(31), Q => 
                           A_ADD_31_port);
   A_ADD_reg_30_inst : DLH_X1 port map( G => n215_port, D => OP1(30), Q => 
                           A_ADD_30_port);
   A_ADD_reg_29_inst : DLH_X1 port map( G => n215_port, D => OP1(29), Q => 
                           A_ADD_29_port);
   A_ADD_reg_28_inst : DLH_X1 port map( G => n215_port, D => OP1(28), Q => 
                           A_ADD_28_port);
   A_ADD_reg_27_inst : DLH_X1 port map( G => n215_port, D => OP1(27), Q => 
                           A_ADD_27_port);
   A_ADD_reg_26_inst : DLH_X1 port map( G => n215_port, D => OP1(26), Q => 
                           A_ADD_26_port);
   A_ADD_reg_25_inst : DLH_X1 port map( G => n215_port, D => OP1(25), Q => 
                           A_ADD_25_port);
   A_ADD_reg_24_inst : DLH_X1 port map( G => n215_port, D => OP1(24), Q => 
                           A_ADD_24_port);
   A_ADD_reg_23_inst : DLH_X1 port map( G => n215_port, D => OP1(23), Q => 
                           A_ADD_23_port);
   A_ADD_reg_22_inst : DLH_X1 port map( G => n215_port, D => OP1(22), Q => 
                           A_ADD_22_port);
   A_ADD_reg_21_inst : DLH_X1 port map( G => n215_port, D => OP1(21), Q => 
                           A_ADD_21_port);
   A_ADD_reg_20_inst : DLH_X1 port map( G => n215_port, D => OP1(20), Q => 
                           A_ADD_20_port);
   A_ADD_reg_19_inst : DLH_X1 port map( G => n215_port, D => OP1(19), Q => 
                           A_ADD_19_port);
   A_ADD_reg_18_inst : DLH_X1 port map( G => n219_port, D => OP1(18), Q => 
                           A_ADD_18_port);
   A_ADD_reg_17_inst : DLH_X1 port map( G => n218_port, D => OP1(17), Q => 
                           A_ADD_17_port);
   A_ADD_reg_16_inst : DLH_X1 port map( G => n218_port, D => OP1(16), Q => 
                           A_ADD_16_port);
   A_ADD_reg_15_inst : DLH_X1 port map( G => n218_port, D => OP1(15), Q => 
                           A_ADD_15_port);
   A_ADD_reg_14_inst : DLH_X1 port map( G => n218_port, D => OP1(14), Q => 
                           A_ADD_14_port);
   A_ADD_reg_13_inst : DLH_X1 port map( G => n218_port, D => OP1(13), Q => 
                           A_ADD_13_port);
   A_ADD_reg_12_inst : DLH_X1 port map( G => n218_port, D => OP1(12), Q => 
                           A_ADD_12_port);
   A_ADD_reg_11_inst : DLH_X1 port map( G => n218_port, D => OP1(11), Q => 
                           A_ADD_11_port);
   A_ADD_reg_10_inst : DLH_X1 port map( G => n218_port, D => OP1(10), Q => 
                           A_ADD_10_port);
   A_ADD_reg_9_inst : DLH_X1 port map( G => n218_port, D => OP1(9), Q => 
                           A_ADD_9_port);
   A_ADD_reg_8_inst : DLH_X1 port map( G => n218_port, D => OP1(8), Q => 
                           A_ADD_8_port);
   A_ADD_reg_7_inst : DLH_X1 port map( G => n218_port, D => OP1(7), Q => 
                           A_ADD_7_port);
   A_ADD_reg_6_inst : DLH_X1 port map( G => n218_port, D => OP1(6), Q => 
                           A_ADD_6_port);
   A_ADD_reg_5_inst : DLH_X1 port map( G => n218_port, D => OP1(5), Q => 
                           A_ADD_5_port);
   A_ADD_reg_4_inst : DLH_X1 port map( G => n218_port, D => OP1(4), Q => 
                           A_ADD_4_port);
   A_ADD_reg_3_inst : DLH_X1 port map( G => n219_port, D => OP1(3), Q => 
                           A_ADD_3_port);
   A_ADD_reg_2_inst : DLH_X1 port map( G => n217_port, D => OP1(2), Q => 
                           A_ADD_2_port);
   A_ADD_reg_1_inst : DLH_X1 port map( G => n217_port, D => OP1(1), Q => 
                           A_ADD_1_port);
   A_ADD_reg_0_inst : DLH_X1 port map( G => n217_port, D => OP1(0), Q => 
                           A_ADD_0_port);
   B_ADD_reg_31_inst : DLH_X1 port map( G => n218_port, D => N210, Q => 
                           B_ADD_31_port);
   B_ADD_reg_30_inst : DLH_X1 port map( G => n218_port, D => N209, Q => 
                           B_ADD_30_port);
   B_ADD_reg_29_inst : DLH_X1 port map( G => n217_port, D => N208, Q => 
                           B_ADD_29_port);
   B_ADD_reg_28_inst : DLH_X1 port map( G => n217_port, D => N207, Q => 
                           B_ADD_28_port);
   B_ADD_reg_27_inst : DLH_X1 port map( G => n217_port, D => N206, Q => 
                           B_ADD_27_port);
   B_ADD_reg_26_inst : DLH_X1 port map( G => n217_port, D => N205, Q => 
                           B_ADD_26_port);
   B_ADD_reg_25_inst : DLH_X1 port map( G => n217_port, D => N204, Q => 
                           B_ADD_25_port);
   B_ADD_reg_24_inst : DLH_X1 port map( G => n217_port, D => N203, Q => 
                           B_ADD_24_port);
   B_ADD_reg_23_inst : DLH_X1 port map( G => n217_port, D => N202, Q => 
                           B_ADD_23_port);
   B_ADD_reg_22_inst : DLH_X1 port map( G => n217_port, D => N201, Q => 
                           B_ADD_22_port);
   B_ADD_reg_21_inst : DLH_X1 port map( G => n217_port, D => N200, Q => 
                           B_ADD_21_port);
   B_ADD_reg_20_inst : DLH_X1 port map( G => n217_port, D => N199, Q => 
                           B_ADD_20_port);
   B_ADD_reg_19_inst : DLH_X1 port map( G => n217_port, D => N198, Q => 
                           B_ADD_19_port);
   B_ADD_reg_18_inst : DLH_X1 port map( G => n217_port, D => N197, Q => 
                           B_ADD_18_port);
   B_ADD_reg_17_inst : DLH_X1 port map( G => n217_port, D => N196, Q => 
                           B_ADD_17_port);
   B_ADD_reg_16_inst : DLH_X1 port map( G => n216_port, D => N195, Q => 
                           B_ADD_16_port);
   B_ADD_reg_15_inst : DLH_X1 port map( G => n216_port, D => N194, Q => 
                           B_ADD_15_port);
   B_ADD_reg_14_inst : DLH_X1 port map( G => n216_port, D => N193, Q => 
                           B_ADD_14_port);
   B_ADD_reg_13_inst : DLH_X1 port map( G => n216_port, D => N192, Q => 
                           B_ADD_13_port);
   B_ADD_reg_12_inst : DLH_X1 port map( G => n216_port, D => N191, Q => 
                           B_ADD_12_port);
   B_ADD_reg_11_inst : DLH_X1 port map( G => n216_port, D => N190, Q => 
                           B_ADD_11_port);
   B_ADD_reg_10_inst : DLH_X1 port map( G => n216_port, D => N189, Q => 
                           B_ADD_10_port);
   B_ADD_reg_9_inst : DLH_X1 port map( G => n216_port, D => N188, Q => 
                           B_ADD_9_port);
   B_ADD_reg_8_inst : DLH_X1 port map( G => n216_port, D => N187, Q => 
                           B_ADD_8_port);
   B_ADD_reg_7_inst : DLH_X1 port map( G => n216_port, D => N186, Q => 
                           B_ADD_7_port);
   B_ADD_reg_6_inst : DLH_X1 port map( G => n216_port, D => N185, Q => 
                           B_ADD_6_port);
   B_ADD_reg_5_inst : DLH_X1 port map( G => n216_port, D => N184, Q => 
                           B_ADD_5_port);
   B_ADD_reg_4_inst : DLH_X1 port map( G => n216_port, D => N183, Q => 
                           B_ADD_4_port);
   B_ADD_reg_3_inst : DLH_X1 port map( G => n216_port, D => N182, Q => 
                           B_ADD_3_port);
   B_ADD_reg_2_inst : DLH_X1 port map( G => n216_port, D => N181, Q => 
                           B_ADD_2_port);
   B_ADD_reg_1_inst : DLH_X1 port map( G => n216_port, D => N180, Q => 
                           B_ADD_1_port);
   B_ADD_reg_0_inst : DLH_X1 port map( G => n215_port, D => N179, Q => 
                           B_ADD_0_port);
   LOGIC_RES_reg_31_inst : DLH_X1 port map( G => n213_port, D => N243, Q => 
                           LOGIC_RES_31_port);
   LOGIC_RES_reg_30_inst : DLH_X1 port map( G => n213_port, D => N242, Q => 
                           LOGIC_RES_30_port);
   LOGIC_RES_reg_29_inst : DLH_X1 port map( G => n213_port, D => N241, Q => 
                           LOGIC_RES_29_port);
   LOGIC_RES_reg_28_inst : DLH_X1 port map( G => n213_port, D => N240, Q => 
                           LOGIC_RES_28_port);
   LOGIC_RES_reg_27_inst : DLH_X1 port map( G => n213_port, D => N239, Q => 
                           LOGIC_RES_27_port);
   LOGIC_RES_reg_26_inst : DLH_X1 port map( G => n213_port, D => N238, Q => 
                           LOGIC_RES_26_port);
   LOGIC_RES_reg_25_inst : DLH_X1 port map( G => n213_port, D => N237, Q => 
                           LOGIC_RES_25_port);
   LOGIC_RES_reg_24_inst : DLH_X1 port map( G => n213_port, D => N236, Q => 
                           LOGIC_RES_24_port);
   LOGIC_RES_reg_23_inst : DLH_X1 port map( G => n213_port, D => N235, Q => 
                           LOGIC_RES_23_port);
   LOGIC_RES_reg_22_inst : DLH_X1 port map( G => n213_port, D => N234, Q => 
                           LOGIC_RES_22_port);
   LOGIC_RES_reg_21_inst : DLH_X1 port map( G => n213_port, D => N233, Q => 
                           LOGIC_RES_21_port);
   LOGIC_RES_reg_20_inst : DLH_X1 port map( G => n213_port, D => N232, Q => 
                           LOGIC_RES_20_port);
   LOGIC_RES_reg_19_inst : DLH_X1 port map( G => n213_port, D => N231, Q => 
                           LOGIC_RES_19_port);
   LOGIC_RES_reg_18_inst : DLH_X1 port map( G => n213_port, D => N230, Q => 
                           LOGIC_RES_18_port);
   LOGIC_RES_reg_17_inst : DLH_X1 port map( G => n213_port, D => N229, Q => 
                           LOGIC_RES_17_port);
   LOGIC_RES_reg_16_inst : DLH_X1 port map( G => n214_port, D => N228, Q => 
                           LOGIC_RES_16_port);
   LOGIC_RES_reg_15_inst : DLH_X1 port map( G => n214_port, D => N227, Q => 
                           LOGIC_RES_15_port);
   LOGIC_RES_reg_14_inst : DLH_X1 port map( G => n214_port, D => N226, Q => 
                           LOGIC_RES_14_port);
   LOGIC_RES_reg_13_inst : DLH_X1 port map( G => n214_port, D => N225, Q => 
                           LOGIC_RES_13_port);
   LOGIC_RES_reg_12_inst : DLH_X1 port map( G => n214_port, D => N224, Q => 
                           LOGIC_RES_12_port);
   LOGIC_RES_reg_11_inst : DLH_X1 port map( G => n214_port, D => N223, Q => 
                           LOGIC_RES_11_port);
   LOGIC_RES_reg_10_inst : DLH_X1 port map( G => n214_port, D => N222, Q => 
                           LOGIC_RES_10_port);
   LOGIC_RES_reg_9_inst : DLH_X1 port map( G => n214_port, D => N221, Q => 
                           LOGIC_RES_9_port);
   LOGIC_RES_reg_8_inst : DLH_X1 port map( G => n214_port, D => N220, Q => 
                           LOGIC_RES_8_port);
   LOGIC_RES_reg_7_inst : DLH_X1 port map( G => n214_port, D => N219, Q => 
                           LOGIC_RES_7_port);
   LOGIC_RES_reg_6_inst : DLH_X1 port map( G => n214_port, D => N218, Q => 
                           LOGIC_RES_6_port);
   LOGIC_RES_reg_5_inst : DLH_X1 port map( G => n214_port, D => N217, Q => 
                           LOGIC_RES_5_port);
   LOGIC_RES_reg_4_inst : DLH_X1 port map( G => n214_port, D => N216, Q => 
                           LOGIC_RES_4_port);
   LOGIC_RES_reg_3_inst : DLH_X1 port map( G => n214_port, D => N215, Q => 
                           LOGIC_RES_3_port);
   LOGIC_RES_reg_2_inst : DLH_X1 port map( G => n214_port, D => N214, Q => 
                           LOGIC_RES_2_port);
   LOGIC_RES_reg_1_inst : DLH_X1 port map( G => n214_port, D => N213, Q => 
                           LOGIC_RES_1_port);
   LOGIC_RES_reg_0_inst : DLH_X1 port map( G => N211, D => N212, Q => 
                           LOGIC_RES_0_port);
   LEFT_RIGHT_reg : DLH_X1 port map( G => n208_port, D => n149, Q => LEFT_RIGHT
                           );
   A_SHF_reg_31_inst : DLH_X1 port map( G => n211_port, D => OP1(31), Q => 
                           A_SHF_31_port);
   A_SHF_reg_30_inst : DLH_X1 port map( G => n211_port, D => OP1(30), Q => 
                           A_SHF_30_port);
   A_SHF_reg_29_inst : DLH_X1 port map( G => n211_port, D => OP1(29), Q => 
                           A_SHF_29_port);
   A_SHF_reg_28_inst : DLH_X1 port map( G => n211_port, D => OP1(28), Q => 
                           A_SHF_28_port);
   A_SHF_reg_27_inst : DLH_X1 port map( G => n211_port, D => OP1(27), Q => 
                           A_SHF_27_port);
   A_SHF_reg_26_inst : DLH_X1 port map( G => n211_port, D => OP1(26), Q => 
                           A_SHF_26_port);
   A_SHF_reg_25_inst : DLH_X1 port map( G => n211_port, D => OP1(25), Q => 
                           A_SHF_25_port);
   A_SHF_reg_24_inst : DLH_X1 port map( G => n211_port, D => OP1(24), Q => 
                           A_SHF_24_port);
   A_SHF_reg_23_inst : DLH_X1 port map( G => n211_port, D => OP1(23), Q => 
                           A_SHF_23_port);
   A_SHF_reg_22_inst : DLH_X1 port map( G => n211_port, D => OP1(22), Q => 
                           A_SHF_22_port);
   A_SHF_reg_21_inst : DLH_X1 port map( G => n211_port, D => OP1(21), Q => 
                           A_SHF_21_port);
   A_SHF_reg_20_inst : DLH_X1 port map( G => n212_port, D => OP1(20), Q => 
                           A_SHF_20_port);
   A_SHF_reg_19_inst : DLH_X1 port map( G => n212_port, D => OP1(19), Q => 
                           A_SHF_19_port);
   A_SHF_reg_18_inst : DLH_X1 port map( G => n212_port, D => OP1(18), Q => 
                           A_SHF_18_port);
   A_SHF_reg_17_inst : DLH_X1 port map( G => n210_port, D => OP1(17), Q => 
                           A_SHF_17_port);
   A_SHF_reg_16_inst : DLH_X1 port map( G => n208_port, D => OP1(16), Q => 
                           A_SHF_16_port);
   A_SHF_reg_15_inst : DLH_X1 port map( G => n208_port, D => OP1(15), Q => 
                           A_SHF_15_port);
   A_SHF_reg_14_inst : DLH_X1 port map( G => n208_port, D => OP1(14), Q => 
                           A_SHF_14_port);
   A_SHF_reg_13_inst : DLH_X1 port map( G => n208_port, D => OP1(13), Q => 
                           A_SHF_13_port);
   A_SHF_reg_12_inst : DLH_X1 port map( G => n208_port, D => OP1(12), Q => 
                           A_SHF_12_port);
   A_SHF_reg_11_inst : DLH_X1 port map( G => n208_port, D => OP1(11), Q => 
                           A_SHF_11_port);
   A_SHF_reg_10_inst : DLH_X1 port map( G => n208_port, D => OP1(10), Q => 
                           A_SHF_10_port);
   A_SHF_reg_9_inst : DLH_X1 port map( G => n208_port, D => OP1(9), Q => 
                           A_SHF_9_port);
   A_SHF_reg_8_inst : DLH_X1 port map( G => n208_port, D => OP1(8), Q => 
                           A_SHF_8_port);
   A_SHF_reg_7_inst : DLH_X1 port map( G => n208_port, D => OP1(7), Q => 
                           A_SHF_7_port);
   A_SHF_reg_6_inst : DLH_X1 port map( G => n208_port, D => OP1(6), Q => 
                           A_SHF_6_port);
   A_SHF_reg_5_inst : DLH_X1 port map( G => n208_port, D => OP1(5), Q => 
                           A_SHF_5_port);
   A_SHF_reg_4_inst : DLH_X1 port map( G => n208_port, D => OP1(4), Q => 
                           A_SHF_4_port);
   A_SHF_reg_3_inst : DLH_X1 port map( G => n209_port, D => OP1(3), Q => 
                           A_SHF_3_port);
   A_SHF_reg_2_inst : DLH_X1 port map( G => n209_port, D => OP1(2), Q => 
                           A_SHF_2_port);
   A_SHF_reg_1_inst : DLH_X1 port map( G => n210_port, D => OP1(1), Q => 
                           A_SHF_1_port);
   A_SHF_reg_0_inst : DLH_X1 port map( G => n210_port, D => OP1(0), Q => 
                           A_SHF_0_port);
   B_SHF_reg_31_inst : DLH_X1 port map( G => n209_port, D => OP2(31), Q => 
                           B_SHF_31_port);
   B_SHF_reg_30_inst : DLH_X1 port map( G => n209_port, D => OP2(30), Q => 
                           B_SHF_30_port);
   B_SHF_reg_29_inst : DLH_X1 port map( G => n209_port, D => OP2(29), Q => 
                           B_SHF_29_port);
   B_SHF_reg_28_inst : DLH_X1 port map( G => n209_port, D => OP2(28), Q => 
                           B_SHF_28_port);
   B_SHF_reg_27_inst : DLH_X1 port map( G => n209_port, D => OP2(27), Q => 
                           B_SHF_27_port);
   B_SHF_reg_26_inst : DLH_X1 port map( G => n209_port, D => OP2(26), Q => 
                           B_SHF_26_port);
   B_SHF_reg_25_inst : DLH_X1 port map( G => n209_port, D => OP2(25), Q => 
                           B_SHF_25_port);
   B_SHF_reg_24_inst : DLH_X1 port map( G => n209_port, D => OP2(24), Q => 
                           B_SHF_24_port);
   B_SHF_reg_23_inst : DLH_X1 port map( G => n209_port, D => OP2(23), Q => 
                           B_SHF_23_port);
   B_SHF_reg_22_inst : DLH_X1 port map( G => n209_port, D => OP2(22), Q => 
                           B_SHF_22_port);
   B_SHF_reg_21_inst : DLH_X1 port map( G => n209_port, D => OP2(21), Q => 
                           B_SHF_21_port);
   B_SHF_reg_20_inst : DLH_X1 port map( G => n209_port, D => OP2(20), Q => 
                           B_SHF_20_port);
   B_SHF_reg_19_inst : DLH_X1 port map( G => n209_port, D => OP2(19), Q => 
                           B_SHF_19_port);
   B_SHF_reg_18_inst : DLH_X1 port map( G => n209_port, D => OP2(18), Q => 
                           B_SHF_18_port);
   B_SHF_reg_17_inst : DLH_X1 port map( G => n210_port, D => OP2(17), Q => 
                           B_SHF_17_port);
   B_SHF_reg_16_inst : DLH_X1 port map( G => n210_port, D => OP2(16), Q => 
                           B_SHF_16_port);
   B_SHF_reg_15_inst : DLH_X1 port map( G => n210_port, D => OP2(15), Q => 
                           B_SHF_15_port);
   B_SHF_reg_14_inst : DLH_X1 port map( G => n210_port, D => OP2(14), Q => 
                           B_SHF_14_port);
   B_SHF_reg_13_inst : DLH_X1 port map( G => n210_port, D => OP2(13), Q => 
                           B_SHF_13_port);
   B_SHF_reg_12_inst : DLH_X1 port map( G => n210_port, D => OP2(12), Q => 
                           B_SHF_12_port);
   B_SHF_reg_11_inst : DLH_X1 port map( G => n210_port, D => OP2(11), Q => 
                           B_SHF_11_port);
   B_SHF_reg_10_inst : DLH_X1 port map( G => n210_port, D => OP2(10), Q => 
                           B_SHF_10_port);
   B_SHF_reg_9_inst : DLH_X1 port map( G => n210_port, D => OP2(9), Q => 
                           B_SHF_9_port);
   B_SHF_reg_8_inst : DLH_X1 port map( G => n210_port, D => OP2(8), Q => 
                           B_SHF_8_port);
   B_SHF_reg_7_inst : DLH_X1 port map( G => n211_port, D => OP2(7), Q => 
                           B_SHF_7_port);
   B_SHF_reg_6_inst : DLH_X1 port map( G => n210_port, D => OP2(6), Q => 
                           B_SHF_6_port);
   B_SHF_reg_5_inst : DLH_X1 port map( G => n210_port, D => OP2(5), Q => 
                           B_SHF_5_port);
   B_SHF_reg_4_inst : DLH_X1 port map( G => n210_port, D => OP2(4), Q => 
                           B_SHF_4_port);
   B_SHF_reg_3_inst : DLH_X1 port map( G => n211_port, D => OP2(3), Q => 
                           B_SHF_3_port);
   B_SHF_reg_2_inst : DLH_X1 port map( G => n211_port, D => OP2(2), Q => 
                           B_SHF_2_port);
   B_SHF_reg_1_inst : DLH_X1 port map( G => n211_port, D => OP2(1), Q => 
                           B_SHF_1_port);
   B_SHF_reg_0_inst : DLH_X1 port map( G => n211_port, D => OP2(0), Q => 
                           B_SHF_0_port);
   OPSel_reg_2_inst : DLH_X1 port map( G => n205_port, D => n146, Q => 
                           OPSel_2_port);
   OPSel_reg_1_inst : DLH_X1 port map( G => n205_port, D => n145, Q => 
                           OPSel_1_port);
   A_CMP_reg_31_inst : DLH_X1 port map( G => n206_port, D => OP1(31), Q => 
                           A_CMP_31_port);
   A_CMP_reg_30_inst : DLH_X1 port map( G => n206_port, D => OP1(30), Q => 
                           A_CMP_30_port);
   A_CMP_reg_29_inst : DLH_X1 port map( G => n206_port, D => OP1(29), Q => 
                           A_CMP_29_port);
   A_CMP_reg_28_inst : DLH_X1 port map( G => n206_port, D => OP1(28), Q => 
                           A_CMP_28_port);
   A_CMP_reg_27_inst : DLH_X1 port map( G => n206_port, D => OP1(27), Q => 
                           A_CMP_27_port);
   A_CMP_reg_26_inst : DLH_X1 port map( G => n205_port, D => OP1(26), Q => 
                           A_CMP_26_port);
   A_CMP_reg_25_inst : DLH_X1 port map( G => n205_port, D => OP1(25), Q => 
                           A_CMP_25_port);
   A_CMP_reg_24_inst : DLH_X1 port map( G => n205_port, D => OP1(24), Q => 
                           A_CMP_24_port);
   A_CMP_reg_23_inst : DLH_X1 port map( G => n205_port, D => OP1(23), Q => 
                           A_CMP_23_port);
   A_CMP_reg_22_inst : DLH_X1 port map( G => n205_port, D => OP1(22), Q => 
                           A_CMP_22_port);
   A_CMP_reg_21_inst : DLH_X1 port map( G => n205_port, D => OP1(21), Q => 
                           A_CMP_21_port);
   A_CMP_reg_20_inst : DLH_X1 port map( G => n205_port, D => OP1(20), Q => 
                           A_CMP_20_port);
   A_CMP_reg_19_inst : DLH_X1 port map( G => n205_port, D => OP1(19), Q => 
                           A_CMP_19_port);
   A_CMP_reg_18_inst : DLH_X1 port map( G => n205_port, D => OP1(18), Q => 
                           A_CMP_18_port);
   A_CMP_reg_17_inst : DLH_X1 port map( G => n205_port, D => OP1(17), Q => 
                           A_CMP_17_port);
   A_CMP_reg_16_inst : DLH_X1 port map( G => n205_port, D => OP1(16), Q => 
                           A_CMP_16_port);
   A_CMP_reg_15_inst : DLH_X1 port map( G => n204_port, D => OP1(15), Q => 
                           A_CMP_15_port);
   A_CMP_reg_14_inst : DLH_X1 port map( G => n204_port, D => OP1(14), Q => 
                           A_CMP_14_port);
   A_CMP_reg_13_inst : DLH_X1 port map( G => n204_port, D => OP1(13), Q => 
                           A_CMP_13_port);
   A_CMP_reg_12_inst : DLH_X1 port map( G => n204_port, D => OP1(12), Q => 
                           A_CMP_12_port);
   A_CMP_reg_11_inst : DLH_X1 port map( G => n204_port, D => OP1(11), Q => 
                           A_CMP_11_port);
   A_CMP_reg_10_inst : DLH_X1 port map( G => n204_port, D => OP1(10), Q => 
                           A_CMP_10_port);
   A_CMP_reg_9_inst : DLH_X1 port map( G => n204_port, D => OP1(9), Q => 
                           A_CMP_9_port);
   A_CMP_reg_8_inst : DLH_X1 port map( G => n204_port, D => OP1(8), Q => 
                           A_CMP_8_port);
   A_CMP_reg_7_inst : DLH_X1 port map( G => n204_port, D => OP1(7), Q => 
                           A_CMP_7_port);
   A_CMP_reg_6_inst : DLH_X1 port map( G => n204_port, D => OP1(6), Q => 
                           A_CMP_6_port);
   A_CMP_reg_5_inst : DLH_X1 port map( G => n204_port, D => OP1(5), Q => 
                           A_CMP_5_port);
   A_CMP_reg_4_inst : DLH_X1 port map( G => n204_port, D => OP1(4), Q => 
                           A_CMP_4_port);
   A_CMP_reg_3_inst : DLH_X1 port map( G => n204_port, D => OP1(3), Q => 
                           A_CMP_3_port);
   A_CMP_reg_2_inst : DLH_X1 port map( G => n204_port, D => OP1(2), Q => 
                           A_CMP_2_port);
   A_CMP_reg_1_inst : DLH_X1 port map( G => n204_port, D => OP1(1), Q => 
                           A_CMP_1_port);
   A_CMP_reg_0_inst : DLH_X1 port map( G => n204_port, D => OP1(0), Q => 
                           A_CMP_0_port);
   OPSel_0_port <= '1';
   U188 : NAND3_X1 port map( A1 => n198_port, A2 => n284, A3 => OP2(31), ZN => 
                           n74);
   U189 : NAND3_X1 port map( A1 => n200_port, A2 => n283, A3 => OP2(30), ZN => 
                           n79);
   U190 : NAND3_X1 port map( A1 => n200_port, A2 => n282, A3 => OP2(29), ZN => 
                           n81);
   U191 : NAND3_X1 port map( A1 => n200_port, A2 => n281, A3 => OP2(28), ZN => 
                           n83);
   U192 : NAND3_X1 port map( A1 => n200_port, A2 => n280, A3 => OP2(27), ZN => 
                           n85);
   U193 : NAND3_X1 port map( A1 => n200_port, A2 => n279, A3 => OP2(26), ZN => 
                           n87);
   U194 : NAND3_X1 port map( A1 => n200_port, A2 => n278, A3 => OP2(25), ZN => 
                           n89);
   U195 : NAND3_X1 port map( A1 => n200_port, A2 => n277, A3 => OP2(24), ZN => 
                           n91);
   U196 : NAND3_X1 port map( A1 => n199_port, A2 => n276, A3 => OP2(23), ZN => 
                           n93);
   U197 : NAND3_X1 port map( A1 => n199_port, A2 => n275, A3 => OP2(22), ZN => 
                           n95);
   U198 : NAND3_X1 port map( A1 => n199_port, A2 => n274, A3 => OP2(21), ZN => 
                           n97);
   U199 : NAND3_X1 port map( A1 => n199_port, A2 => n273, A3 => OP2(20), ZN => 
                           n99);
   U200 : NAND3_X1 port map( A1 => n199_port, A2 => n272, A3 => OP2(19), ZN => 
                           n101);
   U201 : NAND3_X1 port map( A1 => n199_port, A2 => n271, A3 => OP2(18), ZN => 
                           n103);
   U202 : NAND3_X1 port map( A1 => n199_port, A2 => n270, A3 => OP2(17), ZN => 
                           n105);
   U203 : NAND3_X1 port map( A1 => n199_port, A2 => n269, A3 => OP2(16), ZN => 
                           n107);
   U204 : NAND3_X1 port map( A1 => n199_port, A2 => n268, A3 => OP2(15), ZN => 
                           n109);
   U205 : NAND3_X1 port map( A1 => n199_port, A2 => n267, A3 => OP2(14), ZN => 
                           n111);
   U206 : NAND3_X1 port map( A1 => n199_port, A2 => n266, A3 => OP2(13), ZN => 
                           n113);
   U207 : NAND3_X1 port map( A1 => n199_port, A2 => n265, A3 => OP2(12), ZN => 
                           n115);
   U208 : NAND3_X1 port map( A1 => n199_port, A2 => n264, A3 => OP2(11), ZN => 
                           n117);
   U209 : NAND3_X1 port map( A1 => n200_port, A2 => n263, A3 => OP2(10), ZN => 
                           n119);
   U210 : NAND3_X1 port map( A1 => n199_port, A2 => n262, A3 => OP2(9), ZN => 
                           n121);
   U211 : NAND3_X1 port map( A1 => n199_port, A2 => n261, A3 => OP2(8), ZN => 
                           n123);
   U212 : NAND3_X1 port map( A1 => n199_port, A2 => n260, A3 => OP2(7), ZN => 
                           n125);
   U213 : NAND3_X1 port map( A1 => n199_port, A2 => n259, A3 => OP2(6), ZN => 
                           n127);
   U214 : NAND3_X1 port map( A1 => n199_port, A2 => n258, A3 => OP2(5), ZN => 
                           n129);
   U215 : NAND3_X1 port map( A1 => n199_port, A2 => n257, A3 => OP2(4), ZN => 
                           n131);
   U216 : NAND3_X1 port map( A1 => n199_port, A2 => n256, A3 => OP2(3), ZN => 
                           n133);
   U217 : NAND3_X1 port map( A1 => n198_port, A2 => n255, A3 => OP2(2), ZN => 
                           n135);
   U218 : NAND3_X1 port map( A1 => n198_port, A2 => n254, A3 => OP2(1), ZN => 
                           n137);
   U219 : NAND3_X1 port map( A1 => n198_port, A2 => n253, A3 => OP2(0), ZN => 
                           n139);
   U220 : NAND3_X1 port map( A1 => ALU_OPC(2), A2 => n318, A3 => ALU_OPC(0), ZN
                           => n71);
   U221 : NAND3_X1 port map( A1 => n319, A2 => n318, A3 => n320, ZN => n144);
   Comp : comparator_NBIT32 port map( A(31) => A_CMP_31_port, A(30) => 
                           A_CMP_30_port, A(29) => A_CMP_29_port, A(28) => 
                           A_CMP_28_port, A(27) => A_CMP_27_port, A(26) => 
                           A_CMP_26_port, A(25) => A_CMP_25_port, A(24) => 
                           A_CMP_24_port, A(23) => A_CMP_23_port, A(22) => 
                           A_CMP_22_port, A(21) => A_CMP_21_port, A(20) => 
                           A_CMP_20_port, A(19) => A_CMP_19_port, A(18) => 
                           A_CMP_18_port, A(17) => A_CMP_17_port, A(16) => 
                           A_CMP_16_port, A(15) => A_CMP_15_port, A(14) => 
                           A_CMP_14_port, A(13) => A_CMP_13_port, A(12) => 
                           A_CMP_12_port, A(11) => A_CMP_11_port, A(10) => 
                           A_CMP_10_port, A(9) => A_CMP_9_port, A(8) => 
                           A_CMP_8_port, A(7) => A_CMP_7_port, A(6) => 
                           A_CMP_6_port, A(5) => A_CMP_5_port, A(4) => 
                           A_CMP_4_port, A(3) => A_CMP_3_port, A(2) => 
                           A_CMP_2_port, A(1) => A_CMP_1_port, A(0) => 
                           A_CMP_0_port, B(31) => B_CMP_31_port, B(30) => 
                           B_CMP_30_port, B(29) => B_CMP_29_port, B(28) => 
                           B_CMP_28_port, B(27) => B_CMP_27_port, B(26) => 
                           B_CMP_26_port, B(25) => B_CMP_25_port, B(24) => 
                           B_CMP_24_port, B(23) => B_CMP_23_port, B(22) => 
                           B_CMP_22_port, B(21) => B_CMP_21_port, B(20) => 
                           B_CMP_20_port, B(19) => B_CMP_19_port, B(18) => 
                           B_CMP_18_port, B(17) => B_CMP_17_port, B(16) => 
                           B_CMP_16_port, B(15) => B_CMP_15_port, B(14) => 
                           B_CMP_14_port, B(13) => B_CMP_13_port, B(12) => 
                           B_CMP_12_port, B(11) => B_CMP_11_port, B(10) => 
                           B_CMP_10_port, B(9) => B_CMP_9_port, B(8) => 
                           B_CMP_8_port, B(7) => B_CMP_7_port, B(6) => 
                           B_CMP_6_port, B(5) => B_CMP_5_port, B(4) => 
                           B_CMP_4_port, B(3) => B_CMP_3_port, B(2) => 
                           B_CMP_2_port, B(1) => B_CMP_1_port, B(0) => 
                           B_CMP_0_port, OPSel(0) => OPSel_2_port, OPSel(1) => 
                           OPSel_1_port, OPSel(2) => OPSel_0_port, RES(31) => 
                           n_1072, RES(30) => n_1073, RES(29) => n_1074, 
                           RES(28) => n_1075, RES(27) => n_1076, RES(26) => 
                           n_1077, RES(25) => n_1078, RES(24) => n_1079, 
                           RES(23) => n_1080, RES(22) => n_1081, RES(21) => 
                           n_1082, RES(20) => n_1083, RES(19) => n_1084, 
                           RES(18) => n_1085, RES(17) => n_1086, RES(16) => 
                           n_1087, RES(15) => n_1088, RES(14) => n_1089, 
                           RES(13) => n_1090, RES(12) => n_1091, RES(11) => 
                           n_1092, RES(10) => n_1093, RES(9) => n_1094, RES(8) 
                           => n_1095, RES(7) => n_1096, RES(6) => n_1097, 
                           RES(5) => n_1098, RES(4) => n_1099, RES(3) => n_1100
                           , RES(2) => n_1101, RES(1) => n_1102, RES(0) => 
                           COMP_RES_0_port);
   Shift : shifter port map( A(31) => A_SHF_31_port, A(30) => A_SHF_30_port, 
                           A(29) => A_SHF_29_port, A(28) => A_SHF_28_port, 
                           A(27) => A_SHF_27_port, A(26) => A_SHF_26_port, 
                           A(25) => A_SHF_25_port, A(24) => A_SHF_24_port, 
                           A(23) => A_SHF_23_port, A(22) => A_SHF_22_port, 
                           A(21) => A_SHF_21_port, A(20) => A_SHF_20_port, 
                           A(19) => A_SHF_19_port, A(18) => A_SHF_18_port, 
                           A(17) => A_SHF_17_port, A(16) => A_SHF_16_port, 
                           A(15) => A_SHF_15_port, A(14) => A_SHF_14_port, 
                           A(13) => A_SHF_13_port, A(12) => A_SHF_12_port, 
                           A(11) => A_SHF_11_port, A(10) => A_SHF_10_port, A(9)
                           => A_SHF_9_port, A(8) => A_SHF_8_port, A(7) => 
                           A_SHF_7_port, A(6) => A_SHF_6_port, A(5) => 
                           A_SHF_5_port, A(4) => A_SHF_4_port, A(3) => 
                           A_SHF_3_port, A(2) => A_SHF_2_port, A(1) => 
                           A_SHF_1_port, A(0) => A_SHF_0_port, B(31) => 
                           B_SHF_31_port, B(30) => B_SHF_30_port, B(29) => 
                           B_SHF_29_port, B(28) => B_SHF_28_port, B(27) => 
                           B_SHF_27_port, B(26) => B_SHF_26_port, B(25) => 
                           B_SHF_25_port, B(24) => B_SHF_24_port, B(23) => 
                           B_SHF_23_port, B(22) => B_SHF_22_port, B(21) => 
                           B_SHF_21_port, B(20) => B_SHF_20_port, B(19) => 
                           B_SHF_19_port, B(18) => B_SHF_18_port, B(17) => 
                           B_SHF_17_port, B(16) => B_SHF_16_port, B(15) => 
                           B_SHF_15_port, B(14) => B_SHF_14_port, B(13) => 
                           B_SHF_13_port, B(12) => B_SHF_12_port, B(11) => 
                           B_SHF_11_port, B(10) => B_SHF_10_port, B(9) => 
                           B_SHF_9_port, B(8) => B_SHF_8_port, B(7) => 
                           B_SHF_7_port, B(6) => B_SHF_6_port, B(5) => 
                           B_SHF_5_port, B(4) => B_SHF_4_port, B(3) => 
                           B_SHF_3_port, B(2) => B_SHF_2_port, B(1) => 
                           B_SHF_1_port, B(0) => B_SHF_0_port, LOGIC_ARITH => 
                           n252, LEFT_RIGHT => LEFT_RIGHT, RES(31) => 
                           SHIFT_RES_31_port, RES(30) => SHIFT_RES_30_port, 
                           RES(29) => SHIFT_RES_29_port, RES(28) => 
                           SHIFT_RES_28_port, RES(27) => SHIFT_RES_27_port, 
                           RES(26) => SHIFT_RES_26_port, RES(25) => 
                           SHIFT_RES_25_port, RES(24) => SHIFT_RES_24_port, 
                           RES(23) => SHIFT_RES_23_port, RES(22) => 
                           SHIFT_RES_22_port, RES(21) => SHIFT_RES_21_port, 
                           RES(20) => SHIFT_RES_20_port, RES(19) => 
                           SHIFT_RES_19_port, RES(18) => SHIFT_RES_18_port, 
                           RES(17) => SHIFT_RES_17_port, RES(16) => 
                           SHIFT_RES_16_port, RES(15) => SHIFT_RES_15_port, 
                           RES(14) => SHIFT_RES_14_port, RES(13) => 
                           SHIFT_RES_13_port, RES(12) => SHIFT_RES_12_port, 
                           RES(11) => SHIFT_RES_11_port, RES(10) => 
                           SHIFT_RES_10_port, RES(9) => SHIFT_RES_9_port, 
                           RES(8) => SHIFT_RES_8_port, RES(7) => 
                           SHIFT_RES_7_port, RES(6) => SHIFT_RES_6_port, RES(5)
                           => SHIFT_RES_5_port, RES(4) => SHIFT_RES_4_port, 
                           RES(3) => SHIFT_RES_3_port, RES(2) => 
                           SHIFT_RES_2_port, RES(1) => SHIFT_RES_1_port, RES(0)
                           => SHIFT_RES_0_port);
   Add_Sub_unit : P4Adder_NBIT32 port map( A(31) => A_ADD_31_port, A(30) => 
                           A_ADD_30_port, A(29) => A_ADD_29_port, A(28) => 
                           A_ADD_28_port, A(27) => A_ADD_27_port, A(26) => 
                           A_ADD_26_port, A(25) => A_ADD_25_port, A(24) => 
                           A_ADD_24_port, A(23) => A_ADD_23_port, A(22) => 
                           A_ADD_22_port, A(21) => A_ADD_21_port, A(20) => 
                           A_ADD_20_port, A(19) => A_ADD_19_port, A(18) => 
                           A_ADD_18_port, A(17) => A_ADD_17_port, A(16) => 
                           A_ADD_16_port, A(15) => A_ADD_15_port, A(14) => 
                           A_ADD_14_port, A(13) => A_ADD_13_port, A(12) => 
                           A_ADD_12_port, A(11) => A_ADD_11_port, A(10) => 
                           A_ADD_10_port, A(9) => A_ADD_9_port, A(8) => 
                           A_ADD_8_port, A(7) => A_ADD_7_port, A(6) => 
                           A_ADD_6_port, A(5) => A_ADD_5_port, A(4) => 
                           A_ADD_4_port, A(3) => A_ADD_3_port, A(2) => 
                           A_ADD_2_port, A(1) => A_ADD_1_port, A(0) => 
                           A_ADD_0_port, B(31) => B_ADD_31_port, B(30) => 
                           B_ADD_30_port, B(29) => B_ADD_29_port, B(28) => 
                           B_ADD_28_port, B(27) => B_ADD_27_port, B(26) => 
                           B_ADD_26_port, B(25) => B_ADD_25_port, B(24) => 
                           B_ADD_24_port, B(23) => B_ADD_23_port, B(22) => 
                           B_ADD_22_port, B(21) => B_ADD_21_port, B(20) => 
                           B_ADD_20_port, B(19) => B_ADD_19_port, B(18) => 
                           B_ADD_18_port, B(17) => B_ADD_17_port, B(16) => 
                           B_ADD_16_port, B(15) => B_ADD_15_port, B(14) => 
                           B_ADD_14_port, B(13) => B_ADD_13_port, B(12) => 
                           B_ADD_12_port, B(11) => B_ADD_11_port, B(10) => 
                           B_ADD_10_port, B(9) => B_ADD_9_port, B(8) => 
                           B_ADD_8_port, B(7) => B_ADD_7_port, B(6) => 
                           B_ADD_6_port, B(5) => B_ADD_5_port, B(4) => 
                           B_ADD_4_port, B(3) => B_ADD_3_port, B(2) => 
                           B_ADD_2_port, B(1) => B_ADD_1_port, B(0) => 
                           B_ADD_0_port, Cin => ADD_SUB, S(31) => 
                           ADD_SUB_RES_31_port, S(30) => ADD_SUB_RES_30_port, 
                           S(29) => ADD_SUB_RES_29_port, S(28) => 
                           ADD_SUB_RES_28_port, S(27) => ADD_SUB_RES_27_port, 
                           S(26) => ADD_SUB_RES_26_port, S(25) => 
                           ADD_SUB_RES_25_port, S(24) => ADD_SUB_RES_24_port, 
                           S(23) => ADD_SUB_RES_23_port, S(22) => 
                           ADD_SUB_RES_22_port, S(21) => ADD_SUB_RES_21_port, 
                           S(20) => ADD_SUB_RES_20_port, S(19) => 
                           ADD_SUB_RES_19_port, S(18) => ADD_SUB_RES_18_port, 
                           S(17) => ADD_SUB_RES_17_port, S(16) => 
                           ADD_SUB_RES_16_port, S(15) => ADD_SUB_RES_15_port, 
                           S(14) => ADD_SUB_RES_14_port, S(13) => 
                           ADD_SUB_RES_13_port, S(12) => ADD_SUB_RES_12_port, 
                           S(11) => ADD_SUB_RES_11_port, S(10) => 
                           ADD_SUB_RES_10_port, S(9) => ADD_SUB_RES_9_port, 
                           S(8) => ADD_SUB_RES_8_port, S(7) => 
                           ADD_SUB_RES_7_port, S(6) => ADD_SUB_RES_6_port, S(5)
                           => ADD_SUB_RES_5_port, S(4) => ADD_SUB_RES_4_port, 
                           S(3) => ADD_SUB_RES_3_port, S(2) => 
                           ADD_SUB_RES_2_port, S(1) => ADD_SUB_RES_1_port, S(0)
                           => ADD_SUB_RES_0_port, Cout => n_1103);
   Res_mux : mux41_NBIT32_1 port map( A(31) => ADD_SUB_RES_31_port, A(30) => 
                           ADD_SUB_RES_30_port, A(29) => ADD_SUB_RES_29_port, 
                           A(28) => ADD_SUB_RES_28_port, A(27) => 
                           ADD_SUB_RES_27_port, A(26) => ADD_SUB_RES_26_port, 
                           A(25) => ADD_SUB_RES_25_port, A(24) => 
                           ADD_SUB_RES_24_port, A(23) => ADD_SUB_RES_23_port, 
                           A(22) => ADD_SUB_RES_22_port, A(21) => 
                           ADD_SUB_RES_21_port, A(20) => ADD_SUB_RES_20_port, 
                           A(19) => ADD_SUB_RES_19_port, A(18) => 
                           ADD_SUB_RES_18_port, A(17) => ADD_SUB_RES_17_port, 
                           A(16) => ADD_SUB_RES_16_port, A(15) => 
                           ADD_SUB_RES_15_port, A(14) => ADD_SUB_RES_14_port, 
                           A(13) => ADD_SUB_RES_13_port, A(12) => 
                           ADD_SUB_RES_12_port, A(11) => ADD_SUB_RES_11_port, 
                           A(10) => ADD_SUB_RES_10_port, A(9) => 
                           ADD_SUB_RES_9_port, A(8) => ADD_SUB_RES_8_port, A(7)
                           => ADD_SUB_RES_7_port, A(6) => ADD_SUB_RES_6_port, 
                           A(5) => ADD_SUB_RES_5_port, A(4) => 
                           ADD_SUB_RES_4_port, A(3) => ADD_SUB_RES_3_port, A(2)
                           => ADD_SUB_RES_2_port, A(1) => ADD_SUB_RES_1_port, 
                           A(0) => ADD_SUB_RES_0_port, B(31) => 
                           LOGIC_RES_31_port, B(30) => LOGIC_RES_30_port, B(29)
                           => LOGIC_RES_29_port, B(28) => LOGIC_RES_28_port, 
                           B(27) => LOGIC_RES_27_port, B(26) => 
                           LOGIC_RES_26_port, B(25) => LOGIC_RES_25_port, B(24)
                           => LOGIC_RES_24_port, B(23) => LOGIC_RES_23_port, 
                           B(22) => LOGIC_RES_22_port, B(21) => 
                           LOGIC_RES_21_port, B(20) => LOGIC_RES_20_port, B(19)
                           => LOGIC_RES_19_port, B(18) => LOGIC_RES_18_port, 
                           B(17) => LOGIC_RES_17_port, B(16) => 
                           LOGIC_RES_16_port, B(15) => LOGIC_RES_15_port, B(14)
                           => LOGIC_RES_14_port, B(13) => LOGIC_RES_13_port, 
                           B(12) => LOGIC_RES_12_port, B(11) => 
                           LOGIC_RES_11_port, B(10) => LOGIC_RES_10_port, B(9) 
                           => LOGIC_RES_9_port, B(8) => LOGIC_RES_8_port, B(7) 
                           => LOGIC_RES_7_port, B(6) => LOGIC_RES_6_port, B(5) 
                           => LOGIC_RES_5_port, B(4) => LOGIC_RES_4_port, B(3) 
                           => LOGIC_RES_3_port, B(2) => LOGIC_RES_2_port, B(1) 
                           => LOGIC_RES_1_port, B(0) => LOGIC_RES_0_port, C(31)
                           => SHIFT_RES_31_port, C(30) => SHIFT_RES_30_port, 
                           C(29) => SHIFT_RES_29_port, C(28) => 
                           SHIFT_RES_28_port, C(27) => SHIFT_RES_27_port, C(26)
                           => SHIFT_RES_26_port, C(25) => SHIFT_RES_25_port, 
                           C(24) => SHIFT_RES_24_port, C(23) => 
                           SHIFT_RES_23_port, C(22) => SHIFT_RES_22_port, C(21)
                           => SHIFT_RES_21_port, C(20) => SHIFT_RES_20_port, 
                           C(19) => SHIFT_RES_19_port, C(18) => 
                           SHIFT_RES_18_port, C(17) => SHIFT_RES_17_port, C(16)
                           => SHIFT_RES_16_port, C(15) => SHIFT_RES_15_port, 
                           C(14) => SHIFT_RES_14_port, C(13) => 
                           SHIFT_RES_13_port, C(12) => SHIFT_RES_12_port, C(11)
                           => SHIFT_RES_11_port, C(10) => SHIFT_RES_10_port, 
                           C(9) => SHIFT_RES_9_port, C(8) => SHIFT_RES_8_port, 
                           C(7) => SHIFT_RES_7_port, C(6) => SHIFT_RES_6_port, 
                           C(5) => SHIFT_RES_5_port, C(4) => SHIFT_RES_4_port, 
                           C(3) => SHIFT_RES_3_port, C(2) => SHIFT_RES_2_port, 
                           C(1) => SHIFT_RES_1_port, C(0) => SHIFT_RES_0_port, 
                           D(31) => n244_port, D(30) => n243_port, D(29) => 
                           n241_port, D(28) => n240_port, D(27) => n239_port, 
                           D(26) => n238_port, D(25) => n237_port, D(24) => 
                           n236_port, D(23) => n235_port, D(22) => n234_port, 
                           D(21) => n233_port, D(20) => n232_port, D(19) => 
                           n230_port, D(18) => n229_port, D(17) => n228_port, 
                           D(16) => n227_port, D(15) => n226_port, D(14) => 
                           n225_port, D(13) => n224_port, D(12) => n223_port, 
                           D(11) => n222_port, D(10) => n221_port, D(9) => n251
                           , D(8) => n250, D(7) => n249, D(6) => n248, D(5) => 
                           n247, D(4) => n246, D(3) => n245_port, D(2) => 
                           n242_port, D(1) => n231_port, D(0) => 
                           COMP_RES_0_port, S(1) => select_type_sig_1_port, 
                           S(0) => select_type_sig_0_port, Z(31) => 
                           sig_intraMux_31_port, Z(30) => sig_intraMux_30_port,
                           Z(29) => sig_intraMux_29_port, Z(28) => 
                           sig_intraMux_28_port, Z(27) => sig_intraMux_27_port,
                           Z(26) => sig_intraMux_26_port, Z(25) => 
                           sig_intraMux_25_port, Z(24) => sig_intraMux_24_port,
                           Z(23) => sig_intraMux_23_port, Z(22) => 
                           sig_intraMux_22_port, Z(21) => sig_intraMux_21_port,
                           Z(20) => sig_intraMux_20_port, Z(19) => 
                           sig_intraMux_19_port, Z(18) => sig_intraMux_18_port,
                           Z(17) => sig_intraMux_17_port, Z(16) => 
                           sig_intraMux_16_port, Z(15) => sig_intraMux_15_port,
                           Z(14) => sig_intraMux_14_port, Z(13) => 
                           sig_intraMux_13_port, Z(12) => sig_intraMux_12_port,
                           Z(11) => sig_intraMux_11_port, Z(10) => 
                           sig_intraMux_10_port, Z(9) => sig_intraMux_9_port, 
                           Z(8) => sig_intraMux_8_port, Z(7) => 
                           sig_intraMux_7_port, Z(6) => sig_intraMux_6_port, 
                           Z(5) => sig_intraMux_5_port, Z(4) => 
                           sig_intraMux_4_port, Z(3) => sig_intraMux_3_port, 
                           Z(2) => sig_intraMux_2_port, Z(1) => 
                           sig_intraMux_1_port, Z(0) => sig_intraMux_0_port);
   Zeros_mux : mux21_NBIT32_1 port map( A(31) => sig_intraMux_31_port, A(30) =>
                           sig_intraMux_30_port, A(29) => sig_intraMux_29_port,
                           A(28) => sig_intraMux_28_port, A(27) => 
                           sig_intraMux_27_port, A(26) => sig_intraMux_26_port,
                           A(25) => sig_intraMux_25_port, A(24) => 
                           sig_intraMux_24_port, A(23) => sig_intraMux_23_port,
                           A(22) => sig_intraMux_22_port, A(21) => 
                           sig_intraMux_21_port, A(20) => sig_intraMux_20_port,
                           A(19) => sig_intraMux_19_port, A(18) => 
                           sig_intraMux_18_port, A(17) => sig_intraMux_17_port,
                           A(16) => sig_intraMux_16_port, A(15) => 
                           sig_intraMux_15_port, A(14) => sig_intraMux_14_port,
                           A(13) => sig_intraMux_13_port, A(12) => 
                           sig_intraMux_12_port, A(11) => sig_intraMux_11_port,
                           A(10) => sig_intraMux_10_port, A(9) => 
                           sig_intraMux_9_port, A(8) => sig_intraMux_8_port, 
                           A(7) => sig_intraMux_7_port, A(6) => 
                           sig_intraMux_6_port, A(5) => sig_intraMux_5_port, 
                           A(4) => sig_intraMux_4_port, A(3) => 
                           sig_intraMux_3_port, A(2) => sig_intraMux_2_port, 
                           A(1) => sig_intraMux_1_port, A(0) => 
                           sig_intraMux_0_port, B(31) => n220_port, B(30) => 
                           n220_port, B(29) => n220_port, B(28) => n220_port, 
                           B(27) => n220_port, B(26) => n220_port, B(25) => 
                           n220_port, B(24) => n220_port, B(23) => n220_port, 
                           B(22) => n220_port, B(21) => n220_port, B(20) => 
                           n220_port, B(19) => n220_port, B(18) => n220_port, 
                           B(17) => n220_port, B(16) => n220_port, B(15) => 
                           n220_port, B(14) => n220_port, B(13) => n220_port, 
                           B(12) => n220_port, B(11) => n220_port, B(10) => 
                           n220_port, B(9) => n220_port, B(8) => n220_port, 
                           B(7) => n220_port, B(6) => n220_port, B(5) => 
                           n220_port, B(4) => n220_port, B(3) => n220_port, 
                           B(2) => n220_port, B(1) => n220_port, B(0) => 
                           n220_port, S => select_zero_sig, Z(31) => 
                           ALU_RES(31), Z(30) => ALU_RES(30), Z(29) => 
                           ALU_RES(29), Z(28) => ALU_RES(28), Z(27) => 
                           ALU_RES(27), Z(26) => ALU_RES(26), Z(25) => 
                           ALU_RES(25), Z(24) => ALU_RES(24), Z(23) => 
                           ALU_RES(23), Z(22) => ALU_RES(22), Z(21) => 
                           ALU_RES(21), Z(20) => ALU_RES(20), Z(19) => 
                           ALU_RES(19), Z(18) => ALU_RES(18), Z(17) => 
                           ALU_RES(17), Z(16) => ALU_RES(16), Z(15) => 
                           ALU_RES(15), Z(14) => ALU_RES(14), Z(13) => 
                           ALU_RES(13), Z(12) => ALU_RES(12), Z(11) => 
                           ALU_RES(11), Z(10) => ALU_RES(10), Z(9) => 
                           ALU_RES(9), Z(8) => ALU_RES(8), Z(7) => ALU_RES(7), 
                           Z(6) => ALU_RES(6), Z(5) => ALU_RES(5), Z(4) => 
                           ALU_RES(4), Z(3) => ALU_RES(3), Z(2) => ALU_RES(2), 
                           Z(1) => ALU_RES(1), Z(0) => ALU_RES(0));
   U4 : BUF_X1 port map( A => N211, Z => n213_port);
   U5 : BUF_X1 port map( A => N178, Z => n215_port);
   U6 : INV_X1 port map( A => n184_port, ZN => n201_port);
   U7 : BUF_X1 port map( A => n77, Z => n188_port);
   U8 : BUF_X1 port map( A => n77, Z => n189_port);
   U9 : INV_X1 port map( A => n184_port, ZN => n202_port);
   U10 : BUF_X1 port map( A => n195_port, Z => n199_port);
   U11 : BUF_X1 port map( A => n194_port, Z => n197_port);
   U12 : BUF_X1 port map( A => n194_port, Z => n196_port);
   U13 : BUF_X1 port map( A => n77, Z => n190_port);
   U14 : BUF_X1 port map( A => n194_port, Z => n198_port);
   U15 : BUF_X1 port map( A => n195_port, Z => n200_port);
   U16 : NAND2_X1 port map( A1 => n201_port, A2 => n185_port, ZN => N178);
   U17 : OR2_X1 port map( A1 => n198_port, A2 => n193_port, ZN => N211);
   U18 : OR2_X1 port map( A1 => n213_port, A2 => n203_port, ZN => 
                           select_type_sig_0_port);
   U19 : OR2_X1 port map( A1 => n208_port, A2 => n203_port, ZN => 
                           select_type_sig_1_port);
   U20 : BUF_X1 port map( A => n76, Z => n192_port);
   U21 : BUF_X1 port map( A => n76, Z => n191_port);
   U22 : BUF_X1 port map( A => n140, Z => n185_port);
   U23 : BUF_X1 port map( A => n76, Z => n193_port);
   U24 : BUF_X1 port map( A => n140, Z => n186_port);
   U25 : BUF_X1 port map( A => N244, Z => n208_port);
   U26 : BUF_X1 port map( A => n140, Z => n187_port);
   U27 : BUF_X1 port map( A => N245, Z => n203_port);
   U28 : AND2_X1 port map( A1 => n142, A2 => n320, ZN => n184_port);
   U29 : OR4_X1 port map( A1 => N177, A2 => n215_port, A3 => n149, A4 => 
                           select_type_sig_0_port, ZN => N176);
   U30 : AND2_X1 port map( A1 => n198_port, A2 => n320, ZN => n77);
   U31 : NOR2_X1 port map( A1 => n320, A2 => n71, ZN => n146);
   U32 : BUF_X1 port map( A => n75, Z => n194_port);
   U33 : BUF_X1 port map( A => n75, Z => n195_port);
   U34 : AND2_X1 port map( A1 => n208_port, A2 => n320, ZN => n149);
   U35 : NOR3_X1 port map( A1 => n319, A2 => ALU_OPC(0), A3 => n318, ZN => N244
                           );
   U36 : NOR3_X1 port map( A1 => ALU_OPC(1), A2 => ALU_OPC(0), A3 => n319, ZN 
                           => n142);
   U37 : NAND4_X1 port map( A1 => ALU_OPC(3), A2 => n319, A3 => n318, A4 => 
                           n317, ZN => n140);
   U38 : NOR3_X1 port map( A1 => ALU_OPC(2), A2 => ALU_OPC(0), A3 => n318, ZN 
                           => n75);
   U39 : INV_X1 port map( A => ALU_OPC(2), ZN => n319);
   U40 : OAI22_X1 port map( A1 => OP2(0), A2 => n202_port, B1 => n285, B2 => 
                           n185_port, ZN => N179);
   U41 : OAI22_X1 port map( A1 => OP2(1), A2 => n202_port, B1 => n286, B2 => 
                           n185_port, ZN => N180);
   U42 : OAI22_X1 port map( A1 => OP2(2), A2 => n201_port, B1 => n287, B2 => 
                           n185_port, ZN => N181);
   U43 : OAI22_X1 port map( A1 => OP2(3), A2 => n202_port, B1 => n288, B2 => 
                           n185_port, ZN => N182);
   U44 : OAI22_X1 port map( A1 => OP2(4), A2 => n201_port, B1 => n289, B2 => 
                           n185_port, ZN => N183);
   U45 : OAI22_X1 port map( A1 => OP2(5), A2 => n202_port, B1 => n290, B2 => 
                           n185_port, ZN => N184);
   U46 : OAI22_X1 port map( A1 => OP2(6), A2 => n201_port, B1 => n291, B2 => 
                           n185_port, ZN => N185);
   U47 : OAI22_X1 port map( A1 => OP2(7), A2 => n202_port, B1 => n292, B2 => 
                           n185_port, ZN => N186);
   U48 : OAI22_X1 port map( A1 => OP2(8), A2 => n202_port, B1 => n293, B2 => 
                           n185_port, ZN => N187);
   U49 : OAI22_X1 port map( A1 => OP2(9), A2 => n202_port, B1 => n294, B2 => 
                           n185_port, ZN => N188);
   U50 : OAI22_X1 port map( A1 => OP2(10), A2 => n202_port, B1 => n295, B2 => 
                           n185_port, ZN => N189);
   U51 : OAI22_X1 port map( A1 => OP2(11), A2 => n202_port, B1 => n296, B2 => 
                           n186_port, ZN => N190);
   U52 : OAI22_X1 port map( A1 => OP2(12), A2 => n202_port, B1 => n297, B2 => 
                           n186_port, ZN => N191);
   U53 : OAI22_X1 port map( A1 => OP2(13), A2 => n202_port, B1 => n298, B2 => 
                           n186_port, ZN => N192);
   U54 : OAI22_X1 port map( A1 => OP2(14), A2 => n202_port, B1 => n299, B2 => 
                           n186_port, ZN => N193);
   U55 : OAI22_X1 port map( A1 => OP2(15), A2 => n202_port, B1 => n300, B2 => 
                           n186_port, ZN => N194);
   U56 : OAI22_X1 port map( A1 => OP2(16), A2 => n202_port, B1 => n301, B2 => 
                           n186_port, ZN => N195);
   U57 : OAI22_X1 port map( A1 => OP2(17), A2 => n202_port, B1 => n302, B2 => 
                           n186_port, ZN => N196);
   U58 : OAI22_X1 port map( A1 => OP2(18), A2 => n202_port, B1 => n303, B2 => 
                           n186_port, ZN => N197);
   U59 : OAI22_X1 port map( A1 => OP2(19), A2 => n202_port, B1 => n304, B2 => 
                           n186_port, ZN => N198);
   U60 : OAI22_X1 port map( A1 => OP2(20), A2 => n201_port, B1 => n305, B2 => 
                           n186_port, ZN => N199);
   U61 : OAI22_X1 port map( A1 => OP2(21), A2 => n201_port, B1 => n306, B2 => 
                           n186_port, ZN => N200);
   U62 : OAI22_X1 port map( A1 => OP2(22), A2 => n201_port, B1 => n307, B2 => 
                           n186_port, ZN => N201);
   U63 : OAI22_X1 port map( A1 => OP2(23), A2 => n201_port, B1 => n308, B2 => 
                           n187_port, ZN => N202);
   U64 : OAI22_X1 port map( A1 => OP2(24), A2 => n201_port, B1 => n309, B2 => 
                           n187_port, ZN => N203);
   U65 : OAI22_X1 port map( A1 => OP2(25), A2 => n201_port, B1 => n310, B2 => 
                           n187_port, ZN => N204);
   U66 : OAI22_X1 port map( A1 => OP2(26), A2 => n201_port, B1 => n311, B2 => 
                           n187_port, ZN => N205);
   U67 : OAI22_X1 port map( A1 => OP2(27), A2 => n201_port, B1 => n312, B2 => 
                           n187_port, ZN => N206);
   U68 : OAI22_X1 port map( A1 => OP2(28), A2 => n201_port, B1 => n313, B2 => 
                           n187_port, ZN => N207);
   U69 : OAI22_X1 port map( A1 => OP2(29), A2 => n201_port, B1 => n314, B2 => 
                           n187_port, ZN => N208);
   U70 : OAI22_X1 port map( A1 => OP2(30), A2 => n201_port, B1 => n315, B2 => 
                           n187_port, ZN => N209);
   U71 : OAI22_X1 port map( A1 => OP2(31), A2 => n201_port, B1 => n316, B2 => 
                           n187_port, ZN => N210);
   U72 : INV_X1 port map( A => ALU_OPC(3), ZN => n320);
   U73 : INV_X1 port map( A => ALU_OPC(1), ZN => n318);
   U74 : OAI21_X1 port map( B1 => n143, B2 => n317, A => n144, ZN => N177);
   U75 : AOI22_X1 port map( A1 => ALU_OPC(3), A2 => n319, B1 => ALU_OPC(1), B2 
                           => ALU_OPC(2), ZN => n143);
   U76 : NAND2_X1 port map( A1 => n71, A2 => n141, ZN => N245);
   U77 : NAND4_X1 port map( A1 => ALU_OPC(0), A2 => ALU_OPC(1), A3 => n320, A4 
                           => n319, ZN => n141);
   U78 : INV_X1 port map( A => ALU_OPC(0), ZN => n317);
   U79 : AND2_X1 port map( A1 => ALU_OPC(3), A2 => n142, ZN => n76);
   U80 : OAI21_X1 port map( B1 => n122, B2 => n261, A => n123, ZN => N220);
   U81 : AOI221_X1 port map( B1 => n197_port, B2 => n293, C1 => OP2(8), C2 => 
                           n192_port, A => n188_port, ZN => n122);
   U82 : INV_X1 port map( A => OP1(8), ZN => n261);
   U83 : OAI21_X1 port map( B1 => n120, B2 => n262, A => n121, ZN => N221);
   U84 : AOI221_X1 port map( B1 => n197_port, B2 => n294, C1 => OP2(9), C2 => 
                           n192_port, A => n188_port, ZN => n120);
   U85 : INV_X1 port map( A => OP1(9), ZN => n262);
   U86 : OAI21_X1 port map( B1 => n118, B2 => n263, A => n119, ZN => N222);
   U87 : AOI221_X1 port map( B1 => n197_port, B2 => n295, C1 => OP2(10), C2 => 
                           n192_port, A => n188_port, ZN => n118);
   U88 : INV_X1 port map( A => OP1(10), ZN => n263);
   U89 : OAI21_X1 port map( B1 => n116, B2 => n264, A => n117, ZN => N223);
   U90 : AOI221_X1 port map( B1 => n197_port, B2 => n296, C1 => OP2(11), C2 => 
                           n192_port, A => n188_port, ZN => n116);
   U91 : INV_X1 port map( A => OP1(11), ZN => n264);
   U92 : OAI21_X1 port map( B1 => n114, B2 => n265, A => n115, ZN => N224);
   U93 : AOI221_X1 port map( B1 => n197_port, B2 => n297, C1 => OP2(12), C2 => 
                           n192_port, A => n189_port, ZN => n114);
   U94 : INV_X1 port map( A => OP1(12), ZN => n265);
   U95 : OAI21_X1 port map( B1 => n112, B2 => n266, A => n113, ZN => N225);
   U96 : AOI221_X1 port map( B1 => n197_port, B2 => n298, C1 => OP2(13), C2 => 
                           n192_port, A => n189_port, ZN => n112);
   U97 : INV_X1 port map( A => OP1(13), ZN => n266);
   U98 : OAI21_X1 port map( B1 => n110, B2 => n267, A => n111, ZN => N226);
   U99 : AOI221_X1 port map( B1 => n197_port, B2 => n299, C1 => OP2(14), C2 => 
                           n192_port, A => n189_port, ZN => n110);
   U100 : INV_X1 port map( A => OP1(14), ZN => n267);
   U101 : OAI21_X1 port map( B1 => n108, B2 => n268, A => n109, ZN => N227);
   U102 : AOI221_X1 port map( B1 => n197_port, B2 => n300, C1 => OP2(15), C2 =>
                           n192_port, A => n189_port, ZN => n108);
   U103 : INV_X1 port map( A => OP1(15), ZN => n268);
   U104 : OAI21_X1 port map( B1 => n106, B2 => n269, A => n107, ZN => N228);
   U105 : AOI221_X1 port map( B1 => n197_port, B2 => n301, C1 => OP2(16), C2 =>
                           n192_port, A => n189_port, ZN => n106);
   U106 : INV_X1 port map( A => OP1(16), ZN => n269);
   U107 : OAI21_X1 port map( B1 => n104, B2 => n270, A => n105, ZN => N229);
   U108 : AOI221_X1 port map( B1 => n197_port, B2 => n302, C1 => OP2(17), C2 =>
                           n192_port, A => n189_port, ZN => n104);
   U109 : INV_X1 port map( A => OP1(17), ZN => n270);
   U110 : OAI21_X1 port map( B1 => n102, B2 => n271, A => n103, ZN => N230);
   U111 : AOI221_X1 port map( B1 => n197_port, B2 => n303, C1 => OP2(18), C2 =>
                           n191_port, A => n189_port, ZN => n102);
   U112 : INV_X1 port map( A => OP1(18), ZN => n271);
   U113 : OAI21_X1 port map( B1 => n100, B2 => n272, A => n101, ZN => N231);
   U114 : AOI221_X1 port map( B1 => n197_port, B2 => n304, C1 => OP2(19), C2 =>
                           n191_port, A => n189_port, ZN => n100);
   U115 : INV_X1 port map( A => OP1(19), ZN => n272);
   U116 : OAI21_X1 port map( B1 => n98, B2 => n273, A => n99, ZN => N232);
   U117 : AOI221_X1 port map( B1 => n196_port, B2 => n305, C1 => OP2(20), C2 =>
                           n191_port, A => n189_port, ZN => n98);
   U118 : INV_X1 port map( A => OP1(20), ZN => n273);
   U119 : OAI21_X1 port map( B1 => n96, B2 => n274, A => n97, ZN => N233);
   U120 : AOI221_X1 port map( B1 => n196_port, B2 => n306, C1 => OP2(21), C2 =>
                           n191_port, A => n189_port, ZN => n96);
   U121 : INV_X1 port map( A => OP1(21), ZN => n274);
   U122 : OAI21_X1 port map( B1 => n94, B2 => n275, A => n95, ZN => N234);
   U123 : AOI221_X1 port map( B1 => n196_port, B2 => n307, C1 => OP2(22), C2 =>
                           n191_port, A => n189_port, ZN => n94);
   U124 : INV_X1 port map( A => OP1(22), ZN => n275);
   U125 : OAI21_X1 port map( B1 => n92, B2 => n276, A => n93, ZN => N235);
   U126 : AOI221_X1 port map( B1 => n196_port, B2 => n308, C1 => OP2(23), C2 =>
                           n192_port, A => n189_port, ZN => n92);
   U127 : INV_X1 port map( A => OP1(23), ZN => n276);
   U128 : OAI21_X1 port map( B1 => n90, B2 => n277, A => n91, ZN => N236);
   U129 : AOI221_X1 port map( B1 => n196_port, B2 => n309, C1 => OP2(24), C2 =>
                           n191_port, A => n190_port, ZN => n90);
   U130 : INV_X1 port map( A => OP1(24), ZN => n277);
   U131 : OAI21_X1 port map( B1 => n88, B2 => n278, A => n89, ZN => N237);
   U132 : AOI221_X1 port map( B1 => n196_port, B2 => n310, C1 => OP2(25), C2 =>
                           n191_port, A => n190_port, ZN => n88);
   U133 : INV_X1 port map( A => OP1(25), ZN => n278);
   U134 : OAI21_X1 port map( B1 => n86, B2 => n279, A => n87, ZN => N238);
   U135 : AOI221_X1 port map( B1 => n196_port, B2 => n311, C1 => OP2(26), C2 =>
                           n191_port, A => n190_port, ZN => n86);
   U136 : INV_X1 port map( A => OP1(26), ZN => n279);
   U137 : OAI21_X1 port map( B1 => n84, B2 => n280, A => n85, ZN => N239);
   U138 : AOI221_X1 port map( B1 => n196_port, B2 => n312, C1 => OP2(27), C2 =>
                           n191_port, A => n190_port, ZN => n84);
   U139 : INV_X1 port map( A => OP1(27), ZN => n280);
   U140 : OAI21_X1 port map( B1 => n82, B2 => n281, A => n83, ZN => N240);
   U141 : AOI221_X1 port map( B1 => n196_port, B2 => n313, C1 => OP2(28), C2 =>
                           n191_port, A => n190_port, ZN => n82);
   U142 : INV_X1 port map( A => OP1(28), ZN => n281);
   U143 : OAI21_X1 port map( B1 => n80, B2 => n282, A => n81, ZN => N241);
   U144 : AOI221_X1 port map( B1 => n196_port, B2 => n314, C1 => OP2(29), C2 =>
                           n191_port, A => n190_port, ZN => n80);
   U145 : INV_X1 port map( A => OP1(29), ZN => n282);
   U146 : OAI21_X1 port map( B1 => n78, B2 => n283, A => n79, ZN => N242);
   U147 : AOI221_X1 port map( B1 => n196_port, B2 => n315, C1 => OP2(30), C2 =>
                           n191_port, A => n190_port, ZN => n78);
   U148 : INV_X1 port map( A => OP1(30), ZN => n283);
   U149 : OAI21_X1 port map( B1 => n73, B2 => n284, A => n74, ZN => N243);
   U150 : AOI221_X1 port map( B1 => n196_port, B2 => n316, C1 => n193_port, C2 
                           => OP2(31), A => n190_port, ZN => n73);
   U151 : INV_X1 port map( A => OP1(31), ZN => n284);
   U152 : OAI21_X1 port map( B1 => n138, B2 => n253, A => n139, ZN => N212);
   U153 : AOI221_X1 port map( B1 => n198_port, B2 => n285, C1 => OP2(0), C2 => 
                           n193_port, A => n188_port, ZN => n138);
   U154 : INV_X1 port map( A => OP1(0), ZN => n253);
   U155 : OAI21_X1 port map( B1 => n136, B2 => n254, A => n137, ZN => N213);
   U156 : AOI221_X1 port map( B1 => n198_port, B2 => n286, C1 => OP2(1), C2 => 
                           n193_port, A => n188_port, ZN => n136);
   U157 : INV_X1 port map( A => OP1(1), ZN => n254);
   U158 : OAI21_X1 port map( B1 => n134, B2 => n255, A => n135, ZN => N214);
   U159 : AOI221_X1 port map( B1 => n198_port, B2 => n287, C1 => OP2(2), C2 => 
                           n193_port, A => n188_port, ZN => n134);
   U160 : INV_X1 port map( A => OP1(2), ZN => n255);
   U161 : OAI21_X1 port map( B1 => n132, B2 => n256, A => n133, ZN => N215);
   U162 : AOI221_X1 port map( B1 => n198_port, B2 => n288, C1 => OP2(3), C2 => 
                           n193_port, A => n188_port, ZN => n132);
   U163 : INV_X1 port map( A => OP1(3), ZN => n256);
   U164 : OAI21_X1 port map( B1 => n130, B2 => n257, A => n131, ZN => N216);
   U165 : AOI221_X1 port map( B1 => n198_port, B2 => n289, C1 => OP2(4), C2 => 
                           n193_port, A => n188_port, ZN => n130);
   U166 : INV_X1 port map( A => OP1(4), ZN => n257);
   U167 : OAI21_X1 port map( B1 => n128, B2 => n258, A => n129, ZN => N217);
   U168 : AOI221_X1 port map( B1 => n198_port, B2 => n290, C1 => OP2(5), C2 => 
                           n193_port, A => n188_port, ZN => n128);
   U169 : INV_X1 port map( A => OP1(5), ZN => n258);
   U170 : OAI21_X1 port map( B1 => n126, B2 => n259, A => n127, ZN => N218);
   U171 : AOI221_X1 port map( B1 => n198_port, B2 => n291, C1 => OP2(6), C2 => 
                           n193_port, A => n188_port, ZN => n126);
   U172 : INV_X1 port map( A => OP1(6), ZN => n259);
   U173 : OAI21_X1 port map( B1 => n124, B2 => n260, A => n125, ZN => N219);
   U174 : AOI221_X1 port map( B1 => n198_port, B2 => n292, C1 => OP2(7), C2 => 
                           n192_port, A => n188_port, ZN => n124);
   U175 : INV_X1 port map( A => OP1(7), ZN => n260);
   U176 : NOR2_X1 port map( A1 => ALU_OPC(3), A2 => n71, ZN => n145);
   U177 : INV_X1 port map( A => OP2(0), ZN => n285);
   U178 : INV_X1 port map( A => OP2(1), ZN => n286);
   U179 : INV_X1 port map( A => OP2(2), ZN => n287);
   U180 : INV_X1 port map( A => OP2(3), ZN => n288);
   U181 : INV_X1 port map( A => OP2(4), ZN => n289);
   U182 : INV_X1 port map( A => OP2(5), ZN => n290);
   U183 : INV_X1 port map( A => OP2(6), ZN => n291);
   U184 : INV_X1 port map( A => OP2(7), ZN => n292);
   U185 : INV_X1 port map( A => OP2(8), ZN => n293);
   U186 : INV_X1 port map( A => OP2(9), ZN => n294);
   U187 : INV_X1 port map( A => OP2(10), ZN => n295);
   U222 : INV_X1 port map( A => OP2(11), ZN => n296);
   U223 : INV_X1 port map( A => OP2(12), ZN => n297);
   U224 : INV_X1 port map( A => OP2(13), ZN => n298);
   U225 : INV_X1 port map( A => OP2(14), ZN => n299);
   U226 : INV_X1 port map( A => OP2(15), ZN => n300);
   U227 : INV_X1 port map( A => OP2(16), ZN => n301);
   U228 : INV_X1 port map( A => OP2(17), ZN => n302);
   U229 : INV_X1 port map( A => OP2(18), ZN => n303);
   U230 : INV_X1 port map( A => OP2(19), ZN => n304);
   U231 : INV_X1 port map( A => OP2(20), ZN => n305);
   U232 : INV_X1 port map( A => OP2(21), ZN => n306);
   U233 : INV_X1 port map( A => OP2(22), ZN => n307);
   U234 : INV_X1 port map( A => OP2(23), ZN => n308);
   U235 : INV_X1 port map( A => OP2(24), ZN => n309);
   U236 : INV_X1 port map( A => OP2(25), ZN => n310);
   U237 : INV_X1 port map( A => OP2(26), ZN => n311);
   U238 : INV_X1 port map( A => OP2(27), ZN => n312);
   U239 : INV_X1 port map( A => OP2(28), ZN => n313);
   U240 : INV_X1 port map( A => OP2(29), ZN => n314);
   U241 : INV_X1 port map( A => OP2(30), ZN => n315);
   U242 : INV_X1 port map( A => OP2(31), ZN => n316);
   U243 : CLKBUF_X1 port map( A => N245, Z => n204_port);
   U244 : CLKBUF_X1 port map( A => N245, Z => n205_port);
   U245 : CLKBUF_X1 port map( A => N245, Z => n206_port);
   U246 : CLKBUF_X1 port map( A => N245, Z => n207_port);
   U247 : CLKBUF_X1 port map( A => N244, Z => n209_port);
   U248 : CLKBUF_X1 port map( A => N244, Z => n210_port);
   U249 : CLKBUF_X1 port map( A => N244, Z => n211_port);
   U250 : CLKBUF_X1 port map( A => N244, Z => n212_port);
   U251 : CLKBUF_X1 port map( A => N211, Z => n214_port);
   U252 : CLKBUF_X1 port map( A => N178, Z => n216_port);
   U253 : CLKBUF_X1 port map( A => N178, Z => n217_port);
   U254 : CLKBUF_X1 port map( A => N178, Z => n218_port);
   U255 : CLKBUF_X1 port map( A => N178, Z => n219_port);
   n220_port <= '0';
   n221_port <= '0';
   n222_port <= '0';
   n223_port <= '0';
   n224_port <= '0';
   n225_port <= '0';
   n226_port <= '0';
   n227_port <= '0';
   n228_port <= '0';
   n229_port <= '0';
   n230_port <= '0';
   n231_port <= '0';
   n232_port <= '0';
   n233_port <= '0';
   n234_port <= '0';
   n235_port <= '0';
   n236_port <= '0';
   n237_port <= '0';
   n238_port <= '0';
   n239_port <= '0';
   n240_port <= '0';
   n241_port <= '0';
   n242_port <= '0';
   n243_port <= '0';
   n244_port <= '0';
   n245_port <= '0';
   n246 <= '0';
   n247 <= '0';
   n248 <= '0';
   n249 <= '0';
   n250 <= '0';
   n251 <= '0';
   n252 <= '1';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FWD_Unit is

   port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB : in 
         std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;  
         FWDA, FWDB : out std_logic_vector (1 downto 0));

end FWD_Unit;

architecture SYN_bhv of FWD_Unit is

   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n43, n44, n45, n46 : std_logic;

begin
   
   U38 : XOR2_X1 port map( A => ADD_WR_WB(4), B => ADD_RS2(4), Z => n13);
   U39 : XOR2_X1 port map( A => ADD_WR_WB(0), B => ADD_RS2(0), Z => n12);
   U40 : XOR2_X1 port map( A => ADD_WR_MEM(4), B => ADD_RS2(4), Z => n19);
   U41 : XOR2_X1 port map( A => ADD_WR_MEM(3), B => ADD_RS2(3), Z => n18);
   U42 : XOR2_X1 port map( A => ADD_WR_WB(1), B => ADD_RS1(1), Z => n33);
   U43 : XOR2_X1 port map( A => ADD_WR_WB(0), B => ADD_RS1(0), Z => n32);
   U44 : XOR2_X1 port map( A => ADD_WR_MEM(4), B => ADD_RS1(4), Z => n39);
   U45 : XOR2_X1 port map( A => ADD_WR_MEM(3), B => ADD_RS1(3), Z => n38);
   U3 : OAI22_X1 port map( A1 => n46, A2 => n6, B1 => n5, B2 => n7, ZN => 
                           FWDB(0));
   U4 : INV_X1 port map( A => n5, ZN => n46);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n21, B1 => n20, B2 => n7, ZN => 
                           FWDA(0));
   U6 : INV_X1 port map( A => n20, ZN => n45);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n5, B1 => n43, B2 => n6, ZN => 
                           FWDB(1));
   U8 : OAI22_X1 port map( A1 => n44, A2 => n20, B1 => n43, B2 => n21, ZN => 
                           FWDA(1));
   U9 : INV_X1 port map( A => RST, ZN => n44);
   U10 : NOR3_X1 port map( A1 => n12, A2 => n44, A3 => n13, ZN => n11);
   U11 : NOR3_X1 port map( A1 => n32, A2 => n44, A3 => n33, ZN => n31);
   U12 : NAND4_X1 port map( A1 => n14, A2 => n15, A3 => n16, A4 => n17, ZN => 
                           n5);
   U13 : NOR2_X1 port map( A1 => n18, A2 => n19, ZN => n17);
   U14 : XNOR2_X1 port map( A => ADD_RS2(0), B => ADD_WR_MEM(0), ZN => n14);
   U15 : XNOR2_X1 port map( A => ADD_RS2(1), B => ADD_WR_MEM(1), ZN => n15);
   U16 : NAND4_X1 port map( A1 => n34, A2 => n35, A3 => n36, A4 => n37, ZN => 
                           n20);
   U17 : NOR2_X1 port map( A1 => n38, A2 => n39, ZN => n37);
   U18 : XNOR2_X1 port map( A => ADD_RS1(0), B => ADD_WR_MEM(0), ZN => n34);
   U19 : XNOR2_X1 port map( A => ADD_RS1(1), B => ADD_WR_MEM(1), ZN => n35);
   U20 : NAND4_X1 port map( A1 => n8, A2 => n9, A3 => n10, A4 => n11, ZN => n6)
                           ;
   U21 : XNOR2_X1 port map( A => ADD_RS2(3), B => ADD_WR_WB(3), ZN => n8);
   U22 : XNOR2_X1 port map( A => ADD_RS2(1), B => ADD_WR_WB(1), ZN => n9);
   U23 : XNOR2_X1 port map( A => ADD_RS2(2), B => ADD_WR_WB(2), ZN => n10);
   U24 : NAND4_X1 port map( A1 => n28, A2 => n29, A3 => n30, A4 => n31, ZN => 
                           n21);
   U25 : XNOR2_X1 port map( A => ADD_RS1(4), B => ADD_WR_WB(4), ZN => n28);
   U26 : XNOR2_X1 port map( A => ADD_RS1(3), B => ADD_WR_WB(3), ZN => n29);
   U27 : XNOR2_X1 port map( A => ADD_RS1(2), B => ADD_WR_WB(2), ZN => n30);
   U28 : XNOR2_X1 port map( A => ADD_RS2(2), B => ADD_WR_MEM(2), ZN => n16);
   U29 : XNOR2_X1 port map( A => ADD_RS1(2), B => ADD_WR_MEM(2), ZN => n36);
   U30 : NAND2_X1 port map( A1 => RST, A2 => n25, ZN => n7);
   U31 : OAI21_X1 port map( B1 => n26, B2 => n27, A => RF_WE_MEM, ZN => n25);
   U32 : OR2_X1 port map( A1 => ADD_WR_MEM(0), A2 => ADD_WR_MEM(1), ZN => n27);
   U33 : OR3_X1 port map( A1 => ADD_WR_MEM(3), A2 => ADD_WR_MEM(4), A3 => 
                           ADD_WR_MEM(2), ZN => n26);
   U34 : INV_X1 port map( A => n22, ZN => n43);
   U35 : OAI21_X1 port map( B1 => n23, B2 => n24, A => RF_WE_WB, ZN => n22);
   U36 : OR2_X1 port map( A1 => ADD_WR_WB(0), A2 => ADD_WR_WB(1), ZN => n24);
   U37 : OR3_X1 port map( A1 => ADD_WR_WB(3), A2 => ADD_WR_WB(4), A3 => 
                           ADD_WR_WB(2), ZN => n23);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N2 is

   port( DIN : in std_logic_vector (1 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (1 downto 0));

end regn_N2;

architecture SYN_bhv of regn_N2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n1, n2 : std_logic;

begin
   
   DOUT_reg_1_inst : DFFR_X1 port map( D => n6, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n4);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n5, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n3);
   U2 : OAI21_X1 port map( B1 => n3, B2 => EN, A => n2, ZN => n5);
   U3 : NAND2_X1 port map( A1 => DIN(0), A2 => EN, ZN => n2);
   U4 : OAI21_X1 port map( B1 => n4, B2 => EN, A => n1, ZN => n6);
   U5 : NAND2_X1 port map( A1 => EN, A2 => DIN(1), ZN => n1);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Branch_Cond_Unit_NBIT32 is

   port( RST : in std_logic;  A : in std_logic_vector (31 downto 0);  ALU_OPC :
         in std_logic_vector (0 to 3);  JUMP_TYPE : in std_logic_vector (1 
         downto 0);  PC_SEL : out std_logic_vector (1 downto 0);  ZERO : out 
         std_logic);

end Branch_Cond_Unit_NBIT32;

architecture SYN_bhv of Branch_Cond_Unit_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => ZERO);
   U4 : NOR4_X1 port map( A1 => A(23), A2 => A(22), A3 => A(21), A4 => A(20), 
                           ZN => n12);
   U5 : NOR4_X1 port map( A1 => A(9), A2 => A(8), A3 => A(7), A4 => A(6), ZN =>
                           n16);
   U6 : NAND4_X1 port map( A1 => ALU_OPC(0), A2 => RST, A3 => JUMP_TYPE(0), A4 
                           => n4, ZN => n2);
   U7 : NOR3_X1 port map( A1 => n5, A2 => ALU_OPC(1), A3 => ALU_OPC(2), ZN => 
                           n4);
   U8 : XNOR2_X1 port map( A => ALU_OPC(3), B => n6, ZN => n5);
   U9 : NOR2_X1 port map( A1 => n7, A2 => n8, ZN => n6);
   U10 : NAND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => n8
                           );
   U11 : NOR4_X1 port map( A1 => A(12), A2 => A(11), A3 => A(10), A4 => A(0), 
                           ZN => n9);
   U12 : NOR4_X1 port map( A1 => A(16), A2 => A(15), A3 => A(14), A4 => A(13), 
                           ZN => n10);
   U13 : NOR4_X1 port map( A1 => A(1), A2 => A(19), A3 => A(18), A4 => A(17), 
                           ZN => n11);
   U14 : NAND4_X1 port map( A1 => n13, A2 => n14, A3 => n15, A4 => n16, ZN => 
                           n7);
   U15 : NOR4_X1 port map( A1 => A(27), A2 => A(26), A3 => A(25), A4 => A(24), 
                           ZN => n13);
   U16 : NOR4_X1 port map( A1 => A(30), A2 => A(2), A3 => A(29), A4 => A(28), 
                           ZN => n14);
   U17 : NOR4_X1 port map( A1 => A(5), A2 => A(4), A3 => A(3), A4 => A(31), ZN 
                           => n15);
   U18 : NAND2_X1 port map( A1 => RST, A2 => JUMP_TYPE(1), ZN => n3);
   U19 : OAI22_X1 port map( A1 => JUMP_TYPE(1), A2 => n2, B1 => JUMP_TYPE(0), 
                           B2 => n3, ZN => PC_SEL(0));
   U20 : NOR2_X1 port map( A1 => n17, A2 => n3, ZN => PC_SEL(1));
   U21 : INV_X1 port map( A => JUMP_TYPE(0), ZN => n17);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity register_file_NBIT_ADD5_NBIT_DATA32 is

   port( CLK, RST, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RS1, 
         ADD_RS2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_NBIT_ADD5_NBIT_DATA32;

architecture SYN_bhv of register_file_NBIT_ADD5_NBIT_DATA32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
      n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, 
      n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, 
      n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, 
      n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, 
      n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, 
      n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, 
      n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, 
      n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, 
      n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, 
      n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, 
      n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, 
      n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, 
      n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, 
      n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, 
      n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, 
      n3143, n3144, n3145, n3146, n3174, n3175, n3176, n3177, n3178, n3206, 
      n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, 
      n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, 
      n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, 
      n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, 
      n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, 
      n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, 
      n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, 
      n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, 
      n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, 
      n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, 
      n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, 
      n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, 
      n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, 
      n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, 
      n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, 
      n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, 
      n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, 
      n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, 
      n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, 
      n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, 
      n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, 
      n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, 
      n3427, n3428, n3429, n3430, n938, n939, n950, n955, n956, n966, n971, 
      n972, n982, n987, n988, n998, n2623, n2624, n2625, n2626, n2627, n2628, 
      n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, 
      n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, 
      n2649, n2650, n2651, n2652, n2653, n2655, n2656, n2657, n2658, n2659, 
      n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, 
      n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, 
      n2680, n2681, n2682, n2683, n2684, n2685, n2690, n2691, n2692, n2693, 
      n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, 
      n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, 
      n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, 
      n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, 
      n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, 
      n2744, n2745, n2746, n2747, n2748, n2749, n2850, n2851, n2852, n2853, 
      n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, 
      n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, 
      n2874, n2875, n2876, n2877, n2910, n2911, n2912, n2913, n2914, n2915, 
      n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, 
      n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, 
      n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, 
      n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, 
      n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, 
      n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, 
      n2976, n2977, n2978, n2979, n2980, n2981, n2982, n3559, n3560, n3561, 
      n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, 
      n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, 
      n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, 
      n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, 
      n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, 
      n3676, n3677, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, 
      n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, 
      n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, 
      n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, 
      n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, 
      n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, 
      n3800, n3801, n3802, n3803, n3804, n3805, n3870, n3871, n3872, n3873, 
      n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, 
      n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, 
      n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, 
      n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, 
      n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, 
      n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, 
      n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, 
      n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, 
      n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, 
      n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, 
      n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, 
      n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, 
      n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, 
      n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, 
      n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, 
      n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, 
      n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, 
      n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, 
      n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, 
      n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, 
      n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, 
      n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, 
      n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, 
      n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, 
      n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, 
      n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, 
      n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, 
      n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, 
      n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, 
      n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, 
      n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, 
      n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, 
      n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, 
      n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, 
      n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, 
      n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, 
      n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, 
      n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, 
      n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, 
      n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, 
      n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, 
      n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, 
      n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, 
      n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, 
      n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, 
      n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, 
      n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, 
      n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, 
      n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, 
      n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, 
      n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, 
      n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, 
      n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, 
      n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, 
      n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, 
      n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, 
      n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, 
      n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, 
      n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, 
      n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, 
      n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, 
      n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, 
      n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, 
      n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, 
      n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, 
      n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, 
      n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n749, n824, n825,
      n826, n834, n835, n836, n837, n838, n840, n841, n842, n843, n844, n845, 
      n847, n848, n849, n871, n872, n873, n876, n877, n878, n888, n889, n890, 
      n893, n894, n895, n905, n906, n907, n910, n911, n912, n922, n923, n924, 
      n927, n928, n929, n941, n942, n943, n946, n947, n948, n961, n962, n963, 
      n967, n968, n969, n981, n983, n984, n989, n990, n991, n1002, n1003, n1004
      , n1007, n1008, n1009, n1019, n1020, n1021, n1024, n1025, n1026, n1036, 
      n1037, n1038, n1041, n1042, n1043, n1053, n1054, n1055, n1058, n1059, 
      n1060, n1070, n1071, n1072, n1075, n1076, n1077, n1087, n1088, n1089, 
      n1092, n1093, n1094, n1104, n1105, n1106, n1109, n1110, n1111, n1121, 
      n1122, n1123, n1126, n1127, n1128, n1138, n1139, n1140, n1143, n1144, 
      n1145, n1155, n1156, n1157, n1160, n1161, n1162, n1172, n1173, n1174, 
      n1177, n1178, n1179, n1189, n1190, n1191, n1194, n1195, n1196, n1206, 
      n1207, n1208, n1211, n1212, n1213, n1223, n1224, n1225, n1228, n1229, 
      n1230, n1240, n1241, n1242, n1245, n1246, n1247, n1257, n1258, n1259, 
      n1262, n1263, n1264, n1274, n1275, n1276, n1279, n1280, n1281, n1291, 
      n1292, n1293, n1296, n1297, n1298, n1308, n1309, n1310, n1313, n1314, 
      n1315, n1325, n1326, n1327, n1330, n1331, n1332, n1342, n1343, n1344, 
      n1347, n1348, n1349, n1359, n1360, n1361, n1364, n1365, n1366, n1376, 
      n1377, n1378, n1381, n1382, n1383, n1393, n1394, n1397, n1398, n1399, 
      n1400, n1401, n1402, n1406, n1412, n1413, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1427, n1437, n1438, n1439, n1447, n1448, n1449, 
      n1450, n1451, n1453, n1454, n1455, n1456, n1457, n1458, n1460, n1461, 
      n1462, n1481, n1482, n1483, n1486, n1487, n1488, n1498, n1499, n1500, 
      n1503, n1504, n1505, n1515, n1516, n1517, n1520, n1521, n1522, n1532, 
      n1533, n1534, n1537, n1538, n1539, n1549, n1550, n1551, n1554, n1555, 
      n1556, n1566, n1567, n1568, n1571, n1572, n1573, n1583, n1584, n1585, 
      n1588, n1589, n1590, n1600, n1601, n1602, n1605, n1606, n1607, n1617, 
      n1618, n1619, n1622, n1623, n1624, n1634, n1635, n1636, n1639, n1640, 
      n1641, n1651, n1652, n1653, n1656, n1657, n1658, n1668, n1669, n1670, 
      n1673, n1674, n1675, n1685, n1686, n1687, n1690, n1691, n1692, n1702, 
      n1703, n1704, n1707, n1708, n1709, n1719, n1720, n1721, n1724, n1725, 
      n1726, n1736, n1737, n1738, n1741, n1742, n1743, n1753, n1754, n1755, 
      n1758, n1759, n1760, n1770, n1771, n1772, n1775, n1776, n1777, n1787, 
      n1788, n1789, n1792, n1793, n1794, n1804, n1805, n1806, n1809, n1810, 
      n1811, n1821, n1822, n1823, n1826, n1827, n1828, n1838, n1839, n1840, 
      n1843, n1844, n1845, n1855, n1856, n1857, n1860, n1861, n1862, n1872, 
      n1873, n1874, n1877, n1878, n1879, n1889, n1890, n1891, n1894, n1895, 
      n1896, n1906, n1907, n1908, n1911, n1912, n1913, n1923, n1924, n1925, 
      n1928, n1929, n1930, n1940, n1941, n1942, n1945, n1946, n1947, n1957, 
      n1958, n1959, n1962, n1963, n1964, n1974, n1975, n1976, n1979, n1980, 
      n1981, n1993, n1994, n1997, n1998, n1999, n2000, n2001, n2002, n2006, 
      n2012, n2013, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2027, 
      n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, 
      n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, 
      n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, 
      n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, 
      n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
      n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, 
      n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, 
      n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, 
      n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
      n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, 
      n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, 
      n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, 
      n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, 
      n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, 
      n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, 
      n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, 
      n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, 
      n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, 
      n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, 
      n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, 
      n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, 
      n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, 
      n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, 
      n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, 
      n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, 
      n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, 
      n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, 
      n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, 
      n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, 
      n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, 
      n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, 
      n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, 
      n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, 
      n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, 
      n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, 
      n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, 
      n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, 
      n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, 
      n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, 
      n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, 
      n2438, n2439, n2440, n2441, n2442, n2443, n4606, n4607, n4608, n4609, 
      n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, 
      n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, 
      n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, 
      n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, 
      n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, 
      n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, 
      n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, 
      n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, 
      n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, 
      n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, 
      n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, 
      n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, 
      n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, 
      n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, 
      n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, 
      n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, 
      n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, 
      n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, 
      n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, 
      n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, 
      n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, 
      n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, 
      n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, 
      n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, 
      n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, 
      n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, 
      n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, 
      n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, 
      n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, 
      n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, 
      n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, 
      n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, 
      n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, 
      n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, 
      n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, 
      n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, 
      n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, 
      n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, 
      n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, 
      n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, 
      n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, 
      n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, 
      n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, 
      n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, 
      n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, 
      n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, 
      n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, 
      n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, 
      n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, 
      n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, 
      n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, 
      n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, 
      n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, 
      n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, 
      n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, 
      n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, 
      n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, 
      n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, 
      n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, 
      n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, 
      n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, 
      n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, 
      n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, 
      n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, 
      n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, 
      n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, 
      n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, 
      n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, 
      n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, 
      n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, 
      n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, 
      n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, 
      n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, 
      n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, 
      n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, 
      n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, 
      n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, 
      n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, 
      n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, 
      n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, 
      n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, 
      n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, 
      n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, 
      n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, 
      n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, 
      n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, 
      n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, 
      n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, 
      n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, 
      n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, 
      n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, 
      n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, 
      n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, 
      n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, 
      n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, 
      n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, 
      n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, 
      n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, 
      n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, 
      n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, 
      n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, 
      n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, 
      n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, 
      n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, 
      n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, 
      n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, 
      n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, 
      n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, 
      n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, 
      n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, 
      n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, 
      n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, 
      n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, 
      n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, 
      n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, 
      n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, 
      n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, 
      n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, 
      n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, 
      n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, 
      n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, 
      n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, 
      n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, 
      n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, 
      n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, 
      n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, 
      n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, 
      n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, 
      n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, 
      n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, 
      n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, 
      n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, 
      n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, 
      n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, 
      n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, 
      n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, 
      n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, 
      n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, 
      n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, 
      n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, 
      n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, 
      n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, 
      n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, 
      n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, 
      n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, 
      n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, 
      n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, 
      n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, 
      n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, 
      n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, 
      n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, 
      n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, 
      n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, 
      n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, 
      n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, 
      n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, 
      n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, 
      n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, 
      n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, 
      n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, 
      n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, 
      n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, 
      n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, 
      n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, 
      n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, 
      n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, 
      n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, 
      n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, 
      n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, 
      n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, 
      n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, 
      n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, 
      n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, 
      n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, 
      n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, 
      n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, 
      n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, 
      n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, 
      n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, 
      n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, 
      n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, 
      n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, 
      n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, 
      n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, 
      n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, 
      n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, 
      n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, 
      n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, 
      n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, 
      n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, 
      n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, 
      n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, 
      n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, 
      n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, 
      n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, 
      n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, 
      n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, 
      n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, 
      n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, 
      n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, 
      n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, 
      n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, 
      n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, 
      n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, 
      n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, 
      n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, 
      n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, 
      n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, 
      n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, 
      n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, 
      n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, 
      n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, 
      n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, 
      n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, 
      n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, 
      n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, 
      n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, 
      n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, 
      n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, 
      n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, 
      n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, 
      n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, 
      n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, 
      n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, 
      n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, 
      n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, 
      n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, 
      n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, 
      n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, 
      n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, 
      n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, 
      n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, 
      n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, 
      n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, 
      n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, 
      n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, 
      n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, 
      n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, 
      n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, 
      n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, 
      n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, 
      n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, 
      n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, 
      n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, 
      n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, 
      n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, 
      n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, 
      n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, 
      n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, 
      n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, 
      n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, 
      n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, 
      n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, 
      n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, 
      n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, 
      n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, 
      n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, 
      n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, 
      n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, 
      n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, 
      n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, 
      n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, 
      n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, 
      n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, 
      n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, 
      n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, 
      n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, 
      n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, 
      n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, 
      n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, 
      n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, 
      n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, 
      n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, 
      n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, 
      n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, 
      n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, 
      n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, 
      n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, 
      n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, 
      n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, 
      n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, 
      n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, 
      n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, 
      n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, 
      n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, 
      n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, 
      n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, 
      n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, 
      n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, 
      n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, 
      n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, 
      n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, 
      n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, 
      n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, 
      n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, 
      n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, 
      n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, 
      n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, 
      n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, 
      n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, 
      n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, 
      n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, 
      n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, 
      n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, 
      n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, 
      n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, 
      n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, 
      n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, 
      n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, 
      n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, 
      n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, 
      n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, 
      n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, 
      n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, 
      n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, 
      n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, 
      n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, 
      n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, 
      n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, 
      n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, 
      n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, 
      n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, 
      n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, 
      n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, 
      n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, 
      n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, 
      n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, 
      n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, 
      n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, 
      n7900, n7901, n7902, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135 : 
      std_logic;

begin
   
   REGISTERS_reg_10_31_inst : DFFR_X1 port map( D => n3430, CK => CLK, RN => 
                           n6444, Q => n5712, QN => n2318);
   REGISTERS_reg_10_30_inst : DFFR_X1 port map( D => n3429, CK => CLK, RN => 
                           n6444, Q => n5713, QN => n2322);
   REGISTERS_reg_10_29_inst : DFFR_X1 port map( D => n3428, CK => CLK, RN => 
                           n6444, Q => n5714, QN => n2326);
   REGISTERS_reg_10_28_inst : DFFR_X1 port map( D => n3427, CK => CLK, RN => 
                           n6444, Q => n5715, QN => n2330);
   REGISTERS_reg_10_27_inst : DFFR_X1 port map( D => n3426, CK => CLK, RN => 
                           n6445, Q => n5716, QN => n2334);
   REGISTERS_reg_10_26_inst : DFFR_X1 port map( D => n3425, CK => CLK, RN => 
                           n6445, Q => n5717, QN => n2338);
   REGISTERS_reg_10_25_inst : DFFR_X1 port map( D => n3424, CK => CLK, RN => 
                           n6445, Q => n5718, QN => n2342);
   REGISTERS_reg_10_24_inst : DFFR_X1 port map( D => n3423, CK => CLK, RN => 
                           n6445, Q => n5719, QN => n2346);
   REGISTERS_reg_10_23_inst : DFFR_X1 port map( D => n3422, CK => CLK, RN => 
                           n6445, Q => n5720, QN => n2350);
   REGISTERS_reg_10_22_inst : DFFR_X1 port map( D => n3421, CK => CLK, RN => 
                           n6445, Q => n5721, QN => n2354);
   REGISTERS_reg_10_21_inst : DFFR_X1 port map( D => n3420, CK => CLK, RN => 
                           n6445, Q => n5722, QN => n2358);
   REGISTERS_reg_10_20_inst : DFFR_X1 port map( D => n3419, CK => CLK, RN => 
                           n6445, Q => n5723, QN => n2362);
   REGISTERS_reg_10_19_inst : DFFR_X1 port map( D => n3418, CK => CLK, RN => 
                           n6443, Q => n5724, QN => n2366);
   REGISTERS_reg_10_18_inst : DFFR_X1 port map( D => n3417, CK => CLK, RN => 
                           n6443, Q => n5725, QN => n2370);
   REGISTERS_reg_10_17_inst : DFFR_X1 port map( D => n3416, CK => CLK, RN => 
                           n6443, Q => n5726, QN => n2374);
   REGISTERS_reg_10_16_inst : DFFR_X1 port map( D => n3415, CK => CLK, RN => 
                           n6443, Q => n5727, QN => n2378);
   REGISTERS_reg_10_15_inst : DFFR_X1 port map( D => n3414, CK => CLK, RN => 
                           n6444, Q => n5728, QN => n2382);
   REGISTERS_reg_10_14_inst : DFFR_X1 port map( D => n3413, CK => CLK, RN => 
                           n6444, Q => n5729, QN => n2386);
   REGISTERS_reg_10_13_inst : DFFR_X1 port map( D => n3412, CK => CLK, RN => 
                           n6444, Q => n5730, QN => n2390);
   REGISTERS_reg_10_12_inst : DFFR_X1 port map( D => n3411, CK => CLK, RN => 
                           n6444, Q => n5731, QN => n2394);
   REGISTERS_reg_10_11_inst : DFFR_X1 port map( D => n3410, CK => CLK, RN => 
                           n6444, Q => n5732, QN => n2398);
   REGISTERS_reg_10_10_inst : DFFR_X1 port map( D => n3409, CK => CLK, RN => 
                           n6444, Q => n5733, QN => n2402);
   REGISTERS_reg_10_9_inst : DFFR_X1 port map( D => n3408, CK => CLK, RN => 
                           n6444, Q => n5734, QN => n2406);
   REGISTERS_reg_10_8_inst : DFFR_X1 port map( D => n3407, CK => CLK, RN => 
                           n6444, Q => n5735, QN => n2410);
   REGISTERS_reg_10_7_inst : DFFR_X1 port map( D => n3406, CK => CLK, RN => 
                           n6443, Q => n5736, QN => n2414);
   REGISTERS_reg_10_6_inst : DFFR_X1 port map( D => n3405, CK => CLK, RN => 
                           n6443, Q => n5737, QN => n2418);
   REGISTERS_reg_10_5_inst : DFFR_X1 port map( D => n3404, CK => CLK, RN => 
                           n6443, Q => n5738, QN => n2422);
   REGISTERS_reg_10_4_inst : DFFR_X1 port map( D => n3403, CK => CLK, RN => 
                           n6443, Q => n5739, QN => n2426);
   REGISTERS_reg_10_3_inst : DFFR_X1 port map( D => n3402, CK => CLK, RN => 
                           n6443, Q => n5740, QN => n2430);
   REGISTERS_reg_10_2_inst : DFFR_X1 port map( D => n3401, CK => CLK, RN => 
                           n6443, Q => n5741, QN => n2434);
   REGISTERS_reg_10_1_inst : DFFR_X1 port map( D => n3400, CK => CLK, RN => 
                           n6443, Q => n5742, QN => n2438);
   REGISTERS_reg_10_0_inst : DFFR_X1 port map( D => n3399, CK => CLK, RN => 
                           n6443, Q => n5743, QN => n2442);
   REGISTERS_reg_11_31_inst : DFFR_X1 port map( D => n3398, CK => CLK, RN => 
                           n6442, Q => n5548, QN => n2319);
   REGISTERS_reg_11_30_inst : DFFR_X1 port map( D => n3397, CK => CLK, RN => 
                           n6442, Q => n5549, QN => n2323);
   REGISTERS_reg_11_29_inst : DFFR_X1 port map( D => n3396, CK => CLK, RN => 
                           n6442, Q => n5550, QN => n2327);
   REGISTERS_reg_11_28_inst : DFFR_X1 port map( D => n3395, CK => CLK, RN => 
                           n6442, Q => n5551, QN => n2331);
   REGISTERS_reg_11_27_inst : DFFR_X1 port map( D => n3394, CK => CLK, RN => 
                           n6441, Q => n5552, QN => n2335);
   REGISTERS_reg_11_26_inst : DFFR_X1 port map( D => n3393, CK => CLK, RN => 
                           n6441, Q => n5553, QN => n2339);
   REGISTERS_reg_11_25_inst : DFFR_X1 port map( D => n3392, CK => CLK, RN => 
                           n6441, Q => n5554, QN => n2343);
   REGISTERS_reg_11_24_inst : DFFR_X1 port map( D => n3391, CK => CLK, RN => 
                           n6441, Q => n5555, QN => n2347);
   REGISTERS_reg_11_23_inst : DFFR_X1 port map( D => n3390, CK => CLK, RN => 
                           n6442, Q => n5556, QN => n2351);
   REGISTERS_reg_11_22_inst : DFFR_X1 port map( D => n3389, CK => CLK, RN => 
                           n6442, Q => n5557, QN => n2355);
   REGISTERS_reg_11_21_inst : DFFR_X1 port map( D => n3388, CK => CLK, RN => 
                           n6442, Q => n5558, QN => n2359);
   REGISTERS_reg_11_20_inst : DFFR_X1 port map( D => n3387, CK => CLK, RN => 
                           n6442, Q => n5559, QN => n2363);
   REGISTERS_reg_11_19_inst : DFFR_X1 port map( D => n3386, CK => CLK, RN => 
                           n6442, Q => n5560, QN => n2367);
   REGISTERS_reg_11_18_inst : DFFR_X1 port map( D => n3385, CK => CLK, RN => 
                           n6442, Q => n5561, QN => n2371);
   REGISTERS_reg_11_17_inst : DFFR_X1 port map( D => n3384, CK => CLK, RN => 
                           n6442, Q => n5562, QN => n2375);
   REGISTERS_reg_11_16_inst : DFFR_X1 port map( D => n3383, CK => CLK, RN => 
                           n6442, Q => n5563, QN => n2379);
   REGISTERS_reg_11_15_inst : DFFR_X1 port map( D => n3382, CK => CLK, RN => 
                           n6440, Q => n5564, QN => n2383);
   REGISTERS_reg_11_14_inst : DFFR_X1 port map( D => n3381, CK => CLK, RN => 
                           n6440, Q => n5565, QN => n2387);
   REGISTERS_reg_11_13_inst : DFFR_X1 port map( D => n3380, CK => CLK, RN => 
                           n6440, Q => n5566, QN => n2391);
   REGISTERS_reg_11_12_inst : DFFR_X1 port map( D => n3379, CK => CLK, RN => 
                           n6440, Q => n5567, QN => n2395);
   REGISTERS_reg_11_11_inst : DFFR_X1 port map( D => n3378, CK => CLK, RN => 
                           n6441, Q => n5568, QN => n2399);
   REGISTERS_reg_11_10_inst : DFFR_X1 port map( D => n3377, CK => CLK, RN => 
                           n6441, Q => n5569, QN => n2403);
   REGISTERS_reg_11_9_inst : DFFR_X1 port map( D => n3376, CK => CLK, RN => 
                           n6441, Q => n5570, QN => n2407);
   REGISTERS_reg_11_8_inst : DFFR_X1 port map( D => n3375, CK => CLK, RN => 
                           n6441, Q => n5571, QN => n2411);
   REGISTERS_reg_11_7_inst : DFFR_X1 port map( D => n3374, CK => CLK, RN => 
                           n6441, Q => n5572, QN => n2415);
   REGISTERS_reg_11_6_inst : DFFR_X1 port map( D => n3373, CK => CLK, RN => 
                           n6441, Q => n5573, QN => n2419);
   REGISTERS_reg_11_5_inst : DFFR_X1 port map( D => n3372, CK => CLK, RN => 
                           n6441, Q => n5574, QN => n2423);
   REGISTERS_reg_11_4_inst : DFFR_X1 port map( D => n3371, CK => CLK, RN => 
                           n6441, Q => n5575, QN => n2427);
   REGISTERS_reg_11_3_inst : DFFR_X1 port map( D => n3370, CK => CLK, RN => 
                           n6452, Q => n5576, QN => n2431);
   REGISTERS_reg_11_2_inst : DFFR_X1 port map( D => n3369, CK => CLK, RN => 
                           n6452, Q => n5577, QN => n2435);
   REGISTERS_reg_11_1_inst : DFFR_X1 port map( D => n3368, CK => CLK, RN => 
                           n6452, Q => n5578, QN => n2439);
   REGISTERS_reg_11_0_inst : DFFR_X1 port map( D => n3367, CK => CLK, RN => 
                           n6452, Q => n5579, QN => n2443);
   REGISTERS_reg_14_31_inst : DFFR_X1 port map( D => n3366, CK => CLK, RN => 
                           n6447, Q => n5236, QN => n2316);
   REGISTERS_reg_14_30_inst : DFFR_X1 port map( D => n3365, CK => CLK, RN => 
                           n6447, Q => n5238, QN => n2320);
   REGISTERS_reg_14_29_inst : DFFR_X1 port map( D => n3364, CK => CLK, RN => 
                           n6447, Q => n5239, QN => n2324);
   REGISTERS_reg_14_28_inst : DFFR_X1 port map( D => n3363, CK => CLK, RN => 
                           n6447, Q => n5240, QN => n2328);
   REGISTERS_reg_14_27_inst : DFFR_X1 port map( D => n3362, CK => CLK, RN => 
                           n6457, Q => n5241, QN => n2332);
   REGISTERS_reg_14_26_inst : DFFR_X1 port map( D => n3361, CK => CLK, RN => 
                           n6457, Q => n5242, QN => n2336);
   REGISTERS_reg_14_25_inst : DFFR_X1 port map( D => n3360, CK => CLK, RN => 
                           n6457, Q => n5243, QN => n2340);
   REGISTERS_reg_14_24_inst : DFFR_X1 port map( D => n3359, CK => CLK, RN => 
                           n6457, Q => n5244, QN => n2344);
   REGISTERS_reg_14_23_inst : DFFR_X1 port map( D => n3358, CK => CLK, RN => 
                           n6458, Q => n5245, QN => n2348);
   REGISTERS_reg_14_22_inst : DFFR_X1 port map( D => n3357, CK => CLK, RN => 
                           n6458, Q => n5246, QN => n2352);
   REGISTERS_reg_14_21_inst : DFFR_X1 port map( D => n3356, CK => CLK, RN => 
                           n6458, Q => n5247, QN => n2356);
   REGISTERS_reg_14_20_inst : DFFR_X1 port map( D => n3355, CK => CLK, RN => 
                           n6458, Q => n5248, QN => n2360);
   REGISTERS_reg_14_19_inst : DFFR_X1 port map( D => n3354, CK => CLK, RN => 
                           n6458, Q => n5249, QN => n2364);
   REGISTERS_reg_14_18_inst : DFFR_X1 port map( D => n3353, CK => CLK, RN => 
                           n6458, Q => n5250, QN => n2368);
   REGISTERS_reg_14_17_inst : DFFR_X1 port map( D => n3352, CK => CLK, RN => 
                           n6458, Q => n5251, QN => n2372);
   REGISTERS_reg_14_16_inst : DFFR_X1 port map( D => n3351, CK => CLK, RN => 
                           n6458, Q => n5252, QN => n2376);
   REGISTERS_reg_14_15_inst : DFFR_X1 port map( D => n3350, CK => CLK, RN => 
                           n6456, Q => n5253, QN => n2380);
   REGISTERS_reg_14_14_inst : DFFR_X1 port map( D => n3349, CK => CLK, RN => 
                           n6456, Q => n5254, QN => n2384);
   REGISTERS_reg_14_13_inst : DFFR_X1 port map( D => n3348, CK => CLK, RN => 
                           n6456, Q => n5255, QN => n2388);
   REGISTERS_reg_14_12_inst : DFFR_X1 port map( D => n3347, CK => CLK, RN => 
                           n6456, Q => n5256, QN => n2392);
   REGISTERS_reg_14_11_inst : DFFR_X1 port map( D => n3346, CK => CLK, RN => 
                           n6457, Q => n5257, QN => n2396);
   REGISTERS_reg_14_10_inst : DFFR_X1 port map( D => n3345, CK => CLK, RN => 
                           n6457, Q => n5258, QN => n2400);
   REGISTERS_reg_14_9_inst : DFFR_X1 port map( D => n3344, CK => CLK, RN => 
                           n6457, Q => n5259, QN => n2404);
   REGISTERS_reg_14_8_inst : DFFR_X1 port map( D => n3343, CK => CLK, RN => 
                           n6457, Q => n5260, QN => n2408);
   REGISTERS_reg_14_7_inst : DFFR_X1 port map( D => n3342, CK => CLK, RN => 
                           n6457, Q => n5261, QN => n2412);
   REGISTERS_reg_14_6_inst : DFFR_X1 port map( D => n3341, CK => CLK, RN => 
                           n6457, Q => n5262, QN => n2416);
   REGISTERS_reg_14_5_inst : DFFR_X1 port map( D => n3340, CK => CLK, RN => 
                           n6457, Q => n5263, QN => n2420);
   REGISTERS_reg_14_4_inst : DFFR_X1 port map( D => n3339, CK => CLK, RN => 
                           n6457, Q => n5264, QN => n2424);
   REGISTERS_reg_14_3_inst : DFFR_X1 port map( D => n3338, CK => CLK, RN => 
                           n6456, Q => n5265, QN => n2428);
   REGISTERS_reg_14_2_inst : DFFR_X1 port map( D => n3337, CK => CLK, RN => 
                           n6456, Q => n5266, QN => n2432);
   REGISTERS_reg_14_1_inst : DFFR_X1 port map( D => n3336, CK => CLK, RN => 
                           n6456, Q => n5267, QN => n2436);
   REGISTERS_reg_14_0_inst : DFFR_X1 port map( D => n3335, CK => CLK, RN => 
                           n6456, Q => n5237, QN => n2440);
   REGISTERS_reg_15_31_inst : DFFR_X1 port map( D => n3334, CK => CLK, RN => 
                           n6455, Q => n5745, QN => n2317);
   REGISTERS_reg_15_30_inst : DFFR_X1 port map( D => n3333, CK => CLK, RN => 
                           n6455, Q => n5746, QN => n2321);
   REGISTERS_reg_15_29_inst : DFFR_X1 port map( D => n3332, CK => CLK, RN => 
                           n6455, Q => n5747, QN => n2325);
   REGISTERS_reg_15_28_inst : DFFR_X1 port map( D => n3331, CK => CLK, RN => 
                           n6455, Q => n5748, QN => n2329);
   REGISTERS_reg_15_27_inst : DFFR_X1 port map( D => n3330, CK => CLK, RN => 
                           n6456, Q => n5749, QN => n2333);
   REGISTERS_reg_15_26_inst : DFFR_X1 port map( D => n3329, CK => CLK, RN => 
                           n6456, Q => n5750, QN => n2337);
   REGISTERS_reg_15_25_inst : DFFR_X1 port map( D => n3328, CK => CLK, RN => 
                           n6456, Q => n5751, QN => n2341);
   REGISTERS_reg_15_24_inst : DFFR_X1 port map( D => n3327, CK => CLK, RN => 
                           n6456, Q => n5752, QN => n2345);
   REGISTERS_reg_15_23_inst : DFFR_X1 port map( D => n3326, CK => CLK, RN => 
                           n6454, Q => n5753, QN => n2349);
   REGISTERS_reg_15_22_inst : DFFR_X1 port map( D => n3325, CK => CLK, RN => 
                           n6454, Q => n5754, QN => n2353);
   REGISTERS_reg_15_21_inst : DFFR_X1 port map( D => n3324, CK => CLK, RN => 
                           n6454, Q => n5755, QN => n2357);
   REGISTERS_reg_15_20_inst : DFFR_X1 port map( D => n3323, CK => CLK, RN => 
                           n6454, Q => n5756, QN => n2361);
   REGISTERS_reg_15_19_inst : DFFR_X1 port map( D => n3322, CK => CLK, RN => 
                           n6455, Q => n5757, QN => n2365);
   REGISTERS_reg_15_18_inst : DFFR_X1 port map( D => n3321, CK => CLK, RN => 
                           n6455, Q => n5758, QN => n2369);
   REGISTERS_reg_15_17_inst : DFFR_X1 port map( D => n3320, CK => CLK, RN => 
                           n6455, Q => n5759, QN => n2373);
   REGISTERS_reg_15_16_inst : DFFR_X1 port map( D => n3319, CK => CLK, RN => 
                           n6455, Q => n5760, QN => n2377);
   REGISTERS_reg_15_15_inst : DFFR_X1 port map( D => n3318, CK => CLK, RN => 
                           n6455, Q => n5761, QN => n2381);
   REGISTERS_reg_15_14_inst : DFFR_X1 port map( D => n3317, CK => CLK, RN => 
                           n6455, Q => n5762, QN => n2385);
   REGISTERS_reg_15_13_inst : DFFR_X1 port map( D => n3316, CK => CLK, RN => 
                           n6455, Q => n5763, QN => n2389);
   REGISTERS_reg_15_12_inst : DFFR_X1 port map( D => n3315, CK => CLK, RN => 
                           n6455, Q => n5764, QN => n2393);
   REGISTERS_reg_15_11_inst : DFFR_X1 port map( D => n3314, CK => CLK, RN => 
                           n6453, Q => n5765, QN => n2397);
   REGISTERS_reg_15_10_inst : DFFR_X1 port map( D => n3313, CK => CLK, RN => 
                           n6453, Q => n5766, QN => n2401);
   REGISTERS_reg_15_9_inst : DFFR_X1 port map( D => n3312, CK => CLK, RN => 
                           n6453, Q => n5767, QN => n2405);
   REGISTERS_reg_15_8_inst : DFFR_X1 port map( D => n3311, CK => CLK, RN => 
                           n6453, Q => n5768, QN => n2409);
   REGISTERS_reg_15_7_inst : DFFR_X1 port map( D => n3310, CK => CLK, RN => 
                           n6454, Q => n5769, QN => n2413);
   REGISTERS_reg_15_6_inst : DFFR_X1 port map( D => n3309, CK => CLK, RN => 
                           n6454, Q => n5770, QN => n2417);
   REGISTERS_reg_15_5_inst : DFFR_X1 port map( D => n3308, CK => CLK, RN => 
                           n6454, Q => n5771, QN => n2421);
   REGISTERS_reg_15_4_inst : DFFR_X1 port map( D => n3307, CK => CLK, RN => 
                           n6454, Q => n5772, QN => n2425);
   REGISTERS_reg_15_3_inst : DFFR_X1 port map( D => n3306, CK => CLK, RN => 
                           n6454, Q => n5773, QN => n2429);
   REGISTERS_reg_15_2_inst : DFFR_X1 port map( D => n3305, CK => CLK, RN => 
                           n6454, Q => n5774, QN => n2433);
   REGISTERS_reg_15_1_inst : DFFR_X1 port map( D => n3304, CK => CLK, RN => 
                           n6454, Q => n5775, QN => n2437);
   REGISTERS_reg_15_0_inst : DFFR_X1 port map( D => n3303, CK => CLK, RN => 
                           n6454, Q => n5776, QN => n2441);
   REGISTERS_reg_18_30_inst : DFFR_X1 port map( D => n3301, CK => CLK, RN => 
                           n6460, Q => n5453, QN => n2250);
   REGISTERS_reg_18_29_inst : DFFR_X1 port map( D => n3300, CK => CLK, RN => 
                           n6460, Q => n5454, QN => n2249);
   REGISTERS_reg_18_28_inst : DFFR_X1 port map( D => n3299, CK => CLK, RN => 
                           n6460, Q => n5455, QN => n2248);
   REGISTERS_reg_18_27_inst : DFFR_X1 port map( D => n3298, CK => CLK, RN => 
                           n6460, Q => n5456, QN => n2247);
   REGISTERS_reg_18_26_inst : DFFR_X1 port map( D => n3297, CK => CLK, RN => 
                           n6460, Q => n5457, QN => n2246);
   REGISTERS_reg_18_25_inst : DFFR_X1 port map( D => n3296, CK => CLK, RN => 
                           n6460, Q => n5458, QN => n2245);
   REGISTERS_reg_18_24_inst : DFFR_X1 port map( D => n3295, CK => CLK, RN => 
                           n6460, Q => n5459, QN => n2244);
   REGISTERS_reg_18_23_inst : DFFR_X1 port map( D => n3294, CK => CLK, RN => 
                           n6458, Q => n5460, QN => n2243);
   REGISTERS_reg_18_22_inst : DFFR_X1 port map( D => n3293, CK => CLK, RN => 
                           n6458, Q => n5461, QN => n2242);
   REGISTERS_reg_18_21_inst : DFFR_X1 port map( D => n3292, CK => CLK, RN => 
                           n6458, Q => n5462, QN => n2241);
   REGISTERS_reg_18_20_inst : DFFR_X1 port map( D => n3291, CK => CLK, RN => 
                           n6458, Q => n5463, QN => n2240);
   REGISTERS_reg_18_19_inst : DFFR_X1 port map( D => n3290, CK => CLK, RN => 
                           n6459, Q => n5464, QN => n2239);
   REGISTERS_reg_18_18_inst : DFFR_X1 port map( D => n3289, CK => CLK, RN => 
                           n6459, Q => n5465, QN => n2238);
   REGISTERS_reg_18_17_inst : DFFR_X1 port map( D => n3288, CK => CLK, RN => 
                           n6459, Q => n5466, QN => n2237);
   REGISTERS_reg_18_16_inst : DFFR_X1 port map( D => n3287, CK => CLK, RN => 
                           n6459, Q => n5467, QN => n2236);
   REGISTERS_reg_18_15_inst : DFFR_X1 port map( D => n3286, CK => CLK, RN => 
                           n6459, Q => n5468, QN => n2235);
   REGISTERS_reg_18_14_inst : DFFR_X1 port map( D => n3285, CK => CLK, RN => 
                           n6459, Q => n5469, QN => n2234);
   REGISTERS_reg_18_13_inst : DFFR_X1 port map( D => n3284, CK => CLK, RN => 
                           n6459, Q => n5470, QN => n2233);
   REGISTERS_reg_18_12_inst : DFFR_X1 port map( D => n3283, CK => CLK, RN => 
                           n6459, Q => n5471, QN => n2232);
   REGISTERS_reg_18_11_inst : DFFR_X1 port map( D => n3282, CK => CLK, RN => 
                           n6387, Q => n5472, QN => n2231);
   REGISTERS_reg_18_10_inst : DFFR_X1 port map( D => n3281, CK => CLK, RN => 
                           n6387, Q => n5473, QN => n2230);
   REGISTERS_reg_18_9_inst : DFFR_X1 port map( D => n3280, CK => CLK, RN => 
                           n6387, Q => n5474, QN => n2229);
   REGISTERS_reg_18_8_inst : DFFR_X1 port map( D => n3279, CK => CLK, RN => 
                           n6387, Q => n5475, QN => n2228);
   REGISTERS_reg_18_7_inst : DFFR_X1 port map( D => n3278, CK => CLK, RN => 
                           n6387, Q => n5476, QN => n2227);
   REGISTERS_reg_18_6_inst : DFFR_X1 port map( D => n3277, CK => CLK, RN => 
                           n6387, Q => n5477, QN => n2226);
   REGISTERS_reg_18_5_inst : DFFR_X1 port map( D => n3276, CK => CLK, RN => 
                           n6387, Q => n5478, QN => n2225);
   REGISTERS_reg_18_4_inst : DFFR_X1 port map( D => n3275, CK => CLK, RN => 
                           n6387, Q => n5479, QN => n2224);
   REGISTERS_reg_18_3_inst : DFFR_X1 port map( D => n3274, CK => CLK, RN => 
                           n6387, Q => n5480, QN => n2223);
   REGISTERS_reg_18_2_inst : DFFR_X1 port map( D => n3273, CK => CLK, RN => 
                           n6387, Q => n5481, QN => n2222);
   REGISTERS_reg_18_1_inst : DFFR_X1 port map( D => n3272, CK => CLK, RN => 
                           n6388, Q => n5482, QN => n2221);
   REGISTERS_reg_18_0_inst : DFFR_X1 port map( D => n3271, CK => CLK, RN => 
                           n6388, Q => n5486, QN => n2220);
   REGISTERS_reg_19_31_inst : DFFR_X1 port map( D => n3270, CK => CLK, RN => 
                           n6386, Q => n5515, QN => n2219);
   REGISTERS_reg_19_30_inst : DFFR_X1 port map( D => n3269, CK => CLK, RN => 
                           n6386, Q => n5516, QN => n2218);
   REGISTERS_reg_19_29_inst : DFFR_X1 port map( D => n3268, CK => CLK, RN => 
                           n6386, Q => n5517, QN => n2217);
   REGISTERS_reg_19_28_inst : DFFR_X1 port map( D => n3267, CK => CLK, RN => 
                           n6386, Q => n5518, QN => n2216);
   REGISTERS_reg_19_27_inst : DFFR_X1 port map( D => n3266, CK => CLK, RN => 
                           n6386, Q => n5519, QN => n2215);
   REGISTERS_reg_19_26_inst : DFFR_X1 port map( D => n3265, CK => CLK, RN => 
                           n6386, Q => n5520, QN => n2214);
   REGISTERS_reg_19_25_inst : DFFR_X1 port map( D => n3264, CK => CLK, RN => 
                           n6386, Q => n5521, QN => n2213);
   REGISTERS_reg_19_24_inst : DFFR_X1 port map( D => n3263, CK => CLK, RN => 
                           n6386, Q => n5522, QN => n2212);
   REGISTERS_reg_19_23_inst : DFFR_X1 port map( D => n3262, CK => CLK, RN => 
                           n6386, Q => n5523, QN => n2211);
   REGISTERS_reg_19_22_inst : DFFR_X1 port map( D => n3261, CK => CLK, RN => 
                           n6386, Q => n5524, QN => n2210);
   REGISTERS_reg_19_21_inst : DFFR_X1 port map( D => n3260, CK => CLK, RN => 
                           n6387, Q => n5525, QN => n2209);
   REGISTERS_reg_19_20_inst : DFFR_X1 port map( D => n3259, CK => CLK, RN => 
                           n6387, Q => n5526, QN => n2208);
   REGISTERS_reg_19_19_inst : DFFR_X1 port map( D => n3258, CK => CLK, RN => 
                           n6385, Q => n5527, QN => n2207);
   REGISTERS_reg_19_18_inst : DFFR_X1 port map( D => n3257, CK => CLK, RN => 
                           n6385, Q => n5528, QN => n2206);
   REGISTERS_reg_19_17_inst : DFFR_X1 port map( D => n3256, CK => CLK, RN => 
                           n6385, Q => n5529, QN => n2205);
   REGISTERS_reg_19_16_inst : DFFR_X1 port map( D => n3255, CK => CLK, RN => 
                           n6385, Q => n5530, QN => n2204);
   REGISTERS_reg_19_15_inst : DFFR_X1 port map( D => n3254, CK => CLK, RN => 
                           n6385, Q => n5531, QN => n2203);
   REGISTERS_reg_19_14_inst : DFFR_X1 port map( D => n3253, CK => CLK, RN => 
                           n6385, Q => n5532, QN => n2202);
   REGISTERS_reg_19_13_inst : DFFR_X1 port map( D => n3252, CK => CLK, RN => 
                           n6385, Q => n5533, QN => n2201);
   REGISTERS_reg_19_12_inst : DFFR_X1 port map( D => n3251, CK => CLK, RN => 
                           n6385, Q => n5534, QN => n2200);
   REGISTERS_reg_19_11_inst : DFFR_X1 port map( D => n3250, CK => CLK, RN => 
                           n6385, Q => n5535, QN => n2199);
   REGISTERS_reg_19_10_inst : DFFR_X1 port map( D => n3249, CK => CLK, RN => 
                           n6385, Q => n5536, QN => n2198);
   REGISTERS_reg_19_9_inst : DFFR_X1 port map( D => n3248, CK => CLK, RN => 
                           n6386, Q => n5537, QN => n2197);
   REGISTERS_reg_19_8_inst : DFFR_X1 port map( D => n3247, CK => CLK, RN => 
                           n6386, Q => n5538, QN => n2196);
   REGISTERS_reg_19_7_inst : DFFR_X1 port map( D => n3246, CK => CLK, RN => 
                           n6385, Q => n5539, QN => n2195);
   REGISTERS_reg_19_6_inst : DFFR_X1 port map( D => n3245, CK => CLK, RN => 
                           n6384, Q => n5540, QN => n2194);
   REGISTERS_reg_19_5_inst : DFFR_X1 port map( D => n3244, CK => CLK, RN => 
                           n6384, Q => n5541, QN => n2193);
   REGISTERS_reg_19_4_inst : DFFR_X1 port map( D => n3243, CK => CLK, RN => 
                           n6384, Q => n5542, QN => n2192);
   REGISTERS_reg_19_3_inst : DFFR_X1 port map( D => n3242, CK => CLK, RN => 
                           n6384, Q => n5543, QN => n2191);
   REGISTERS_reg_19_2_inst : DFFR_X1 port map( D => n3241, CK => CLK, RN => 
                           n6384, Q => n5544, QN => n2190);
   REGISTERS_reg_19_1_inst : DFFR_X1 port map( D => n3240, CK => CLK, RN => 
                           n6384, Q => n5545, QN => n2189);
   REGISTERS_reg_19_0_inst : DFFR_X1 port map( D => n3239, CK => CLK, RN => 
                           n6385, Q => n5680, QN => n2188);
   REGISTERS_reg_25_31_inst : DFFR_X1 port map( D => n3142, CK => CLK, RN => 
                           n6394, Q => n5137, QN => n2187);
   REGISTERS_reg_25_30_inst : DFFR_X1 port map( D => n3141, CK => CLK, RN => 
                           n6394, Q => n5138, QN => n2186);
   REGISTERS_reg_25_29_inst : DFFR_X1 port map( D => n3140, CK => CLK, RN => 
                           n6394, Q => n5139, QN => n2185);
   REGISTERS_reg_25_28_inst : DFFR_X1 port map( D => n3139, CK => CLK, RN => 
                           n6394, Q => n5140, QN => n2184);
   REGISTERS_reg_25_27_inst : DFFR_X1 port map( D => n3138, CK => CLK, RN => 
                           n6394, Q => n5141, QN => n2183);
   REGISTERS_reg_25_26_inst : DFFR_X1 port map( D => n3137, CK => CLK, RN => 
                           n6394, Q => n5142, QN => n2182);
   REGISTERS_reg_25_25_inst : DFFR_X1 port map( D => n3136, CK => CLK, RN => 
                           n6394, Q => n5143, QN => n2181);
   REGISTERS_reg_25_24_inst : DFFR_X1 port map( D => n3135, CK => CLK, RN => 
                           n6394, Q => n5144, QN => n2180);
   REGISTERS_reg_25_23_inst : DFFR_X1 port map( D => n3134, CK => CLK, RN => 
                           n6394, Q => n5145, QN => n2179);
   REGISTERS_reg_25_22_inst : DFFR_X1 port map( D => n3133, CK => CLK, RN => 
                           n6394, Q => n5146, QN => n2178);
   REGISTERS_reg_25_21_inst : DFFR_X1 port map( D => n3132, CK => CLK, RN => 
                           n6395, Q => n5147, QN => n2177);
   REGISTERS_reg_25_20_inst : DFFR_X1 port map( D => n3131, CK => CLK, RN => 
                           n6395, Q => n5148, QN => n2176);
   REGISTERS_reg_25_19_inst : DFFR_X1 port map( D => n3130, CK => CLK, RN => 
                           n6405, Q => n5149, QN => n2175);
   REGISTERS_reg_25_18_inst : DFFR_X1 port map( D => n3129, CK => CLK, RN => 
                           n6405, Q => n5150, QN => n2174);
   REGISTERS_reg_25_17_inst : DFFR_X1 port map( D => n3128, CK => CLK, RN => 
                           n6405, Q => n5151, QN => n2173);
   REGISTERS_reg_25_16_inst : DFFR_X1 port map( D => n3127, CK => CLK, RN => 
                           n6405, Q => n5152, QN => n2172);
   REGISTERS_reg_25_15_inst : DFFR_X1 port map( D => n3126, CK => CLK, RN => 
                           n6405, Q => n5153, QN => n2171);
   REGISTERS_reg_25_14_inst : DFFR_X1 port map( D => n3125, CK => CLK, RN => 
                           n6405, Q => n5154, QN => n2170);
   REGISTERS_reg_25_13_inst : DFFR_X1 port map( D => n3124, CK => CLK, RN => 
                           n6405, Q => n5155, QN => n2169);
   REGISTERS_reg_25_12_inst : DFFR_X1 port map( D => n3123, CK => CLK, RN => 
                           n6405, Q => n5156, QN => n2168);
   REGISTERS_reg_25_11_inst : DFFR_X1 port map( D => n3122, CK => CLK, RN => 
                           n6405, Q => n5157, QN => n2167);
   REGISTERS_reg_25_10_inst : DFFR_X1 port map( D => n3121, CK => CLK, RN => 
                           n6405, Q => n5158, QN => n2166);
   REGISTERS_reg_25_9_inst : DFFR_X1 port map( D => n3120, CK => CLK, RN => 
                           n6405, Q => n5159, QN => n2165);
   REGISTERS_reg_25_8_inst : DFFR_X1 port map( D => n3119, CK => CLK, RN => 
                           n6405, Q => n5160, QN => n2164);
   REGISTERS_reg_25_7_inst : DFFR_X1 port map( D => n3118, CK => CLK, RN => 
                           n6404, Q => n5161, QN => n2163);
   REGISTERS_reg_25_6_inst : DFFR_X1 port map( D => n3117, CK => CLK, RN => 
                           n6404, Q => n5162, QN => n2162);
   REGISTERS_reg_25_5_inst : DFFR_X1 port map( D => n3116, CK => CLK, RN => 
                           n6404, Q => n5163, QN => n2161);
   REGISTERS_reg_25_4_inst : DFFR_X1 port map( D => n3115, CK => CLK, RN => 
                           n6404, Q => n5164, QN => n2160);
   REGISTERS_reg_25_3_inst : DFFR_X1 port map( D => n3114, CK => CLK, RN => 
                           n6404, Q => n5165, QN => n2159);
   REGISTERS_reg_25_2_inst : DFFR_X1 port map( D => n3113, CK => CLK, RN => 
                           n6404, Q => n5166, QN => n2158);
   REGISTERS_reg_25_1_inst : DFFR_X1 port map( D => n3112, CK => CLK, RN => 
                           n6404, Q => n5167, QN => n2157);
   REGISTERS_reg_25_0_inst : DFFR_X1 port map( D => n3111, CK => CLK, RN => 
                           n6404, Q => n5171, QN => n2156);
   REGISTERS_reg_29_31_inst : DFFR_X1 port map( D => n3078, CK => CLK, RN => 
                           n6408, Q => n5234, QN => n2059);
   REGISTERS_reg_29_30_inst : DFFR_X1 port map( D => n3077, CK => CLK, RN => 
                           n6408, Q => n5268, QN => n2058);
   REGISTERS_reg_29_29_inst : DFFR_X1 port map( D => n3076, CK => CLK, RN => 
                           n6408, Q => n5269, QN => n2057);
   REGISTERS_reg_29_28_inst : DFFR_X1 port map( D => n3075, CK => CLK, RN => 
                           n6408, Q => n5270, QN => n2056);
   REGISTERS_reg_29_27_inst : DFFR_X1 port map( D => n3074, CK => CLK, RN => 
                           n6407, Q => n5271, QN => n2055);
   REGISTERS_reg_29_26_inst : DFFR_X1 port map( D => n3073, CK => CLK, RN => 
                           n6407, Q => n5272, QN => n2054);
   REGISTERS_reg_29_25_inst : DFFR_X1 port map( D => n3072, CK => CLK, RN => 
                           n6407, Q => n5273, QN => n2053);
   REGISTERS_reg_29_24_inst : DFFR_X1 port map( D => n3071, CK => CLK, RN => 
                           n6407, Q => n5274, QN => n2052);
   REGISTERS_reg_29_23_inst : DFFR_X1 port map( D => n3070, CK => CLK, RN => 
                           n6407, Q => n5275, QN => n2051);
   REGISTERS_reg_29_22_inst : DFFR_X1 port map( D => n3069, CK => CLK, RN => 
                           n6407, Q => n5276, QN => n2050);
   REGISTERS_reg_29_21_inst : DFFR_X1 port map( D => n3068, CK => CLK, RN => 
                           n6407, Q => n5277, QN => n2049);
   REGISTERS_reg_29_20_inst : DFFR_X1 port map( D => n3067, CK => CLK, RN => 
                           n6407, Q => n5278, QN => n2048);
   REGISTERS_reg_29_19_inst : DFFR_X1 port map( D => n3066, CK => CLK, RN => 
                           n6407, Q => n5279, QN => n2047);
   REGISTERS_reg_29_18_inst : DFFR_X1 port map( D => n3065, CK => CLK, RN => 
                           n6407, Q => n5280, QN => n2046);
   REGISTERS_reg_29_17_inst : DFFR_X1 port map( D => n3064, CK => CLK, RN => 
                           n6407, Q => n5281, QN => n2045);
   REGISTERS_reg_29_16_inst : DFFR_X1 port map( D => n3063, CK => CLK, RN => 
                           n6407, Q => n5282, QN => n2044);
   REGISTERS_reg_29_15_inst : DFFR_X1 port map( D => n3062, CK => CLK, RN => 
                           n6406, Q => n5283, QN => n2043);
   REGISTERS_reg_29_14_inst : DFFR_X1 port map( D => n3061, CK => CLK, RN => 
                           n6406, Q => n5284, QN => n2042);
   REGISTERS_reg_29_13_inst : DFFR_X1 port map( D => n3060, CK => CLK, RN => 
                           n6406, Q => n5285, QN => n2041);
   REGISTERS_reg_29_12_inst : DFFR_X1 port map( D => n3059, CK => CLK, RN => 
                           n6406, Q => n5286, QN => n2040);
   REGISTERS_reg_29_11_inst : DFFR_X1 port map( D => n3058, CK => CLK, RN => 
                           n6406, Q => n5287, QN => n2039);
   REGISTERS_reg_29_10_inst : DFFR_X1 port map( D => n3057, CK => CLK, RN => 
                           n6406, Q => n5288, QN => n2038);
   REGISTERS_reg_29_9_inst : DFFR_X1 port map( D => n3056, CK => CLK, RN => 
                           n6406, Q => n5289, QN => n2037);
   REGISTERS_reg_29_8_inst : DFFR_X1 port map( D => n3055, CK => CLK, RN => 
                           n6406, Q => n5290, QN => n2036);
   REGISTERS_reg_29_7_inst : DFFR_X1 port map( D => n3054, CK => CLK, RN => 
                           n6406, Q => n5291, QN => n2035);
   REGISTERS_reg_29_6_inst : DFFR_X1 port map( D => n3053, CK => CLK, RN => 
                           n6406, Q => n5292, QN => n2034);
   REGISTERS_reg_29_5_inst : DFFR_X1 port map( D => n3052, CK => CLK, RN => 
                           n6406, Q => n5293, QN => n2033);
   REGISTERS_reg_29_4_inst : DFFR_X1 port map( D => n3051, CK => CLK, RN => 
                           n6406, Q => n5294, QN => n2032);
   REGISTERS_reg_29_3_inst : DFFR_X1 port map( D => n3050, CK => CLK, RN => 
                           n6416, Q => n5295, QN => n2031);
   REGISTERS_reg_29_2_inst : DFFR_X1 port map( D => n3049, CK => CLK, RN => 
                           n6416, Q => n5296, QN => n2030);
   REGISTERS_reg_29_1_inst : DFFR_X1 port map( D => n3048, CK => CLK, RN => 
                           n6416, Q => n5297, QN => n2029);
   REGISTERS_reg_29_0_inst : DFFR_X1 port map( D => n3047, CK => CLK, RN => 
                           n6416, Q => n5235, QN => n2028);
   OUT2_reg_31_inst : DFF_X1 port map( D => n3015, CK => CLK, Q => OUT2(31), QN
                           => n7551);
   OUT2_reg_30_inst : DFF_X1 port map( D => n3016, CK => CLK, Q => OUT2(30), QN
                           => n2655);
   OUT2_reg_29_inst : DFF_X1 port map( D => n3017, CK => CLK, Q => OUT2(29), QN
                           => n2656);
   OUT2_reg_28_inst : DFF_X1 port map( D => n3018, CK => CLK, Q => OUT2(28), QN
                           => n2657);
   OUT2_reg_27_inst : DFF_X1 port map( D => n3019, CK => CLK, Q => OUT2(27), QN
                           => n2658);
   OUT2_reg_26_inst : DFF_X1 port map( D => n3020, CK => CLK, Q => OUT2(26), QN
                           => n2659);
   OUT2_reg_25_inst : DFF_X1 port map( D => n3021, CK => CLK, Q => OUT2(25), QN
                           => n2660);
   OUT2_reg_24_inst : DFF_X1 port map( D => n3022, CK => CLK, Q => OUT2(24), QN
                           => n2661);
   OUT2_reg_23_inst : DFF_X1 port map( D => n3023, CK => CLK, Q => OUT2(23), QN
                           => n2662);
   OUT2_reg_22_inst : DFF_X1 port map( D => n3024, CK => CLK, Q => OUT2(22), QN
                           => n2663);
   OUT2_reg_21_inst : DFF_X1 port map( D => n3025, CK => CLK, Q => OUT2(21), QN
                           => n2664);
   OUT2_reg_20_inst : DFF_X1 port map( D => n3026, CK => CLK, Q => OUT2(20), QN
                           => n2665);
   OUT2_reg_19_inst : DFF_X1 port map( D => n3027, CK => CLK, Q => OUT2(19), QN
                           => n2666);
   OUT2_reg_18_inst : DFF_X1 port map( D => n3028, CK => CLK, Q => OUT2(18), QN
                           => n2667);
   OUT2_reg_17_inst : DFF_X1 port map( D => n3029, CK => CLK, Q => OUT2(17), QN
                           => n2668);
   OUT2_reg_16_inst : DFF_X1 port map( D => n3030, CK => CLK, Q => OUT2(16), QN
                           => n2669);
   OUT2_reg_15_inst : DFF_X1 port map( D => n3031, CK => CLK, Q => OUT2(15), QN
                           => n2670);
   OUT2_reg_14_inst : DFF_X1 port map( D => n3032, CK => CLK, Q => OUT2(14), QN
                           => n2671);
   OUT2_reg_13_inst : DFF_X1 port map( D => n3033, CK => CLK, Q => OUT2(13), QN
                           => n2672);
   OUT2_reg_12_inst : DFF_X1 port map( D => n3034, CK => CLK, Q => OUT2(12), QN
                           => n2673);
   OUT2_reg_11_inst : DFF_X1 port map( D => n3035, CK => CLK, Q => OUT2(11), QN
                           => n2674);
   OUT2_reg_10_inst : DFF_X1 port map( D => n3036, CK => CLK, Q => OUT2(10), QN
                           => n2675);
   OUT2_reg_9_inst : DFF_X1 port map( D => n3037, CK => CLK, Q => OUT2(9), QN 
                           => n2676);
   OUT2_reg_8_inst : DFF_X1 port map( D => n3038, CK => CLK, Q => OUT2(8), QN 
                           => n2677);
   OUT2_reg_7_inst : DFF_X1 port map( D => n3039, CK => CLK, Q => OUT2(7), QN 
                           => n2678);
   OUT2_reg_6_inst : DFF_X1 port map( D => n3040, CK => CLK, Q => OUT2(6), QN 
                           => n2679);
   OUT2_reg_5_inst : DFF_X1 port map( D => n3041, CK => CLK, Q => OUT2(5), QN 
                           => n2680);
   OUT2_reg_4_inst : DFF_X1 port map( D => n3042, CK => CLK, Q => OUT2(4), QN 
                           => n2681);
   OUT2_reg_3_inst : DFF_X1 port map( D => n3043, CK => CLK, Q => OUT2(3), QN 
                           => n2682);
   OUT2_reg_2_inst : DFF_X1 port map( D => n3044, CK => CLK, Q => OUT2(2), QN 
                           => n2683);
   OUT2_reg_1_inst : DFF_X1 port map( D => n3045, CK => CLK, Q => OUT2(1), QN 
                           => n2684);
   OUT2_reg_0_inst : DFF_X1 port map( D => n3046, CK => CLK, Q => OUT2(0), QN 
                           => n2685);
   OUT1_reg_31_inst : DFF_X1 port map( D => n3014, CK => CLK, Q => OUT1(31), QN
                           => n2653);
   OUT1_reg_30_inst : DFF_X1 port map( D => n3013, CK => CLK, Q => OUT1(30), QN
                           => n2652);
   OUT1_reg_29_inst : DFF_X1 port map( D => n3012, CK => CLK, Q => OUT1(29), QN
                           => n2651);
   OUT1_reg_28_inst : DFF_X1 port map( D => n3011, CK => CLK, Q => OUT1(28), QN
                           => n2650);
   OUT1_reg_27_inst : DFF_X1 port map( D => n3010, CK => CLK, Q => OUT1(27), QN
                           => n2649);
   OUT1_reg_26_inst : DFF_X1 port map( D => n3009, CK => CLK, Q => OUT1(26), QN
                           => n2648);
   OUT1_reg_25_inst : DFF_X1 port map( D => n3008, CK => CLK, Q => OUT1(25), QN
                           => n2647);
   OUT1_reg_24_inst : DFF_X1 port map( D => n3007, CK => CLK, Q => OUT1(24), QN
                           => n2646);
   OUT1_reg_23_inst : DFF_X1 port map( D => n3006, CK => CLK, Q => OUT1(23), QN
                           => n2645);
   OUT1_reg_22_inst : DFF_X1 port map( D => n3005, CK => CLK, Q => OUT1(22), QN
                           => n2644);
   OUT1_reg_21_inst : DFF_X1 port map( D => n3004, CK => CLK, Q => OUT1(21), QN
                           => n2643);
   OUT1_reg_20_inst : DFF_X1 port map( D => n3003, CK => CLK, Q => OUT1(20), QN
                           => n2642);
   OUT1_reg_19_inst : DFF_X1 port map( D => n3002, CK => CLK, Q => OUT1(19), QN
                           => n2641);
   OUT1_reg_18_inst : DFF_X1 port map( D => n3001, CK => CLK, Q => OUT1(18), QN
                           => n2640);
   OUT1_reg_17_inst : DFF_X1 port map( D => n3000, CK => CLK, Q => OUT1(17), QN
                           => n2639);
   OUT1_reg_16_inst : DFF_X1 port map( D => n2999, CK => CLK, Q => OUT1(16), QN
                           => n2638);
   OUT1_reg_15_inst : DFF_X1 port map( D => n2998, CK => CLK, Q => OUT1(15), QN
                           => n2637);
   OUT1_reg_14_inst : DFF_X1 port map( D => n2997, CK => CLK, Q => OUT1(14), QN
                           => n2636);
   OUT1_reg_13_inst : DFF_X1 port map( D => n2996, CK => CLK, Q => OUT1(13), QN
                           => n2635);
   OUT1_reg_12_inst : DFF_X1 port map( D => n2995, CK => CLK, Q => OUT1(12), QN
                           => n2634);
   OUT1_reg_11_inst : DFF_X1 port map( D => n2994, CK => CLK, Q => OUT1(11), QN
                           => n2633);
   OUT1_reg_10_inst : DFF_X1 port map( D => n2993, CK => CLK, Q => OUT1(10), QN
                           => n2632);
   OUT1_reg_9_inst : DFF_X1 port map( D => n2992, CK => CLK, Q => OUT1(9), QN 
                           => n2631);
   OUT1_reg_8_inst : DFF_X1 port map( D => n2991, CK => CLK, Q => OUT1(8), QN 
                           => n2630);
   OUT1_reg_7_inst : DFF_X1 port map( D => n2990, CK => CLK, Q => OUT1(7), QN 
                           => n2629);
   OUT1_reg_6_inst : DFF_X1 port map( D => n2989, CK => CLK, Q => OUT1(6), QN 
                           => n2628);
   OUT1_reg_5_inst : DFF_X1 port map( D => n2988, CK => CLK, Q => OUT1(5), QN 
                           => n2627);
   OUT1_reg_4_inst : DFF_X1 port map( D => n2987, CK => CLK, Q => OUT1(4), QN 
                           => n2626);
   OUT1_reg_3_inst : DFF_X1 port map( D => n2986, CK => CLK, Q => OUT1(3), QN 
                           => n2625);
   OUT1_reg_2_inst : DFF_X1 port map( D => n2985, CK => CLK, Q => OUT1(2), QN 
                           => n2624);
   OUT1_reg_1_inst : DFF_X1 port map( D => n2984, CK => CLK, Q => OUT1(1), QN 
                           => n2623);
   OUT1_reg_0_inst : DFF_X1 port map( D => n2983, CK => CLK, Q => OUT1(0), QN 
                           => n6512);
   REGISTERS_reg_24_31_inst : DFFR_X1 port map( D => n3174, CK => CLK, RN => 
                           n6382, Q => n2877, QN => n5880);
   REGISTERS_reg_24_30_inst : DFFR_X1 port map( D => n7656, CK => CLK, RN => 
                           n6398, Q => n2876, QN => n5881);
   REGISTERS_reg_24_29_inst : DFFR_X1 port map( D => n7657, CK => CLK, RN => 
                           n6397, Q => n2875, QN => n5882);
   REGISTERS_reg_24_28_inst : DFFR_X1 port map( D => n7658, CK => CLK, RN => 
                           n6397, Q => n2874, QN => n5883);
   REGISTERS_reg_24_27_inst : DFFR_X1 port map( D => n7659, CK => CLK, RN => 
                           n6397, Q => n2873, QN => n5884);
   REGISTERS_reg_24_26_inst : DFFR_X1 port map( D => n7660, CK => CLK, RN => 
                           n6397, Q => n2872, QN => n5885);
   REGISTERS_reg_24_25_inst : DFFR_X1 port map( D => n7661, CK => CLK, RN => 
                           n6397, Q => n2871, QN => n5886);
   REGISTERS_reg_24_24_inst : DFFR_X1 port map( D => n7662, CK => CLK, RN => 
                           n6397, Q => n2870, QN => n5887);
   REGISTERS_reg_24_23_inst : DFFR_X1 port map( D => n7663, CK => CLK, RN => 
                           n6397, Q => n2869, QN => n5888);
   REGISTERS_reg_24_22_inst : DFFR_X1 port map( D => n7664, CK => CLK, RN => 
                           n6397, Q => n2868, QN => n5889);
   REGISTERS_reg_24_21_inst : DFFR_X1 port map( D => n7665, CK => CLK, RN => 
                           n6396, Q => n2867, QN => n5890);
   REGISTERS_reg_24_20_inst : DFFR_X1 port map( D => n7666, CK => CLK, RN => 
                           n6396, Q => n2866, QN => n5891);
   REGISTERS_reg_24_19_inst : DFFR_X1 port map( D => n7667, CK => CLK, RN => 
                           n6396, Q => n2865, QN => n5892);
   REGISTERS_reg_24_18_inst : DFFR_X1 port map( D => n7668, CK => CLK, RN => 
                           n6396, Q => n2864, QN => n5893);
   REGISTERS_reg_24_17_inst : DFFR_X1 port map( D => n7669, CK => CLK, RN => 
                           n6396, Q => n2863, QN => n5894);
   REGISTERS_reg_24_16_inst : DFFR_X1 port map( D => n7670, CK => CLK, RN => 
                           n6396, Q => n2862, QN => n5895);
   REGISTERS_reg_24_15_inst : DFFR_X1 port map( D => n7671, CK => CLK, RN => 
                           n6396, Q => n2861, QN => n5896);
   REGISTERS_reg_24_14_inst : DFFR_X1 port map( D => n7672, CK => CLK, RN => 
                           n6396, Q => n2860, QN => n5897);
   REGISTERS_reg_24_13_inst : DFFR_X1 port map( D => n7673, CK => CLK, RN => 
                           n6396, Q => n2859, QN => n5898);
   REGISTERS_reg_24_12_inst : DFFR_X1 port map( D => n7674, CK => CLK, RN => 
                           n6396, Q => n2858, QN => n5899);
   REGISTERS_reg_24_11_inst : DFFR_X1 port map( D => n7675, CK => CLK, RN => 
                           n6396, Q => n2857, QN => n5900);
   REGISTERS_reg_24_10_inst : DFFR_X1 port map( D => n7676, CK => CLK, RN => 
                           n6396, Q => n2856, QN => n5901);
   REGISTERS_reg_24_9_inst : DFFR_X1 port map( D => n7677, CK => CLK, RN => 
                           n6395, Q => n2855, QN => n5902);
   REGISTERS_reg_24_8_inst : DFFR_X1 port map( D => n7678, CK => CLK, RN => 
                           n6395, Q => n2854, QN => n5903);
   REGISTERS_reg_24_7_inst : DFFR_X1 port map( D => n7679, CK => CLK, RN => 
                           n6395, Q => n2853, QN => n5904);
   REGISTERS_reg_24_6_inst : DFFR_X1 port map( D => n7680, CK => CLK, RN => 
                           n6395, Q => n2852, QN => n5905);
   REGISTERS_reg_24_5_inst : DFFR_X1 port map( D => n7681, CK => CLK, RN => 
                           n6395, Q => n2851, QN => n5906);
   REGISTERS_reg_24_4_inst : DFFR_X1 port map( D => n7682, CK => CLK, RN => 
                           n6395, Q => n2850, QN => n5907);
   REGISTERS_reg_24_3_inst : DFFR_X1 port map( D => n3146, CK => CLK, RN => 
                           n6395, Q => n5483, QN => n987);
   REGISTERS_reg_24_2_inst : DFFR_X1 port map( D => n3145, CK => CLK, RN => 
                           n6395, Q => n5484, QN => n971);
   REGISTERS_reg_24_1_inst : DFFR_X1 port map( D => n3144, CK => CLK, RN => 
                           n6395, Q => n5485, QN => n955);
   REGISTERS_reg_24_0_inst : DFFR_X1 port map( D => n3143, CK => CLK, RN => 
                           n6395, Q => n5583, QN => n938);
   REGISTERS_reg_23_3_inst : DFFR_X1 port map( D => n3178, CK => CLK, RN => 
                           n6397, Q => n5580, QN => n988);
   REGISTERS_reg_23_2_inst : DFFR_X1 port map( D => n3177, CK => CLK, RN => 
                           n6397, Q => n5581, QN => n972);
   REGISTERS_reg_23_1_inst : DFFR_X1 port map( D => n3176, CK => CLK, RN => 
                           n6397, Q => n5582, QN => n956);
   REGISTERS_reg_23_0_inst : DFFR_X1 port map( D => n3175, CK => CLK, RN => 
                           n6397, Q => n5647, QN => n939);
   REGISTERS_reg_3_26_inst : DFFR_X1 port map( D => n7779, CK => CLK, RN => 
                           n6428, Q => n4056, QN => n5915);
   REGISTERS_reg_3_25_inst : DFFR_X1 port map( D => n7780, CK => CLK, RN => 
                           n6428, Q => n4055, QN => n5916);
   REGISTERS_reg_3_24_inst : DFFR_X1 port map( D => n7781, CK => CLK, RN => 
                           n6428, Q => n4054, QN => n5917);
   REGISTERS_reg_3_23_inst : DFFR_X1 port map( D => n7782, CK => CLK, RN => 
                           n6427, Q => n4053, QN => n5918);
   REGISTERS_reg_3_22_inst : DFFR_X1 port map( D => n7783, CK => CLK, RN => 
                           n6427, Q => n4052, QN => n5919);
   REGISTERS_reg_3_21_inst : DFFR_X1 port map( D => n7784, CK => CLK, RN => 
                           n6427, Q => n4051, QN => n5920);
   REGISTERS_reg_3_20_inst : DFFR_X1 port map( D => n7785, CK => CLK, RN => 
                           n6427, Q => n4050, QN => n5921);
   REGISTERS_reg_3_19_inst : DFFR_X1 port map( D => n7786, CK => CLK, RN => 
                           n6427, Q => n4049, QN => n5922);
   REGISTERS_reg_3_18_inst : DFFR_X1 port map( D => n7787, CK => CLK, RN => 
                           n6427, Q => n4048, QN => n5923);
   REGISTERS_reg_3_17_inst : DFFR_X1 port map( D => n7788, CK => CLK, RN => 
                           n6427, Q => n4047, QN => n5924);
   REGISTERS_reg_3_16_inst : DFFR_X1 port map( D => n7789, CK => CLK, RN => 
                           n6427, Q => n4046, QN => n5925);
   REGISTERS_reg_3_15_inst : DFFR_X1 port map( D => n7790, CK => CLK, RN => 
                           n6426, Q => n4045, QN => n5926);
   REGISTERS_reg_3_14_inst : DFFR_X1 port map( D => n7791, CK => CLK, RN => 
                           n6426, Q => n4044, QN => n5927);
   REGISTERS_reg_3_13_inst : DFFR_X1 port map( D => n7792, CK => CLK, RN => 
                           n6426, Q => n4043, QN => n5928);
   REGISTERS_reg_3_12_inst : DFFR_X1 port map( D => n7793, CK => CLK, RN => 
                           n6426, Q => n4042, QN => n5929);
   REGISTERS_reg_3_11_inst : DFFR_X1 port map( D => n7794, CK => CLK, RN => 
                           n6426, Q => n4041, QN => n5930);
   REGISTERS_reg_3_10_inst : DFFR_X1 port map( D => n7795, CK => CLK, RN => 
                           n6426, Q => n4040, QN => n5931);
   REGISTERS_reg_3_9_inst : DFFR_X1 port map( D => n7796, CK => CLK, RN => 
                           n6426, Q => n4039, QN => n5932);
   REGISTERS_reg_3_8_inst : DFFR_X1 port map( D => n7797, CK => CLK, RN => 
                           n6426, Q => n4038, QN => n5933);
   REGISTERS_reg_3_7_inst : DFFR_X1 port map( D => n7798, CK => CLK, RN => 
                           n6426, Q => n4037, QN => n5934);
   REGISTERS_reg_3_6_inst : DFFR_X1 port map( D => n7799, CK => CLK, RN => 
                           n6426, Q => n4036, QN => n5935);
   REGISTERS_reg_3_5_inst : DFFR_X1 port map( D => n7800, CK => CLK, RN => 
                           n6426, Q => n4035, QN => n5936);
   REGISTERS_reg_3_4_inst : DFFR_X1 port map( D => n7801, CK => CLK, RN => 
                           n6426, Q => n4034, QN => n5937);
   REGISTERS_reg_3_3_inst : DFFR_X1 port map( D => n7802, CK => CLK, RN => 
                           n6425, Q => n4033, QN => n5938);
   REGISTERS_reg_3_2_inst : DFFR_X1 port map( D => n7803, CK => CLK, RN => 
                           n6425, Q => n4032, QN => n5939);
   REGISTERS_reg_3_1_inst : DFFR_X1 port map( D => n7804, CK => CLK, RN => 
                           n6425, Q => n4031, QN => n5940);
   REGISTERS_reg_3_0_inst : DFFR_X1 port map( D => n7805, CK => CLK, RN => 
                           n6425, Q => n4030, QN => n5910);
   REGISTERS_reg_2_31_inst : DFFR_X1 port map( D => n7806, CK => CLK, RN => 
                           n6420, Q => n4093, QN => n5973);
   REGISTERS_reg_2_30_inst : DFFR_X1 port map( D => n7807, CK => CLK, RN => 
                           n6420, Q => n4092, QN => n5975);
   REGISTERS_reg_2_29_inst : DFFR_X1 port map( D => n7808, CK => CLK, RN => 
                           n6420, Q => n4091, QN => n5976);
   REGISTERS_reg_2_28_inst : DFFR_X1 port map( D => n7809, CK => CLK, RN => 
                           n6420, Q => n4090, QN => n5977);
   REGISTERS_reg_2_27_inst : DFFR_X1 port map( D => n7810, CK => CLK, RN => 
                           n6419, Q => n4089, QN => n5978);
   REGISTERS_reg_2_26_inst : DFFR_X1 port map( D => n7811, CK => CLK, RN => 
                           n6419, Q => n4088, QN => n5979);
   REGISTERS_reg_2_25_inst : DFFR_X1 port map( D => n7812, CK => CLK, RN => 
                           n6419, Q => n4087, QN => n5980);
   REGISTERS_reg_2_24_inst : DFFR_X1 port map( D => n7813, CK => CLK, RN => 
                           n6419, Q => n4086, QN => n5981);
   REGISTERS_reg_2_23_inst : DFFR_X1 port map( D => n7814, CK => CLK, RN => 
                           n6419, Q => n4085, QN => n5982);
   REGISTERS_reg_2_22_inst : DFFR_X1 port map( D => n7815, CK => CLK, RN => 
                           n6419, Q => n4084, QN => n5983);
   REGISTERS_reg_2_21_inst : DFFR_X1 port map( D => n7816, CK => CLK, RN => 
                           n6419, Q => n4083, QN => n5984);
   REGISTERS_reg_2_20_inst : DFFR_X1 port map( D => n7817, CK => CLK, RN => 
                           n6419, Q => n4082, QN => n5985);
   REGISTERS_reg_2_19_inst : DFFR_X1 port map( D => n7818, CK => CLK, RN => 
                           n6418, Q => n4081, QN => n5986);
   REGISTERS_reg_2_18_inst : DFFR_X1 port map( D => n7819, CK => CLK, RN => 
                           n6418, Q => n4080, QN => n5987);
   REGISTERS_reg_2_17_inst : DFFR_X1 port map( D => n7820, CK => CLK, RN => 
                           n6418, Q => n4079, QN => n5988);
   REGISTERS_reg_2_16_inst : DFFR_X1 port map( D => n7821, CK => CLK, RN => 
                           n6418, Q => n4078, QN => n5989);
   REGISTERS_reg_2_15_inst : DFFR_X1 port map( D => n7822, CK => CLK, RN => 
                           n6418, Q => n4077, QN => n5990);
   REGISTERS_reg_2_14_inst : DFFR_X1 port map( D => n7823, CK => CLK, RN => 
                           n6418, Q => n4076, QN => n5991);
   REGISTERS_reg_2_13_inst : DFFR_X1 port map( D => n7824, CK => CLK, RN => 
                           n6418, Q => n4075, QN => n5992);
   REGISTERS_reg_2_12_inst : DFFR_X1 port map( D => n7825, CK => CLK, RN => 
                           n6418, Q => n4074, QN => n5993);
   REGISTERS_reg_2_11_inst : DFFR_X1 port map( D => n7826, CK => CLK, RN => 
                           n6418, Q => n4073, QN => n5994);
   REGISTERS_reg_2_10_inst : DFFR_X1 port map( D => n7827, CK => CLK, RN => 
                           n6418, Q => n4072, QN => n5995);
   REGISTERS_reg_2_9_inst : DFFR_X1 port map( D => n7828, CK => CLK, RN => 
                           n6418, Q => n4071, QN => n5996);
   REGISTERS_reg_2_8_inst : DFFR_X1 port map( D => n7829, CK => CLK, RN => 
                           n6418, Q => n4070, QN => n5997);
   REGISTERS_reg_2_7_inst : DFFR_X1 port map( D => n7830, CK => CLK, RN => 
                           n6417, Q => n4069, QN => n5998);
   REGISTERS_reg_2_6_inst : DFFR_X1 port map( D => n7831, CK => CLK, RN => 
                           n6417, Q => n4068, QN => n5999);
   REGISTERS_reg_2_5_inst : DFFR_X1 port map( D => n7832, CK => CLK, RN => 
                           n6417, Q => n4067, QN => n6000);
   REGISTERS_reg_2_4_inst : DFFR_X1 port map( D => n7833, CK => CLK, RN => 
                           n6417, Q => n4066, QN => n6001);
   REGISTERS_reg_2_3_inst : DFFR_X1 port map( D => n7834, CK => CLK, RN => 
                           n6427, Q => n4065, QN => n6002);
   REGISTERS_reg_2_2_inst : DFFR_X1 port map( D => n7835, CK => CLK, RN => 
                           n6427, Q => n4064, QN => n6003);
   REGISTERS_reg_2_1_inst : DFFR_X1 port map( D => n7836, CK => CLK, RN => 
                           n6427, Q => n4063, QN => n6004);
   REGISTERS_reg_2_0_inst : DFFR_X1 port map( D => n7837, CK => CLK, RN => 
                           n6427, Q => n4062, QN => n5974);
   REGISTERS_reg_28_31_inst : DFFR_X1 port map( D => n3110, CK => CLK, RN => 
                           n6410, Q => n5681, QN => n2091);
   REGISTERS_reg_28_30_inst : DFFR_X1 port map( D => n3109, CK => CLK, RN => 
                           n6410, Q => n5682, QN => n2090);
   REGISTERS_reg_28_29_inst : DFFR_X1 port map( D => n3108, CK => CLK, RN => 
                           n6410, Q => n5683, QN => n2089);
   REGISTERS_reg_28_28_inst : DFFR_X1 port map( D => n3107, CK => CLK, RN => 
                           n6410, Q => n5684, QN => n2088);
   REGISTERS_reg_28_27_inst : DFFR_X1 port map( D => n3106, CK => CLK, RN => 
                           n6410, Q => n5685, QN => n2087);
   REGISTERS_reg_28_26_inst : DFFR_X1 port map( D => n3105, CK => CLK, RN => 
                           n6410, Q => n5686, QN => n2086);
   REGISTERS_reg_28_25_inst : DFFR_X1 port map( D => n3104, CK => CLK, RN => 
                           n6410, Q => n5687, QN => n2085);
   REGISTERS_reg_28_24_inst : DFFR_X1 port map( D => n3103, CK => CLK, RN => 
                           n6410, Q => n5688, QN => n2084);
   REGISTERS_reg_28_23_inst : DFFR_X1 port map( D => n3102, CK => CLK, RN => 
                           n6410, Q => n5689, QN => n2083);
   REGISTERS_reg_28_22_inst : DFFR_X1 port map( D => n3101, CK => CLK, RN => 
                           n6410, Q => n5690, QN => n2082);
   REGISTERS_reg_28_21_inst : DFFR_X1 port map( D => n3100, CK => CLK, RN => 
                           n6410, Q => n5691, QN => n2081);
   REGISTERS_reg_28_20_inst : DFFR_X1 port map( D => n3099, CK => CLK, RN => 
                           n6410, Q => n5692, QN => n2080);
   REGISTERS_reg_28_19_inst : DFFR_X1 port map( D => n3098, CK => CLK, RN => 
                           n6409, Q => n5693, QN => n2079);
   REGISTERS_reg_28_18_inst : DFFR_X1 port map( D => n3097, CK => CLK, RN => 
                           n6409, Q => n5694, QN => n2078);
   REGISTERS_reg_28_17_inst : DFFR_X1 port map( D => n3096, CK => CLK, RN => 
                           n6409, Q => n5695, QN => n2077);
   REGISTERS_reg_28_16_inst : DFFR_X1 port map( D => n3095, CK => CLK, RN => 
                           n6409, Q => n5696, QN => n2076);
   REGISTERS_reg_28_15_inst : DFFR_X1 port map( D => n3094, CK => CLK, RN => 
                           n6409, Q => n5697, QN => n2075);
   REGISTERS_reg_28_14_inst : DFFR_X1 port map( D => n3093, CK => CLK, RN => 
                           n6409, Q => n5698, QN => n2074);
   REGISTERS_reg_28_13_inst : DFFR_X1 port map( D => n3092, CK => CLK, RN => 
                           n6409, Q => n5699, QN => n2073);
   REGISTERS_reg_28_12_inst : DFFR_X1 port map( D => n3091, CK => CLK, RN => 
                           n6409, Q => n5700, QN => n2072);
   REGISTERS_reg_28_11_inst : DFFR_X1 port map( D => n3090, CK => CLK, RN => 
                           n6409, Q => n5701, QN => n2071);
   REGISTERS_reg_28_10_inst : DFFR_X1 port map( D => n3089, CK => CLK, RN => 
                           n6409, Q => n5702, QN => n2070);
   REGISTERS_reg_28_9_inst : DFFR_X1 port map( D => n3088, CK => CLK, RN => 
                           n6409, Q => n5703, QN => n2069);
   REGISTERS_reg_28_8_inst : DFFR_X1 port map( D => n3087, CK => CLK, RN => 
                           n6409, Q => n5704, QN => n2068);
   REGISTERS_reg_28_7_inst : DFFR_X1 port map( D => n3086, CK => CLK, RN => 
                           n6408, Q => n5705, QN => n2067);
   REGISTERS_reg_28_6_inst : DFFR_X1 port map( D => n3085, CK => CLK, RN => 
                           n6408, Q => n5706, QN => n2066);
   REGISTERS_reg_28_5_inst : DFFR_X1 port map( D => n3084, CK => CLK, RN => 
                           n6408, Q => n5707, QN => n2065);
   REGISTERS_reg_28_4_inst : DFFR_X1 port map( D => n3083, CK => CLK, RN => 
                           n6408, Q => n5708, QN => n2064);
   REGISTERS_reg_28_3_inst : DFFR_X1 port map( D => n3082, CK => CLK, RN => 
                           n6408, Q => n5709, QN => n2063);
   REGISTERS_reg_28_2_inst : DFFR_X1 port map( D => n3081, CK => CLK, RN => 
                           n6408, Q => n5710, QN => n2062);
   REGISTERS_reg_28_1_inst : DFFR_X1 port map( D => n3080, CK => CLK, RN => 
                           n6408, Q => n5711, QN => n2061);
   REGISTERS_reg_28_0_inst : DFFR_X1 port map( D => n3079, CK => CLK, RN => 
                           n6408, Q => n5358, QN => n2060);
   REGISTERS_reg_18_31_inst : DFFR_X1 port map( D => n3302, CK => CLK, RN => 
                           n6460, Q => n5744, QN => n2251);
   REGISTERS_reg_27_31_inst : DFFR_X1 port map( D => n4541, CK => CLK, RN => 
                           n6382, Q => n5391, QN => n2123);
   REGISTERS_reg_27_30_inst : DFFR_X1 port map( D => n4540, CK => CLK, RN => 
                           n6401, Q => n5392, QN => n2122);
   REGISTERS_reg_27_29_inst : DFFR_X1 port map( D => n4539, CK => CLK, RN => 
                           n6401, Q => n5393, QN => n2121);
   REGISTERS_reg_27_28_inst : DFFR_X1 port map( D => n4538, CK => CLK, RN => 
                           n6401, Q => n5394, QN => n2120);
   REGISTERS_reg_27_27_inst : DFFR_X1 port map( D => n4537, CK => CLK, RN => 
                           n6401, Q => n5395, QN => n2119);
   REGISTERS_reg_27_26_inst : DFFR_X1 port map( D => n4536, CK => CLK, RN => 
                           n6401, Q => n5396, QN => n2118);
   REGISTERS_reg_27_25_inst : DFFR_X1 port map( D => n4535, CK => CLK, RN => 
                           n6401, Q => n5397, QN => n2117);
   REGISTERS_reg_27_24_inst : DFFR_X1 port map( D => n4534, CK => CLK, RN => 
                           n6401, Q => n5398, QN => n2116);
   REGISTERS_reg_27_23_inst : DFFR_X1 port map( D => n4533, CK => CLK, RN => 
                           n6401, Q => n5399, QN => n2115);
   REGISTERS_reg_27_22_inst : DFFR_X1 port map( D => n4532, CK => CLK, RN => 
                           n6400, Q => n5400, QN => n2114);
   REGISTERS_reg_27_21_inst : DFFR_X1 port map( D => n4531, CK => CLK, RN => 
                           n6400, Q => n5401, QN => n2113);
   REGISTERS_reg_27_20_inst : DFFR_X1 port map( D => n4530, CK => CLK, RN => 
                           n6400, Q => n5402, QN => n2112);
   REGISTERS_reg_27_19_inst : DFFR_X1 port map( D => n4529, CK => CLK, RN => 
                           n6400, Q => n5403, QN => n2111);
   REGISTERS_reg_27_18_inst : DFFR_X1 port map( D => n4528, CK => CLK, RN => 
                           n6400, Q => n5404, QN => n2110);
   REGISTERS_reg_27_17_inst : DFFR_X1 port map( D => n4527, CK => CLK, RN => 
                           n6400, Q => n5405, QN => n2109);
   REGISTERS_reg_27_16_inst : DFFR_X1 port map( D => n4526, CK => CLK, RN => 
                           n6400, Q => n5406, QN => n2108);
   REGISTERS_reg_27_15_inst : DFFR_X1 port map( D => n4525, CK => CLK, RN => 
                           n6400, Q => n5407, QN => n2107);
   REGISTERS_reg_27_14_inst : DFFR_X1 port map( D => n4524, CK => CLK, RN => 
                           n6400, Q => n5408, QN => n2106);
   REGISTERS_reg_27_13_inst : DFFR_X1 port map( D => n4523, CK => CLK, RN => 
                           n6400, Q => n5409, QN => n2105);
   REGISTERS_reg_27_12_inst : DFFR_X1 port map( D => n4522, CK => CLK, RN => 
                           n6400, Q => n5410, QN => n2104);
   REGISTERS_reg_27_11_inst : DFFR_X1 port map( D => n4521, CK => CLK, RN => 
                           n6411, Q => n5411, QN => n2103);
   REGISTERS_reg_27_10_inst : DFFR_X1 port map( D => n4520, CK => CLK, RN => 
                           n6411, Q => n5412, QN => n2102);
   REGISTERS_reg_27_9_inst : DFFR_X1 port map( D => n4519, CK => CLK, RN => 
                           n6411, Q => n5413, QN => n2101);
   REGISTERS_reg_27_8_inst : DFFR_X1 port map( D => n4518, CK => CLK, RN => 
                           n6411, Q => n5414, QN => n2100);
   REGISTERS_reg_27_7_inst : DFFR_X1 port map( D => n4517, CK => CLK, RN => 
                           n6411, Q => n5415, QN => n2099);
   REGISTERS_reg_27_6_inst : DFFR_X1 port map( D => n4516, CK => CLK, RN => 
                           n6411, Q => n5416, QN => n2098);
   REGISTERS_reg_27_5_inst : DFFR_X1 port map( D => n4515, CK => CLK, RN => 
                           n6411, Q => n5417, QN => n2097);
   REGISTERS_reg_27_4_inst : DFFR_X1 port map( D => n4514, CK => CLK, RN => 
                           n6411, Q => n5418, QN => n2096);
   REGISTERS_reg_27_3_inst : DFFR_X1 port map( D => n4513, CK => CLK, RN => 
                           n6411, Q => n5419, QN => n2095);
   REGISTERS_reg_27_2_inst : DFFR_X1 port map( D => n4512, CK => CLK, RN => 
                           n6411, Q => n5420, QN => n2094);
   REGISTERS_reg_27_1_inst : DFFR_X1 port map( D => n4511, CK => CLK, RN => 
                           n6411, Q => n5421, QN => n2093);
   REGISTERS_reg_27_0_inst : DFFR_X1 port map( D => n4510, CK => CLK, RN => 
                           n6411, Q => n5546, QN => n2092);
   REGISTERS_reg_4_31_inst : DFFR_X1 port map( D => n4317, CK => CLK, RN => 
                           n6425, Q => n5875, QN => n2315);
   REGISTERS_reg_4_30_inst : DFFR_X1 port map( D => n4316, CK => CLK, RN => 
                           n6425, Q => n5298, QN => n2314);
   REGISTERS_reg_4_29_inst : DFFR_X1 port map( D => n4315, CK => CLK, RN => 
                           n6425, Q => n5299, QN => n2313);
   REGISTERS_reg_4_28_inst : DFFR_X1 port map( D => n4314, CK => CLK, RN => 
                           n6425, Q => n5300, QN => n2312);
   REGISTERS_reg_4_27_inst : DFFR_X1 port map( D => n4313, CK => CLK, RN => 
                           n6425, Q => n5301, QN => n2311);
   REGISTERS_reg_4_26_inst : DFFR_X1 port map( D => n4312, CK => CLK, RN => 
                           n6425, Q => n5302, QN => n2310);
   REGISTERS_reg_4_25_inst : DFFR_X1 port map( D => n4311, CK => CLK, RN => 
                           n6425, Q => n5303, QN => n2309);
   REGISTERS_reg_4_24_inst : DFFR_X1 port map( D => n4310, CK => CLK, RN => 
                           n6425, Q => n5304, QN => n2308);
   REGISTERS_reg_4_23_inst : DFFR_X1 port map( D => n4309, CK => CLK, RN => 
                           n6424, Q => n5305, QN => n2307);
   REGISTERS_reg_4_22_inst : DFFR_X1 port map( D => n4308, CK => CLK, RN => 
                           n6424, Q => n5306, QN => n2306);
   REGISTERS_reg_4_21_inst : DFFR_X1 port map( D => n4307, CK => CLK, RN => 
                           n6424, Q => n5307, QN => n2305);
   REGISTERS_reg_4_20_inst : DFFR_X1 port map( D => n4306, CK => CLK, RN => 
                           n6424, Q => n5308, QN => n2304);
   REGISTERS_reg_4_19_inst : DFFR_X1 port map( D => n4305, CK => CLK, RN => 
                           n6424, Q => n5309, QN => n2303);
   REGISTERS_reg_4_18_inst : DFFR_X1 port map( D => n4304, CK => CLK, RN => 
                           n6424, Q => n5310, QN => n2302);
   REGISTERS_reg_4_17_inst : DFFR_X1 port map( D => n4303, CK => CLK, RN => 
                           n6424, Q => n5311, QN => n2301);
   REGISTERS_reg_4_16_inst : DFFR_X1 port map( D => n4302, CK => CLK, RN => 
                           n6424, Q => n5312, QN => n2300);
   REGISTERS_reg_4_15_inst : DFFR_X1 port map( D => n4301, CK => CLK, RN => 
                           n6424, Q => n5313, QN => n2299);
   REGISTERS_reg_4_14_inst : DFFR_X1 port map( D => n4300, CK => CLK, RN => 
                           n6424, Q => n5314, QN => n2298);
   REGISTERS_reg_4_13_inst : DFFR_X1 port map( D => n4299, CK => CLK, RN => 
                           n6424, Q => n5315, QN => n2297);
   REGISTERS_reg_4_12_inst : DFFR_X1 port map( D => n4298, CK => CLK, RN => 
                           n6424, Q => n5316, QN => n2296);
   REGISTERS_reg_4_11_inst : DFFR_X1 port map( D => n4297, CK => CLK, RN => 
                           n6423, Q => n5317, QN => n2295);
   REGISTERS_reg_4_10_inst : DFFR_X1 port map( D => n4296, CK => CLK, RN => 
                           n6423, Q => n5318, QN => n2294);
   REGISTERS_reg_4_9_inst : DFFR_X1 port map( D => n4295, CK => CLK, RN => 
                           n6423, Q => n5319, QN => n2293);
   REGISTERS_reg_4_8_inst : DFFR_X1 port map( D => n4294, CK => CLK, RN => 
                           n6423, Q => n5320, QN => n2292);
   REGISTERS_reg_4_7_inst : DFFR_X1 port map( D => n4293, CK => CLK, RN => 
                           n6423, Q => n5321, QN => n2291);
   REGISTERS_reg_4_6_inst : DFFR_X1 port map( D => n4292, CK => CLK, RN => 
                           n6423, Q => n5322, QN => n2290);
   REGISTERS_reg_4_5_inst : DFFR_X1 port map( D => n4291, CK => CLK, RN => 
                           n6423, Q => n5323, QN => n2289);
   REGISTERS_reg_4_4_inst : DFFR_X1 port map( D => n4290, CK => CLK, RN => 
                           n6423, Q => n5324, QN => n2288);
   REGISTERS_reg_4_3_inst : DFFR_X1 port map( D => n4289, CK => CLK, RN => 
                           n6423, Q => n5325, QN => n2287);
   REGISTERS_reg_4_2_inst : DFFR_X1 port map( D => n4288, CK => CLK, RN => 
                           n6423, Q => n5326, QN => n2286);
   REGISTERS_reg_4_1_inst : DFFR_X1 port map( D => n4287, CK => CLK, RN => 
                           n6423, Q => n5327, QN => n2285);
   REGISTERS_reg_4_0_inst : DFFR_X1 port map( D => n4286, CK => CLK, RN => 
                           n6423, Q => n5876, QN => n2284);
   REGISTERS_reg_26_31_inst : DFFR_X1 port map( D => n4509, CK => CLK, RN => 
                           n6404, Q => n5649, QN => n2155);
   REGISTERS_reg_26_30_inst : DFFR_X1 port map( D => n4508, CK => CLK, RN => 
                           n6404, Q => n5650, QN => n2154);
   REGISTERS_reg_26_29_inst : DFFR_X1 port map( D => n4507, CK => CLK, RN => 
                           n6404, Q => n5651, QN => n2153);
   REGISTERS_reg_26_28_inst : DFFR_X1 port map( D => n4506, CK => CLK, RN => 
                           n6404, Q => n5652, QN => n2152);
   REGISTERS_reg_26_27_inst : DFFR_X1 port map( D => n4505, CK => CLK, RN => 
                           n6403, Q => n5653, QN => n2151);
   REGISTERS_reg_26_26_inst : DFFR_X1 port map( D => n4504, CK => CLK, RN => 
                           n6403, Q => n5654, QN => n2150);
   REGISTERS_reg_26_25_inst : DFFR_X1 port map( D => n4503, CK => CLK, RN => 
                           n6403, Q => n5655, QN => n2149);
   REGISTERS_reg_26_24_inst : DFFR_X1 port map( D => n4502, CK => CLK, RN => 
                           n6403, Q => n5656, QN => n2148);
   REGISTERS_reg_26_23_inst : DFFR_X1 port map( D => n4501, CK => CLK, RN => 
                           n6403, Q => n5657, QN => n2147);
   REGISTERS_reg_26_22_inst : DFFR_X1 port map( D => n4500, CK => CLK, RN => 
                           n6403, Q => n5658, QN => n2146);
   REGISTERS_reg_26_21_inst : DFFR_X1 port map( D => n4499, CK => CLK, RN => 
                           n6403, Q => n5659, QN => n2145);
   REGISTERS_reg_26_20_inst : DFFR_X1 port map( D => n4498, CK => CLK, RN => 
                           n6403, Q => n5660, QN => n2144);
   REGISTERS_reg_26_19_inst : DFFR_X1 port map( D => n4497, CK => CLK, RN => 
                           n6403, Q => n5661, QN => n2143);
   REGISTERS_reg_26_18_inst : DFFR_X1 port map( D => n4496, CK => CLK, RN => 
                           n6403, Q => n5662, QN => n2142);
   REGISTERS_reg_26_17_inst : DFFR_X1 port map( D => n4495, CK => CLK, RN => 
                           n6403, Q => n5663, QN => n2141);
   REGISTERS_reg_26_16_inst : DFFR_X1 port map( D => n4494, CK => CLK, RN => 
                           n6403, Q => n5664, QN => n2140);
   REGISTERS_reg_26_15_inst : DFFR_X1 port map( D => n4493, CK => CLK, RN => 
                           n6402, Q => n5665, QN => n2139);
   REGISTERS_reg_26_14_inst : DFFR_X1 port map( D => n4492, CK => CLK, RN => 
                           n6402, Q => n5666, QN => n2138);
   REGISTERS_reg_26_13_inst : DFFR_X1 port map( D => n4491, CK => CLK, RN => 
                           n6402, Q => n5667, QN => n2137);
   REGISTERS_reg_26_12_inst : DFFR_X1 port map( D => n4490, CK => CLK, RN => 
                           n6402, Q => n5668, QN => n2136);
   REGISTERS_reg_26_11_inst : DFFR_X1 port map( D => n4489, CK => CLK, RN => 
                           n6402, Q => n5669, QN => n2135);
   REGISTERS_reg_26_10_inst : DFFR_X1 port map( D => n4488, CK => CLK, RN => 
                           n6402, Q => n5670, QN => n2134);
   REGISTERS_reg_26_9_inst : DFFR_X1 port map( D => n4487, CK => CLK, RN => 
                           n6402, Q => n5671, QN => n2133);
   REGISTERS_reg_26_8_inst : DFFR_X1 port map( D => n4486, CK => CLK, RN => 
                           n6402, Q => n5672, QN => n2132);
   REGISTERS_reg_26_7_inst : DFFR_X1 port map( D => n4485, CK => CLK, RN => 
                           n6402, Q => n5673, QN => n2131);
   REGISTERS_reg_26_6_inst : DFFR_X1 port map( D => n4484, CK => CLK, RN => 
                           n6402, Q => n5674, QN => n2130);
   REGISTERS_reg_26_5_inst : DFFR_X1 port map( D => n4483, CK => CLK, RN => 
                           n6402, Q => n5675, QN => n2129);
   REGISTERS_reg_26_4_inst : DFFR_X1 port map( D => n4482, CK => CLK, RN => 
                           n6402, Q => n5676, QN => n2128);
   REGISTERS_reg_26_3_inst : DFFR_X1 port map( D => n4481, CK => CLK, RN => 
                           n6401, Q => n5677, QN => n2127);
   REGISTERS_reg_26_2_inst : DFFR_X1 port map( D => n4480, CK => CLK, RN => 
                           n6401, Q => n5678, QN => n2126);
   REGISTERS_reg_26_1_inst : DFFR_X1 port map( D => n4479, CK => CLK, RN => 
                           n6401, Q => n5679, QN => n2125);
   REGISTERS_reg_26_0_inst : DFFR_X1 port map( D => n4478, CK => CLK, RN => 
                           n6401, Q => n5648, QN => n2124);
   REGISTERS_reg_17_31_inst : DFFR_X1 port map( D => n4413, CK => CLK, RN => 
                           n6463, Q => n5168, QN => n2283);
   REGISTERS_reg_17_30_inst : DFFR_X1 port map( D => n4412, CK => CLK, RN => 
                           n6463, Q => n5361, QN => n2282);
   REGISTERS_reg_17_29_inst : DFFR_X1 port map( D => n4411, CK => CLK, RN => 
                           n6463, Q => n5362, QN => n2281);
   REGISTERS_reg_17_28_inst : DFFR_X1 port map( D => n4410, CK => CLK, RN => 
                           n6463, Q => n5363, QN => n2280);
   REGISTERS_reg_17_27_inst : DFFR_X1 port map( D => n4409, CK => CLK, RN => 
                           n6462, Q => n5364, QN => n2279);
   REGISTERS_reg_17_26_inst : DFFR_X1 port map( D => n4408, CK => CLK, RN => 
                           n6462, Q => n5365, QN => n2278);
   REGISTERS_reg_17_25_inst : DFFR_X1 port map( D => n4407, CK => CLK, RN => 
                           n6462, Q => n5366, QN => n2277);
   REGISTERS_reg_17_24_inst : DFFR_X1 port map( D => n4406, CK => CLK, RN => 
                           n6462, Q => n5367, QN => n2276);
   REGISTERS_reg_17_23_inst : DFFR_X1 port map( D => n4405, CK => CLK, RN => 
                           n6462, Q => n5368, QN => n2275);
   REGISTERS_reg_17_22_inst : DFFR_X1 port map( D => n4404, CK => CLK, RN => 
                           n6462, Q => n5369, QN => n2274);
   REGISTERS_reg_17_21_inst : DFFR_X1 port map( D => n4403, CK => CLK, RN => 
                           n6462, Q => n5370, QN => n2273);
   REGISTERS_reg_17_20_inst : DFFR_X1 port map( D => n4402, CK => CLK, RN => 
                           n6462, Q => n5371, QN => n2272);
   REGISTERS_reg_17_19_inst : DFFR_X1 port map( D => n4401, CK => CLK, RN => 
                           n6461, Q => n5372, QN => n2271);
   REGISTERS_reg_17_18_inst : DFFR_X1 port map( D => n4400, CK => CLK, RN => 
                           n6461, Q => n5373, QN => n2270);
   REGISTERS_reg_17_17_inst : DFFR_X1 port map( D => n4399, CK => CLK, RN => 
                           n6461, Q => n5374, QN => n2269);
   REGISTERS_reg_17_16_inst : DFFR_X1 port map( D => n4398, CK => CLK, RN => 
                           n6461, Q => n5375, QN => n2268);
   REGISTERS_reg_17_15_inst : DFFR_X1 port map( D => n4397, CK => CLK, RN => 
                           n6461, Q => n5376, QN => n2267);
   REGISTERS_reg_17_14_inst : DFFR_X1 port map( D => n4396, CK => CLK, RN => 
                           n6461, Q => n5377, QN => n2266);
   REGISTERS_reg_17_13_inst : DFFR_X1 port map( D => n4395, CK => CLK, RN => 
                           n6461, Q => n5378, QN => n2265);
   REGISTERS_reg_17_12_inst : DFFR_X1 port map( D => n4394, CK => CLK, RN => 
                           n6461, Q => n5379, QN => n2264);
   REGISTERS_reg_17_11_inst : DFFR_X1 port map( D => n4393, CK => CLK, RN => 
                           n6461, Q => n5380, QN => n2263);
   REGISTERS_reg_17_10_inst : DFFR_X1 port map( D => n4392, CK => CLK, RN => 
                           n6461, Q => n5381, QN => n2262);
   REGISTERS_reg_17_9_inst : DFFR_X1 port map( D => n4391, CK => CLK, RN => 
                           n6461, Q => n5382, QN => n2261);
   REGISTERS_reg_17_8_inst : DFFR_X1 port map( D => n4390, CK => CLK, RN => 
                           n6461, Q => n5383, QN => n2260);
   REGISTERS_reg_17_7_inst : DFFR_X1 port map( D => n4389, CK => CLK, RN => 
                           n6460, Q => n5384, QN => n2259);
   REGISTERS_reg_17_6_inst : DFFR_X1 port map( D => n4388, CK => CLK, RN => 
                           n6460, Q => n5385, QN => n2258);
   REGISTERS_reg_17_5_inst : DFFR_X1 port map( D => n4387, CK => CLK, RN => 
                           n6460, Q => n5386, QN => n2257);
   REGISTERS_reg_17_4_inst : DFFR_X1 port map( D => n4386, CK => CLK, RN => 
                           n6460, Q => n5387, QN => n2256);
   REGISTERS_reg_17_3_inst : DFFR_X1 port map( D => n4385, CK => CLK, RN => 
                           n6459, Q => n5388, QN => n2255);
   REGISTERS_reg_17_2_inst : DFFR_X1 port map( D => n4384, CK => CLK, RN => 
                           n6459, Q => n5389, QN => n2254);
   REGISTERS_reg_17_1_inst : DFFR_X1 port map( D => n4383, CK => CLK, RN => 
                           n6459, Q => n5390, QN => n2253);
   REGISTERS_reg_17_0_inst : DFFR_X1 port map( D => n4382, CK => CLK, RN => 
                           n6459, Q => n5233, QN => n2252);
   REGISTERS_reg_5_31_inst : DFFR_X1 port map( D => n4349, CK => CLK, RN => 
                           n6422, Q => n5809, QN => n4029);
   REGISTERS_reg_5_30_inst : DFFR_X1 port map( D => n4348, CK => CLK, RN => 
                           n6422, Q => n5810, QN => n4028);
   REGISTERS_reg_5_29_inst : DFFR_X1 port map( D => n4347, CK => CLK, RN => 
                           n6422, Q => n5811, QN => n4027);
   REGISTERS_reg_5_28_inst : DFFR_X1 port map( D => n4346, CK => CLK, RN => 
                           n6422, Q => n5812, QN => n4026);
   REGISTERS_reg_5_27_inst : DFFR_X1 port map( D => n4345, CK => CLK, RN => 
                           n6434, Q => n5813, QN => n4025);
   REGISTERS_reg_5_26_inst : DFFR_X1 port map( D => n4344, CK => CLK, RN => 
                           n6434, Q => n5814, QN => n4024);
   REGISTERS_reg_5_25_inst : DFFR_X1 port map( D => n4343, CK => CLK, RN => 
                           n6434, Q => n5815, QN => n4023);
   REGISTERS_reg_5_24_inst : DFFR_X1 port map( D => n4342, CK => CLK, RN => 
                           n6434, Q => n5816, QN => n4022);
   REGISTERS_reg_5_23_inst : DFFR_X1 port map( D => n4341, CK => CLK, RN => 
                           n6434, Q => n5817, QN => n4021);
   REGISTERS_reg_5_22_inst : DFFR_X1 port map( D => n4340, CK => CLK, RN => 
                           n6434, Q => n5818, QN => n4020);
   REGISTERS_reg_5_21_inst : DFFR_X1 port map( D => n4339, CK => CLK, RN => 
                           n6434, Q => n5819, QN => n4019);
   REGISTERS_reg_5_20_inst : DFFR_X1 port map( D => n4338, CK => CLK, RN => 
                           n6434, Q => n5820, QN => n4018);
   REGISTERS_reg_5_19_inst : DFFR_X1 port map( D => n4337, CK => CLK, RN => 
                           n6433, Q => n5821, QN => n4017);
   REGISTERS_reg_5_18_inst : DFFR_X1 port map( D => n4336, CK => CLK, RN => 
                           n6433, Q => n5822, QN => n4016);
   REGISTERS_reg_5_17_inst : DFFR_X1 port map( D => n4335, CK => CLK, RN => 
                           n6433, Q => n5823, QN => n4015);
   REGISTERS_reg_5_16_inst : DFFR_X1 port map( D => n4334, CK => CLK, RN => 
                           n6433, Q => n5824, QN => n4014);
   REGISTERS_reg_5_15_inst : DFFR_X1 port map( D => n4333, CK => CLK, RN => 
                           n6433, Q => n5825, QN => n4013);
   REGISTERS_reg_5_14_inst : DFFR_X1 port map( D => n4332, CK => CLK, RN => 
                           n6433, Q => n5826, QN => n4012);
   REGISTERS_reg_5_13_inst : DFFR_X1 port map( D => n4331, CK => CLK, RN => 
                           n6433, Q => n5827, QN => n4011);
   REGISTERS_reg_5_12_inst : DFFR_X1 port map( D => n4330, CK => CLK, RN => 
                           n6433, Q => n5828, QN => n4010);
   REGISTERS_reg_5_11_inst : DFFR_X1 port map( D => n4329, CK => CLK, RN => 
                           n6433, Q => n5829, QN => n4009);
   REGISTERS_reg_5_10_inst : DFFR_X1 port map( D => n4328, CK => CLK, RN => 
                           n6433, Q => n5830, QN => n4008);
   REGISTERS_reg_5_9_inst : DFFR_X1 port map( D => n4327, CK => CLK, RN => 
                           n6433, Q => n5831, QN => n4007);
   REGISTERS_reg_5_8_inst : DFFR_X1 port map( D => n4326, CK => CLK, RN => 
                           n6433, Q => n5832, QN => n4006);
   REGISTERS_reg_5_7_inst : DFFR_X1 port map( D => n4325, CK => CLK, RN => 
                           n6432, Q => n5833, QN => n4005);
   REGISTERS_reg_5_6_inst : DFFR_X1 port map( D => n4324, CK => CLK, RN => 
                           n6432, Q => n5834, QN => n4004);
   REGISTERS_reg_5_5_inst : DFFR_X1 port map( D => n4323, CK => CLK, RN => 
                           n6432, Q => n5835, QN => n4003);
   REGISTERS_reg_5_4_inst : DFFR_X1 port map( D => n4322, CK => CLK, RN => 
                           n6432, Q => n5836, QN => n4002);
   REGISTERS_reg_5_3_inst : DFFR_X1 port map( D => n4321, CK => CLK, RN => 
                           n6431, Q => n5837, QN => n4001);
   REGISTERS_reg_5_2_inst : DFFR_X1 port map( D => n4320, CK => CLK, RN => 
                           n6431, Q => n5838, QN => n4000);
   REGISTERS_reg_5_1_inst : DFFR_X1 port map( D => n4319, CK => CLK, RN => 
                           n6431, Q => n5839, QN => n3999);
   REGISTERS_reg_5_0_inst : DFFR_X1 port map( D => n4318, CK => CLK, RN => 
                           n6431, Q => n5840, QN => n3998);
   REGISTERS_reg_31_31_inst : DFFR_X1 port map( D => n4605, CK => CLK, RN => 
                           n6413, Q => n5487, QN => n2717);
   REGISTERS_reg_31_30_inst : DFFR_X1 port map( D => n4604, CK => CLK, RN => 
                           n6413, Q => n5488, QN => n2716);
   REGISTERS_reg_31_29_inst : DFFR_X1 port map( D => n4603, CK => CLK, RN => 
                           n6413, Q => n5489, QN => n2715);
   REGISTERS_reg_31_28_inst : DFFR_X1 port map( D => n4602, CK => CLK, RN => 
                           n6413, Q => n5490, QN => n2714);
   REGISTERS_reg_31_27_inst : DFFR_X1 port map( D => n4601, CK => CLK, RN => 
                           n6413, Q => n5491, QN => n2713);
   REGISTERS_reg_31_26_inst : DFFR_X1 port map( D => n4600, CK => CLK, RN => 
                           n6413, Q => n5492, QN => n2712);
   REGISTERS_reg_31_25_inst : DFFR_X1 port map( D => n4599, CK => CLK, RN => 
                           n6413, Q => n5493, QN => n2711);
   REGISTERS_reg_31_24_inst : DFFR_X1 port map( D => n4598, CK => CLK, RN => 
                           n6413, Q => n5494, QN => n2710);
   REGISTERS_reg_31_23_inst : DFFR_X1 port map( D => n4597, CK => CLK, RN => 
                           n6413, Q => n5495, QN => n2709);
   REGISTERS_reg_31_22_inst : DFFR_X1 port map( D => n4596, CK => CLK, RN => 
                           n6413, Q => n5496, QN => n2708);
   REGISTERS_reg_31_21_inst : DFFR_X1 port map( D => n4595, CK => CLK, RN => 
                           n6413, Q => n5497, QN => n2707);
   REGISTERS_reg_31_20_inst : DFFR_X1 port map( D => n4594, CK => CLK, RN => 
                           n6413, Q => n5498, QN => n2706);
   REGISTERS_reg_31_19_inst : DFFR_X1 port map( D => n4593, CK => CLK, RN => 
                           n6412, Q => n5499, QN => n2705);
   REGISTERS_reg_31_18_inst : DFFR_X1 port map( D => n4592, CK => CLK, RN => 
                           n6412, Q => n5500, QN => n2704);
   REGISTERS_reg_31_17_inst : DFFR_X1 port map( D => n4591, CK => CLK, RN => 
                           n6412, Q => n5501, QN => n2703);
   REGISTERS_reg_31_16_inst : DFFR_X1 port map( D => n4590, CK => CLK, RN => 
                           n6412, Q => n5502, QN => n2702);
   REGISTERS_reg_31_15_inst : DFFR_X1 port map( D => n4589, CK => CLK, RN => 
                           n6412, Q => n5503, QN => n2701);
   REGISTERS_reg_31_14_inst : DFFR_X1 port map( D => n4588, CK => CLK, RN => 
                           n6412, Q => n5504, QN => n2700);
   REGISTERS_reg_31_13_inst : DFFR_X1 port map( D => n4587, CK => CLK, RN => 
                           n6412, Q => n5505, QN => n2699);
   REGISTERS_reg_31_12_inst : DFFR_X1 port map( D => n4586, CK => CLK, RN => 
                           n6412, Q => n5506, QN => n2698);
   REGISTERS_reg_31_11_inst : DFFR_X1 port map( D => n4585, CK => CLK, RN => 
                           n6412, Q => n5507, QN => n2697);
   REGISTERS_reg_31_10_inst : DFFR_X1 port map( D => n4584, CK => CLK, RN => 
                           n6412, Q => n5508, QN => n2696);
   REGISTERS_reg_31_9_inst : DFFR_X1 port map( D => n4583, CK => CLK, RN => 
                           n6412, Q => n5509, QN => n2695);
   REGISTERS_reg_31_8_inst : DFFR_X1 port map( D => n4582, CK => CLK, RN => 
                           n6412, Q => n5510, QN => n2694);
   REGISTERS_reg_31_7_inst : DFFR_X1 port map( D => n4581, CK => CLK, RN => 
                           n6417, Q => n5511, QN => n2693);
   REGISTERS_reg_31_6_inst : DFFR_X1 port map( D => n4580, CK => CLK, RN => 
                           n6417, Q => n5512, QN => n2692);
   REGISTERS_reg_31_5_inst : DFFR_X1 port map( D => n4579, CK => CLK, RN => 
                           n6417, Q => n5513, QN => n2691);
   REGISTERS_reg_31_4_inst : DFFR_X1 port map( D => n4578, CK => CLK, RN => 
                           n6417, Q => n5514, QN => n2690);
   REGISTERS_reg_31_3_inst : DFFR_X1 port map( D => n4577, CK => CLK, RN => 
                           n6417, Q => n998, QN => n5877);
   REGISTERS_reg_31_2_inst : DFFR_X1 port map( D => n4576, CK => CLK, RN => 
                           n6417, Q => n982, QN => n5878);
   REGISTERS_reg_31_1_inst : DFFR_X1 port map( D => n4575, CK => CLK, RN => 
                           n6417, Q => n966, QN => n5879);
   REGISTERS_reg_31_0_inst : DFFR_X1 port map( D => n4574, CK => CLK, RN => 
                           n6417, Q => n950, QN => n5908);
   REGISTERS_reg_21_31_inst : DFFR_X1 port map( D => n4477, CK => CLK, RN => 
                           n6394, Q => n5172, QN => n2973);
   REGISTERS_reg_21_30_inst : DFFR_X1 port map( D => n4476, CK => CLK, RN => 
                           n6394, Q => n5173, QN => n2972);
   REGISTERS_reg_21_29_inst : DFFR_X1 port map( D => n4475, CK => CLK, RN => 
                           n6393, Q => n5174, QN => n2971);
   REGISTERS_reg_21_28_inst : DFFR_X1 port map( D => n4474, CK => CLK, RN => 
                           n6393, Q => n5175, QN => n2970);
   REGISTERS_reg_21_27_inst : DFFR_X1 port map( D => n4473, CK => CLK, RN => 
                           n6393, Q => n5176, QN => n2969);
   REGISTERS_reg_21_26_inst : DFFR_X1 port map( D => n4472, CK => CLK, RN => 
                           n6393, Q => n5177, QN => n2968);
   REGISTERS_reg_21_25_inst : DFFR_X1 port map( D => n4471, CK => CLK, RN => 
                           n6393, Q => n5178, QN => n2967);
   REGISTERS_reg_21_24_inst : DFFR_X1 port map( D => n4470, CK => CLK, RN => 
                           n6393, Q => n5179, QN => n2966);
   REGISTERS_reg_21_23_inst : DFFR_X1 port map( D => n4469, CK => CLK, RN => 
                           n6393, Q => n5180, QN => n2965);
   REGISTERS_reg_21_22_inst : DFFR_X1 port map( D => n4468, CK => CLK, RN => 
                           n6393, Q => n5181, QN => n2964);
   REGISTERS_reg_21_21_inst : DFFR_X1 port map( D => n4467, CK => CLK, RN => 
                           n6392, Q => n5182, QN => n2963);
   REGISTERS_reg_21_20_inst : DFFR_X1 port map( D => n4466, CK => CLK, RN => 
                           n6392, Q => n5183, QN => n2962);
   REGISTERS_reg_21_19_inst : DFFR_X1 port map( D => n4465, CK => CLK, RN => 
                           n6392, Q => n5184, QN => n2961);
   REGISTERS_reg_21_18_inst : DFFR_X1 port map( D => n4464, CK => CLK, RN => 
                           n6392, Q => n5185, QN => n2960);
   REGISTERS_reg_21_17_inst : DFFR_X1 port map( D => n4463, CK => CLK, RN => 
                           n6392, Q => n5186, QN => n2959);
   REGISTERS_reg_21_16_inst : DFFR_X1 port map( D => n4462, CK => CLK, RN => 
                           n6392, Q => n5187, QN => n2958);
   REGISTERS_reg_21_15_inst : DFFR_X1 port map( D => n4461, CK => CLK, RN => 
                           n6392, Q => n5188, QN => n2957);
   REGISTERS_reg_21_14_inst : DFFR_X1 port map( D => n4460, CK => CLK, RN => 
                           n6392, Q => n5189, QN => n2956);
   REGISTERS_reg_21_13_inst : DFFR_X1 port map( D => n4459, CK => CLK, RN => 
                           n6392, Q => n5190, QN => n2955);
   REGISTERS_reg_21_12_inst : DFFR_X1 port map( D => n4458, CK => CLK, RN => 
                           n6392, Q => n5191, QN => n2954);
   REGISTERS_reg_21_11_inst : DFFR_X1 port map( D => n4457, CK => CLK, RN => 
                           n6392, Q => n5192, QN => n2953);
   REGISTERS_reg_21_10_inst : DFFR_X1 port map( D => n4456, CK => CLK, RN => 
                           n6392, Q => n5193, QN => n2952);
   REGISTERS_reg_21_9_inst : DFFR_X1 port map( D => n4455, CK => CLK, RN => 
                           n6391, Q => n5194, QN => n2951);
   REGISTERS_reg_21_8_inst : DFFR_X1 port map( D => n4454, CK => CLK, RN => 
                           n6391, Q => n5195, QN => n2950);
   REGISTERS_reg_21_7_inst : DFFR_X1 port map( D => n4453, CK => CLK, RN => 
                           n6391, Q => n5196, QN => n2949);
   REGISTERS_reg_21_6_inst : DFFR_X1 port map( D => n4452, CK => CLK, RN => 
                           n6391, Q => n5197, QN => n2948);
   REGISTERS_reg_21_5_inst : DFFR_X1 port map( D => n4451, CK => CLK, RN => 
                           n6391, Q => n5198, QN => n2947);
   REGISTERS_reg_21_4_inst : DFFR_X1 port map( D => n4450, CK => CLK, RN => 
                           n6391, Q => n5199, QN => n2946);
   REGISTERS_reg_21_3_inst : DFFR_X1 port map( D => n4449, CK => CLK, RN => 
                           n6391, Q => n5200, QN => n2945);
   REGISTERS_reg_21_2_inst : DFFR_X1 port map( D => n4448, CK => CLK, RN => 
                           n6391, Q => n5201, QN => n2944);
   REGISTERS_reg_21_1_inst : DFFR_X1 port map( D => n4447, CK => CLK, RN => 
                           n6391, Q => n5202, QN => n2943);
   REGISTERS_reg_21_0_inst : DFFR_X1 port map( D => n4446, CK => CLK, RN => 
                           n6391, Q => n5359, QN => n2942);
   REGISTERS_reg_12_31_inst : DFFR_X1 port map( D => n4221, CK => CLK, RN => 
                           n6452, Q => n5615, QN => n3805);
   REGISTERS_reg_12_30_inst : DFFR_X1 port map( D => n4220, CK => CLK, RN => 
                           n6452, Q => n5616, QN => n3804);
   REGISTERS_reg_12_29_inst : DFFR_X1 port map( D => n4219, CK => CLK, RN => 
                           n6452, Q => n5617, QN => n3803);
   REGISTERS_reg_12_28_inst : DFFR_X1 port map( D => n4218, CK => CLK, RN => 
                           n6452, Q => n5618, QN => n3802);
   REGISTERS_reg_12_27_inst : DFFR_X1 port map( D => n4217, CK => CLK, RN => 
                           n6451, Q => n5619, QN => n3801);
   REGISTERS_reg_12_26_inst : DFFR_X1 port map( D => n4216, CK => CLK, RN => 
                           n6451, Q => n5620, QN => n3800);
   REGISTERS_reg_12_25_inst : DFFR_X1 port map( D => n4215, CK => CLK, RN => 
                           n6451, Q => n5621, QN => n3799);
   REGISTERS_reg_12_24_inst : DFFR_X1 port map( D => n4214, CK => CLK, RN => 
                           n6451, Q => n5622, QN => n3798);
   REGISTERS_reg_12_23_inst : DFFR_X1 port map( D => n4213, CK => CLK, RN => 
                           n6451, Q => n5623, QN => n3797);
   REGISTERS_reg_12_22_inst : DFFR_X1 port map( D => n4212, CK => CLK, RN => 
                           n6451, Q => n5624, QN => n3796);
   REGISTERS_reg_12_21_inst : DFFR_X1 port map( D => n4211, CK => CLK, RN => 
                           n6451, Q => n5625, QN => n3795);
   REGISTERS_reg_12_20_inst : DFFR_X1 port map( D => n4210, CK => CLK, RN => 
                           n6451, Q => n5626, QN => n3794);
   REGISTERS_reg_12_19_inst : DFFR_X1 port map( D => n4209, CK => CLK, RN => 
                           n6451, Q => n5627, QN => n3793);
   REGISTERS_reg_12_18_inst : DFFR_X1 port map( D => n4208, CK => CLK, RN => 
                           n6451, Q => n5628, QN => n3792);
   REGISTERS_reg_12_17_inst : DFFR_X1 port map( D => n4207, CK => CLK, RN => 
                           n6451, Q => n5629, QN => n3791);
   REGISTERS_reg_12_16_inst : DFFR_X1 port map( D => n4206, CK => CLK, RN => 
                           n6451, Q => n5630, QN => n3790);
   REGISTERS_reg_12_15_inst : DFFR_X1 port map( D => n4205, CK => CLK, RN => 
                           n6450, Q => n5631, QN => n3789);
   REGISTERS_reg_12_14_inst : DFFR_X1 port map( D => n4204, CK => CLK, RN => 
                           n6450, Q => n5632, QN => n3788);
   REGISTERS_reg_12_13_inst : DFFR_X1 port map( D => n4203, CK => CLK, RN => 
                           n6450, Q => n5633, QN => n3787);
   REGISTERS_reg_12_12_inst : DFFR_X1 port map( D => n4202, CK => CLK, RN => 
                           n6450, Q => n5634, QN => n3786);
   REGISTERS_reg_12_11_inst : DFFR_X1 port map( D => n4201, CK => CLK, RN => 
                           n6450, Q => n5635, QN => n3785);
   REGISTERS_reg_12_10_inst : DFFR_X1 port map( D => n4200, CK => CLK, RN => 
                           n6450, Q => n5636, QN => n3784);
   REGISTERS_reg_12_9_inst : DFFR_X1 port map( D => n4199, CK => CLK, RN => 
                           n6450, Q => n5637, QN => n3783);
   REGISTERS_reg_12_8_inst : DFFR_X1 port map( D => n4198, CK => CLK, RN => 
                           n6450, Q => n5638, QN => n3782);
   REGISTERS_reg_12_7_inst : DFFR_X1 port map( D => n4197, CK => CLK, RN => 
                           n6450, Q => n5639, QN => n3781);
   REGISTERS_reg_12_6_inst : DFFR_X1 port map( D => n4196, CK => CLK, RN => 
                           n6450, Q => n5640, QN => n3780);
   REGISTERS_reg_12_5_inst : DFFR_X1 port map( D => n4195, CK => CLK, RN => 
                           n6450, Q => n5641, QN => n3779);
   REGISTERS_reg_12_4_inst : DFFR_X1 port map( D => n4194, CK => CLK, RN => 
                           n6450, Q => n5642, QN => n3778);
   REGISTERS_reg_12_3_inst : DFFR_X1 port map( D => n4193, CK => CLK, RN => 
                           n6449, Q => n5643, QN => n3777);
   REGISTERS_reg_12_2_inst : DFFR_X1 port map( D => n4192, CK => CLK, RN => 
                           n6449, Q => n5644, QN => n3776);
   REGISTERS_reg_12_1_inst : DFFR_X1 port map( D => n4191, CK => CLK, RN => 
                           n6449, Q => n5645, QN => n3775);
   REGISTERS_reg_12_0_inst : DFFR_X1 port map( D => n4190, CK => CLK, RN => 
                           n6449, Q => n5646, QN => n3774);
   REGISTERS_reg_8_31_inst : DFFR_X1 port map( D => n4157, CK => CLK, RN => 
                           n6438, Q => n5777, QN => n3933);
   REGISTERS_reg_8_30_inst : DFFR_X1 port map( D => n4156, CK => CLK, RN => 
                           n6438, Q => n5778, QN => n3932);
   REGISTERS_reg_8_29_inst : DFFR_X1 port map( D => n4155, CK => CLK, RN => 
                           n6438, Q => n5779, QN => n3931);
   REGISTERS_reg_8_28_inst : DFFR_X1 port map( D => n4154, CK => CLK, RN => 
                           n6438, Q => n5780, QN => n3930);
   REGISTERS_reg_8_27_inst : DFFR_X1 port map( D => n4153, CK => CLK, RN => 
                           n6438, Q => n5781, QN => n3929);
   REGISTERS_reg_8_26_inst : DFFR_X1 port map( D => n4152, CK => CLK, RN => 
                           n6438, Q => n5782, QN => n3928);
   REGISTERS_reg_8_25_inst : DFFR_X1 port map( D => n4151, CK => CLK, RN => 
                           n6438, Q => n5783, QN => n3927);
   REGISTERS_reg_8_24_inst : DFFR_X1 port map( D => n4150, CK => CLK, RN => 
                           n6438, Q => n5784, QN => n3926);
   REGISTERS_reg_8_23_inst : DFFR_X1 port map( D => n4149, CK => CLK, RN => 
                           n6438, Q => n5785, QN => n3925);
   REGISTERS_reg_8_22_inst : DFFR_X1 port map( D => n4148, CK => CLK, RN => 
                           n6438, Q => n5786, QN => n3924);
   REGISTERS_reg_8_21_inst : DFFR_X1 port map( D => n4147, CK => CLK, RN => 
                           n6438, Q => n5787, QN => n3923);
   REGISTERS_reg_8_20_inst : DFFR_X1 port map( D => n4146, CK => CLK, RN => 
                           n6438, Q => n5788, QN => n3922);
   REGISTERS_reg_8_19_inst : DFFR_X1 port map( D => n4145, CK => CLK, RN => 
                           n6437, Q => n5789, QN => n3921);
   REGISTERS_reg_8_18_inst : DFFR_X1 port map( D => n4144, CK => CLK, RN => 
                           n6437, Q => n5790, QN => n3920);
   REGISTERS_reg_8_17_inst : DFFR_X1 port map( D => n4143, CK => CLK, RN => 
                           n6437, Q => n5791, QN => n3919);
   REGISTERS_reg_8_16_inst : DFFR_X1 port map( D => n4142, CK => CLK, RN => 
                           n6437, Q => n5792, QN => n3918);
   REGISTERS_reg_8_15_inst : DFFR_X1 port map( D => n4141, CK => CLK, RN => 
                           n6437, Q => n5793, QN => n3917);
   REGISTERS_reg_8_14_inst : DFFR_X1 port map( D => n4140, CK => CLK, RN => 
                           n6437, Q => n5794, QN => n3916);
   REGISTERS_reg_8_13_inst : DFFR_X1 port map( D => n4139, CK => CLK, RN => 
                           n6437, Q => n5795, QN => n3915);
   REGISTERS_reg_8_12_inst : DFFR_X1 port map( D => n4138, CK => CLK, RN => 
                           n6437, Q => n5796, QN => n3914);
   REGISTERS_reg_8_11_inst : DFFR_X1 port map( D => n4137, CK => CLK, RN => 
                           n6437, Q => n5797, QN => n3913);
   REGISTERS_reg_8_10_inst : DFFR_X1 port map( D => n4136, CK => CLK, RN => 
                           n6437, Q => n5798, QN => n3912);
   REGISTERS_reg_8_9_inst : DFFR_X1 port map( D => n4135, CK => CLK, RN => 
                           n6437, Q => n5799, QN => n3911);
   REGISTERS_reg_8_8_inst : DFFR_X1 port map( D => n4134, CK => CLK, RN => 
                           n6437, Q => n5800, QN => n3910);
   REGISTERS_reg_8_7_inst : DFFR_X1 port map( D => n4133, CK => CLK, RN => 
                           n6436, Q => n5801, QN => n3909);
   REGISTERS_reg_8_6_inst : DFFR_X1 port map( D => n4132, CK => CLK, RN => 
                           n6436, Q => n5802, QN => n3908);
   REGISTERS_reg_8_5_inst : DFFR_X1 port map( D => n4131, CK => CLK, RN => 
                           n6436, Q => n5803, QN => n3907);
   REGISTERS_reg_8_4_inst : DFFR_X1 port map( D => n4130, CK => CLK, RN => 
                           n6436, Q => n5804, QN => n3906);
   REGISTERS_reg_8_3_inst : DFFR_X1 port map( D => n4129, CK => CLK, RN => 
                           n6436, Q => n5805, QN => n3905);
   REGISTERS_reg_8_2_inst : DFFR_X1 port map( D => n4128, CK => CLK, RN => 
                           n6436, Q => n5806, QN => n3904);
   REGISTERS_reg_8_1_inst : DFFR_X1 port map( D => n4127, CK => CLK, RN => 
                           n6436, Q => n5807, QN => n3903);
   REGISTERS_reg_8_0_inst : DFFR_X1 port map( D => n4126, CK => CLK, RN => 
                           n6436, Q => n5808, QN => n3902);
   REGISTERS_reg_30_31_inst : DFFR_X1 port map( D => n4573, CK => CLK, RN => 
                           n6416, Q => n5584, QN => n2749);
   REGISTERS_reg_30_30_inst : DFFR_X1 port map( D => n4572, CK => CLK, RN => 
                           n6416, Q => n5585, QN => n2748);
   REGISTERS_reg_30_29_inst : DFFR_X1 port map( D => n4571, CK => CLK, RN => 
                           n6416, Q => n5586, QN => n2747);
   REGISTERS_reg_30_28_inst : DFFR_X1 port map( D => n4570, CK => CLK, RN => 
                           n6416, Q => n5587, QN => n2746);
   REGISTERS_reg_30_27_inst : DFFR_X1 port map( D => n4569, CK => CLK, RN => 
                           n6416, Q => n5588, QN => n2745);
   REGISTERS_reg_30_26_inst : DFFR_X1 port map( D => n4568, CK => CLK, RN => 
                           n6416, Q => n5589, QN => n2744);
   REGISTERS_reg_30_25_inst : DFFR_X1 port map( D => n4567, CK => CLK, RN => 
                           n6416, Q => n5590, QN => n2743);
   REGISTERS_reg_30_24_inst : DFFR_X1 port map( D => n4566, CK => CLK, RN => 
                           n6416, Q => n5591, QN => n2742);
   REGISTERS_reg_30_23_inst : DFFR_X1 port map( D => n4565, CK => CLK, RN => 
                           n6415, Q => n5592, QN => n2741);
   REGISTERS_reg_30_22_inst : DFFR_X1 port map( D => n4564, CK => CLK, RN => 
                           n6415, Q => n5593, QN => n2740);
   REGISTERS_reg_30_21_inst : DFFR_X1 port map( D => n4563, CK => CLK, RN => 
                           n6415, Q => n5594, QN => n2739);
   REGISTERS_reg_30_20_inst : DFFR_X1 port map( D => n4562, CK => CLK, RN => 
                           n6415, Q => n5595, QN => n2738);
   REGISTERS_reg_30_19_inst : DFFR_X1 port map( D => n4561, CK => CLK, RN => 
                           n6415, Q => n5596, QN => n2737);
   REGISTERS_reg_30_18_inst : DFFR_X1 port map( D => n4560, CK => CLK, RN => 
                           n6415, Q => n5597, QN => n2736);
   REGISTERS_reg_30_17_inst : DFFR_X1 port map( D => n4559, CK => CLK, RN => 
                           n6415, Q => n5598, QN => n2735);
   REGISTERS_reg_30_16_inst : DFFR_X1 port map( D => n4558, CK => CLK, RN => 
                           n6415, Q => n5599, QN => n2734);
   REGISTERS_reg_30_15_inst : DFFR_X1 port map( D => n4557, CK => CLK, RN => 
                           n6415, Q => n5600, QN => n2733);
   REGISTERS_reg_30_14_inst : DFFR_X1 port map( D => n4556, CK => CLK, RN => 
                           n6415, Q => n5601, QN => n2732);
   REGISTERS_reg_30_13_inst : DFFR_X1 port map( D => n4555, CK => CLK, RN => 
                           n6415, Q => n5602, QN => n2731);
   REGISTERS_reg_30_12_inst : DFFR_X1 port map( D => n4554, CK => CLK, RN => 
                           n6415, Q => n5603, QN => n2730);
   REGISTERS_reg_30_11_inst : DFFR_X1 port map( D => n4553, CK => CLK, RN => 
                           n6414, Q => n5604, QN => n2729);
   REGISTERS_reg_30_10_inst : DFFR_X1 port map( D => n4552, CK => CLK, RN => 
                           n6414, Q => n5605, QN => n2728);
   REGISTERS_reg_30_9_inst : DFFR_X1 port map( D => n4551, CK => CLK, RN => 
                           n6414, Q => n5606, QN => n2727);
   REGISTERS_reg_30_8_inst : DFFR_X1 port map( D => n4550, CK => CLK, RN => 
                           n6414, Q => n5607, QN => n2726);
   REGISTERS_reg_30_7_inst : DFFR_X1 port map( D => n4549, CK => CLK, RN => 
                           n6414, Q => n5608, QN => n2725);
   REGISTERS_reg_30_6_inst : DFFR_X1 port map( D => n4548, CK => CLK, RN => 
                           n6414, Q => n5609, QN => n2724);
   REGISTERS_reg_30_5_inst : DFFR_X1 port map( D => n4547, CK => CLK, RN => 
                           n6414, Q => n5610, QN => n2723);
   REGISTERS_reg_30_4_inst : DFFR_X1 port map( D => n4546, CK => CLK, RN => 
                           n6414, Q => n5611, QN => n2722);
   REGISTERS_reg_30_3_inst : DFFR_X1 port map( D => n4545, CK => CLK, RN => 
                           n6414, Q => n5612, QN => n2721);
   REGISTERS_reg_30_2_inst : DFFR_X1 port map( D => n4544, CK => CLK, RN => 
                           n6414, Q => n5613, QN => n2720);
   REGISTERS_reg_30_1_inst : DFFR_X1 port map( D => n4543, CK => CLK, RN => 
                           n6414, Q => n5614, QN => n2719);
   REGISTERS_reg_30_0_inst : DFFR_X1 port map( D => n4542, CK => CLK, RN => 
                           n6414, Q => n5360, QN => n2718);
   REGISTERS_reg_20_31_inst : DFFR_X1 port map( D => n4445, CK => CLK, RN => 
                           n6384, Q => n5105, QN => n3581);
   REGISTERS_reg_20_30_inst : DFFR_X1 port map( D => n4444, CK => CLK, RN => 
                           n6384, Q => n5106, QN => n3580);
   REGISTERS_reg_20_29_inst : DFFR_X1 port map( D => n4443, CK => CLK, RN => 
                           n6384, Q => n5107, QN => n3579);
   REGISTERS_reg_20_28_inst : DFFR_X1 port map( D => n4442, CK => CLK, RN => 
                           n6384, Q => n5108, QN => n3578);
   REGISTERS_reg_20_27_inst : DFFR_X1 port map( D => n4441, CK => CLK, RN => 
                           n6384, Q => n5109, QN => n3577);
   REGISTERS_reg_20_26_inst : DFFR_X1 port map( D => n4440, CK => CLK, RN => 
                           n6384, Q => n5110, QN => n3576);
   REGISTERS_reg_20_25_inst : DFFR_X1 port map( D => n4439, CK => CLK, RN => 
                           n6383, Q => n5111, QN => n3575);
   REGISTERS_reg_20_24_inst : DFFR_X1 port map( D => n4438, CK => CLK, RN => 
                           n6383, Q => n5112, QN => n3574);
   REGISTERS_reg_20_23_inst : DFFR_X1 port map( D => n4437, CK => CLK, RN => 
                           n6383, Q => n5113, QN => n3573);
   REGISTERS_reg_20_22_inst : DFFR_X1 port map( D => n4436, CK => CLK, RN => 
                           n6383, Q => n5114, QN => n3572);
   REGISTERS_reg_20_21_inst : DFFR_X1 port map( D => n4435, CK => CLK, RN => 
                           n6383, Q => n5115, QN => n3571);
   REGISTERS_reg_20_20_inst : DFFR_X1 port map( D => n4434, CK => CLK, RN => 
                           n6383, Q => n5116, QN => n3570);
   REGISTERS_reg_20_19_inst : DFFR_X1 port map( D => n4433, CK => CLK, RN => 
                           n6383, Q => n5117, QN => n3569);
   REGISTERS_reg_20_18_inst : DFFR_X1 port map( D => n4432, CK => CLK, RN => 
                           n6383, Q => n5118, QN => n3568);
   REGISTERS_reg_20_17_inst : DFFR_X1 port map( D => n4431, CK => CLK, RN => 
                           n6383, Q => n5119, QN => n3567);
   REGISTERS_reg_20_16_inst : DFFR_X1 port map( D => n4430, CK => CLK, RN => 
                           n6383, Q => n5120, QN => n3566);
   REGISTERS_reg_20_15_inst : DFFR_X1 port map( D => n4429, CK => CLK, RN => 
                           n6383, Q => n5121, QN => n3565);
   REGISTERS_reg_20_14_inst : DFFR_X1 port map( D => n4428, CK => CLK, RN => 
                           n6383, Q => n5122, QN => n3564);
   REGISTERS_reg_20_13_inst : DFFR_X1 port map( D => n4427, CK => CLK, RN => 
                           n6382, Q => n5123, QN => n3563);
   REGISTERS_reg_20_12_inst : DFFR_X1 port map( D => n4426, CK => CLK, RN => 
                           n6382, Q => n5124, QN => n3562);
   REGISTERS_reg_20_11_inst : DFFR_X1 port map( D => n4425, CK => CLK, RN => 
                           n6382, Q => n5125, QN => n3561);
   REGISTERS_reg_20_10_inst : DFFR_X1 port map( D => n4424, CK => CLK, RN => 
                           n6382, Q => n5126, QN => n3560);
   REGISTERS_reg_20_9_inst : DFFR_X1 port map( D => n4423, CK => CLK, RN => 
                           n6382, Q => n5127, QN => n3559);
   REGISTERS_reg_20_8_inst : DFFR_X1 port map( D => n4422, CK => CLK, RN => 
                           n6382, Q => n5128, QN => n2982);
   REGISTERS_reg_20_7_inst : DFFR_X1 port map( D => n4421, CK => CLK, RN => 
                           n6382, Q => n5129, QN => n2981);
   REGISTERS_reg_20_6_inst : DFFR_X1 port map( D => n4420, CK => CLK, RN => 
                           n6382, Q => n5130, QN => n2980);
   REGISTERS_reg_20_5_inst : DFFR_X1 port map( D => n4419, CK => CLK, RN => 
                           n6382, Q => n5131, QN => n2979);
   REGISTERS_reg_20_4_inst : DFFR_X1 port map( D => n4418, CK => CLK, RN => 
                           n6382, Q => n5132, QN => n2978);
   REGISTERS_reg_20_3_inst : DFFR_X1 port map( D => n4417, CK => CLK, RN => 
                           n6393, Q => n5133, QN => n2977);
   REGISTERS_reg_20_2_inst : DFFR_X1 port map( D => n4416, CK => CLK, RN => 
                           n6393, Q => n5134, QN => n2976);
   REGISTERS_reg_20_1_inst : DFFR_X1 port map( D => n4415, CK => CLK, RN => 
                           n6393, Q => n5135, QN => n2975);
   REGISTERS_reg_20_0_inst : DFFR_X1 port map( D => n4414, CK => CLK, RN => 
                           n6393, Q => n5136, QN => n2974);
   REGISTERS_reg_16_31_inst : DFFR_X1 port map( D => n4381, CK => CLK, RN => 
                           n6453, Q => n5422, QN => n3677);
   REGISTERS_reg_16_30_inst : DFFR_X1 port map( D => n4380, CK => CLK, RN => 
                           n6453, Q => n5423, QN => n3676);
   REGISTERS_reg_16_29_inst : DFFR_X1 port map( D => n4379, CK => CLK, RN => 
                           n6453, Q => n5424, QN => n3675);
   REGISTERS_reg_16_28_inst : DFFR_X1 port map( D => n4378, CK => CLK, RN => 
                           n6453, Q => n5425, QN => n3674);
   REGISTERS_reg_16_27_inst : DFFR_X1 port map( D => n4377, CK => CLK, RN => 
                           n6453, Q => n5426, QN => n3673);
   REGISTERS_reg_16_26_inst : DFFR_X1 port map( D => n4376, CK => CLK, RN => 
                           n6453, Q => n5427, QN => n3672);
   REGISTERS_reg_16_25_inst : DFFR_X1 port map( D => n4375, CK => CLK, RN => 
                           n6453, Q => n5428, QN => n3671);
   REGISTERS_reg_16_24_inst : DFFR_X1 port map( D => n4374, CK => CLK, RN => 
                           n6453, Q => n5429, QN => n3670);
   REGISTERS_reg_16_23_inst : DFFR_X1 port map( D => n4373, CK => CLK, RN => 
                           n6452, Q => n5430, QN => n3669);
   REGISTERS_reg_16_22_inst : DFFR_X1 port map( D => n4372, CK => CLK, RN => 
                           n6452, Q => n5431, QN => n3668);
   REGISTERS_reg_16_21_inst : DFFR_X1 port map( D => n4371, CK => CLK, RN => 
                           n6452, Q => n5432, QN => n3667);
   REGISTERS_reg_16_20_inst : DFFR_X1 port map( D => n4370, CK => CLK, RN => 
                           n6452, Q => n5433, QN => n3666);
   REGISTERS_reg_16_19_inst : DFFR_X1 port map( D => n4369, CK => CLK, RN => 
                           n6464, Q => n5434, QN => n3665);
   REGISTERS_reg_16_18_inst : DFFR_X1 port map( D => n4368, CK => CLK, RN => 
                           n6464, Q => n5435, QN => n3664);
   REGISTERS_reg_16_17_inst : DFFR_X1 port map( D => n4367, CK => CLK, RN => 
                           n6464, Q => n5436, QN => n3663);
   REGISTERS_reg_16_16_inst : DFFR_X1 port map( D => n4366, CK => CLK, RN => 
                           n6464, Q => n5437, QN => n3662);
   REGISTERS_reg_16_15_inst : DFFR_X1 port map( D => n4365, CK => CLK, RN => 
                           n6464, Q => n5438, QN => n3661);
   REGISTERS_reg_16_14_inst : DFFR_X1 port map( D => n4364, CK => CLK, RN => 
                           n6464, Q => n5439, QN => n3660);
   REGISTERS_reg_16_13_inst : DFFR_X1 port map( D => n4363, CK => CLK, RN => 
                           n6464, Q => n5440, QN => n3659);
   REGISTERS_reg_16_12_inst : DFFR_X1 port map( D => n4362, CK => CLK, RN => 
                           n6464, Q => n5441, QN => n3658);
   REGISTERS_reg_16_11_inst : DFFR_X1 port map( D => n4361, CK => CLK, RN => 
                           n6463, Q => n5442, QN => n3657);
   REGISTERS_reg_16_10_inst : DFFR_X1 port map( D => n4360, CK => CLK, RN => 
                           n6463, Q => n5443, QN => n3656);
   REGISTERS_reg_16_9_inst : DFFR_X1 port map( D => n4359, CK => CLK, RN => 
                           n6463, Q => n5444, QN => n3655);
   REGISTERS_reg_16_8_inst : DFFR_X1 port map( D => n4358, CK => CLK, RN => 
                           n6463, Q => n5445, QN => n3654);
   REGISTERS_reg_16_7_inst : DFFR_X1 port map( D => n4357, CK => CLK, RN => 
                           n6463, Q => n5446, QN => n3653);
   REGISTERS_reg_16_6_inst : DFFR_X1 port map( D => n4356, CK => CLK, RN => 
                           n6463, Q => n5447, QN => n3652);
   REGISTERS_reg_16_5_inst : DFFR_X1 port map( D => n4355, CK => CLK, RN => 
                           n6463, Q => n5448, QN => n3651);
   REGISTERS_reg_16_4_inst : DFFR_X1 port map( D => n4354, CK => CLK, RN => 
                           n6463, Q => n5449, QN => n3650);
   REGISTERS_reg_16_3_inst : DFFR_X1 port map( D => n4353, CK => CLK, RN => 
                           n6462, Q => n5450, QN => n3649);
   REGISTERS_reg_16_2_inst : DFFR_X1 port map( D => n4352, CK => CLK, RN => 
                           n6462, Q => n5451, QN => n3648);
   REGISTERS_reg_16_1_inst : DFFR_X1 port map( D => n4351, CK => CLK, RN => 
                           n6462, Q => n5452, QN => n3647);
   REGISTERS_reg_16_0_inst : DFFR_X1 port map( D => n4350, CK => CLK, RN => 
                           n6462, Q => n5547, QN => n3646);
   REGISTERS_reg_13_31_inst : DFFR_X1 port map( D => n4253, CK => CLK, RN => 
                           n6449, Q => n5873, QN => n3773);
   REGISTERS_reg_13_30_inst : DFFR_X1 port map( D => n4252, CK => CLK, RN => 
                           n6449, Q => n5328, QN => n3772);
   REGISTERS_reg_13_29_inst : DFFR_X1 port map( D => n4251, CK => CLK, RN => 
                           n6449, Q => n5329, QN => n3771);
   REGISTERS_reg_13_28_inst : DFFR_X1 port map( D => n4250, CK => CLK, RN => 
                           n6449, Q => n5330, QN => n3770);
   REGISTERS_reg_13_27_inst : DFFR_X1 port map( D => n4249, CK => CLK, RN => 
                           n6449, Q => n5331, QN => n3769);
   REGISTERS_reg_13_26_inst : DFFR_X1 port map( D => n4248, CK => CLK, RN => 
                           n6449, Q => n5332, QN => n3768);
   REGISTERS_reg_13_25_inst : DFFR_X1 port map( D => n4247, CK => CLK, RN => 
                           n6449, Q => n5333, QN => n3767);
   REGISTERS_reg_13_24_inst : DFFR_X1 port map( D => n4246, CK => CLK, RN => 
                           n6449, Q => n5334, QN => n3766);
   REGISTERS_reg_13_23_inst : DFFR_X1 port map( D => n4245, CK => CLK, RN => 
                           n6448, Q => n5335, QN => n3765);
   REGISTERS_reg_13_22_inst : DFFR_X1 port map( D => n4244, CK => CLK, RN => 
                           n6448, Q => n5336, QN => n3764);
   REGISTERS_reg_13_21_inst : DFFR_X1 port map( D => n4243, CK => CLK, RN => 
                           n6448, Q => n5337, QN => n3763);
   REGISTERS_reg_13_20_inst : DFFR_X1 port map( D => n4242, CK => CLK, RN => 
                           n6448, Q => n5338, QN => n3762);
   REGISTERS_reg_13_19_inst : DFFR_X1 port map( D => n4241, CK => CLK, RN => 
                           n6448, Q => n5339, QN => n3761);
   REGISTERS_reg_13_18_inst : DFFR_X1 port map( D => n4240, CK => CLK, RN => 
                           n6448, Q => n5340, QN => n3760);
   REGISTERS_reg_13_17_inst : DFFR_X1 port map( D => n4239, CK => CLK, RN => 
                           n6448, Q => n5341, QN => n3759);
   REGISTERS_reg_13_16_inst : DFFR_X1 port map( D => n4238, CK => CLK, RN => 
                           n6448, Q => n5342, QN => n3758);
   REGISTERS_reg_13_15_inst : DFFR_X1 port map( D => n4237, CK => CLK, RN => 
                           n6448, Q => n5343, QN => n3757);
   REGISTERS_reg_13_14_inst : DFFR_X1 port map( D => n4236, CK => CLK, RN => 
                           n6448, Q => n5344, QN => n3756);
   REGISTERS_reg_13_13_inst : DFFR_X1 port map( D => n4235, CK => CLK, RN => 
                           n6448, Q => n5345, QN => n3755);
   REGISTERS_reg_13_12_inst : DFFR_X1 port map( D => n4234, CK => CLK, RN => 
                           n6448, Q => n5346, QN => n3754);
   REGISTERS_reg_13_11_inst : DFFR_X1 port map( D => n4233, CK => CLK, RN => 
                           n6447, Q => n5347, QN => n3753);
   REGISTERS_reg_13_10_inst : DFFR_X1 port map( D => n4232, CK => CLK, RN => 
                           n6447, Q => n5348, QN => n3752);
   REGISTERS_reg_13_9_inst : DFFR_X1 port map( D => n4231, CK => CLK, RN => 
                           n6447, Q => n5349, QN => n3751);
   REGISTERS_reg_13_8_inst : DFFR_X1 port map( D => n4230, CK => CLK, RN => 
                           n6447, Q => n5350, QN => n3750);
   REGISTERS_reg_13_7_inst : DFFR_X1 port map( D => n4229, CK => CLK, RN => 
                           n6447, Q => n5351, QN => n3749);
   REGISTERS_reg_13_6_inst : DFFR_X1 port map( D => n4228, CK => CLK, RN => 
                           n6447, Q => n5352, QN => n3748);
   REGISTERS_reg_13_5_inst : DFFR_X1 port map( D => n4227, CK => CLK, RN => 
                           n6447, Q => n5353, QN => n3747);
   REGISTERS_reg_13_4_inst : DFFR_X1 port map( D => n4226, CK => CLK, RN => 
                           n6447, Q => n5354, QN => n3746);
   REGISTERS_reg_13_3_inst : DFFR_X1 port map( D => n4225, CK => CLK, RN => 
                           n6446, Q => n5355, QN => n3745);
   REGISTERS_reg_13_2_inst : DFFR_X1 port map( D => n4224, CK => CLK, RN => 
                           n6446, Q => n5356, QN => n3744);
   REGISTERS_reg_13_1_inst : DFFR_X1 port map( D => n4223, CK => CLK, RN => 
                           n6446, Q => n5357, QN => n3743);
   REGISTERS_reg_13_0_inst : DFFR_X1 port map( D => n4222, CK => CLK, RN => 
                           n6446, Q => n5874, QN => n3742);
   REGISTERS_reg_9_31_inst : DFFR_X1 port map( D => n4189, CK => CLK, RN => 
                           n6436, Q => n5841, QN => n3901);
   REGISTERS_reg_9_30_inst : DFFR_X1 port map( D => n4188, CK => CLK, RN => 
                           n6436, Q => n5842, QN => n3900);
   REGISTERS_reg_9_29_inst : DFFR_X1 port map( D => n4187, CK => CLK, RN => 
                           n6436, Q => n5843, QN => n3899);
   REGISTERS_reg_9_28_inst : DFFR_X1 port map( D => n4186, CK => CLK, RN => 
                           n6436, Q => n5844, QN => n3898);
   REGISTERS_reg_9_27_inst : DFFR_X1 port map( D => n4185, CK => CLK, RN => 
                           n6435, Q => n5845, QN => n3897);
   REGISTERS_reg_9_26_inst : DFFR_X1 port map( D => n4184, CK => CLK, RN => 
                           n6435, Q => n5846, QN => n3896);
   REGISTERS_reg_9_25_inst : DFFR_X1 port map( D => n4183, CK => CLK, RN => 
                           n6435, Q => n5847, QN => n3895);
   REGISTERS_reg_9_24_inst : DFFR_X1 port map( D => n4182, CK => CLK, RN => 
                           n6435, Q => n5848, QN => n3894);
   REGISTERS_reg_9_23_inst : DFFR_X1 port map( D => n4181, CK => CLK, RN => 
                           n6435, Q => n5849, QN => n3893);
   REGISTERS_reg_9_22_inst : DFFR_X1 port map( D => n4180, CK => CLK, RN => 
                           n6435, Q => n5850, QN => n3892);
   REGISTERS_reg_9_21_inst : DFFR_X1 port map( D => n4179, CK => CLK, RN => 
                           n6435, Q => n5851, QN => n3891);
   REGISTERS_reg_9_20_inst : DFFR_X1 port map( D => n4178, CK => CLK, RN => 
                           n6435, Q => n5852, QN => n3890);
   REGISTERS_reg_9_19_inst : DFFR_X1 port map( D => n4177, CK => CLK, RN => 
                           n6435, Q => n5853, QN => n3889);
   REGISTERS_reg_9_18_inst : DFFR_X1 port map( D => n4176, CK => CLK, RN => 
                           n6435, Q => n5854, QN => n3888);
   REGISTERS_reg_9_17_inst : DFFR_X1 port map( D => n4175, CK => CLK, RN => 
                           n6435, Q => n5855, QN => n3887);
   REGISTERS_reg_9_16_inst : DFFR_X1 port map( D => n4174, CK => CLK, RN => 
                           n6435, Q => n5856, QN => n3886);
   REGISTERS_reg_9_15_inst : DFFR_X1 port map( D => n4173, CK => CLK, RN => 
                           n6434, Q => n5857, QN => n3885);
   REGISTERS_reg_9_14_inst : DFFR_X1 port map( D => n4172, CK => CLK, RN => 
                           n6434, Q => n5858, QN => n3884);
   REGISTERS_reg_9_13_inst : DFFR_X1 port map( D => n4171, CK => CLK, RN => 
                           n6434, Q => n5859, QN => n3883);
   REGISTERS_reg_9_12_inst : DFFR_X1 port map( D => n4170, CK => CLK, RN => 
                           n6434, Q => n5860, QN => n3882);
   REGISTERS_reg_9_11_inst : DFFR_X1 port map( D => n4169, CK => CLK, RN => 
                           n6446, Q => n5861, QN => n3881);
   REGISTERS_reg_9_10_inst : DFFR_X1 port map( D => n4168, CK => CLK, RN => 
                           n6446, Q => n5862, QN => n3880);
   REGISTERS_reg_9_9_inst : DFFR_X1 port map( D => n4167, CK => CLK, RN => 
                           n6446, Q => n5863, QN => n3879);
   REGISTERS_reg_9_8_inst : DFFR_X1 port map( D => n4166, CK => CLK, RN => 
                           n6446, Q => n5864, QN => n3878);
   REGISTERS_reg_9_7_inst : DFFR_X1 port map( D => n4165, CK => CLK, RN => 
                           n6446, Q => n5865, QN => n3877);
   REGISTERS_reg_9_6_inst : DFFR_X1 port map( D => n4164, CK => CLK, RN => 
                           n6446, Q => n5866, QN => n3876);
   REGISTERS_reg_9_5_inst : DFFR_X1 port map( D => n4163, CK => CLK, RN => 
                           n6446, Q => n5867, QN => n3875);
   REGISTERS_reg_9_4_inst : DFFR_X1 port map( D => n4162, CK => CLK, RN => 
                           n6446, Q => n5868, QN => n3874);
   REGISTERS_reg_9_3_inst : DFFR_X1 port map( D => n4161, CK => CLK, RN => 
                           n6445, Q => n5869, QN => n3873);
   REGISTERS_reg_9_2_inst : DFFR_X1 port map( D => n4160, CK => CLK, RN => 
                           n6445, Q => n5870, QN => n3872);
   REGISTERS_reg_9_1_inst : DFFR_X1 port map( D => n4159, CK => CLK, RN => 
                           n6445, Q => n5871, QN => n3871);
   REGISTERS_reg_9_0_inst : DFFR_X1 port map( D => n4158, CK => CLK, RN => 
                           n6445, Q => n5872, QN => n3870);
   REGISTERS_reg_1_31_inst : DFFR_X1 port map( D => n4285, CK => CLK, RN => 
                           n6422, Q => n5169, QN => n4094);
   REGISTERS_reg_1_30_inst : DFFR_X1 port map( D => n4284, CK => CLK, RN => 
                           n6422, Q => n5203, QN => n4095);
   REGISTERS_reg_1_29_inst : DFFR_X1 port map( D => n4283, CK => CLK, RN => 
                           n6422, Q => n5204, QN => n4096);
   REGISTERS_reg_1_28_inst : DFFR_X1 port map( D => n4282, CK => CLK, RN => 
                           n6422, Q => n5205, QN => n4097);
   REGISTERS_reg_1_27_inst : DFFR_X1 port map( D => n4281, CK => CLK, RN => 
                           n6422, Q => n5206, QN => n4098);
   REGISTERS_reg_1_26_inst : DFFR_X1 port map( D => n4280, CK => CLK, RN => 
                           n6422, Q => n5207, QN => n4099);
   REGISTERS_reg_1_25_inst : DFFR_X1 port map( D => n4279, CK => CLK, RN => 
                           n6422, Q => n5208, QN => n4100);
   REGISTERS_reg_1_24_inst : DFFR_X1 port map( D => n4278, CK => CLK, RN => 
                           n6422, Q => n5209, QN => n4101);
   REGISTERS_reg_1_23_inst : DFFR_X1 port map( D => n4277, CK => CLK, RN => 
                           n6421, Q => n5210, QN => n4102);
   REGISTERS_reg_1_22_inst : DFFR_X1 port map( D => n4276, CK => CLK, RN => 
                           n6421, Q => n5211, QN => n4103);
   REGISTERS_reg_1_21_inst : DFFR_X1 port map( D => n4275, CK => CLK, RN => 
                           n6421, Q => n5212, QN => n4104);
   REGISTERS_reg_1_20_inst : DFFR_X1 port map( D => n4274, CK => CLK, RN => 
                           n6421, Q => n5213, QN => n4105);
   REGISTERS_reg_1_19_inst : DFFR_X1 port map( D => n4273, CK => CLK, RN => 
                           n6421, Q => n5214, QN => n4106);
   REGISTERS_reg_1_18_inst : DFFR_X1 port map( D => n4272, CK => CLK, RN => 
                           n6421, Q => n5215, QN => n4107);
   REGISTERS_reg_1_17_inst : DFFR_X1 port map( D => n4271, CK => CLK, RN => 
                           n6421, Q => n5216, QN => n4108);
   REGISTERS_reg_1_16_inst : DFFR_X1 port map( D => n4270, CK => CLK, RN => 
                           n6421, Q => n5217, QN => n4109);
   REGISTERS_reg_1_15_inst : DFFR_X1 port map( D => n4269, CK => CLK, RN => 
                           n6421, Q => n5218, QN => n4110);
   REGISTERS_reg_1_14_inst : DFFR_X1 port map( D => n4268, CK => CLK, RN => 
                           n6421, Q => n5219, QN => n4111);
   REGISTERS_reg_1_13_inst : DFFR_X1 port map( D => n4267, CK => CLK, RN => 
                           n6421, Q => n5220, QN => n4112);
   REGISTERS_reg_1_12_inst : DFFR_X1 port map( D => n4266, CK => CLK, RN => 
                           n6421, Q => n5221, QN => n4113);
   REGISTERS_reg_1_11_inst : DFFR_X1 port map( D => n4265, CK => CLK, RN => 
                           n6420, Q => n5222, QN => n4114);
   REGISTERS_reg_1_10_inst : DFFR_X1 port map( D => n4264, CK => CLK, RN => 
                           n6420, Q => n5223, QN => n4115);
   REGISTERS_reg_1_9_inst : DFFR_X1 port map( D => n4263, CK => CLK, RN => 
                           n6420, Q => n5224, QN => n4116);
   REGISTERS_reg_1_8_inst : DFFR_X1 port map( D => n4262, CK => CLK, RN => 
                           n6420, Q => n5225, QN => n4117);
   REGISTERS_reg_1_7_inst : DFFR_X1 port map( D => n4261, CK => CLK, RN => 
                           n6420, Q => n5226, QN => n4118);
   REGISTERS_reg_1_6_inst : DFFR_X1 port map( D => n4260, CK => CLK, RN => 
                           n6420, Q => n5227, QN => n4119);
   REGISTERS_reg_1_5_inst : DFFR_X1 port map( D => n4259, CK => CLK, RN => 
                           n6420, Q => n5228, QN => n4120);
   REGISTERS_reg_1_4_inst : DFFR_X1 port map( D => n4258, CK => CLK, RN => 
                           n6420, Q => n5229, QN => n4121);
   REGISTERS_reg_1_3_inst : DFFR_X1 port map( D => n4257, CK => CLK, RN => 
                           n6419, Q => n5230, QN => n4122);
   REGISTERS_reg_1_2_inst : DFFR_X1 port map( D => n4256, CK => CLK, RN => 
                           n6419, Q => n5231, QN => n4123);
   REGISTERS_reg_1_1_inst : DFFR_X1 port map( D => n4255, CK => CLK, RN => 
                           n6419, Q => n5232, QN => n4124);
   REGISTERS_reg_1_0_inst : DFFR_X1 port map( D => n4254, CK => CLK, RN => 
                           n6419, Q => n5170, QN => n4125);
   REGISTERS_reg_23_31_inst : DFFR_X1 port map( D => n3206, CK => CLK, RN => 
                           RST, Q => n4750, QN => n7521);
   REGISTERS_reg_23_30_inst : DFFR_X1 port map( D => n7683, CK => CLK, RN => 
                           n6389, Q => n4748, QN => n7498);
   REGISTERS_reg_23_29_inst : DFFR_X1 port map( D => n7684, CK => CLK, RN => 
                           n6388, Q => n4742, QN => n7479);
   REGISTERS_reg_23_28_inst : DFFR_X1 port map( D => n7685, CK => CLK, RN => 
                           n6388, Q => n4744, QN => n7460);
   REGISTERS_reg_23_27_inst : DFFR_X1 port map( D => n7686, CK => CLK, RN => 
                           n6400, Q => n4746, QN => n7441);
   REGISTERS_reg_23_26_inst : DFFR_X1 port map( D => n7687, CK => CLK, RN => 
                           n6399, Q => n4736, QN => n7422);
   REGISTERS_reg_23_25_inst : DFFR_X1 port map( D => n7688, CK => CLK, RN => 
                           n6399, Q => n4738, QN => n7403);
   REGISTERS_reg_23_24_inst : DFFR_X1 port map( D => n7689, CK => CLK, RN => 
                           n6399, Q => n4740, QN => n7384);
   REGISTERS_reg_23_23_inst : DFFR_X1 port map( D => n7690, CK => CLK, RN => 
                           n6399, Q => n4730, QN => n7365);
   REGISTERS_reg_23_22_inst : DFFR_X1 port map( D => n7691, CK => CLK, RN => 
                           n6399, Q => n4732, QN => n7346);
   REGISTERS_reg_23_21_inst : DFFR_X1 port map( D => n7692, CK => CLK, RN => 
                           n6399, Q => n4734, QN => n7327);
   REGISTERS_reg_23_20_inst : DFFR_X1 port map( D => n7693, CK => CLK, RN => 
                           n6399, Q => n4724, QN => n7308);
   REGISTERS_reg_23_19_inst : DFFR_X1 port map( D => n7694, CK => CLK, RN => 
                           n6399, Q => n4726, QN => n7289);
   REGISTERS_reg_23_18_inst : DFFR_X1 port map( D => n7695, CK => CLK, RN => 
                           n6399, Q => n4728, QN => n7270);
   REGISTERS_reg_23_17_inst : DFFR_X1 port map( D => n7696, CK => CLK, RN => 
                           n6399, Q => n4718, QN => n7251);
   REGISTERS_reg_23_16_inst : DFFR_X1 port map( D => n7697, CK => CLK, RN => 
                           n6399, Q => n4720, QN => n7232);
   REGISTERS_reg_23_15_inst : DFFR_X1 port map( D => n7698, CK => CLK, RN => 
                           n6399, Q => n4722, QN => n7213);
   REGISTERS_reg_23_14_inst : DFFR_X1 port map( D => n7699, CK => CLK, RN => 
                           n6398, Q => n4712, QN => n7194);
   REGISTERS_reg_23_13_inst : DFFR_X1 port map( D => n7700, CK => CLK, RN => 
                           n6398, Q => n4714, QN => n7175);
   REGISTERS_reg_23_12_inst : DFFR_X1 port map( D => n7701, CK => CLK, RN => 
                           n6398, Q => n4716, QN => n7156);
   REGISTERS_reg_23_11_inst : DFFR_X1 port map( D => n7702, CK => CLK, RN => 
                           n6398, Q => n4706, QN => n7137);
   REGISTERS_reg_23_10_inst : DFFR_X1 port map( D => n7703, CK => CLK, RN => 
                           n6398, Q => n4708, QN => n7118);
   REGISTERS_reg_23_9_inst : DFFR_X1 port map( D => n7704, CK => CLK, RN => 
                           n6398, Q => n4710, QN => n7099);
   REGISTERS_reg_23_8_inst : DFFR_X1 port map( D => n7705, CK => CLK, RN => 
                           n6398, Q => n4700, QN => n7080);
   REGISTERS_reg_23_7_inst : DFFR_X1 port map( D => n7706, CK => CLK, RN => 
                           n6398, Q => n4702, QN => n7061);
   REGISTERS_reg_23_6_inst : DFFR_X1 port map( D => n7707, CK => CLK, RN => 
                           n6398, Q => n4704, QN => n7042);
   REGISTERS_reg_23_5_inst : DFFR_X1 port map( D => n7708, CK => CLK, RN => 
                           n6398, Q => n4696, QN => n7023);
   REGISTERS_reg_23_4_inst : DFFR_X1 port map( D => n7709, CK => CLK, RN => 
                           n6398, Q => n4698, QN => n7004);
   REGISTERS_reg_22_31_inst : DFFR_X1 port map( D => n3238, CK => CLK, RN => 
                           n6391, Q => n2941, QN => n5941);
   REGISTERS_reg_22_30_inst : DFFR_X1 port map( D => n3237, CK => CLK, RN => 
                           n6391, Q => n2940, QN => n5942);
   REGISTERS_reg_22_29_inst : DFFR_X1 port map( D => n3236, CK => CLK, RN => 
                           n6390, Q => n2939, QN => n5943);
   REGISTERS_reg_22_28_inst : DFFR_X1 port map( D => n3235, CK => CLK, RN => 
                           n6390, Q => n2938, QN => n5944);
   REGISTERS_reg_22_27_inst : DFFR_X1 port map( D => n3234, CK => CLK, RN => 
                           n6390, Q => n2937, QN => n5945);
   REGISTERS_reg_22_26_inst : DFFR_X1 port map( D => n3233, CK => CLK, RN => 
                           n6390, Q => n2936, QN => n5946);
   REGISTERS_reg_22_25_inst : DFFR_X1 port map( D => n3232, CK => CLK, RN => 
                           n6390, Q => n2935, QN => n5947);
   REGISTERS_reg_22_24_inst : DFFR_X1 port map( D => n3231, CK => CLK, RN => 
                           n6390, Q => n2934, QN => n5948);
   REGISTERS_reg_22_23_inst : DFFR_X1 port map( D => n3230, CK => CLK, RN => 
                           n6390, Q => n2933, QN => n5949);
   REGISTERS_reg_22_22_inst : DFFR_X1 port map( D => n3229, CK => CLK, RN => 
                           n6390, Q => n2932, QN => n5950);
   REGISTERS_reg_22_21_inst : DFFR_X1 port map( D => n3228, CK => CLK, RN => 
                           n6390, Q => n2931, QN => n5951);
   REGISTERS_reg_22_20_inst : DFFR_X1 port map( D => n3227, CK => CLK, RN => 
                           n6390, Q => n2930, QN => n5952);
   REGISTERS_reg_22_19_inst : DFFR_X1 port map( D => n3226, CK => CLK, RN => 
                           n6390, Q => n2929, QN => n5953);
   REGISTERS_reg_22_18_inst : DFFR_X1 port map( D => n3225, CK => CLK, RN => 
                           n6390, Q => n2928, QN => n5954);
   REGISTERS_reg_22_17_inst : DFFR_X1 port map( D => n3224, CK => CLK, RN => 
                           n6389, Q => n2927, QN => n5955);
   REGISTERS_reg_22_16_inst : DFFR_X1 port map( D => n3223, CK => CLK, RN => 
                           n6389, Q => n2926, QN => n5956);
   REGISTERS_reg_22_15_inst : DFFR_X1 port map( D => n3222, CK => CLK, RN => 
                           n6389, Q => n2925, QN => n5957);
   REGISTERS_reg_22_14_inst : DFFR_X1 port map( D => n3221, CK => CLK, RN => 
                           n6389, Q => n2924, QN => n5958);
   REGISTERS_reg_22_13_inst : DFFR_X1 port map( D => n3220, CK => CLK, RN => 
                           n6389, Q => n2923, QN => n5959);
   REGISTERS_reg_22_12_inst : DFFR_X1 port map( D => n3219, CK => CLK, RN => 
                           n6389, Q => n2922, QN => n5960);
   REGISTERS_reg_22_11_inst : DFFR_X1 port map( D => n3218, CK => CLK, RN => 
                           n6389, Q => n2921, QN => n5961);
   REGISTERS_reg_22_10_inst : DFFR_X1 port map( D => n3217, CK => CLK, RN => 
                           n6389, Q => n2920, QN => n5962);
   REGISTERS_reg_22_9_inst : DFFR_X1 port map( D => n3216, CK => CLK, RN => 
                           n6389, Q => n2919, QN => n5963);
   REGISTERS_reg_22_8_inst : DFFR_X1 port map( D => n3215, CK => CLK, RN => 
                           n6389, Q => n2918, QN => n5964);
   REGISTERS_reg_22_7_inst : DFFR_X1 port map( D => n3214, CK => CLK, RN => 
                           n6388, Q => n2917, QN => n5965);
   REGISTERS_reg_22_6_inst : DFFR_X1 port map( D => n3213, CK => CLK, RN => 
                           n6388, Q => n2916, QN => n5966);
   REGISTERS_reg_22_5_inst : DFFR_X1 port map( D => n3212, CK => CLK, RN => 
                           n6388, Q => n2915, QN => n5967);
   REGISTERS_reg_22_4_inst : DFFR_X1 port map( D => n3211, CK => CLK, RN => 
                           n6388, Q => n2914, QN => n5968);
   REGISTERS_reg_22_3_inst : DFFR_X1 port map( D => n3210, CK => CLK, RN => 
                           n6388, Q => n2913, QN => n5969);
   REGISTERS_reg_22_2_inst : DFFR_X1 port map( D => n3209, CK => CLK, RN => 
                           n6388, Q => n2912, QN => n5970);
   REGISTERS_reg_22_1_inst : DFFR_X1 port map( D => n3208, CK => CLK, RN => 
                           n6388, Q => n2911, QN => n5971);
   REGISTERS_reg_22_0_inst : DFFR_X1 port map( D => n3207, CK => CLK, RN => 
                           n6388, Q => n2910, QN => n5972);
   REGISTERS_reg_7_31_inst : DFFR_X1 port map( D => n7710, CK => CLK, RN => 
                           n6429, Q => n4814, QN => n7535);
   REGISTERS_reg_7_30_inst : DFFR_X1 port map( D => n7711, CK => CLK, RN => 
                           n6429, Q => n4780, QN => n7505);
   REGISTERS_reg_7_29_inst : DFFR_X1 port map( D => n7712, CK => CLK, RN => 
                           n6429, Q => n4776, QN => n7486);
   REGISTERS_reg_7_28_inst : DFFR_X1 port map( D => n7713, CK => CLK, RN => 
                           n6429, Q => n4778, QN => n7467);
   REGISTERS_reg_7_27_inst : DFFR_X1 port map( D => n7714, CK => CLK, RN => 
                           n6429, Q => n4754, QN => n7448);
   REGISTERS_reg_7_26_inst : DFFR_X1 port map( D => n7715, CK => CLK, RN => 
                           n6429, Q => n4772, QN => n7429);
   REGISTERS_reg_7_25_inst : DFFR_X1 port map( D => n7716, CK => CLK, RN => 
                           n6429, Q => n4774, QN => n7410);
   REGISTERS_reg_7_24_inst : DFFR_X1 port map( D => n7717, CK => CLK, RN => 
                           n6429, Q => n4766, QN => n7391);
   REGISTERS_reg_7_23_inst : DFFR_X1 port map( D => n7718, CK => CLK, RN => 
                           n6428, Q => n4770, QN => n7372);
   REGISTERS_reg_7_22_inst : DFFR_X1 port map( D => n7719, CK => CLK, RN => 
                           n6428, Q => n4764, QN => n7353);
   REGISTERS_reg_7_21_inst : DFFR_X1 port map( D => n7720, CK => CLK, RN => 
                           n6428, Q => n4760, QN => n7334);
   REGISTERS_reg_7_20_inst : DFFR_X1 port map( D => n7721, CK => CLK, RN => 
                           n6428, Q => n4768, QN => n7315);
   REGISTERS_reg_7_19_inst : DFFR_X1 port map( D => n7722, CK => CLK, RN => 
                           n6440, Q => n4758, QN => n7296);
   REGISTERS_reg_7_18_inst : DFFR_X1 port map( D => n7723, CK => CLK, RN => 
                           n6440, Q => n4756, QN => n7277);
   REGISTERS_reg_7_17_inst : DFFR_X1 port map( D => n7724, CK => CLK, RN => 
                           n6440, Q => n4762, QN => n7258);
   REGISTERS_reg_7_16_inst : DFFR_X1 port map( D => n7725, CK => CLK, RN => 
                           n6440, Q => n4752, QN => n7239);
   REGISTERS_reg_7_15_inst : DFFR_X1 port map( D => n7726, CK => CLK, RN => 
                           n6440, Q => n4782, QN => n7220);
   REGISTERS_reg_7_14_inst : DFFR_X1 port map( D => n7727, CK => CLK, RN => 
                           n6440, Q => n4784, QN => n7201);
   REGISTERS_reg_7_13_inst : DFFR_X1 port map( D => n7728, CK => CLK, RN => 
                           n6440, Q => n4786, QN => n7182);
   REGISTERS_reg_7_12_inst : DFFR_X1 port map( D => n7729, CK => CLK, RN => 
                           n6440, Q => n4788, QN => n7163);
   REGISTERS_reg_7_11_inst : DFFR_X1 port map( D => n7730, CK => CLK, RN => 
                           n6439, Q => n4790, QN => n7144);
   REGISTERS_reg_7_10_inst : DFFR_X1 port map( D => n7731, CK => CLK, RN => 
                           n6439, Q => n4792, QN => n7125);
   REGISTERS_reg_7_9_inst : DFFR_X1 port map( D => n7732, CK => CLK, RN => 
                           n6439, Q => n4794, QN => n7106);
   REGISTERS_reg_7_8_inst : DFFR_X1 port map( D => n7733, CK => CLK, RN => 
                           n6439, Q => n4796, QN => n7087);
   REGISTERS_reg_7_7_inst : DFFR_X1 port map( D => n7734, CK => CLK, RN => 
                           n6439, Q => n4798, QN => n7068);
   REGISTERS_reg_7_6_inst : DFFR_X1 port map( D => n7735, CK => CLK, RN => 
                           n6439, Q => n4800, QN => n7049);
   REGISTERS_reg_7_5_inst : DFFR_X1 port map( D => n7736, CK => CLK, RN => 
                           n6439, Q => n4802, QN => n7030);
   REGISTERS_reg_7_4_inst : DFFR_X1 port map( D => n7737, CK => CLK, RN => 
                           n6439, Q => n4804, QN => n7011);
   REGISTERS_reg_7_3_inst : DFFR_X1 port map( D => n7738, CK => CLK, RN => 
                           n6439, Q => n4806, QN => n6992);
   REGISTERS_reg_7_2_inst : DFFR_X1 port map( D => n7739, CK => CLK, RN => 
                           n6439, Q => n4808, QN => n6974);
   REGISTERS_reg_7_1_inst : DFFR_X1 port map( D => n7740, CK => CLK, RN => 
                           n6439, Q => n4810, QN => n6956);
   REGISTERS_reg_7_0_inst : DFFR_X1 port map( D => n7741, CK => CLK, RN => 
                           n6439, Q => n4812, QN => n6937);
   REGISTERS_reg_6_31_inst : DFFR_X1 port map( D => n7742, CK => CLK, RN => 
                           n6432, Q => n_1104, QN => n7534);
   REGISTERS_reg_6_30_inst : DFFR_X1 port map( D => n7743, CK => CLK, RN => 
                           n6432, Q => n_1105, QN => n7504);
   REGISTERS_reg_6_29_inst : DFFR_X1 port map( D => n7744, CK => CLK, RN => 
                           n6432, Q => n_1106, QN => n7485);
   REGISTERS_reg_6_28_inst : DFFR_X1 port map( D => n7745, CK => CLK, RN => 
                           n6432, Q => n_1107, QN => n7466);
   REGISTERS_reg_6_27_inst : DFFR_X1 port map( D => n7746, CK => CLK, RN => 
                           n6432, Q => n_1108, QN => n7447);
   REGISTERS_reg_6_26_inst : DFFR_X1 port map( D => n7747, CK => CLK, RN => 
                           n6432, Q => n_1109, QN => n7428);
   REGISTERS_reg_6_25_inst : DFFR_X1 port map( D => n7748, CK => CLK, RN => 
                           n6432, Q => n_1110, QN => n7409);
   REGISTERS_reg_6_24_inst : DFFR_X1 port map( D => n7749, CK => CLK, RN => 
                           n6432, Q => n_1111, QN => n7390);
   REGISTERS_reg_6_23_inst : DFFR_X1 port map( D => n7750, CK => CLK, RN => 
                           n6431, Q => n_1112, QN => n7371);
   REGISTERS_reg_6_22_inst : DFFR_X1 port map( D => n7751, CK => CLK, RN => 
                           n6431, Q => n_1113, QN => n7352);
   REGISTERS_reg_6_21_inst : DFFR_X1 port map( D => n7752, CK => CLK, RN => 
                           n6431, Q => n_1114, QN => n7333);
   REGISTERS_reg_6_20_inst : DFFR_X1 port map( D => n7753, CK => CLK, RN => 
                           n6431, Q => n_1115, QN => n7314);
   REGISTERS_reg_6_19_inst : DFFR_X1 port map( D => n7754, CK => CLK, RN => 
                           n6431, Q => n_1116, QN => n7295);
   REGISTERS_reg_6_18_inst : DFFR_X1 port map( D => n7755, CK => CLK, RN => 
                           n6431, Q => n_1117, QN => n7276);
   REGISTERS_reg_6_17_inst : DFFR_X1 port map( D => n7756, CK => CLK, RN => 
                           n6431, Q => n_1118, QN => n7257);
   REGISTERS_reg_6_16_inst : DFFR_X1 port map( D => n7757, CK => CLK, RN => 
                           n6431, Q => n_1119, QN => n7238);
   REGISTERS_reg_6_15_inst : DFFR_X1 port map( D => n7758, CK => CLK, RN => 
                           n6430, Q => n_1120, QN => n7219);
   REGISTERS_reg_6_14_inst : DFFR_X1 port map( D => n7759, CK => CLK, RN => 
                           n6430, Q => n_1121, QN => n7200);
   REGISTERS_reg_6_13_inst : DFFR_X1 port map( D => n7760, CK => CLK, RN => 
                           n6430, Q => n_1122, QN => n7181);
   REGISTERS_reg_6_12_inst : DFFR_X1 port map( D => n7761, CK => CLK, RN => 
                           n6430, Q => n_1123, QN => n7162);
   REGISTERS_reg_6_11_inst : DFFR_X1 port map( D => n7762, CK => CLK, RN => 
                           n6430, Q => n_1124, QN => n7143);
   REGISTERS_reg_6_10_inst : DFFR_X1 port map( D => n7763, CK => CLK, RN => 
                           n6430, Q => n_1125, QN => n7124);
   REGISTERS_reg_6_9_inst : DFFR_X1 port map( D => n7764, CK => CLK, RN => 
                           n6430, Q => n_1126, QN => n7105);
   REGISTERS_reg_6_8_inst : DFFR_X1 port map( D => n7765, CK => CLK, RN => 
                           n6430, Q => n_1127, QN => n7086);
   REGISTERS_reg_6_7_inst : DFFR_X1 port map( D => n7766, CK => CLK, RN => 
                           n6430, Q => n_1128, QN => n7067);
   REGISTERS_reg_6_6_inst : DFFR_X1 port map( D => n7767, CK => CLK, RN => 
                           n6430, Q => n_1129, QN => n7048);
   REGISTERS_reg_6_5_inst : DFFR_X1 port map( D => n7768, CK => CLK, RN => 
                           n6430, Q => n_1130, QN => n7029);
   REGISTERS_reg_6_4_inst : DFFR_X1 port map( D => n7769, CK => CLK, RN => 
                           n6430, Q => n_1131, QN => n7010);
   REGISTERS_reg_6_3_inst : DFFR_X1 port map( D => n7770, CK => CLK, RN => 
                           n6429, Q => n_1132, QN => n6991);
   REGISTERS_reg_6_2_inst : DFFR_X1 port map( D => n7771, CK => CLK, RN => 
                           n6429, Q => n_1133, QN => n6973);
   REGISTERS_reg_6_1_inst : DFFR_X1 port map( D => n7772, CK => CLK, RN => 
                           n6429, Q => n_1134, QN => n6955);
   REGISTERS_reg_6_0_inst : DFFR_X1 port map( D => n7773, CK => CLK, RN => 
                           n6429, Q => n_1135, QN => n6936);
   REGISTERS_reg_3_31_inst : DFFR_X1 port map( D => n7774, CK => CLK, RN => 
                           n6428, Q => n4061, QN => n5909);
   REGISTERS_reg_3_30_inst : DFFR_X1 port map( D => n7775, CK => CLK, RN => 
                           n6428, Q => n4060, QN => n5911);
   REGISTERS_reg_3_29_inst : DFFR_X1 port map( D => n7776, CK => CLK, RN => 
                           n6428, Q => n4059, QN => n5912);
   REGISTERS_reg_3_28_inst : DFFR_X1 port map( D => n7777, CK => CLK, RN => 
                           n6428, Q => n4058, QN => n5913);
   REGISTERS_reg_3_27_inst : DFFR_X1 port map( D => n7778, CK => CLK, RN => 
                           n6428, Q => n4057, QN => n5914);
   U2 : AND2_X1 port map( A1 => n4662, A2 => ADD_WR(3), ZN => n4606);
   U3 : AND2_X1 port map( A1 => n4662, A2 => n7590, ZN => n4607);
   U4 : AND2_X1 port map( A1 => n6480, A2 => n7898, ZN => n4608);
   U5 : AND3_X1 port map( A1 => n749, A2 => ADD_WR(3), A3 => n7589, ZN => n4609
                           );
   U6 : AND3_X1 port map( A1 => ADD_RS1(0), A2 => ADD_RS1(4), A3 => n7592, ZN 
                           => n4610);
   U7 : AND2_X1 port map( A1 => n4663, A2 => ADD_WR(0), ZN => n4611);
   U8 : AND3_X1 port map( A1 => ADD_RS1(3), A2 => ADD_RS1(4), A3 => n7593, ZN 
                           => n4612);
   U9 : AND2_X1 port map( A1 => n6479, A2 => n7900, ZN => n4613);
   U10 : AND2_X1 port map( A1 => n4663, A2 => n6485, ZN => n4614);
   U11 : AND4_X1 port map( A1 => ADD_RS2(3), A2 => ADD_RS2(4), A3 => n6237, A4 
                           => n7595, ZN => n4615);
   U12 : AND4_X1 port map( A1 => n1999, A2 => n1997, A3 => n6173, A4 => n1998, 
                           ZN => n4616);
   U13 : AND4_X1 port map( A1 => ADD_RS2(0), A2 => ADD_RS2(4), A3 => n6237, A4 
                           => n7594, ZN => n4617);
   U14 : AND2_X1 port map( A1 => n2013, A2 => n6163, ZN => n4618);
   U15 : AND3_X1 port map( A1 => ADD_WR(1), A2 => n7591, A3 => n6485, ZN => 
                           n4619);
   U16 : AND3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n7591, ZN =>
                           n4620);
   U17 : AND2_X1 port map( A1 => n6163, A2 => n4613, ZN => n4621);
   U18 : AND3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(2), A3 => n6482, ZN =>
                           n4622);
   U19 : AND3_X1 port map( A1 => ADD_WR(0), A2 => n7591, A3 => n6482, ZN => 
                           n4623);
   U20 : AND3_X1 port map( A1 => ADD_WR(2), A2 => n6485, A3 => n6482, ZN => 
                           n4624);
   U21 : AND3_X1 port map( A1 => n7591, A2 => n6485, A3 => n6482, ZN => n4625);
   U22 : AND2_X1 port map( A1 => n2012, A2 => n6163, ZN => n4626);
   U23 : AND3_X1 port map( A1 => n1406, A2 => n4608, A3 => n6236, ZN => n4627);
   U24 : AND3_X1 port map( A1 => n1406, A2 => n1413, A3 => n6236, ZN => n4628);
   U25 : AND3_X1 port map( A1 => n1393, A2 => n4608, A3 => n6236, ZN => n4629);
   U26 : AND2_X1 port map( A1 => n1394, A2 => n4617, ZN => n4630);
   U27 : AND2_X1 port map( A1 => n2019, A2 => n4613, ZN => n4631);
   U28 : AND2_X1 port map( A1 => n1419, A2 => n4608, ZN => n4632);
   U29 : AND2_X1 port map( A1 => n2006, A2 => n4621, ZN => n4633);
   U30 : AND2_X1 port map( A1 => n2006, A2 => n4626, ZN => n4634);
   U31 : AND2_X1 port map( A1 => n4609, A2 => n4619, ZN => n4635);
   U32 : AND2_X1 port map( A1 => n4606, A2 => n4614, ZN => n4636);
   U33 : AND2_X1 port map( A1 => n4606, A2 => n4619, ZN => n4637);
   U34 : AND2_X1 port map( A1 => n4606, A2 => n4620, ZN => n4638);
   U35 : AND2_X1 port map( A1 => n4607, A2 => n4620, ZN => n4639);
   U36 : AND2_X1 port map( A1 => n4607, A2 => n4619, ZN => n4640);
   U37 : AND2_X1 port map( A1 => n6489, A2 => n4623, ZN => n4641);
   U38 : AND2_X1 port map( A1 => n6489, A2 => n4622, ZN => n4642);
   U39 : AND2_X1 port map( A1 => n4623, A2 => n4609, ZN => n4643);
   U40 : AND2_X1 port map( A1 => n4622, A2 => n4609, ZN => n4644);
   U41 : AND2_X1 port map( A1 => n4625, A2 => n4609, ZN => n4645);
   U42 : AND2_X1 port map( A1 => n4624, A2 => n4609, ZN => n4646);
   U43 : AND2_X1 port map( A1 => n4611, A2 => n4609, ZN => n4647);
   U44 : AND2_X1 port map( A1 => n4614, A2 => n4609, ZN => n4648);
   U45 : AND2_X1 port map( A1 => n4620, A2 => n4609, ZN => n4649);
   U46 : AND2_X1 port map( A1 => n4625, A2 => n4607, ZN => n4650);
   U47 : AND2_X1 port map( A1 => n4624, A2 => n4607, ZN => n4651);
   U48 : AND2_X1 port map( A1 => n4622, A2 => n4607, ZN => n4652);
   U49 : AND2_X1 port map( A1 => n4623, A2 => n4607, ZN => n4653);
   U50 : AND2_X1 port map( A1 => n4624, A2 => n4606, ZN => n4654);
   U51 : AND2_X1 port map( A1 => n4622, A2 => n4606, ZN => n4655);
   U52 : AND2_X1 port map( A1 => n4623, A2 => n4606, ZN => n4656);
   U53 : AND2_X1 port map( A1 => ENABLE, A2 => n6464, ZN => n4657);
   U54 : AND2_X1 port map( A1 => n4624, A2 => n6489, ZN => n4658);
   U55 : AND2_X1 port map( A1 => n4621, A2 => n4610, ZN => n4659);
   U56 : AND2_X1 port map( A1 => RD1, A2 => n4657, ZN => n4660);
   U57 : AND2_X1 port map( A1 => n1994, A2 => n6163, ZN => n4661);
   U58 : AND2_X1 port map( A1 => n749, A2 => ADD_WR(4), ZN => n4662);
   U59 : AND2_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), ZN => n4663);
   U60 : INV_X1 port map( A => n2877, ZN => n4664);
   U61 : INV_X1 port map( A => n2876, ZN => n4665);
   U62 : INV_X1 port map( A => n2875, ZN => n4666);
   U63 : INV_X1 port map( A => n2874, ZN => n4667);
   U64 : INV_X1 port map( A => n2873, ZN => n4668);
   U65 : INV_X1 port map( A => n2872, ZN => n4669);
   U66 : INV_X1 port map( A => n2871, ZN => n4670);
   U67 : INV_X1 port map( A => n2870, ZN => n4671);
   U68 : INV_X1 port map( A => n2869, ZN => n4672);
   U69 : INV_X1 port map( A => n2868, ZN => n4673);
   U70 : INV_X1 port map( A => n2867, ZN => n4674);
   U71 : INV_X1 port map( A => n2866, ZN => n4675);
   U72 : INV_X1 port map( A => n2865, ZN => n4676);
   U73 : INV_X1 port map( A => n2864, ZN => n4677);
   U74 : INV_X1 port map( A => n2863, ZN => n4678);
   U75 : INV_X1 port map( A => n2862, ZN => n4679);
   U76 : INV_X1 port map( A => n2861, ZN => n4680);
   U77 : INV_X1 port map( A => n2860, ZN => n4681);
   U78 : INV_X1 port map( A => n2859, ZN => n4682);
   U79 : INV_X1 port map( A => n2858, ZN => n4683);
   U80 : INV_X1 port map( A => n2857, ZN => n4684);
   U81 : INV_X1 port map( A => n2856, ZN => n4685);
   U82 : INV_X1 port map( A => n2855, ZN => n4686);
   U83 : INV_X1 port map( A => n2854, ZN => n4687);
   U84 : INV_X1 port map( A => n2853, ZN => n4688);
   U85 : INV_X1 port map( A => n2852, ZN => n4689);
   U86 : INV_X1 port map( A => n2851, ZN => n4690);
   U87 : INV_X1 port map( A => n2850, ZN => n4691);
   U88 : INV_X1 port map( A => n998, ZN => n4692);
   U89 : INV_X1 port map( A => n982, ZN => n4693);
   U90 : INV_X1 port map( A => n966, ZN => n4694);
   U91 : INV_X1 port map( A => n950, ZN => n4695);
   U92 : INV_X1 port map( A => n4696, ZN => n4697);
   U93 : INV_X1 port map( A => n4698, ZN => n4699);
   U94 : INV_X1 port map( A => n4700, ZN => n4701);
   U95 : INV_X1 port map( A => n4702, ZN => n4703);
   U96 : INV_X1 port map( A => n4704, ZN => n4705);
   U97 : INV_X1 port map( A => n4706, ZN => n4707);
   U98 : INV_X1 port map( A => n4708, ZN => n4709);
   U99 : INV_X1 port map( A => n4710, ZN => n4711);
   U100 : INV_X1 port map( A => n4712, ZN => n4713);
   U101 : INV_X1 port map( A => n4714, ZN => n4715);
   U102 : INV_X1 port map( A => n4716, ZN => n4717);
   U103 : INV_X1 port map( A => n4718, ZN => n4719);
   U104 : INV_X1 port map( A => n4720, ZN => n4721);
   U105 : INV_X1 port map( A => n4722, ZN => n4723);
   U106 : INV_X1 port map( A => n4724, ZN => n4725);
   U107 : INV_X1 port map( A => n4726, ZN => n4727);
   U108 : INV_X1 port map( A => n4728, ZN => n4729);
   U109 : INV_X1 port map( A => n4730, ZN => n4731);
   U110 : INV_X1 port map( A => n4732, ZN => n4733);
   U111 : INV_X1 port map( A => n4734, ZN => n4735);
   U112 : INV_X1 port map( A => n4736, ZN => n4737);
   U113 : INV_X1 port map( A => n4738, ZN => n4739);
   U114 : INV_X1 port map( A => n4740, ZN => n4741);
   U115 : INV_X1 port map( A => n4742, ZN => n4743);
   U116 : INV_X1 port map( A => n4744, ZN => n4745);
   U117 : INV_X1 port map( A => n4746, ZN => n4747);
   U118 : INV_X1 port map( A => n4748, ZN => n4749);
   U119 : INV_X1 port map( A => n4750, ZN => n4751);
   U120 : INV_X1 port map( A => n4752, ZN => n4753);
   U121 : INV_X1 port map( A => n4754, ZN => n4755);
   U122 : INV_X1 port map( A => n4756, ZN => n4757);
   U123 : INV_X1 port map( A => n4758, ZN => n4759);
   U124 : INV_X1 port map( A => n4760, ZN => n4761);
   U125 : INV_X1 port map( A => n4762, ZN => n4763);
   U126 : INV_X1 port map( A => n4764, ZN => n4765);
   U127 : INV_X1 port map( A => n4766, ZN => n4767);
   U128 : INV_X1 port map( A => n4768, ZN => n4769);
   U129 : INV_X1 port map( A => n4770, ZN => n4771);
   U130 : INV_X1 port map( A => n4772, ZN => n4773);
   U131 : INV_X1 port map( A => n4774, ZN => n4775);
   U132 : INV_X1 port map( A => n4776, ZN => n4777);
   U133 : INV_X1 port map( A => n4778, ZN => n4779);
   U134 : INV_X1 port map( A => n4780, ZN => n4781);
   U135 : INV_X1 port map( A => n4782, ZN => n4783);
   U136 : INV_X1 port map( A => n4784, ZN => n4785);
   U137 : INV_X1 port map( A => n4786, ZN => n4787);
   U138 : INV_X1 port map( A => n4788, ZN => n4789);
   U139 : INV_X1 port map( A => n4790, ZN => n4791);
   U140 : INV_X1 port map( A => n4792, ZN => n4793);
   U141 : INV_X1 port map( A => n4794, ZN => n4795);
   U142 : INV_X1 port map( A => n4796, ZN => n4797);
   U143 : INV_X1 port map( A => n4798, ZN => n4799);
   U144 : INV_X1 port map( A => n4800, ZN => n4801);
   U145 : INV_X1 port map( A => n4802, ZN => n4803);
   U146 : INV_X1 port map( A => n4804, ZN => n4805);
   U147 : INV_X1 port map( A => n4806, ZN => n4807);
   U148 : INV_X1 port map( A => n4808, ZN => n4809);
   U149 : INV_X1 port map( A => n4810, ZN => n4811);
   U150 : INV_X1 port map( A => n4812, ZN => n4813);
   U151 : INV_X1 port map( A => n4814, ZN => n4815);
   U152 : BUF_X1 port map( A => n4641, Z => n6007);
   U153 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n6006, ZN => n4844);
   U154 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n6007, ZN => n4826);
   U155 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n6007, ZN => n4824);
   U156 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n6007, ZN => n4822);
   U157 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n6007, ZN => n4820);
   U158 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n6007, ZN => n4818);
   U159 : NAND2_X1 port map( A1 => n5205, A2 => n4816, ZN => n4817);
   U160 : NAND2_X1 port map( A1 => n4817, A2 => n4818, ZN => n4282);
   U161 : INV_X1 port map( A => n6007, ZN => n4816);
   U162 : NAND2_X1 port map( A1 => n5206, A2 => n4836, ZN => n4819);
   U163 : NAND2_X1 port map( A1 => n4819, A2 => n4820, ZN => n4281);
   U164 : NAND2_X1 port map( A1 => n5207, A2 => n4833, ZN => n4821);
   U165 : NAND2_X1 port map( A1 => n4821, A2 => n4822, ZN => n4280);
   U166 : NAND2_X1 port map( A1 => n5208, A2 => n4830, ZN => n4823);
   U167 : NAND2_X1 port map( A1 => n4823, A2 => n4824, ZN => n4279);
   U168 : NAND2_X1 port map( A1 => n5209, A2 => n4827, ZN => n4825);
   U169 : NAND2_X1 port map( A1 => n4825, A2 => n4826, ZN => n4278);
   U170 : BUF_X1 port map( A => n4641, Z => n6006);
   U171 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n6006, ZN => n4853);
   U172 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n6006, ZN => n4841);
   U173 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n6006, ZN => n4838);
   U174 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n6006, ZN => n4835);
   U175 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n6006, ZN => n4832);
   U176 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n6006, ZN => n4829);
   U177 : NAND2_X1 port map( A1 => n5211, A2 => n4827, ZN => n4828);
   U178 : NAND2_X1 port map( A1 => n4828, A2 => n4829, ZN => n4276);
   U179 : INV_X1 port map( A => n6006, ZN => n4827);
   U180 : NAND2_X1 port map( A1 => n5212, A2 => n4830, ZN => n4831);
   U181 : NAND2_X1 port map( A1 => n4831, A2 => n4832, ZN => n4275);
   U182 : INV_X1 port map( A => n6006, ZN => n4830);
   U183 : NAND2_X1 port map( A1 => n5213, A2 => n4833, ZN => n4834);
   U184 : NAND2_X1 port map( A1 => n4834, A2 => n4835, ZN => n4274);
   U185 : INV_X1 port map( A => n6006, ZN => n4833);
   U186 : NAND2_X1 port map( A1 => n5214, A2 => n4836, ZN => n4837);
   U187 : NAND2_X1 port map( A1 => n4837, A2 => n4838, ZN => n4273);
   U188 : INV_X1 port map( A => n6006, ZN => n4836);
   U189 : NAND2_X1 port map( A1 => n5215, A2 => n4839, ZN => n4840);
   U190 : NAND2_X1 port map( A1 => n4840, A2 => n4841, ZN => n4272);
   U191 : INV_X1 port map( A => n6006, ZN => n4839);
   U192 : NAND2_X1 port map( A1 => n5216, A2 => n4842, ZN => n4843);
   U193 : NAND2_X1 port map( A1 => n4843, A2 => n4844, ZN => n4271);
   U194 : INV_X1 port map( A => n6006, ZN => n4842);
   U195 : BUF_X1 port map( A => n4641, Z => n6005);
   U196 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n6005, ZN => n4871);
   U197 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n6006, ZN => n4850);
   U198 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n6006, ZN => n4847);
   U199 : NAND2_X1 port map( A1 => n5217, A2 => n4845, ZN => n4846);
   U200 : NAND2_X1 port map( A1 => n4846, A2 => n4847, ZN => n4270);
   U201 : INV_X1 port map( A => n6006, ZN => n4845);
   U202 : NAND2_X1 port map( A1 => n5218, A2 => n4848, ZN => n4849);
   U203 : NAND2_X1 port map( A1 => n4849, A2 => n4850, ZN => n4269);
   U204 : INV_X1 port map( A => n6006, ZN => n4848);
   U205 : NAND2_X1 port map( A1 => n5219, A2 => n4851, ZN => n4852);
   U206 : NAND2_X1 port map( A1 => n4852, A2 => n4853, ZN => n4268);
   U207 : INV_X1 port map( A => n6006, ZN => n4851);
   U208 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n6005, ZN => n4877);
   U209 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n6005, ZN => n4868);
   U210 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n6005, ZN => n4865);
   U211 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n6005, ZN => n4862);
   U212 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n6006, ZN => n4859);
   U213 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n6006, ZN => n4856);
   U214 : NAND2_X1 port map( A1 => n5220, A2 => n4854, ZN => n4855);
   U215 : NAND2_X1 port map( A1 => n4855, A2 => n4856, ZN => n4267);
   U216 : INV_X1 port map( A => n6006, ZN => n4854);
   U217 : NAND2_X1 port map( A1 => n5221, A2 => n4857, ZN => n4858);
   U218 : NAND2_X1 port map( A1 => n4858, A2 => n4859, ZN => n4266);
   U219 : INV_X1 port map( A => n6006, ZN => n4857);
   U220 : NAND2_X1 port map( A1 => n5222, A2 => n4860, ZN => n4861);
   U221 : NAND2_X1 port map( A1 => n4861, A2 => n4862, ZN => n4265);
   U222 : INV_X1 port map( A => n6005, ZN => n4860);
   U223 : NAND2_X1 port map( A1 => n5223, A2 => n4863, ZN => n4864);
   U224 : NAND2_X1 port map( A1 => n4864, A2 => n4865, ZN => n4264);
   U225 : INV_X1 port map( A => n6005, ZN => n4863);
   U226 : NAND2_X1 port map( A1 => n5224, A2 => n4866, ZN => n4867);
   U227 : NAND2_X1 port map( A1 => n4867, A2 => n4868, ZN => n4263);
   U228 : INV_X1 port map( A => n6005, ZN => n4866);
   U229 : NAND2_X1 port map( A1 => n5225, A2 => n4869, ZN => n4870);
   U230 : NAND2_X1 port map( A1 => n4870, A2 => n4871, ZN => n4262);
   U231 : INV_X1 port map( A => n6005, ZN => n4869);
   U232 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n6005, ZN => n4883);
   U233 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n6005, ZN => n4874);
   U234 : NAND2_X1 port map( A1 => n5226, A2 => n4872, ZN => n4873);
   U235 : NAND2_X1 port map( A1 => n4873, A2 => n4874, ZN => n4261);
   U236 : INV_X1 port map( A => n6005, ZN => n4872);
   U237 : NAND2_X1 port map( A1 => n5227, A2 => n4875, ZN => n4876);
   U238 : NAND2_X1 port map( A1 => n4876, A2 => n4877, ZN => n4260);
   U239 : INV_X1 port map( A => n6005, ZN => n4875);
   U240 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n6005, ZN => n4889);
   U241 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n6005, ZN => n4880);
   U242 : NAND2_X1 port map( A1 => n5228, A2 => n4878, ZN => n4879);
   U243 : NAND2_X1 port map( A1 => n4879, A2 => n4880, ZN => n4259);
   U244 : INV_X1 port map( A => n6005, ZN => n4878);
   U245 : NAND2_X1 port map( A1 => n5229, A2 => n4881, ZN => n4882);
   U246 : NAND2_X1 port map( A1 => n4882, A2 => n4883, ZN => n4258);
   U247 : INV_X1 port map( A => n6005, ZN => n4881);
   U248 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n6005, ZN => n4895);
   U249 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n6005, ZN => n4886);
   U250 : NAND2_X1 port map( A1 => n5230, A2 => n4884, ZN => n4885);
   U251 : NAND2_X1 port map( A1 => n4885, A2 => n4886, ZN => n4257);
   U252 : INV_X1 port map( A => n6005, ZN => n4884);
   U253 : NAND2_X1 port map( A1 => n5231, A2 => n4887, ZN => n4888);
   U254 : NAND2_X1 port map( A1 => n4888, A2 => n4889, ZN => n4256);
   U255 : INV_X1 port map( A => n6005, ZN => n4887);
   U256 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n6005, ZN => n4892);
   U257 : NAND2_X1 port map( A1 => n5232, A2 => n4890, ZN => n4891);
   U258 : NAND2_X1 port map( A1 => n4891, A2 => n4892, ZN => n4255);
   U259 : INV_X1 port map( A => n6005, ZN => n4890);
   U260 : NAND2_X1 port map( A1 => n5170, A2 => n4893, ZN => n4894);
   U261 : NAND2_X1 port map( A1 => n4894, A2 => n4895, ZN => n4254);
   U262 : INV_X1 port map( A => n6005, ZN => n4893);
   U263 : INV_X1 port map( A => n6075, ZN => n6074);
   U264 : INV_X1 port map( A => n6075, ZN => n6073);
   U265 : INV_X1 port map( A => n6093, ZN => n6091);
   U266 : BUF_X1 port map( A => n6465, Z => n6464);
   U267 : BUF_X1 port map( A => n7511, Z => n6180);
   U268 : BUF_X1 port map( A => n7511, Z => n6179);
   U269 : BUF_X1 port map( A => n6908, Z => n6127);
   U270 : BUF_X1 port map( A => n6911, Z => n6138);
   U271 : BUF_X1 port map( A => n6919, Z => n6167);
   U272 : BUF_X1 port map( A => n6908, Z => n6128);
   U273 : BUF_X1 port map( A => n6911, Z => n6139);
   U274 : BUF_X1 port map( A => n6919, Z => n6168);
   U275 : BUF_X1 port map( A => n7525, Z => n6202);
   U276 : BUF_X1 port map( A => n7525, Z => n6203);
   U277 : BUF_X1 port map( A => n4633, Z => n6124);
   U278 : BUF_X1 port map( A => n4634, Z => n6135);
   U279 : BUF_X1 port map( A => n6910, Z => n6130);
   U280 : BUF_X1 port map( A => n6910, Z => n6131);
   U281 : BUF_X1 port map( A => n4633, Z => n6125);
   U282 : BUF_X1 port map( A => n4634, Z => n6136);
   U283 : BUF_X1 port map( A => n7525, Z => n6204);
   U284 : BUF_X1 port map( A => n6910, Z => n6132);
   U285 : BUF_X1 port map( A => n4633, Z => n6126);
   U286 : BUF_X1 port map( A => n4634, Z => n6137);
   U287 : BUF_X1 port map( A => n6908, Z => n6129);
   U288 : BUF_X1 port map( A => n6911, Z => n6140);
   U289 : BUF_X1 port map( A => n6919, Z => n6169);
   U290 : BUF_X1 port map( A => n7511, Z => n6181);
   U291 : INV_X1 port map( A => n4902, ZN => n6288);
   U292 : INV_X1 port map( A => n4902, ZN => n6289);
   U293 : INV_X1 port map( A => n4901, ZN => n6326);
   U294 : INV_X1 port map( A => n4901, ZN => n6325);
   U295 : INV_X1 port map( A => n4900, ZN => n6271);
   U296 : INV_X1 port map( A => n4900, ZN => n6272);
   U297 : INV_X1 port map( A => n4899, ZN => n6309);
   U298 : INV_X1 port map( A => n4899, ZN => n6308);
   U299 : INV_X1 port map( A => n6102, ZN => n6100);
   U300 : INV_X1 port map( A => n6111, ZN => n6109);
   U301 : INV_X1 port map( A => n6102, ZN => n6101);
   U302 : INV_X1 port map( A => n6111, ZN => n6110);
   U303 : INV_X1 port map( A => n6057, ZN => n6056);
   U304 : INV_X1 port map( A => n6057, ZN => n6055);
   U305 : INV_X1 port map( A => n6066, ZN => n6065);
   U306 : INV_X1 port map( A => n6066, ZN => n6064);
   U307 : INV_X1 port map( A => n6084, ZN => n6082);
   U308 : INV_X1 port map( A => n4897, ZN => n6119);
   U309 : INV_X1 port map( A => n4897, ZN => n6120);
   U310 : INV_X1 port map( A => n4898, ZN => n6133);
   U311 : INV_X1 port map( A => n4898, ZN => n6134);
   U312 : INV_X1 port map( A => n4896, ZN => n6182);
   U313 : INV_X1 port map( A => n4896, ZN => n6183);
   U314 : BUF_X1 port map( A => n1458, Z => n6274);
   U315 : BUF_X1 port map( A => n1458, Z => n6273);
   U316 : BUF_X1 port map( A => n845, Z => n6310);
   U317 : BUF_X1 port map( A => n845, Z => n6311);
   U318 : BUF_X1 port map( A => n1453, Z => n6286);
   U319 : BUF_X1 port map( A => n1453, Z => n6285);
   U320 : BUF_X1 port map( A => n840, Z => n6322);
   U321 : BUF_X1 port map( A => n840, Z => n6323);
   U322 : BUF_X1 port map( A => n845, Z => n6312);
   U323 : BUF_X1 port map( A => n1458, Z => n6275);
   U324 : BUF_X1 port map( A => n1453, Z => n6287);
   U325 : BUF_X1 port map( A => n840, Z => n6324);
   U326 : BUF_X1 port map( A => n4906, Z => n6149);
   U327 : BUF_X1 port map( A => n4906, Z => n6150);
   U328 : BUF_X1 port map( A => n4904, Z => n6223);
   U329 : BUF_X1 port map( A => n4904, Z => n6224);
   U330 : BUF_X1 port map( A => n4629, Z => n6208);
   U331 : BUF_X1 port map( A => n4628, Z => n6196);
   U332 : BUF_X1 port map( A => n4628, Z => n6197);
   U333 : BUF_X1 port map( A => n4629, Z => n6209);
   U334 : BUF_X1 port map( A => n4908, Z => n6229);
   U335 : BUF_X1 port map( A => n4908, Z => n6230);
   U336 : BUF_X1 port map( A => n4905, Z => n6146);
   U337 : BUF_X1 port map( A => n4905, Z => n6147);
   U338 : BUF_X1 port map( A => n4903, Z => n6220);
   U339 : BUF_X1 port map( A => n4903, Z => n6221);
   U340 : BUF_X1 port map( A => n7520, Z => n6187);
   U341 : BUF_X1 port map( A => n7520, Z => n6188);
   U342 : BUF_X1 port map( A => n7529, Z => n6214);
   U343 : BUF_X1 port map( A => n7529, Z => n6215);
   U344 : BUF_X1 port map( A => n4907, Z => n6155);
   U345 : BUF_X1 port map( A => n4907, Z => n6156);
   U346 : BUF_X1 port map( A => n4631, Z => n6159);
   U347 : BUF_X1 port map( A => n4631, Z => n6158);
   U348 : BUF_X1 port map( A => n4632, Z => n6217);
   U349 : BUF_X1 port map( A => n4632, Z => n6218);
   U350 : BUF_X1 port map( A => n7519, Z => n6185);
   U351 : BUF_X1 port map( A => n7519, Z => n6184);
   U352 : BUF_X1 port map( A => n6907, Z => n6121);
   U353 : BUF_X1 port map( A => n6907, Z => n6122);
   U354 : BUF_X1 port map( A => n4659, Z => n6164);
   U355 : BUF_X1 port map( A => n6913, Z => n6141);
   U356 : BUF_X1 port map( A => n6913, Z => n6142);
   U357 : BUF_X1 port map( A => n7528, Z => n6211);
   U358 : BUF_X1 port map( A => n7528, Z => n6212);
   U359 : BUF_X1 port map( A => n7524, Z => n6199);
   U360 : BUF_X1 port map( A => n7524, Z => n6200);
   U361 : BUF_X1 port map( A => n4659, Z => n6165);
   U362 : BUF_X1 port map( A => n4627, Z => n6193);
   U363 : BUF_X1 port map( A => n4630, Z => n6205);
   U364 : BUF_X1 port map( A => n4627, Z => n6194);
   U365 : BUF_X1 port map( A => n4630, Z => n6206);
   U366 : BUF_X1 port map( A => n7522, Z => n6190);
   U367 : BUF_X1 port map( A => n4909, Z => n6152);
   U368 : BUF_X1 port map( A => n4909, Z => n6153);
   U369 : BUF_X1 port map( A => n7522, Z => n6191);
   U370 : BUF_X1 port map( A => n6906, Z => n6116);
   U371 : BUF_X1 port map( A => n6906, Z => n6117);
   U372 : BUF_X1 port map( A => n4910, Z => n6226);
   U373 : BUF_X1 port map( A => n4910, Z => n6227);
   U374 : BUF_X1 port map( A => n6922, Z => n6170);
   U375 : BUF_X1 port map( A => n6922, Z => n6171);
   U376 : BUF_X1 port map( A => n6071, Z => n6075);
   U377 : BUF_X1 port map( A => n6089, Z => n6093);
   U378 : BUF_X1 port map( A => n835, Z => n6334);
   U379 : BUF_X1 port map( A => n1448, Z => n6297);
   U380 : BUF_X1 port map( A => n835, Z => n6333);
   U381 : BUF_X1 port map( A => n1448, Z => n6296);
   U382 : BUF_X1 port map( A => n843, Z => n6317);
   U383 : BUF_X1 port map( A => n843, Z => n6316);
   U384 : BUF_X1 port map( A => n1456, Z => n6280);
   U385 : BUF_X1 port map( A => n1456, Z => n6279);
   U386 : BUF_X1 port map( A => n838, Z => n6328);
   U387 : BUF_X1 port map( A => n838, Z => n6327);
   U388 : BUF_X1 port map( A => n1451, Z => n6291);
   U389 : BUF_X1 port map( A => n1462, Z => n6266);
   U390 : BUF_X1 port map( A => n849, Z => n6303);
   U391 : BUF_X1 port map( A => n849, Z => n6302);
   U392 : BUF_X1 port map( A => n1462, Z => n6265);
   U393 : BUF_X1 port map( A => n1451, Z => n6290);
   U394 : BUF_X1 port map( A => n842, Z => n6320);
   U395 : BUF_X1 port map( A => n842, Z => n6319);
   U396 : BUF_X1 port map( A => n1455, Z => n6283);
   U397 : BUF_X1 port map( A => n1455, Z => n6282);
   U398 : BUF_X1 port map( A => n4904, Z => n6225);
   U399 : BUF_X1 port map( A => n4906, Z => n6151);
   U400 : BUF_X1 port map( A => n4629, Z => n6210);
   U401 : BUF_X1 port map( A => n4628, Z => n6198);
   U402 : BUF_X1 port map( A => n1461, Z => n6269);
   U403 : BUF_X1 port map( A => n848, Z => n6306);
   U404 : BUF_X1 port map( A => n848, Z => n6305);
   U405 : BUF_X1 port map( A => n1461, Z => n6268);
   U406 : BUF_X1 port map( A => n837, Z => n6331);
   U407 : BUF_X1 port map( A => n837, Z => n6330);
   U408 : BUF_X1 port map( A => n1450, Z => n6294);
   U409 : BUF_X1 port map( A => n1450, Z => n6293);
   U410 : BUF_X1 port map( A => n834, Z => n6337);
   U411 : BUF_X1 port map( A => n1447, Z => n6300);
   U412 : BUF_X1 port map( A => n834, Z => n6336);
   U413 : BUF_X1 port map( A => n1447, Z => n6299);
   U414 : BUF_X1 port map( A => n844, Z => n6314);
   U415 : BUF_X1 port map( A => n844, Z => n6313);
   U416 : BUF_X1 port map( A => n1457, Z => n6277);
   U417 : BUF_X1 port map( A => n1457, Z => n6276);
   U418 : BUF_X1 port map( A => n4908, Z => n6231);
   U419 : BUF_X1 port map( A => n835, Z => n6335);
   U420 : BUF_X1 port map( A => n1448, Z => n6298);
   U421 : BUF_X1 port map( A => n7520, Z => n6189);
   U422 : BUF_X1 port map( A => n4903, Z => n6222);
   U423 : BUF_X1 port map( A => n4905, Z => n6148);
   U424 : BUF_X1 port map( A => n843, Z => n6318);
   U425 : BUF_X1 port map( A => n1456, Z => n6281);
   U426 : BUF_X1 port map( A => n1462, Z => n6267);
   U427 : BUF_X1 port map( A => n1451, Z => n6292);
   U428 : BUF_X1 port map( A => n838, Z => n6329);
   U429 : BUF_X1 port map( A => n849, Z => n6304);
   U430 : BUF_X1 port map( A => n7529, Z => n6216);
   U431 : BUF_X1 port map( A => n4907, Z => n6157);
   U432 : BUF_X1 port map( A => n6907, Z => n6123);
   U433 : BUF_X1 port map( A => n4632, Z => n6219);
   U434 : BUF_X1 port map( A => n4631, Z => n6160);
   U435 : BUF_X1 port map( A => n842, Z => n6321);
   U436 : BUF_X1 port map( A => n1455, Z => n6284);
   U437 : BUF_X1 port map( A => n6913, Z => n6143);
   U438 : BUF_X1 port map( A => n7519, Z => n6186);
   U439 : BUF_X1 port map( A => n7528, Z => n6213);
   U440 : BUF_X1 port map( A => n7524, Z => n6201);
   U441 : BUF_X1 port map( A => n1461, Z => n6270);
   U442 : BUF_X1 port map( A => n848, Z => n6307);
   U443 : BUF_X1 port map( A => n1450, Z => n6295);
   U444 : BUF_X1 port map( A => n837, Z => n6332);
   U445 : BUF_X1 port map( A => n4627, Z => n6195);
   U446 : BUF_X1 port map( A => n4630, Z => n6207);
   U447 : BUF_X1 port map( A => n4659, Z => n6166);
   U448 : BUF_X1 port map( A => n4909, Z => n6154);
   U449 : BUF_X1 port map( A => n7522, Z => n6192);
   U450 : BUF_X1 port map( A => n834, Z => n6338);
   U451 : BUF_X1 port map( A => n1447, Z => n6301);
   U452 : BUF_X1 port map( A => n6906, Z => n6118);
   U453 : BUF_X1 port map( A => n844, Z => n6315);
   U454 : BUF_X1 port map( A => n1457, Z => n6278);
   U455 : BUF_X1 port map( A => n4910, Z => n6228);
   U456 : BUF_X1 port map( A => n6922, Z => n6172);
   U457 : BUF_X1 port map( A => n6071, Z => n6076);
   U458 : BUF_X1 port map( A => n6071, Z => n6077);
   U459 : BUF_X1 port map( A => n6089, Z => n6094);
   U460 : BUF_X1 port map( A => n6089, Z => n6095);
   U461 : BUF_X1 port map( A => n6072, Z => n6078);
   U462 : BUF_X1 port map( A => n6072, Z => n6079);
   U463 : BUF_X1 port map( A => n6090, Z => n6096);
   U464 : BUF_X1 port map( A => n6090, Z => n6097);
   U465 : BUF_X1 port map( A => n6375, Z => n6465);
   U466 : BUF_X1 port map( A => n6377, Z => n6472);
   U467 : BUF_X1 port map( A => n6377, Z => n6471);
   U468 : BUF_X1 port map( A => n6376, Z => n6470);
   U469 : BUF_X1 port map( A => n6377, Z => n6473);
   U470 : BUF_X1 port map( A => n6378, Z => n6475);
   U471 : BUF_X1 port map( A => n6378, Z => n6474);
   U472 : BUF_X1 port map( A => n6378, Z => n6476);
   U473 : BUF_X1 port map( A => n6375, Z => n6466);
   U474 : BUF_X1 port map( A => n6375, Z => n6467);
   U475 : BUF_X1 port map( A => n6376, Z => n6469);
   U476 : BUF_X1 port map( A => n6376, Z => n6468);
   U477 : BUF_X1 port map( A => n6379, Z => n6477);
   U478 : BUF_X1 port map( A => n6379, Z => n6478);
   U479 : NOR2_X1 port map( A1 => n7898, A2 => n6480, ZN => n1412);
   U480 : NOR2_X1 port map( A1 => n7900, A2 => n6479, ZN => n2012);
   U481 : NOR3_X1 port map( A1 => n7592, A2 => n7593, A3 => n7901, ZN => n2006)
                           ;
   U482 : NOR3_X1 port map( A1 => n7594, A2 => n7595, A3 => n7899, ZN => n1406)
                           ;
   U483 : BUF_X1 port map( A => n6484, Z => n6033);
   U484 : BUF_X1 port map( A => n6484, Z => n6032);
   U485 : BUF_X1 port map( A => n4650, Z => n6014);
   U486 : BUF_X1 port map( A => n4650, Z => n6015);
   U487 : BUF_X1 port map( A => n6916, Z => n6161);
   U488 : BUF_X1 port map( A => n6916, Z => n6162);
   U489 : BUF_X1 port map( A => n7510, Z => n6176);
   U490 : BUF_X1 port map( A => n7510, Z => n6177);
   U491 : NAND2_X1 port map( A1 => n2023, A2 => n2012, ZN => n1462);
   U492 : NAND2_X1 port map( A1 => n2022, A2 => n2013, ZN => n1456);
   U493 : NAND2_X1 port map( A1 => n2023, A2 => n2013, ZN => n1455);
   U494 : NAND2_X1 port map( A1 => n2022, A2 => n1994, ZN => n1457);
   U495 : NAND2_X1 port map( A1 => n2022, A2 => n4613, ZN => n1451);
   U496 : NAND2_X1 port map( A1 => n2023, A2 => n4613, ZN => n1450);
   U497 : NAND2_X1 port map( A1 => n1422, A2 => n1413, ZN => n843);
   U498 : NAND2_X1 port map( A1 => n1423, A2 => n1413, ZN => n842);
   U499 : NAND2_X1 port map( A1 => n1422, A2 => n1394, ZN => n844);
   U500 : NAND2_X1 port map( A1 => n1423, A2 => n1412, ZN => n849);
   U501 : NAND2_X1 port map( A1 => n1422, A2 => n4608, ZN => n838);
   U502 : NAND2_X1 port map( A1 => n1423, A2 => n4608, ZN => n837);
   U503 : NAND2_X1 port map( A1 => n1394, A2 => n1419, ZN => n848);
   U504 : BUF_X1 port map( A => n6916, Z => n6163);
   U505 : NAND2_X1 port map( A1 => n1994, A2 => n2019, ZN => n1461);
   U506 : BUF_X1 port map( A => n4650, Z => n6016);
   U507 : AND2_X1 port map( A1 => n4617, A2 => n4608, ZN => n4896);
   U508 : BUF_X1 port map( A => n6484, Z => n6034);
   U509 : BUF_X1 port map( A => n6232, Z => n6234);
   U510 : BUF_X1 port map( A => n6232, Z => n6235);
   U511 : BUF_X1 port map( A => n6233, Z => n6236);
   U512 : BUF_X1 port map( A => n6053, Z => n6057);
   U513 : BUF_X1 port map( A => n6062, Z => n6066);
   U514 : BUF_X1 port map( A => n6080, Z => n6084);
   U515 : BUF_X1 port map( A => n6098, Z => n6102);
   U516 : BUF_X1 port map( A => n6107, Z => n6111);
   U517 : AND2_X1 port map( A1 => n4612, A2 => n4626, ZN => n4897);
   U518 : AND2_X1 port map( A1 => n4612, A2 => n4661, ZN => n4898);
   U519 : AND2_X1 port map( A1 => n2022, A2 => n2012, ZN => n1453);
   U520 : AND2_X1 port map( A1 => n1422, A2 => n1412, ZN => n840);
   U521 : NAND2_X1 port map( A1 => n1420, A2 => n1394, ZN => n4899);
   U522 : NAND2_X1 port map( A1 => n2020, A2 => n1994, ZN => n4900);
   U523 : NAND2_X1 port map( A1 => n1423, A2 => n1394, ZN => n4901);
   U524 : NAND2_X1 port map( A1 => n2023, A2 => n1994, ZN => n4902);
   U525 : AND2_X1 port map( A1 => n1413, A2 => n1420, ZN => n835);
   U526 : AND2_X1 port map( A1 => n1413, A2 => n1419, ZN => n834);
   U527 : AND2_X1 port map( A1 => n1406, A2 => n1394, ZN => n845);
   U528 : AND2_X1 port map( A1 => n2006, A2 => n1994, ZN => n1458);
   U529 : AND2_X1 port map( A1 => n2013, A2 => n2019, ZN => n1447);
   U530 : AND2_X1 port map( A1 => n2013, A2 => n2020, ZN => n1448);
   U531 : AND2_X1 port map( A1 => n1394, A2 => n1393, ZN => n4903);
   U532 : AND2_X1 port map( A1 => n1412, A2 => n1393, ZN => n4904);
   U533 : AND2_X1 port map( A1 => n1994, A2 => n1993, ZN => n4905);
   U534 : AND2_X1 port map( A1 => n2012, A2 => n1993, ZN => n4906);
   U535 : BUF_X1 port map( A => n6053, Z => n6058);
   U536 : BUF_X1 port map( A => n6053, Z => n6059);
   U537 : BUF_X1 port map( A => n6062, Z => n6067);
   U538 : BUF_X1 port map( A => n6062, Z => n6068);
   U539 : BUF_X1 port map( A => n6080, Z => n6085);
   U540 : BUF_X1 port map( A => n6080, Z => n6086);
   U541 : BUF_X1 port map( A => n6098, Z => n6103);
   U542 : BUF_X1 port map( A => n6098, Z => n6104);
   U543 : BUF_X1 port map( A => n6107, Z => n6112);
   U544 : BUF_X1 port map( A => n6107, Z => n6113);
   U545 : BUF_X1 port map( A => n6054, Z => n6060);
   U546 : BUF_X1 port map( A => n6054, Z => n6061);
   U547 : BUF_X1 port map( A => n6063, Z => n6069);
   U548 : BUF_X1 port map( A => n6063, Z => n6070);
   U549 : BUF_X1 port map( A => n6081, Z => n6087);
   U550 : BUF_X1 port map( A => n6081, Z => n6088);
   U551 : BUF_X1 port map( A => n6099, Z => n6105);
   U552 : BUF_X1 port map( A => n6108, Z => n6114);
   U553 : NAND2_X1 port map( A1 => n2012, A2 => n2019, ZN => n4907);
   U554 : NAND2_X1 port map( A1 => n1412, A2 => n1419, ZN => n4908);
   U555 : NAND2_X1 port map( A1 => n2020, A2 => n2012, ZN => n4909);
   U556 : NAND2_X1 port map( A1 => n1420, A2 => n1412, ZN => n4910);
   U557 : BUF_X1 port map( A => n7510, Z => n6178);
   U558 : BUF_X1 port map( A => n6233, Z => n6237);
   U559 : BUF_X1 port map( A => n6099, Z => n6106);
   U560 : BUF_X1 port map( A => n6108, Z => n6115);
   U561 : BUF_X1 port map( A => n6488, Z => n6071);
   U562 : BUF_X1 port map( A => n6491, Z => n6089);
   U563 : BUF_X1 port map( A => n6380, Z => n6377);
   U564 : BUF_X1 port map( A => n6380, Z => n6378);
   U565 : BUF_X1 port map( A => n6381, Z => n6375);
   U566 : BUF_X1 port map( A => n6381, Z => n6376);
   U567 : BUF_X1 port map( A => n6488, Z => n6072);
   U568 : BUF_X1 port map( A => n6491, Z => n6090);
   U569 : BUF_X1 port map( A => n6380, Z => n6379);
   U570 : NOR3_X1 port map( A1 => ADD_RS1(0), A2 => ADD_RS1(4), A3 => n7592, ZN
                           => n2022);
   U571 : NOR3_X1 port map( A1 => n7593, A2 => ADD_RS1(4), A3 => n7592, ZN => 
                           n2023);
   U572 : NOR3_X1 port map( A1 => ADD_RS2(0), A2 => ADD_RS2(4), A3 => n7594, ZN
                           => n1422);
   U573 : NOR3_X1 port map( A1 => n7595, A2 => ADD_RS2(4), A3 => n7594, ZN => 
                           n1423);
   U574 : NOR2_X1 port map( A1 => n7898, A2 => ADD_RS2(1), ZN => n1394);
   U575 : NOR3_X1 port map( A1 => ADD_RS1(0), A2 => ADD_RS1(3), A3 => n7901, ZN
                           => n1993);
   U576 : NOR3_X1 port map( A1 => ADD_RS2(0), A2 => ADD_RS2(3), A3 => n7899, ZN
                           => n1393);
   U577 : NOR2_X1 port map( A1 => n6480, A2 => ADD_RS2(2), ZN => n1413);
   U578 : NOR2_X1 port map( A1 => n7900, A2 => ADD_RS1(1), ZN => n1994);
   U579 : NOR3_X1 port map( A1 => ADD_RS1(3), A2 => ADD_RS1(4), A3 => n7593, ZN
                           => n2019);
   U580 : NOR3_X1 port map( A1 => ADD_RS2(3), A2 => ADD_RS2(4), A3 => n7595, ZN
                           => n1419);
   U581 : NOR2_X1 port map( A1 => n6479, A2 => ADD_RS1(2), ZN => n2013);
   U582 : NOR3_X1 port map( A1 => ADD_RS1(3), A2 => ADD_RS1(4), A3 => 
                           ADD_RS1(0), ZN => n2020);
   U583 : NOR3_X1 port map( A1 => ADD_RS2(3), A2 => ADD_RS2(4), A3 => 
                           ADD_RS2(0), ZN => n1420);
   U584 : INV_X1 port map( A => n4616, ZN => n6144);
   U585 : INV_X1 port map( A => n4616, ZN => n6145);
   U586 : BUF_X1 port map( A => n4643, Z => n6008);
   U587 : BUF_X1 port map( A => n4643, Z => n6009);
   U588 : BUF_X1 port map( A => n4644, Z => n6011);
   U589 : BUF_X1 port map( A => n4644, Z => n6012);
   U590 : BUF_X1 port map( A => n4651, Z => n6017);
   U591 : BUF_X1 port map( A => n4651, Z => n6018);
   U592 : BUF_X1 port map( A => n4636, Z => n6020);
   U593 : BUF_X1 port map( A => n4636, Z => n6021);
   U594 : BUF_X1 port map( A => n4645, Z => n6023);
   U595 : BUF_X1 port map( A => n4645, Z => n6024);
   U596 : BUF_X1 port map( A => n4646, Z => n6026);
   U597 : BUF_X1 port map( A => n4646, Z => n6027);
   U598 : BUF_X1 port map( A => n4652, Z => n6029);
   U599 : BUF_X1 port map( A => n4652, Z => n6030);
   U600 : BUF_X1 port map( A => n4642, Z => n6035);
   U601 : BUF_X1 port map( A => n4642, Z => n6036);
   U602 : BUF_X1 port map( A => n4653, Z => n6038);
   U603 : BUF_X1 port map( A => n4653, Z => n6039);
   U604 : BUF_X1 port map( A => n4637, Z => n6041);
   U605 : BUF_X1 port map( A => n4637, Z => n6042);
   U606 : BUF_X1 port map( A => n4658, Z => n6044);
   U607 : BUF_X1 port map( A => n4658, Z => n6045);
   U608 : BUF_X1 port map( A => n4638, Z => n6047);
   U609 : BUF_X1 port map( A => n4638, Z => n6048);
   U610 : BUF_X1 port map( A => n4654, Z => n6050);
   U611 : BUF_X1 port map( A => n4654, Z => n6051);
   U612 : BUF_X1 port map( A => n4655, Z => n6241);
   U613 : BUF_X1 port map( A => n4655, Z => n6242);
   U614 : BUF_X1 port map( A => n4656, Z => n6244);
   U615 : BUF_X1 port map( A => n4656, Z => n6245);
   U616 : BUF_X1 port map( A => n4639, Z => n6247);
   U617 : BUF_X1 port map( A => n4639, Z => n6248);
   U618 : BUF_X1 port map( A => n4640, Z => n6250);
   U619 : BUF_X1 port map( A => n4640, Z => n6251);
   U620 : BUF_X1 port map( A => n4647, Z => n6253);
   U621 : BUF_X1 port map( A => n4647, Z => n6254);
   U622 : BUF_X1 port map( A => n4648, Z => n6256);
   U623 : BUF_X1 port map( A => n4648, Z => n6257);
   U624 : BUF_X1 port map( A => n4649, Z => n6259);
   U625 : BUF_X1 port map( A => n4649, Z => n6260);
   U626 : BUF_X1 port map( A => n4635, Z => n6262);
   U627 : BUF_X1 port map( A => n4635, Z => n6263);
   U628 : BUF_X1 port map( A => n7552, Z => n6238);
   U629 : BUF_X1 port map( A => n7552, Z => n6239);
   U630 : BUF_X1 port map( A => n4643, Z => n6010);
   U631 : BUF_X1 port map( A => n4644, Z => n6013);
   U632 : BUF_X1 port map( A => n4651, Z => n6019);
   U633 : BUF_X1 port map( A => n4636, Z => n6022);
   U634 : BUF_X1 port map( A => n4645, Z => n6025);
   U635 : BUF_X1 port map( A => n4646, Z => n6028);
   U636 : BUF_X1 port map( A => n4652, Z => n6031);
   U637 : BUF_X1 port map( A => n4642, Z => n6037);
   U638 : BUF_X1 port map( A => n4653, Z => n6040);
   U639 : BUF_X1 port map( A => n4637, Z => n6043);
   U640 : BUF_X1 port map( A => n4658, Z => n6046);
   U641 : BUF_X1 port map( A => n4638, Z => n6049);
   U642 : BUF_X1 port map( A => n4654, Z => n6052);
   U643 : BUF_X1 port map( A => n4655, Z => n6243);
   U644 : BUF_X1 port map( A => n4656, Z => n6246);
   U645 : BUF_X1 port map( A => n4639, Z => n6249);
   U646 : BUF_X1 port map( A => n4640, Z => n6252);
   U647 : BUF_X1 port map( A => n4647, Z => n6255);
   U648 : BUF_X1 port map( A => n4648, Z => n6258);
   U649 : BUF_X1 port map( A => n4649, Z => n6261);
   U650 : BUF_X1 port map( A => n4635, Z => n6264);
   U651 : BUF_X1 port map( A => n7552, Z => n6240);
   U652 : INV_X1 port map( A => ADD_RS1(2), ZN => n7900);
   U653 : INV_X1 port map( A => ADD_RS2(2), ZN => n7898);
   U654 : BUF_X1 port map( A => n7542, Z => n6232);
   U655 : BUF_X1 port map( A => n7542, Z => n6233);
   U656 : BUF_X1 port map( A => n6493, Z => n6107);
   U657 : BUF_X1 port map( A => n6486, Z => n6053);
   U658 : BUF_X1 port map( A => n6487, Z => n6062);
   U659 : BUF_X1 port map( A => n6490, Z => n6080);
   U660 : BUF_X1 port map( A => n6492, Z => n6098);
   U661 : BUF_X1 port map( A => RST, Z => n6380);
   U662 : BUF_X1 port map( A => n6493, Z => n6108);
   U663 : BUF_X1 port map( A => n6486, Z => n6054);
   U664 : BUF_X1 port map( A => n6487, Z => n6063);
   U665 : BUF_X1 port map( A => n6490, Z => n6081);
   U666 : BUF_X1 port map( A => n6492, Z => n6099);
   U667 : BUF_X1 port map( A => RST, Z => n6381);
   U668 : NOR4_X1 port map( A1 => n7902, A2 => n1400, A3 => n1401, A4 => n1402,
                           ZN => n1399);
   U669 : XNOR2_X1 port map( A => n7590, B => ADD_RS1(3), ZN => n2001);
   U670 : XNOR2_X1 port map( A => n7589, B => ADD_RS1(4), ZN => n2000);
   U671 : XNOR2_X1 port map( A => ADD_RS2(2), B => n7591, ZN => n1402);
   U672 : XNOR2_X1 port map( A => n7589, B => ADD_RS2(4), ZN => n1400);
   U673 : XNOR2_X1 port map( A => n7590, B => ADD_RS2(3), ZN => n1401);
   U674 : XNOR2_X1 port map( A => ADD_RS1(2), B => n7591, ZN => n2002);
   U675 : BUF_X1 port map( A => n4660, Z => n6173);
   U676 : BUF_X1 port map( A => n4660, Z => n6174);
   U677 : AOI21_X1 port map( B1 => n6931, B2 => n6930, A => n6929, ZN => n7542)
                           ;
   U678 : AND2_X1 port map( A1 => n1397, A2 => n1427, ZN => n6931);
   U679 : NOR2_X1 port map( A1 => n1402, A2 => n6928, ZN => n6930);
   U680 : NOR3_X1 port map( A1 => n1401, A2 => n7902, A3 => n1400, ZN => n1427)
                           ;
   U681 : BUF_X1 port map( A => n4660, Z => n6175);
   U682 : NOR4_X1 port map( A1 => n7902, A2 => n2000, A3 => n2001, A4 => n2002,
                           ZN => n1999);
   U683 : NOR3_X1 port map( A1 => n2001, A2 => n7902, A3 => n2000, ZN => n2027)
                           ;
   U684 : INV_X1 port map( A => n1398, ZN => n6928);
   U685 : AOI221_X1 port map( B1 => n6275, B2 => n7655, C1 => n6271, C2 => 
                           n7867, A => n1981, ZN => n1974);
   U686 : AOI221_X1 port map( B1 => n6275, B2 => n7654, C1 => n6271, C2 => 
                           n7866, A => n1964, ZN => n1957);
   U687 : AOI221_X1 port map( B1 => n6275, B2 => n7653, C1 => n6271, C2 => 
                           n7865, A => n1947, ZN => n1940);
   U688 : AOI221_X1 port map( B1 => n6275, B2 => n7652, C1 => n6271, C2 => 
                           n7864, A => n1930, ZN => n1923);
   U689 : AOI221_X1 port map( B1 => n6275, B2 => n7651, C1 => n6271, C2 => 
                           n7863, A => n1913, ZN => n1906);
   U690 : AOI221_X1 port map( B1 => n6275, B2 => n7650, C1 => n6271, C2 => 
                           n7862, A => n1896, ZN => n1889);
   U691 : AOI221_X1 port map( B1 => n6275, B2 => n7649, C1 => n6271, C2 => 
                           n7861, A => n1879, ZN => n1872);
   U692 : AOI221_X1 port map( B1 => n6274, B2 => n7648, C1 => n6271, C2 => 
                           n7860, A => n1862, ZN => n1855);
   U693 : AOI221_X1 port map( B1 => n6274, B2 => n7647, C1 => n6271, C2 => 
                           n7859, A => n1845, ZN => n1838);
   U694 : AOI221_X1 port map( B1 => n6274, B2 => n7646, C1 => n6271, C2 => 
                           n7858, A => n1828, ZN => n1821);
   U695 : AOI221_X1 port map( B1 => n6274, B2 => n7645, C1 => n6271, C2 => 
                           n7857, A => n1811, ZN => n1804);
   U696 : AOI221_X1 port map( B1 => n6274, B2 => n7644, C1 => n6271, C2 => 
                           n7856, A => n1794, ZN => n1787);
   U697 : AOI221_X1 port map( B1 => n6274, B2 => n7643, C1 => n6272, C2 => 
                           n7855, A => n1777, ZN => n1770);
   U698 : AOI221_X1 port map( B1 => n6274, B2 => n7642, C1 => n6272, C2 => 
                           n7854, A => n1760, ZN => n1753);
   U699 : AOI221_X1 port map( B1 => n6274, B2 => n7641, C1 => n6272, C2 => 
                           n7853, A => n1743, ZN => n1736);
   U700 : AOI221_X1 port map( B1 => n6274, B2 => n7640, C1 => n6272, C2 => 
                           n7852, A => n1726, ZN => n1719);
   U701 : AOI221_X1 port map( B1 => n6274, B2 => n7639, C1 => n6272, C2 => 
                           n7851, A => n1709, ZN => n1702);
   U702 : AOI221_X1 port map( B1 => n6274, B2 => n7638, C1 => n6272, C2 => 
                           n7850, A => n1692, ZN => n1685);
   U703 : AOI221_X1 port map( B1 => n6274, B2 => n7637, C1 => n6272, C2 => 
                           n7849, A => n1675, ZN => n1668);
   U704 : AOI221_X1 port map( B1 => n6273, B2 => n7636, C1 => n6272, C2 => 
                           n7848, A => n1658, ZN => n1651);
   U705 : AOI221_X1 port map( B1 => n6273, B2 => n7635, C1 => n6272, C2 => 
                           n7847, A => n1641, ZN => n1634);
   U706 : AOI221_X1 port map( B1 => n6273, B2 => n7634, C1 => n6272, C2 => 
                           n7846, A => n1624, ZN => n1617);
   U707 : AOI221_X1 port map( B1 => n6273, B2 => n7633, C1 => n6272, C2 => 
                           n7845, A => n1607, ZN => n1600);
   U708 : AOI221_X1 port map( B1 => n6273, B2 => n7632, C1 => n6272, C2 => 
                           n7844, A => n1590, ZN => n1583);
   U709 : AOI221_X1 port map( B1 => n6273, B2 => n7631, C1 => n6271, C2 => 
                           n7843, A => n1573, ZN => n1566);
   U710 : AOI221_X1 port map( B1 => n6273, B2 => n7630, C1 => n6272, C2 => 
                           n7842, A => n1556, ZN => n1549);
   U711 : AOI221_X1 port map( B1 => n6273, B2 => n7629, C1 => n6271, C2 => 
                           n7841, A => n1539, ZN => n1532);
   U712 : AOI221_X1 port map( B1 => n6273, B2 => n7628, C1 => n6272, C2 => 
                           n7840, A => n1522, ZN => n1515);
   U713 : AOI221_X1 port map( B1 => n6273, B2 => n7627, C1 => n6271, C2 => 
                           n7839, A => n1505, ZN => n1498);
   U714 : AOI221_X1 port map( B1 => n6273, B2 => n7626, C1 => n6272, C2 => 
                           n7838, A => n1488, ZN => n1481);
   U715 : AOI221_X1 port map( B1 => n6273, B2 => n7587, C1 => n6271, C2 => 
                           n5103, A => n1460, ZN => n1437);
   U716 : AOI221_X1 port map( B1 => n6310, B2 => n7588, C1 => n6309, C2 => 
                           n5104, A => n847, ZN => n824);
   U717 : AOI221_X1 port map( B1 => n6310, B2 => n7655, C1 => n6308, C2 => 
                           n7867, A => n878, ZN => n871);
   U718 : AOI221_X1 port map( B1 => n6310, B2 => n7654, C1 => n6309, C2 => 
                           n7866, A => n895, ZN => n888);
   U719 : AOI221_X1 port map( B1 => n6310, B2 => n7653, C1 => n6308, C2 => 
                           n7865, A => n912, ZN => n905);
   U720 : AOI221_X1 port map( B1 => n6310, B2 => n7652, C1 => n6309, C2 => 
                           n7864, A => n929, ZN => n922);
   U721 : AOI221_X1 port map( B1 => n6310, B2 => n7651, C1 => n6308, C2 => 
                           n7863, A => n948, ZN => n941);
   U722 : AOI221_X1 port map( B1 => n6310, B2 => n7650, C1 => n6309, C2 => 
                           n7862, A => n969, ZN => n961);
   U723 : AOI221_X1 port map( B1 => n6310, B2 => n7649, C1 => n6309, C2 => 
                           n7861, A => n991, ZN => n981);
   U724 : AOI221_X1 port map( B1 => n6310, B2 => n7648, C1 => n6309, C2 => 
                           n7860, A => n1009, ZN => n1002);
   U725 : AOI221_X1 port map( B1 => n6310, B2 => n7647, C1 => n6309, C2 => 
                           n7859, A => n1026, ZN => n1019);
   U726 : AOI221_X1 port map( B1 => n6310, B2 => n7646, C1 => n6309, C2 => 
                           n7858, A => n1043, ZN => n1036);
   U727 : AOI221_X1 port map( B1 => n6310, B2 => n7645, C1 => n6309, C2 => 
                           n7857, A => n1060, ZN => n1053);
   U728 : AOI221_X1 port map( B1 => n6311, B2 => n7644, C1 => n6309, C2 => 
                           n7856, A => n1077, ZN => n1070);
   U729 : AOI221_X1 port map( B1 => n6311, B2 => n7643, C1 => n6309, C2 => 
                           n7855, A => n1094, ZN => n1087);
   U730 : AOI221_X1 port map( B1 => n6311, B2 => n7642, C1 => n6309, C2 => 
                           n7854, A => n1111, ZN => n1104);
   U731 : AOI221_X1 port map( B1 => n6311, B2 => n7641, C1 => n6309, C2 => 
                           n7853, A => n1128, ZN => n1121);
   U732 : AOI221_X1 port map( B1 => n6311, B2 => n7640, C1 => n6309, C2 => 
                           n7852, A => n1145, ZN => n1138);
   U733 : AOI221_X1 port map( B1 => n6311, B2 => n7639, C1 => n6309, C2 => 
                           n7851, A => n1162, ZN => n1155);
   U734 : AOI221_X1 port map( B1 => n6311, B2 => n7638, C1 => n6309, C2 => 
                           n7850, A => n1179, ZN => n1172);
   U735 : AOI221_X1 port map( B1 => n6311, B2 => n7637, C1 => n6308, C2 => 
                           n7849, A => n1196, ZN => n1189);
   U736 : AOI221_X1 port map( B1 => n6311, B2 => n7636, C1 => n6308, C2 => 
                           n7848, A => n1213, ZN => n1206);
   U737 : AOI221_X1 port map( B1 => n6311, B2 => n7635, C1 => n6308, C2 => 
                           n7847, A => n1230, ZN => n1223);
   U738 : AOI221_X1 port map( B1 => n6311, B2 => n7634, C1 => n6308, C2 => 
                           n7846, A => n1247, ZN => n1240);
   U739 : AOI221_X1 port map( B1 => n6311, B2 => n7633, C1 => n6308, C2 => 
                           n7845, A => n1264, ZN => n1257);
   U740 : AOI221_X1 port map( B1 => n6312, B2 => n7632, C1 => n6308, C2 => 
                           n7844, A => n1281, ZN => n1274);
   U741 : AOI221_X1 port map( B1 => n6312, B2 => n7631, C1 => n6308, C2 => 
                           n7843, A => n1298, ZN => n1291);
   U742 : AOI221_X1 port map( B1 => n6312, B2 => n7630, C1 => n6308, C2 => 
                           n7842, A => n1315, ZN => n1308);
   U743 : AOI221_X1 port map( B1 => n6312, B2 => n7629, C1 => n6308, C2 => 
                           n7841, A => n1332, ZN => n1325);
   U744 : AOI221_X1 port map( B1 => n6312, B2 => n7628, C1 => n6308, C2 => 
                           n7840, A => n1349, ZN => n1342);
   U745 : AOI221_X1 port map( B1 => n6312, B2 => n7627, C1 => n6308, C2 => 
                           n7839, A => n1366, ZN => n1359);
   U746 : AOI221_X1 port map( B1 => n6312, B2 => n7626, C1 => n6308, C2 => 
                           n7838, A => n1383, ZN => n1376);
   U747 : AOI221_X1 port map( B1 => n6288, B2 => n7897, C1 => n6287, C2 => 
                           n7625, A => n1980, ZN => n1975);
   U748 : AOI221_X1 port map( B1 => n6288, B2 => n7896, C1 => n6287, C2 => 
                           n7624, A => n1963, ZN => n1958);
   U749 : AOI221_X1 port map( B1 => n6288, B2 => n7895, C1 => n6287, C2 => 
                           n7623, A => n1946, ZN => n1941);
   U750 : AOI221_X1 port map( B1 => n6288, B2 => n7894, C1 => n6287, C2 => 
                           n7622, A => n1929, ZN => n1924);
   U751 : AOI221_X1 port map( B1 => n6288, B2 => n7893, C1 => n6287, C2 => 
                           n7621, A => n1912, ZN => n1907);
   U752 : AOI221_X1 port map( B1 => n6288, B2 => n7892, C1 => n6287, C2 => 
                           n7620, A => n1895, ZN => n1890);
   U753 : AOI221_X1 port map( B1 => n6288, B2 => n7891, C1 => n6287, C2 => 
                           n7619, A => n1878, ZN => n1873);
   U754 : AOI221_X1 port map( B1 => n6288, B2 => n7890, C1 => n6286, C2 => 
                           n7618, A => n1861, ZN => n1856);
   U755 : AOI221_X1 port map( B1 => n6288, B2 => n7889, C1 => n6286, C2 => 
                           n7617, A => n1844, ZN => n1839);
   U756 : AOI221_X1 port map( B1 => n6288, B2 => n7888, C1 => n6286, C2 => 
                           n7616, A => n1827, ZN => n1822);
   U757 : AOI221_X1 port map( B1 => n6288, B2 => n7887, C1 => n6286, C2 => 
                           n7615, A => n1810, ZN => n1805);
   U758 : AOI221_X1 port map( B1 => n6288, B2 => n7886, C1 => n6286, C2 => 
                           n7614, A => n1793, ZN => n1788);
   U759 : AOI221_X1 port map( B1 => n6289, B2 => n7885, C1 => n6286, C2 => 
                           n7613, A => n1776, ZN => n1771);
   U760 : AOI221_X1 port map( B1 => n6289, B2 => n7884, C1 => n6286, C2 => 
                           n7612, A => n1759, ZN => n1754);
   U761 : AOI221_X1 port map( B1 => n6289, B2 => n7883, C1 => n6286, C2 => 
                           n7611, A => n1742, ZN => n1737);
   U762 : AOI221_X1 port map( B1 => n6289, B2 => n7882, C1 => n6286, C2 => 
                           n7610, A => n1725, ZN => n1720);
   U763 : AOI221_X1 port map( B1 => n6289, B2 => n7881, C1 => n6286, C2 => 
                           n7609, A => n1708, ZN => n1703);
   U764 : AOI221_X1 port map( B1 => n6289, B2 => n7880, C1 => n6286, C2 => 
                           n7608, A => n1691, ZN => n1686);
   U765 : AOI221_X1 port map( B1 => n6289, B2 => n7879, C1 => n6286, C2 => 
                           n7607, A => n1674, ZN => n1669);
   U766 : AOI221_X1 port map( B1 => n6289, B2 => n7878, C1 => n6285, C2 => 
                           n7606, A => n1657, ZN => n1652);
   U767 : AOI221_X1 port map( B1 => n6289, B2 => n7877, C1 => n6285, C2 => 
                           n7605, A => n1640, ZN => n1635);
   U768 : AOI221_X1 port map( B1 => n6289, B2 => n7876, C1 => n6285, C2 => 
                           n7604, A => n1623, ZN => n1618);
   U769 : AOI221_X1 port map( B1 => n6289, B2 => n7875, C1 => n6285, C2 => 
                           n7603, A => n1606, ZN => n1601);
   U770 : AOI221_X1 port map( B1 => n6289, B2 => n7874, C1 => n6285, C2 => 
                           n7602, A => n1589, ZN => n1584);
   U771 : AOI221_X1 port map( B1 => n6288, B2 => n7873, C1 => n6285, C2 => 
                           n7601, A => n1572, ZN => n1567);
   U772 : AOI221_X1 port map( B1 => n6289, B2 => n7872, C1 => n6285, C2 => 
                           n7600, A => n1555, ZN => n1550);
   U773 : AOI221_X1 port map( B1 => n6288, B2 => n7871, C1 => n6285, C2 => 
                           n7599, A => n1538, ZN => n1533);
   U774 : AOI221_X1 port map( B1 => n6289, B2 => n7870, C1 => n6285, C2 => 
                           n7598, A => n1521, ZN => n1516);
   U775 : AOI221_X1 port map( B1 => n6288, B2 => n7869, C1 => n6285, C2 => 
                           n7597, A => n1504, ZN => n1499);
   U776 : AOI221_X1 port map( B1 => n6289, B2 => n7868, C1 => n6285, C2 => 
                           n7596, A => n1487, ZN => n1482);
   U777 : AOI221_X1 port map( B1 => n6288, B2 => n5101, C1 => n6285, C2 => 
                           n7585, A => n1454, ZN => n1438);
   U778 : AOI221_X1 port map( B1 => n6326, B2 => n5102, C1 => n6322, C2 => 
                           n7586, A => n841, ZN => n825);
   U779 : AOI221_X1 port map( B1 => n6325, B2 => n7897, C1 => n6322, C2 => 
                           n7625, A => n877, ZN => n872);
   U780 : AOI221_X1 port map( B1 => n6326, B2 => n7896, C1 => n6322, C2 => 
                           n7624, A => n894, ZN => n889);
   U781 : AOI221_X1 port map( B1 => n6325, B2 => n7895, C1 => n6322, C2 => 
                           n7623, A => n911, ZN => n906);
   U782 : AOI221_X1 port map( B1 => n6326, B2 => n7894, C1 => n6322, C2 => 
                           n7622, A => n928, ZN => n923);
   U783 : AOI221_X1 port map( B1 => n6325, B2 => n7893, C1 => n6322, C2 => 
                           n7621, A => n947, ZN => n942);
   U784 : AOI221_X1 port map( B1 => n6326, B2 => n7892, C1 => n6322, C2 => 
                           n7620, A => n968, ZN => n962);
   U785 : AOI221_X1 port map( B1 => n6326, B2 => n7891, C1 => n6322, C2 => 
                           n7619, A => n990, ZN => n983);
   U786 : AOI221_X1 port map( B1 => n6326, B2 => n7890, C1 => n6322, C2 => 
                           n7618, A => n1008, ZN => n1003);
   U787 : AOI221_X1 port map( B1 => n6326, B2 => n7889, C1 => n6322, C2 => 
                           n7617, A => n1025, ZN => n1020);
   U788 : AOI221_X1 port map( B1 => n6326, B2 => n7888, C1 => n6322, C2 => 
                           n7616, A => n1042, ZN => n1037);
   U789 : AOI221_X1 port map( B1 => n6326, B2 => n7887, C1 => n6322, C2 => 
                           n7615, A => n1059, ZN => n1054);
   U790 : AOI221_X1 port map( B1 => n6326, B2 => n7886, C1 => n6323, C2 => 
                           n7614, A => n1076, ZN => n1071);
   U791 : AOI221_X1 port map( B1 => n6326, B2 => n7885, C1 => n6323, C2 => 
                           n7613, A => n1093, ZN => n1088);
   U792 : AOI221_X1 port map( B1 => n6326, B2 => n7884, C1 => n6323, C2 => 
                           n7612, A => n1110, ZN => n1105);
   U793 : AOI221_X1 port map( B1 => n6326, B2 => n7883, C1 => n6323, C2 => 
                           n7611, A => n1127, ZN => n1122);
   U794 : AOI221_X1 port map( B1 => n6326, B2 => n7882, C1 => n6323, C2 => 
                           n7610, A => n1144, ZN => n1139);
   U795 : AOI221_X1 port map( B1 => n6326, B2 => n7881, C1 => n6323, C2 => 
                           n7609, A => n1161, ZN => n1156);
   U796 : AOI221_X1 port map( B1 => n6326, B2 => n7880, C1 => n6323, C2 => 
                           n7608, A => n1178, ZN => n1173);
   U797 : AOI221_X1 port map( B1 => n6325, B2 => n7879, C1 => n6323, C2 => 
                           n7607, A => n1195, ZN => n1190);
   U798 : AOI221_X1 port map( B1 => n6325, B2 => n7878, C1 => n6323, C2 => 
                           n7606, A => n1212, ZN => n1207);
   U799 : AOI221_X1 port map( B1 => n6325, B2 => n7877, C1 => n6323, C2 => 
                           n7605, A => n1229, ZN => n1224);
   U800 : AOI221_X1 port map( B1 => n6325, B2 => n7876, C1 => n6323, C2 => 
                           n7604, A => n1246, ZN => n1241);
   U801 : AOI221_X1 port map( B1 => n6325, B2 => n7875, C1 => n6323, C2 => 
                           n7603, A => n1263, ZN => n1258);
   U802 : AOI221_X1 port map( B1 => n6325, B2 => n7874, C1 => n6324, C2 => 
                           n7602, A => n1280, ZN => n1275);
   U803 : AOI221_X1 port map( B1 => n6325, B2 => n7873, C1 => n6324, C2 => 
                           n7601, A => n1297, ZN => n1292);
   U804 : AOI221_X1 port map( B1 => n6325, B2 => n7872, C1 => n6324, C2 => 
                           n7600, A => n1314, ZN => n1309);
   U805 : AOI221_X1 port map( B1 => n6325, B2 => n7871, C1 => n6324, C2 => 
                           n7599, A => n1331, ZN => n1326);
   U806 : AOI221_X1 port map( B1 => n6325, B2 => n7870, C1 => n6324, C2 => 
                           n7598, A => n1348, ZN => n1343);
   U807 : AOI221_X1 port map( B1 => n6325, B2 => n7869, C1 => n6324, C2 => 
                           n7597, A => n1365, ZN => n1360);
   U808 : AOI221_X1 port map( B1 => n6325, B2 => n7868, C1 => n6324, C2 => 
                           n7596, A => n1382, ZN => n1377);
   U809 : XNOR2_X1 port map( A => ADD_RS2(1), B => ADD_WR(1), ZN => n1398);
   U810 : XNOR2_X1 port map( A => ADD_RS1(0), B => ADD_WR(0), ZN => n1997);
   U811 : XNOR2_X1 port map( A => ADD_RS1(1), B => ADD_WR(1), ZN => n1998);
   U812 : INV_X1 port map( A => WR, ZN => n7902);
   U813 : XNOR2_X1 port map( A => ADD_RS2(0), B => ADD_WR(0), ZN => n1397);
   U814 : AOI221_X1 port map( B1 => n6299, B2 => n4061, C1 => n6296, C2 => 
                           n4093, A => n1449, ZN => n1439);
   U815 : AOI221_X1 port map( B1 => n6336, B2 => n4030, C1 => n6333, C2 => 
                           n4062, A => n836, ZN => n826);
   U816 : INV_X1 port map( A => DATAIN(31), ZN => n6374);
   U817 : INV_X1 port map( A => DATAIN(4), ZN => n6347);
   U818 : INV_X1 port map( A => DATAIN(5), ZN => n6348);
   U819 : INV_X1 port map( A => DATAIN(6), ZN => n6349);
   U820 : INV_X1 port map( A => DATAIN(7), ZN => n6350);
   U821 : INV_X1 port map( A => DATAIN(8), ZN => n6351);
   U822 : INV_X1 port map( A => DATAIN(9), ZN => n6352);
   U823 : INV_X1 port map( A => DATAIN(10), ZN => n6353);
   U824 : INV_X1 port map( A => DATAIN(11), ZN => n6354);
   U825 : INV_X1 port map( A => DATAIN(12), ZN => n6355);
   U826 : INV_X1 port map( A => DATAIN(13), ZN => n6356);
   U827 : INV_X1 port map( A => DATAIN(14), ZN => n6357);
   U828 : INV_X1 port map( A => DATAIN(15), ZN => n6358);
   U829 : INV_X1 port map( A => DATAIN(16), ZN => n6359);
   U830 : INV_X1 port map( A => DATAIN(17), ZN => n6360);
   U831 : INV_X1 port map( A => DATAIN(18), ZN => n6361);
   U832 : INV_X1 port map( A => DATAIN(19), ZN => n6362);
   U833 : INV_X1 port map( A => DATAIN(20), ZN => n6363);
   U834 : INV_X1 port map( A => DATAIN(21), ZN => n6364);
   U835 : INV_X1 port map( A => DATAIN(22), ZN => n6365);
   U836 : INV_X1 port map( A => DATAIN(23), ZN => n6366);
   U837 : INV_X1 port map( A => DATAIN(24), ZN => n6367);
   U838 : INV_X1 port map( A => DATAIN(25), ZN => n6368);
   U839 : INV_X1 port map( A => DATAIN(26), ZN => n6369);
   U840 : INV_X1 port map( A => DATAIN(27), ZN => n6370);
   U841 : INV_X1 port map( A => DATAIN(28), ZN => n6371);
   U842 : INV_X1 port map( A => DATAIN(29), ZN => n6372);
   U843 : INV_X1 port map( A => DATAIN(30), ZN => n6373);
   U844 : INV_X1 port map( A => n2285, ZN => n7867);
   U845 : INV_X1 port map( A => n2436, ZN => n7625);
   U846 : INV_X1 port map( A => n2286, ZN => n7866);
   U847 : INV_X1 port map( A => n2432, ZN => n7624);
   U848 : INV_X1 port map( A => n2287, ZN => n7865);
   U849 : INV_X1 port map( A => n2428, ZN => n7623);
   U850 : INV_X1 port map( A => n2288, ZN => n7864);
   U851 : INV_X1 port map( A => n2424, ZN => n7622);
   U852 : INV_X1 port map( A => n2289, ZN => n7863);
   U853 : INV_X1 port map( A => n2420, ZN => n7621);
   U854 : INV_X1 port map( A => n2290, ZN => n7862);
   U855 : INV_X1 port map( A => n2416, ZN => n7620);
   U856 : INV_X1 port map( A => n2291, ZN => n7861);
   U857 : INV_X1 port map( A => n2412, ZN => n7619);
   U858 : INV_X1 port map( A => n2292, ZN => n7860);
   U859 : INV_X1 port map( A => n2408, ZN => n7618);
   U860 : INV_X1 port map( A => n2293, ZN => n7859);
   U861 : INV_X1 port map( A => n2404, ZN => n7617);
   U862 : INV_X1 port map( A => n2294, ZN => n7858);
   U863 : INV_X1 port map( A => n2400, ZN => n7616);
   U864 : INV_X1 port map( A => n2295, ZN => n7857);
   U865 : INV_X1 port map( A => n2396, ZN => n7615);
   U866 : INV_X1 port map( A => n2296, ZN => n7856);
   U867 : INV_X1 port map( A => n2392, ZN => n7614);
   U868 : INV_X1 port map( A => n2297, ZN => n7855);
   U869 : INV_X1 port map( A => n2388, ZN => n7613);
   U870 : INV_X1 port map( A => n2298, ZN => n7854);
   U871 : INV_X1 port map( A => n2384, ZN => n7612);
   U872 : INV_X1 port map( A => n2299, ZN => n7853);
   U873 : INV_X1 port map( A => n2380, ZN => n7611);
   U874 : INV_X1 port map( A => n2300, ZN => n7852);
   U875 : INV_X1 port map( A => n2376, ZN => n7610);
   U876 : INV_X1 port map( A => n2301, ZN => n7851);
   U877 : INV_X1 port map( A => n2372, ZN => n7609);
   U878 : INV_X1 port map( A => n2302, ZN => n7850);
   U879 : INV_X1 port map( A => n2368, ZN => n7608);
   U880 : INV_X1 port map( A => n2303, ZN => n7849);
   U881 : INV_X1 port map( A => n2364, ZN => n7607);
   U882 : INV_X1 port map( A => n2304, ZN => n7848);
   U883 : INV_X1 port map( A => n2360, ZN => n7606);
   U884 : INV_X1 port map( A => n2305, ZN => n7847);
   U885 : INV_X1 port map( A => n2356, ZN => n7605);
   U886 : INV_X1 port map( A => n2306, ZN => n7846);
   U887 : INV_X1 port map( A => n2352, ZN => n7604);
   U888 : INV_X1 port map( A => n2307, ZN => n7845);
   U889 : INV_X1 port map( A => n2348, ZN => n7603);
   U890 : INV_X1 port map( A => n2308, ZN => n7844);
   U891 : INV_X1 port map( A => n2344, ZN => n7602);
   U892 : INV_X1 port map( A => n2309, ZN => n7843);
   U893 : INV_X1 port map( A => n2340, ZN => n7601);
   U894 : INV_X1 port map( A => n2310, ZN => n7842);
   U895 : INV_X1 port map( A => n2336, ZN => n7600);
   U896 : INV_X1 port map( A => n2311, ZN => n7841);
   U897 : INV_X1 port map( A => n2332, ZN => n7599);
   U898 : INV_X1 port map( A => n2312, ZN => n7840);
   U899 : INV_X1 port map( A => n2328, ZN => n7598);
   U900 : INV_X1 port map( A => n2313, ZN => n7839);
   U901 : INV_X1 port map( A => n2324, ZN => n7597);
   U902 : INV_X1 port map( A => n2314, ZN => n7838);
   U903 : INV_X1 port map( A => n2320, ZN => n7596);
   U904 : INV_X1 port map( A => n2029, ZN => n7655);
   U905 : INV_X1 port map( A => n3743, ZN => n7897);
   U906 : INV_X1 port map( A => n2030, ZN => n7654);
   U907 : INV_X1 port map( A => n3744, ZN => n7896);
   U908 : INV_X1 port map( A => n2031, ZN => n7653);
   U909 : INV_X1 port map( A => n3745, ZN => n7895);
   U910 : INV_X1 port map( A => n2032, ZN => n7652);
   U911 : INV_X1 port map( A => n3746, ZN => n7894);
   U912 : INV_X1 port map( A => n2033, ZN => n7651);
   U913 : INV_X1 port map( A => n3747, ZN => n7893);
   U914 : INV_X1 port map( A => n2034, ZN => n7650);
   U915 : INV_X1 port map( A => n3748, ZN => n7892);
   U916 : INV_X1 port map( A => n2035, ZN => n7649);
   U917 : INV_X1 port map( A => n3749, ZN => n7891);
   U918 : INV_X1 port map( A => n2036, ZN => n7648);
   U919 : INV_X1 port map( A => n3750, ZN => n7890);
   U920 : INV_X1 port map( A => n2037, ZN => n7647);
   U921 : INV_X1 port map( A => n3751, ZN => n7889);
   U922 : INV_X1 port map( A => n2038, ZN => n7646);
   U923 : INV_X1 port map( A => n3752, ZN => n7888);
   U924 : INV_X1 port map( A => n2039, ZN => n7645);
   U925 : INV_X1 port map( A => n3753, ZN => n7887);
   U926 : INV_X1 port map( A => n2040, ZN => n7644);
   U927 : INV_X1 port map( A => n3754, ZN => n7886);
   U928 : INV_X1 port map( A => n2041, ZN => n7643);
   U929 : INV_X1 port map( A => n3755, ZN => n7885);
   U930 : INV_X1 port map( A => n2042, ZN => n7642);
   U931 : INV_X1 port map( A => n3756, ZN => n7884);
   U932 : INV_X1 port map( A => n2043, ZN => n7641);
   U933 : INV_X1 port map( A => n3757, ZN => n7883);
   U934 : INV_X1 port map( A => n2044, ZN => n7640);
   U935 : INV_X1 port map( A => n3758, ZN => n7882);
   U936 : INV_X1 port map( A => n2045, ZN => n7639);
   U937 : INV_X1 port map( A => n3759, ZN => n7881);
   U938 : INV_X1 port map( A => n2046, ZN => n7638);
   U939 : INV_X1 port map( A => n3760, ZN => n7880);
   U940 : INV_X1 port map( A => n2047, ZN => n7637);
   U941 : INV_X1 port map( A => n3761, ZN => n7879);
   U942 : INV_X1 port map( A => n2048, ZN => n7636);
   U943 : INV_X1 port map( A => n3762, ZN => n7878);
   U944 : INV_X1 port map( A => n2049, ZN => n7635);
   U945 : INV_X1 port map( A => n3763, ZN => n7877);
   U946 : INV_X1 port map( A => n2050, ZN => n7634);
   U947 : INV_X1 port map( A => n3764, ZN => n7876);
   U948 : INV_X1 port map( A => n2051, ZN => n7633);
   U949 : INV_X1 port map( A => n3765, ZN => n7875);
   U950 : INV_X1 port map( A => n2052, ZN => n7632);
   U951 : INV_X1 port map( A => n3766, ZN => n7874);
   U952 : INV_X1 port map( A => n2053, ZN => n7631);
   U953 : INV_X1 port map( A => n3767, ZN => n7873);
   U954 : INV_X1 port map( A => n2054, ZN => n7630);
   U955 : INV_X1 port map( A => n3768, ZN => n7872);
   U956 : INV_X1 port map( A => n2055, ZN => n7629);
   U957 : INV_X1 port map( A => n3769, ZN => n7871);
   U958 : INV_X1 port map( A => n2056, ZN => n7628);
   U959 : INV_X1 port map( A => n3770, ZN => n7870);
   U960 : INV_X1 port map( A => n2057, ZN => n7627);
   U961 : INV_X1 port map( A => n3771, ZN => n7869);
   U962 : INV_X1 port map( A => n2058, ZN => n7626);
   U963 : INV_X1 port map( A => n3772, ZN => n7868);
   U964 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n749);
   U965 : INV_X1 port map( A => n2220, ZN => n4911);
   U966 : INV_X1 port map( A => n2060, ZN => n4912);
   U967 : INV_X1 port map( A => n2282, ZN => n4913);
   U968 : INV_X1 port map( A => n2281, ZN => n4914);
   U969 : INV_X1 port map( A => n2280, ZN => n4915);
   U970 : INV_X1 port map( A => n2279, ZN => n4916);
   U971 : INV_X1 port map( A => n2278, ZN => n4917);
   U972 : INV_X1 port map( A => n2277, ZN => n4918);
   U973 : INV_X1 port map( A => n2276, ZN => n4919);
   U974 : INV_X1 port map( A => n2275, ZN => n4920);
   U975 : INV_X1 port map( A => n2274, ZN => n4921);
   U976 : INV_X1 port map( A => n2273, ZN => n4922);
   U977 : INV_X1 port map( A => n2272, ZN => n4923);
   U978 : INV_X1 port map( A => n2271, ZN => n4924);
   U979 : INV_X1 port map( A => n2270, ZN => n4925);
   U980 : INV_X1 port map( A => n2269, ZN => n4926);
   U981 : INV_X1 port map( A => n2268, ZN => n4927);
   U982 : INV_X1 port map( A => n2267, ZN => n4928);
   U983 : INV_X1 port map( A => n2266, ZN => n4929);
   U984 : INV_X1 port map( A => n2265, ZN => n4930);
   U985 : INV_X1 port map( A => n2264, ZN => n4931);
   U986 : INV_X1 port map( A => n2263, ZN => n4932);
   U987 : INV_X1 port map( A => n2262, ZN => n4933);
   U988 : INV_X1 port map( A => n2261, ZN => n4934);
   U989 : INV_X1 port map( A => n2260, ZN => n4935);
   U990 : INV_X1 port map( A => n2259, ZN => n4936);
   U991 : INV_X1 port map( A => n2258, ZN => n4937);
   U992 : INV_X1 port map( A => n2257, ZN => n4938);
   U993 : INV_X1 port map( A => n2256, ZN => n4939);
   U994 : INV_X1 port map( A => n2255, ZN => n4940);
   U995 : INV_X1 port map( A => n2254, ZN => n4941);
   U996 : INV_X1 port map( A => n2253, ZN => n4942);
   U997 : INV_X1 port map( A => n2717, ZN => n4943);
   U998 : INV_X1 port map( A => n2716, ZN => n4944);
   U999 : INV_X1 port map( A => n2715, ZN => n4945);
   U1000 : INV_X1 port map( A => n2714, ZN => n4946);
   U1001 : INV_X1 port map( A => n2713, ZN => n4947);
   U1002 : INV_X1 port map( A => n2712, ZN => n4948);
   U1003 : INV_X1 port map( A => n2711, ZN => n4949);
   U1004 : INV_X1 port map( A => n2710, ZN => n4950);
   U1005 : INV_X1 port map( A => n2709, ZN => n4951);
   U1006 : INV_X1 port map( A => n2708, ZN => n4952);
   U1007 : INV_X1 port map( A => n2707, ZN => n4953);
   U1008 : INV_X1 port map( A => n2706, ZN => n4954);
   U1009 : INV_X1 port map( A => n2705, ZN => n4955);
   U1010 : INV_X1 port map( A => n2704, ZN => n4956);
   U1011 : INV_X1 port map( A => n2703, ZN => n4957);
   U1012 : INV_X1 port map( A => n2702, ZN => n4958);
   U1013 : INV_X1 port map( A => n2701, ZN => n4959);
   U1014 : INV_X1 port map( A => n2700, ZN => n4960);
   U1015 : INV_X1 port map( A => n2699, ZN => n4961);
   U1016 : INV_X1 port map( A => n2698, ZN => n4962);
   U1017 : INV_X1 port map( A => n2697, ZN => n4963);
   U1018 : INV_X1 port map( A => n2696, ZN => n4964);
   U1019 : INV_X1 port map( A => n2695, ZN => n4965);
   U1020 : INV_X1 port map( A => n2694, ZN => n4966);
   U1021 : INV_X1 port map( A => n2693, ZN => n4967);
   U1022 : INV_X1 port map( A => n2692, ZN => n4968);
   U1023 : INV_X1 port map( A => n2691, ZN => n4969);
   U1024 : INV_X1 port map( A => n2690, ZN => n4970);
   U1025 : INV_X1 port map( A => n2942, ZN => n4971);
   U1026 : INV_X1 port map( A => n2718, ZN => n4972);
   U1027 : INV_X1 port map( A => n2250, ZN => n4973);
   U1028 : INV_X1 port map( A => n2249, ZN => n4974);
   U1029 : INV_X1 port map( A => n2248, ZN => n4975);
   U1030 : INV_X1 port map( A => n2247, ZN => n4976);
   U1031 : INV_X1 port map( A => n2246, ZN => n4977);
   U1032 : INV_X1 port map( A => n2245, ZN => n4978);
   U1033 : INV_X1 port map( A => n2244, ZN => n4979);
   U1034 : INV_X1 port map( A => n2243, ZN => n4980);
   U1035 : INV_X1 port map( A => n2242, ZN => n4981);
   U1036 : INV_X1 port map( A => n2241, ZN => n4982);
   U1037 : INV_X1 port map( A => n2240, ZN => n4983);
   U1038 : INV_X1 port map( A => n2239, ZN => n4984);
   U1039 : INV_X1 port map( A => n2238, ZN => n4985);
   U1040 : INV_X1 port map( A => n2237, ZN => n4986);
   U1041 : INV_X1 port map( A => n2236, ZN => n4987);
   U1042 : INV_X1 port map( A => n2235, ZN => n4988);
   U1043 : INV_X1 port map( A => n2234, ZN => n4989);
   U1044 : INV_X1 port map( A => n2233, ZN => n4990);
   U1045 : INV_X1 port map( A => n2232, ZN => n4991);
   U1046 : INV_X1 port map( A => n2231, ZN => n4992);
   U1047 : INV_X1 port map( A => n2230, ZN => n4993);
   U1048 : INV_X1 port map( A => n2229, ZN => n4994);
   U1049 : INV_X1 port map( A => n2228, ZN => n4995);
   U1050 : INV_X1 port map( A => n2227, ZN => n4996);
   U1051 : INV_X1 port map( A => n2226, ZN => n4997);
   U1052 : INV_X1 port map( A => n2225, ZN => n4998);
   U1053 : INV_X1 port map( A => n2224, ZN => n4999);
   U1054 : INV_X1 port map( A => n2223, ZN => n5000);
   U1055 : INV_X1 port map( A => n2222, ZN => n5001);
   U1056 : INV_X1 port map( A => n2221, ZN => n5002);
   U1057 : INV_X1 port map( A => n2219, ZN => n5003);
   U1058 : INV_X1 port map( A => n2218, ZN => n5004);
   U1059 : INV_X1 port map( A => n2217, ZN => n5005);
   U1060 : INV_X1 port map( A => n2216, ZN => n5006);
   U1061 : INV_X1 port map( A => n2215, ZN => n5007);
   U1062 : INV_X1 port map( A => n2214, ZN => n5008);
   U1063 : INV_X1 port map( A => n2213, ZN => n5009);
   U1064 : INV_X1 port map( A => n2212, ZN => n5010);
   U1065 : INV_X1 port map( A => n2211, ZN => n5011);
   U1066 : INV_X1 port map( A => n2210, ZN => n5012);
   U1067 : INV_X1 port map( A => n2209, ZN => n5013);
   U1068 : INV_X1 port map( A => n2208, ZN => n5014);
   U1069 : INV_X1 port map( A => n2207, ZN => n5015);
   U1070 : INV_X1 port map( A => n2206, ZN => n5016);
   U1071 : INV_X1 port map( A => n2205, ZN => n5017);
   U1072 : INV_X1 port map( A => n2204, ZN => n5018);
   U1073 : INV_X1 port map( A => n2203, ZN => n5019);
   U1074 : INV_X1 port map( A => n2202, ZN => n5020);
   U1075 : INV_X1 port map( A => n2201, ZN => n5021);
   U1076 : INV_X1 port map( A => n2200, ZN => n5022);
   U1077 : INV_X1 port map( A => n2199, ZN => n5023);
   U1078 : INV_X1 port map( A => n2198, ZN => n5024);
   U1079 : INV_X1 port map( A => n2197, ZN => n5025);
   U1080 : INV_X1 port map( A => n2196, ZN => n5026);
   U1081 : INV_X1 port map( A => n2195, ZN => n5027);
   U1082 : INV_X1 port map( A => n2194, ZN => n5028);
   U1083 : INV_X1 port map( A => n2193, ZN => n5029);
   U1084 : INV_X1 port map( A => n2192, ZN => n5030);
   U1085 : INV_X1 port map( A => n2191, ZN => n5031);
   U1086 : INV_X1 port map( A => n2190, ZN => n5032);
   U1087 : INV_X1 port map( A => n2189, ZN => n5033);
   U1088 : INV_X1 port map( A => n987, ZN => n5034);
   U1089 : INV_X1 port map( A => n971, ZN => n5035);
   U1090 : INV_X1 port map( A => n955, ZN => n5036);
   U1091 : INV_X1 port map( A => n2123, ZN => n5037);
   U1092 : INV_X1 port map( A => n2122, ZN => n5038);
   U1093 : INV_X1 port map( A => n2121, ZN => n5039);
   U1094 : INV_X1 port map( A => n2120, ZN => n5040);
   U1095 : INV_X1 port map( A => n2119, ZN => n5041);
   U1096 : INV_X1 port map( A => n2118, ZN => n5042);
   U1097 : INV_X1 port map( A => n2117, ZN => n5043);
   U1098 : INV_X1 port map( A => n2116, ZN => n5044);
   U1099 : INV_X1 port map( A => n2115, ZN => n5045);
   U1100 : INV_X1 port map( A => n2114, ZN => n5046);
   U1101 : INV_X1 port map( A => n2113, ZN => n5047);
   U1102 : INV_X1 port map( A => n2112, ZN => n5048);
   U1103 : INV_X1 port map( A => n2111, ZN => n5049);
   U1104 : INV_X1 port map( A => n2110, ZN => n5050);
   U1105 : INV_X1 port map( A => n2109, ZN => n5051);
   U1106 : INV_X1 port map( A => n2108, ZN => n5052);
   U1107 : INV_X1 port map( A => n2107, ZN => n5053);
   U1108 : INV_X1 port map( A => n2106, ZN => n5054);
   U1109 : INV_X1 port map( A => n2105, ZN => n5055);
   U1110 : INV_X1 port map( A => n2104, ZN => n5056);
   U1111 : INV_X1 port map( A => n2103, ZN => n5057);
   U1112 : INV_X1 port map( A => n2102, ZN => n5058);
   U1113 : INV_X1 port map( A => n2101, ZN => n5059);
   U1114 : INV_X1 port map( A => n2100, ZN => n5060);
   U1115 : INV_X1 port map( A => n2099, ZN => n5061);
   U1116 : INV_X1 port map( A => n2098, ZN => n5062);
   U1117 : INV_X1 port map( A => n2097, ZN => n5063);
   U1118 : INV_X1 port map( A => n2096, ZN => n5064);
   U1119 : INV_X1 port map( A => n2095, ZN => n5065);
   U1120 : INV_X1 port map( A => n2094, ZN => n5066);
   U1121 : INV_X1 port map( A => n2093, ZN => n5067);
   U1122 : INV_X1 port map( A => n2092, ZN => n5068);
   U1123 : INV_X1 port map( A => n3677, ZN => n5069);
   U1124 : INV_X1 port map( A => n3676, ZN => n5070);
   U1125 : INV_X1 port map( A => n3675, ZN => n5071);
   U1126 : INV_X1 port map( A => n3674, ZN => n5072);
   U1127 : INV_X1 port map( A => n3673, ZN => n5073);
   U1128 : INV_X1 port map( A => n3672, ZN => n5074);
   U1129 : INV_X1 port map( A => n3671, ZN => n5075);
   U1130 : INV_X1 port map( A => n3670, ZN => n5076);
   U1131 : INV_X1 port map( A => n3669, ZN => n5077);
   U1132 : INV_X1 port map( A => n3668, ZN => n5078);
   U1133 : INV_X1 port map( A => n3667, ZN => n5079);
   U1134 : INV_X1 port map( A => n3666, ZN => n5080);
   U1135 : INV_X1 port map( A => n3665, ZN => n5081);
   U1136 : INV_X1 port map( A => n3664, ZN => n5082);
   U1137 : INV_X1 port map( A => n3663, ZN => n5083);
   U1138 : INV_X1 port map( A => n3662, ZN => n5084);
   U1139 : INV_X1 port map( A => n3661, ZN => n5085);
   U1140 : INV_X1 port map( A => n3660, ZN => n5086);
   U1141 : INV_X1 port map( A => n3659, ZN => n5087);
   U1142 : INV_X1 port map( A => n3658, ZN => n5088);
   U1143 : INV_X1 port map( A => n3657, ZN => n5089);
   U1144 : INV_X1 port map( A => n3656, ZN => n5090);
   U1145 : INV_X1 port map( A => n3655, ZN => n5091);
   U1146 : INV_X1 port map( A => n3654, ZN => n5092);
   U1147 : INV_X1 port map( A => n3653, ZN => n5093);
   U1148 : INV_X1 port map( A => n3652, ZN => n5094);
   U1149 : INV_X1 port map( A => n3651, ZN => n5095);
   U1150 : INV_X1 port map( A => n3650, ZN => n5096);
   U1151 : INV_X1 port map( A => n3649, ZN => n5097);
   U1152 : INV_X1 port map( A => n3648, ZN => n5098);
   U1153 : INV_X1 port map( A => n3647, ZN => n5099);
   U1154 : INV_X1 port map( A => n3646, ZN => n5100);
   U1155 : INV_X1 port map( A => n3773, ZN => n5101);
   U1156 : INV_X1 port map( A => n3742, ZN => n5102);
   U1157 : INV_X1 port map( A => n2315, ZN => n5103);
   U1158 : INV_X1 port map( A => n2284, ZN => n5104);
   U1159 : OAI22_X1 port map( A1 => n4029, A2 => n6305, B1 => n2317, B2 => 
                           n6302, ZN => n1425);
   U1160 : OAI22_X1 port map( A1 => n4029, A2 => n6270, B1 => n2317, B2 => 
                           n6267, ZN => n1460);
   U1161 : OAI22_X1 port map( A1 => n4028, A2 => n6305, B1 => n2321, B2 => 
                           n6302, ZN => n1383);
   U1162 : OAI22_X1 port map( A1 => n4028, A2 => n6270, B1 => n2321, B2 => 
                           n6267, ZN => n1488);
   U1163 : OAI22_X1 port map( A1 => n4027, A2 => n6305, B1 => n2325, B2 => 
                           n6302, ZN => n1366);
   U1164 : OAI22_X1 port map( A1 => n4027, A2 => n6270, B1 => n2325, B2 => 
                           n6267, ZN => n1505);
   U1165 : OAI22_X1 port map( A1 => n4026, A2 => n6305, B1 => n2329, B2 => 
                           n6302, ZN => n1349);
   U1166 : OAI22_X1 port map( A1 => n4026, A2 => n6270, B1 => n2329, B2 => 
                           n6267, ZN => n1522);
   U1167 : OAI22_X1 port map( A1 => n4025, A2 => n6305, B1 => n2333, B2 => 
                           n6302, ZN => n1332);
   U1168 : OAI22_X1 port map( A1 => n4025, A2 => n6270, B1 => n2333, B2 => 
                           n6267, ZN => n1539);
   U1169 : OAI22_X1 port map( A1 => n4024, A2 => n6305, B1 => n2337, B2 => 
                           n6302, ZN => n1315);
   U1170 : OAI22_X1 port map( A1 => n4024, A2 => n6270, B1 => n2337, B2 => 
                           n6267, ZN => n1556);
   U1171 : OAI22_X1 port map( A1 => n4023, A2 => n6305, B1 => n2341, B2 => 
                           n6302, ZN => n1298);
   U1172 : OAI22_X1 port map( A1 => n4023, A2 => n6270, B1 => n2341, B2 => 
                           n6267, ZN => n1573);
   U1173 : OAI22_X1 port map( A1 => n4022, A2 => n6305, B1 => n2345, B2 => 
                           n6302, ZN => n1281);
   U1174 : OAI22_X1 port map( A1 => n4022, A2 => n6270, B1 => n2345, B2 => 
                           n6267, ZN => n1590);
   U1175 : OAI22_X1 port map( A1 => n4021, A2 => n6305, B1 => n2349, B2 => 
                           n6302, ZN => n1264);
   U1176 : OAI22_X1 port map( A1 => n4021, A2 => n6269, B1 => n2349, B2 => 
                           n6266, ZN => n1607);
   U1177 : OAI22_X1 port map( A1 => n4020, A2 => n6305, B1 => n2353, B2 => 
                           n6302, ZN => n1247);
   U1178 : OAI22_X1 port map( A1 => n4020, A2 => n6269, B1 => n2353, B2 => 
                           n6266, ZN => n1624);
   U1179 : OAI22_X1 port map( A1 => n4019, A2 => n6305, B1 => n2357, B2 => 
                           n6302, ZN => n1230);
   U1180 : OAI22_X1 port map( A1 => n4019, A2 => n6269, B1 => n2357, B2 => 
                           n6266, ZN => n1641);
   U1181 : OAI22_X1 port map( A1 => n4018, A2 => n6305, B1 => n2361, B2 => 
                           n6302, ZN => n1213);
   U1182 : OAI22_X1 port map( A1 => n4018, A2 => n6269, B1 => n2361, B2 => 
                           n6266, ZN => n1658);
   U1183 : OAI22_X1 port map( A1 => n4017, A2 => n6306, B1 => n2365, B2 => 
                           n6303, ZN => n1196);
   U1184 : OAI22_X1 port map( A1 => n4017, A2 => n6269, B1 => n2365, B2 => 
                           n6266, ZN => n1675);
   U1185 : OAI22_X1 port map( A1 => n4016, A2 => n6306, B1 => n2369, B2 => 
                           n6303, ZN => n1179);
   U1186 : OAI22_X1 port map( A1 => n4016, A2 => n6269, B1 => n2369, B2 => 
                           n6266, ZN => n1692);
   U1187 : OAI22_X1 port map( A1 => n4015, A2 => n6306, B1 => n2373, B2 => 
                           n6303, ZN => n1162);
   U1188 : OAI22_X1 port map( A1 => n4015, A2 => n6269, B1 => n2373, B2 => 
                           n6266, ZN => n1709);
   U1189 : OAI22_X1 port map( A1 => n4014, A2 => n6306, B1 => n2377, B2 => 
                           n6303, ZN => n1145);
   U1190 : OAI22_X1 port map( A1 => n4014, A2 => n6269, B1 => n2377, B2 => 
                           n6266, ZN => n1726);
   U1191 : OAI22_X1 port map( A1 => n4013, A2 => n6306, B1 => n2381, B2 => 
                           n6303, ZN => n1128);
   U1192 : OAI22_X1 port map( A1 => n4013, A2 => n6269, B1 => n2381, B2 => 
                           n6266, ZN => n1743);
   U1193 : OAI22_X1 port map( A1 => n4012, A2 => n6306, B1 => n2385, B2 => 
                           n6303, ZN => n1111);
   U1194 : OAI22_X1 port map( A1 => n4012, A2 => n6269, B1 => n2385, B2 => 
                           n6266, ZN => n1760);
   U1195 : OAI22_X1 port map( A1 => n4011, A2 => n6306, B1 => n2389, B2 => 
                           n6303, ZN => n1094);
   U1196 : OAI22_X1 port map( A1 => n4011, A2 => n6269, B1 => n2389, B2 => 
                           n6266, ZN => n1777);
   U1197 : OAI22_X1 port map( A1 => n4010, A2 => n6306, B1 => n2393, B2 => 
                           n6303, ZN => n1077);
   U1198 : OAI22_X1 port map( A1 => n4010, A2 => n6269, B1 => n2393, B2 => 
                           n6266, ZN => n1794);
   U1199 : OAI22_X1 port map( A1 => n4009, A2 => n6306, B1 => n2397, B2 => 
                           n6303, ZN => n1060);
   U1200 : OAI22_X1 port map( A1 => n4009, A2 => n6268, B1 => n2397, B2 => 
                           n6265, ZN => n1811);
   U1201 : OAI22_X1 port map( A1 => n4008, A2 => n6306, B1 => n2401, B2 => 
                           n6303, ZN => n1043);
   U1202 : OAI22_X1 port map( A1 => n4008, A2 => n6268, B1 => n2401, B2 => 
                           n6265, ZN => n1828);
   U1203 : OAI22_X1 port map( A1 => n4007, A2 => n6306, B1 => n2405, B2 => 
                           n6303, ZN => n1026);
   U1204 : OAI22_X1 port map( A1 => n4007, A2 => n6268, B1 => n2405, B2 => 
                           n6265, ZN => n1845);
   U1205 : OAI22_X1 port map( A1 => n4006, A2 => n6306, B1 => n2409, B2 => 
                           n6303, ZN => n1009);
   U1206 : OAI22_X1 port map( A1 => n4006, A2 => n6268, B1 => n2409, B2 => 
                           n6265, ZN => n1862);
   U1207 : OAI22_X1 port map( A1 => n4005, A2 => n6307, B1 => n2413, B2 => 
                           n6304, ZN => n991);
   U1208 : OAI22_X1 port map( A1 => n4005, A2 => n6268, B1 => n2413, B2 => 
                           n6265, ZN => n1879);
   U1209 : OAI22_X1 port map( A1 => n4004, A2 => n6307, B1 => n2417, B2 => 
                           n6304, ZN => n969);
   U1210 : OAI22_X1 port map( A1 => n4004, A2 => n6268, B1 => n2417, B2 => 
                           n6265, ZN => n1896);
   U1211 : OAI22_X1 port map( A1 => n4003, A2 => n6307, B1 => n2421, B2 => 
                           n6304, ZN => n948);
   U1212 : OAI22_X1 port map( A1 => n4003, A2 => n6268, B1 => n2421, B2 => 
                           n6265, ZN => n1913);
   U1213 : OAI22_X1 port map( A1 => n4002, A2 => n6307, B1 => n2425, B2 => 
                           n6304, ZN => n929);
   U1214 : OAI22_X1 port map( A1 => n4002, A2 => n6268, B1 => n2425, B2 => 
                           n6265, ZN => n1930);
   U1215 : OAI22_X1 port map( A1 => n4001, A2 => n6307, B1 => n2429, B2 => 
                           n6304, ZN => n912);
   U1216 : OAI22_X1 port map( A1 => n4001, A2 => n6268, B1 => n2429, B2 => 
                           n6265, ZN => n1947);
   U1217 : OAI22_X1 port map( A1 => n4000, A2 => n6307, B1 => n2433, B2 => 
                           n6304, ZN => n895);
   U1218 : OAI22_X1 port map( A1 => n4000, A2 => n6268, B1 => n2433, B2 => 
                           n6265, ZN => n1964);
   U1219 : OAI22_X1 port map( A1 => n3999, A2 => n6307, B1 => n2437, B2 => 
                           n6304, ZN => n878);
   U1220 : OAI22_X1 port map( A1 => n3999, A2 => n6268, B1 => n2437, B2 => 
                           n6265, ZN => n1981);
   U1221 : OAI22_X1 port map( A1 => n3998, A2 => n6307, B1 => n2441, B2 => 
                           n6304, ZN => n847);
   U1222 : OAI22_X1 port map( A1 => n3998, A2 => n6268, B1 => n2441, B2 => 
                           n6265, ZN => n2025);
   U1223 : OAI22_X1 port map( A1 => n3901, A2 => n6330, B1 => n3933, B2 => 
                           n6327, ZN => n1421);
   U1224 : OAI22_X1 port map( A1 => n3901, A2 => n6295, B1 => n3933, B2 => 
                           n6292, ZN => n1449);
   U1225 : OAI22_X1 port map( A1 => n3900, A2 => n6330, B1 => n3932, B2 => 
                           n6327, ZN => n1381);
   U1226 : OAI22_X1 port map( A1 => n3900, A2 => n6295, B1 => n3932, B2 => 
                           n6292, ZN => n1486);
   U1227 : OAI22_X1 port map( A1 => n3899, A2 => n6330, B1 => n3931, B2 => 
                           n6327, ZN => n1364);
   U1228 : OAI22_X1 port map( A1 => n3899, A2 => n6295, B1 => n3931, B2 => 
                           n6292, ZN => n1503);
   U1229 : OAI22_X1 port map( A1 => n3898, A2 => n6330, B1 => n3930, B2 => 
                           n6327, ZN => n1347);
   U1230 : OAI22_X1 port map( A1 => n3898, A2 => n6295, B1 => n3930, B2 => 
                           n6292, ZN => n1520);
   U1231 : OAI22_X1 port map( A1 => n3897, A2 => n6330, B1 => n3929, B2 => 
                           n6327, ZN => n1330);
   U1232 : OAI22_X1 port map( A1 => n3897, A2 => n6295, B1 => n3929, B2 => 
                           n6292, ZN => n1537);
   U1233 : OAI22_X1 port map( A1 => n3896, A2 => n6330, B1 => n3928, B2 => 
                           n6327, ZN => n1313);
   U1234 : OAI22_X1 port map( A1 => n3896, A2 => n6295, B1 => n3928, B2 => 
                           n6292, ZN => n1554);
   U1235 : OAI22_X1 port map( A1 => n3895, A2 => n6330, B1 => n3927, B2 => 
                           n6327, ZN => n1296);
   U1236 : OAI22_X1 port map( A1 => n3895, A2 => n6295, B1 => n3927, B2 => 
                           n6292, ZN => n1571);
   U1237 : OAI22_X1 port map( A1 => n3894, A2 => n6330, B1 => n3926, B2 => 
                           n6327, ZN => n1279);
   U1238 : OAI22_X1 port map( A1 => n3894, A2 => n6295, B1 => n3926, B2 => 
                           n6292, ZN => n1588);
   U1239 : OAI22_X1 port map( A1 => n3893, A2 => n6330, B1 => n3925, B2 => 
                           n6327, ZN => n1262);
   U1240 : OAI22_X1 port map( A1 => n3893, A2 => n6294, B1 => n3925, B2 => 
                           n6291, ZN => n1605);
   U1241 : OAI22_X1 port map( A1 => n3892, A2 => n6330, B1 => n3924, B2 => 
                           n6327, ZN => n1245);
   U1242 : OAI22_X1 port map( A1 => n3892, A2 => n6294, B1 => n3924, B2 => 
                           n6291, ZN => n1622);
   U1243 : OAI22_X1 port map( A1 => n3891, A2 => n6330, B1 => n3923, B2 => 
                           n6327, ZN => n1228);
   U1244 : OAI22_X1 port map( A1 => n3891, A2 => n6294, B1 => n3923, B2 => 
                           n6291, ZN => n1639);
   U1245 : OAI22_X1 port map( A1 => n3890, A2 => n6330, B1 => n3922, B2 => 
                           n6327, ZN => n1211);
   U1246 : OAI22_X1 port map( A1 => n3890, A2 => n6294, B1 => n3922, B2 => 
                           n6291, ZN => n1656);
   U1247 : OAI22_X1 port map( A1 => n3889, A2 => n6331, B1 => n3921, B2 => 
                           n6328, ZN => n1194);
   U1248 : OAI22_X1 port map( A1 => n3889, A2 => n6294, B1 => n3921, B2 => 
                           n6291, ZN => n1673);
   U1249 : OAI22_X1 port map( A1 => n3888, A2 => n6331, B1 => n3920, B2 => 
                           n6328, ZN => n1177);
   U1250 : OAI22_X1 port map( A1 => n3888, A2 => n6294, B1 => n3920, B2 => 
                           n6291, ZN => n1690);
   U1251 : OAI22_X1 port map( A1 => n3887, A2 => n6331, B1 => n3919, B2 => 
                           n6328, ZN => n1160);
   U1252 : OAI22_X1 port map( A1 => n3887, A2 => n6294, B1 => n3919, B2 => 
                           n6291, ZN => n1707);
   U1253 : OAI22_X1 port map( A1 => n3886, A2 => n6331, B1 => n3918, B2 => 
                           n6328, ZN => n1143);
   U1254 : OAI22_X1 port map( A1 => n3886, A2 => n6294, B1 => n3918, B2 => 
                           n6291, ZN => n1724);
   U1255 : OAI22_X1 port map( A1 => n3885, A2 => n6331, B1 => n3917, B2 => 
                           n6328, ZN => n1126);
   U1256 : OAI22_X1 port map( A1 => n3885, A2 => n6294, B1 => n3917, B2 => 
                           n6291, ZN => n1741);
   U1257 : OAI22_X1 port map( A1 => n3884, A2 => n6331, B1 => n3916, B2 => 
                           n6328, ZN => n1109);
   U1258 : OAI22_X1 port map( A1 => n3884, A2 => n6294, B1 => n3916, B2 => 
                           n6291, ZN => n1758);
   U1259 : OAI22_X1 port map( A1 => n3883, A2 => n6331, B1 => n3915, B2 => 
                           n6328, ZN => n1092);
   U1260 : OAI22_X1 port map( A1 => n3883, A2 => n6294, B1 => n3915, B2 => 
                           n6291, ZN => n1775);
   U1261 : OAI22_X1 port map( A1 => n3882, A2 => n6331, B1 => n3914, B2 => 
                           n6328, ZN => n1075);
   U1262 : OAI22_X1 port map( A1 => n3882, A2 => n6294, B1 => n3914, B2 => 
                           n6291, ZN => n1792);
   U1263 : OAI22_X1 port map( A1 => n3881, A2 => n6331, B1 => n3913, B2 => 
                           n6328, ZN => n1058);
   U1264 : OAI22_X1 port map( A1 => n3881, A2 => n6293, B1 => n3913, B2 => 
                           n6290, ZN => n1809);
   U1265 : OAI22_X1 port map( A1 => n3880, A2 => n6331, B1 => n3912, B2 => 
                           n6328, ZN => n1041);
   U1266 : OAI22_X1 port map( A1 => n3880, A2 => n6293, B1 => n3912, B2 => 
                           n6290, ZN => n1826);
   U1267 : OAI22_X1 port map( A1 => n3879, A2 => n6331, B1 => n3911, B2 => 
                           n6328, ZN => n1024);
   U1268 : OAI22_X1 port map( A1 => n3879, A2 => n6293, B1 => n3911, B2 => 
                           n6290, ZN => n1843);
   U1269 : OAI22_X1 port map( A1 => n3878, A2 => n6331, B1 => n3910, B2 => 
                           n6328, ZN => n1007);
   U1270 : OAI22_X1 port map( A1 => n3878, A2 => n6293, B1 => n3910, B2 => 
                           n6290, ZN => n1860);
   U1271 : OAI22_X1 port map( A1 => n3877, A2 => n6332, B1 => n3909, B2 => 
                           n6329, ZN => n989);
   U1272 : OAI22_X1 port map( A1 => n3877, A2 => n6293, B1 => n3909, B2 => 
                           n6290, ZN => n1877);
   U1273 : OAI22_X1 port map( A1 => n3876, A2 => n6332, B1 => n3908, B2 => 
                           n6329, ZN => n967);
   U1274 : OAI22_X1 port map( A1 => n3876, A2 => n6293, B1 => n3908, B2 => 
                           n6290, ZN => n1894);
   U1275 : OAI22_X1 port map( A1 => n3875, A2 => n6332, B1 => n3907, B2 => 
                           n6329, ZN => n946);
   U1276 : OAI22_X1 port map( A1 => n3875, A2 => n6293, B1 => n3907, B2 => 
                           n6290, ZN => n1911);
   U1277 : OAI22_X1 port map( A1 => n3874, A2 => n6332, B1 => n3906, B2 => 
                           n6329, ZN => n927);
   U1278 : OAI22_X1 port map( A1 => n3874, A2 => n6293, B1 => n3906, B2 => 
                           n6290, ZN => n1928);
   U1279 : OAI22_X1 port map( A1 => n3873, A2 => n6332, B1 => n3905, B2 => 
                           n6329, ZN => n910);
   U1280 : OAI22_X1 port map( A1 => n3873, A2 => n6293, B1 => n3905, B2 => 
                           n6290, ZN => n1945);
   U1281 : OAI22_X1 port map( A1 => n3872, A2 => n6332, B1 => n3904, B2 => 
                           n6329, ZN => n893);
   U1282 : OAI22_X1 port map( A1 => n3872, A2 => n6293, B1 => n3904, B2 => 
                           n6290, ZN => n1962);
   U1283 : OAI22_X1 port map( A1 => n3871, A2 => n6332, B1 => n3903, B2 => 
                           n6329, ZN => n876);
   U1284 : OAI22_X1 port map( A1 => n3871, A2 => n6293, B1 => n3903, B2 => 
                           n6290, ZN => n1979);
   U1285 : OAI22_X1 port map( A1 => n3870, A2 => n6332, B1 => n3902, B2 => 
                           n6329, ZN => n836);
   U1286 : OAI22_X1 port map( A1 => n3870, A2 => n6293, B1 => n3902, B2 => 
                           n6290, ZN => n2021);
   U1287 : OAI222_X1 port map( A1 => n2319, A2 => n6319, B1 => n2318, B2 => 
                           n6316, C1 => n3805, C2 => n6313, ZN => n1424);
   U1288 : OAI222_X1 port map( A1 => n2319, A2 => n6284, B1 => n2318, B2 => 
                           n6281, C1 => n3805, C2 => n6278, ZN => n1454);
   U1289 : OAI222_X1 port map( A1 => n2323, A2 => n6319, B1 => n2322, B2 => 
                           n6316, C1 => n3804, C2 => n6313, ZN => n1382);
   U1290 : OAI222_X1 port map( A1 => n2323, A2 => n6284, B1 => n2322, B2 => 
                           n6281, C1 => n3804, C2 => n6278, ZN => n1487);
   U1291 : OAI222_X1 port map( A1 => n2327, A2 => n6319, B1 => n2326, B2 => 
                           n6316, C1 => n3803, C2 => n6313, ZN => n1365);
   U1292 : OAI222_X1 port map( A1 => n2327, A2 => n6284, B1 => n2326, B2 => 
                           n6281, C1 => n3803, C2 => n6278, ZN => n1504);
   U1293 : OAI222_X1 port map( A1 => n2331, A2 => n6319, B1 => n2330, B2 => 
                           n6316, C1 => n3802, C2 => n6313, ZN => n1348);
   U1294 : OAI222_X1 port map( A1 => n2331, A2 => n6284, B1 => n2330, B2 => 
                           n6281, C1 => n3802, C2 => n6278, ZN => n1521);
   U1295 : OAI222_X1 port map( A1 => n2335, A2 => n6319, B1 => n2334, B2 => 
                           n6316, C1 => n3801, C2 => n6313, ZN => n1331);
   U1296 : OAI222_X1 port map( A1 => n2335, A2 => n6284, B1 => n2334, B2 => 
                           n6281, C1 => n3801, C2 => n6278, ZN => n1538);
   U1297 : OAI222_X1 port map( A1 => n2339, A2 => n6319, B1 => n2338, B2 => 
                           n6316, C1 => n3800, C2 => n6313, ZN => n1314);
   U1298 : OAI222_X1 port map( A1 => n2339, A2 => n6284, B1 => n2338, B2 => 
                           n6281, C1 => n3800, C2 => n6278, ZN => n1555);
   U1299 : OAI222_X1 port map( A1 => n2343, A2 => n6319, B1 => n2342, B2 => 
                           n6316, C1 => n3799, C2 => n6313, ZN => n1297);
   U1300 : OAI222_X1 port map( A1 => n2343, A2 => n6284, B1 => n2342, B2 => 
                           n6281, C1 => n3799, C2 => n6278, ZN => n1572);
   U1301 : OAI222_X1 port map( A1 => n2347, A2 => n6319, B1 => n2346, B2 => 
                           n6316, C1 => n3798, C2 => n6313, ZN => n1280);
   U1302 : OAI222_X1 port map( A1 => n2347, A2 => n6284, B1 => n2346, B2 => 
                           n6281, C1 => n3798, C2 => n6278, ZN => n1589);
   U1303 : OAI222_X1 port map( A1 => n2351, A2 => n6319, B1 => n2350, B2 => 
                           n6316, C1 => n3797, C2 => n6313, ZN => n1263);
   U1304 : OAI222_X1 port map( A1 => n2351, A2 => n6283, B1 => n2350, B2 => 
                           n6280, C1 => n3797, C2 => n6277, ZN => n1606);
   U1305 : OAI222_X1 port map( A1 => n2355, A2 => n6319, B1 => n2354, B2 => 
                           n6316, C1 => n3796, C2 => n6313, ZN => n1246);
   U1306 : OAI222_X1 port map( A1 => n2355, A2 => n6283, B1 => n2354, B2 => 
                           n6280, C1 => n3796, C2 => n6277, ZN => n1623);
   U1307 : OAI222_X1 port map( A1 => n2359, A2 => n6319, B1 => n2358, B2 => 
                           n6316, C1 => n3795, C2 => n6313, ZN => n1229);
   U1308 : OAI222_X1 port map( A1 => n2359, A2 => n6283, B1 => n2358, B2 => 
                           n6280, C1 => n3795, C2 => n6277, ZN => n1640);
   U1309 : OAI222_X1 port map( A1 => n2363, A2 => n6319, B1 => n2362, B2 => 
                           n6316, C1 => n3794, C2 => n6313, ZN => n1212);
   U1310 : OAI222_X1 port map( A1 => n2363, A2 => n6283, B1 => n2362, B2 => 
                           n6280, C1 => n3794, C2 => n6277, ZN => n1657);
   U1311 : OAI222_X1 port map( A1 => n2367, A2 => n6320, B1 => n2366, B2 => 
                           n6317, C1 => n3793, C2 => n6314, ZN => n1195);
   U1312 : OAI222_X1 port map( A1 => n2367, A2 => n6283, B1 => n2366, B2 => 
                           n6280, C1 => n3793, C2 => n6277, ZN => n1674);
   U1313 : OAI222_X1 port map( A1 => n2371, A2 => n6320, B1 => n2370, B2 => 
                           n6317, C1 => n3792, C2 => n6314, ZN => n1178);
   U1314 : OAI222_X1 port map( A1 => n2371, A2 => n6283, B1 => n2370, B2 => 
                           n6280, C1 => n3792, C2 => n6277, ZN => n1691);
   U1315 : OAI222_X1 port map( A1 => n2375, A2 => n6320, B1 => n2374, B2 => 
                           n6317, C1 => n3791, C2 => n6314, ZN => n1161);
   U1316 : OAI222_X1 port map( A1 => n2375, A2 => n6283, B1 => n2374, B2 => 
                           n6280, C1 => n3791, C2 => n6277, ZN => n1708);
   U1317 : OAI222_X1 port map( A1 => n2379, A2 => n6320, B1 => n2378, B2 => 
                           n6317, C1 => n3790, C2 => n6314, ZN => n1144);
   U1318 : OAI222_X1 port map( A1 => n2379, A2 => n6283, B1 => n2378, B2 => 
                           n6280, C1 => n3790, C2 => n6277, ZN => n1725);
   U1319 : OAI222_X1 port map( A1 => n2383, A2 => n6320, B1 => n2382, B2 => 
                           n6317, C1 => n3789, C2 => n6314, ZN => n1127);
   U1320 : OAI222_X1 port map( A1 => n2383, A2 => n6283, B1 => n2382, B2 => 
                           n6280, C1 => n3789, C2 => n6277, ZN => n1742);
   U1321 : OAI222_X1 port map( A1 => n2387, A2 => n6320, B1 => n2386, B2 => 
                           n6317, C1 => n3788, C2 => n6314, ZN => n1110);
   U1322 : OAI222_X1 port map( A1 => n2387, A2 => n6283, B1 => n2386, B2 => 
                           n6280, C1 => n3788, C2 => n6277, ZN => n1759);
   U1323 : OAI222_X1 port map( A1 => n2391, A2 => n6320, B1 => n2390, B2 => 
                           n6317, C1 => n3787, C2 => n6314, ZN => n1093);
   U1324 : OAI222_X1 port map( A1 => n2391, A2 => n6283, B1 => n2390, B2 => 
                           n6280, C1 => n3787, C2 => n6277, ZN => n1776);
   U1325 : OAI222_X1 port map( A1 => n2395, A2 => n6320, B1 => n2394, B2 => 
                           n6317, C1 => n3786, C2 => n6314, ZN => n1076);
   U1326 : OAI222_X1 port map( A1 => n2395, A2 => n6283, B1 => n2394, B2 => 
                           n6280, C1 => n3786, C2 => n6277, ZN => n1793);
   U1327 : OAI222_X1 port map( A1 => n2399, A2 => n6320, B1 => n2398, B2 => 
                           n6317, C1 => n3785, C2 => n6314, ZN => n1059);
   U1328 : OAI222_X1 port map( A1 => n2399, A2 => n6282, B1 => n2398, B2 => 
                           n6279, C1 => n3785, C2 => n6276, ZN => n1810);
   U1329 : OAI222_X1 port map( A1 => n2403, A2 => n6320, B1 => n2402, B2 => 
                           n6317, C1 => n3784, C2 => n6314, ZN => n1042);
   U1330 : OAI222_X1 port map( A1 => n2403, A2 => n6282, B1 => n2402, B2 => 
                           n6279, C1 => n3784, C2 => n6276, ZN => n1827);
   U1331 : OAI222_X1 port map( A1 => n2407, A2 => n6320, B1 => n2406, B2 => 
                           n6317, C1 => n3783, C2 => n6314, ZN => n1025);
   U1332 : OAI222_X1 port map( A1 => n2407, A2 => n6282, B1 => n2406, B2 => 
                           n6279, C1 => n3783, C2 => n6276, ZN => n1844);
   U1333 : OAI222_X1 port map( A1 => n2411, A2 => n6320, B1 => n2410, B2 => 
                           n6317, C1 => n3782, C2 => n6314, ZN => n1008);
   U1334 : OAI222_X1 port map( A1 => n2411, A2 => n6282, B1 => n2410, B2 => 
                           n6279, C1 => n3782, C2 => n6276, ZN => n1861);
   U1335 : OAI222_X1 port map( A1 => n2415, A2 => n6321, B1 => n2414, B2 => 
                           n6318, C1 => n3781, C2 => n6315, ZN => n990);
   U1336 : OAI222_X1 port map( A1 => n2415, A2 => n6282, B1 => n2414, B2 => 
                           n6279, C1 => n3781, C2 => n6276, ZN => n1878);
   U1337 : OAI222_X1 port map( A1 => n2419, A2 => n6321, B1 => n2418, B2 => 
                           n6318, C1 => n3780, C2 => n6315, ZN => n968);
   U1338 : OAI222_X1 port map( A1 => n2419, A2 => n6282, B1 => n2418, B2 => 
                           n6279, C1 => n3780, C2 => n6276, ZN => n1895);
   U1339 : OAI222_X1 port map( A1 => n2423, A2 => n6321, B1 => n2422, B2 => 
                           n6318, C1 => n3779, C2 => n6315, ZN => n947);
   U1340 : OAI222_X1 port map( A1 => n2423, A2 => n6282, B1 => n2422, B2 => 
                           n6279, C1 => n3779, C2 => n6276, ZN => n1912);
   U1341 : OAI222_X1 port map( A1 => n2427, A2 => n6321, B1 => n2426, B2 => 
                           n6318, C1 => n3778, C2 => n6315, ZN => n928);
   U1342 : OAI222_X1 port map( A1 => n2427, A2 => n6282, B1 => n2426, B2 => 
                           n6279, C1 => n3778, C2 => n6276, ZN => n1929);
   U1343 : OAI222_X1 port map( A1 => n2431, A2 => n6321, B1 => n2430, B2 => 
                           n6318, C1 => n3777, C2 => n6315, ZN => n911);
   U1344 : OAI222_X1 port map( A1 => n2431, A2 => n6282, B1 => n2430, B2 => 
                           n6279, C1 => n3777, C2 => n6276, ZN => n1946);
   U1345 : OAI222_X1 port map( A1 => n2435, A2 => n6321, B1 => n2434, B2 => 
                           n6318, C1 => n3776, C2 => n6315, ZN => n894);
   U1346 : OAI222_X1 port map( A1 => n2435, A2 => n6282, B1 => n2434, B2 => 
                           n6279, C1 => n3776, C2 => n6276, ZN => n1963);
   U1347 : OAI222_X1 port map( A1 => n2439, A2 => n6321, B1 => n2438, B2 => 
                           n6318, C1 => n3775, C2 => n6315, ZN => n877);
   U1348 : OAI222_X1 port map( A1 => n2439, A2 => n6282, B1 => n2438, B2 => 
                           n6279, C1 => n3775, C2 => n6276, ZN => n1980);
   U1349 : OAI222_X1 port map( A1 => n2443, A2 => n6321, B1 => n2442, B2 => 
                           n6318, C1 => n3774, C2 => n6315, ZN => n841);
   U1350 : OAI222_X1 port map( A1 => n2443, A2 => n6282, B1 => n2442, B2 => 
                           n6279, C1 => n3774, C2 => n6276, ZN => n2024);
   U1351 : AOI221_X1 port map( B1 => n6338, B2 => n4060, C1 => n6335, C2 => 
                           n4092, A => n1381, ZN => n1378);
   U1352 : AOI221_X1 port map( B1 => n6299, B2 => n4060, C1 => n6296, C2 => 
                           n4092, A => n1486, ZN => n1483);
   U1353 : AOI221_X1 port map( B1 => n6338, B2 => n4059, C1 => n6335, C2 => 
                           n4091, A => n1364, ZN => n1361);
   U1354 : AOI221_X1 port map( B1 => n6299, B2 => n4059, C1 => n6296, C2 => 
                           n4091, A => n1503, ZN => n1500);
   U1355 : AOI221_X1 port map( B1 => n6338, B2 => n4058, C1 => n6335, C2 => 
                           n4090, A => n1347, ZN => n1344);
   U1356 : AOI221_X1 port map( B1 => n6299, B2 => n4058, C1 => n6296, C2 => 
                           n4090, A => n1520, ZN => n1517);
   U1357 : AOI221_X1 port map( B1 => n6338, B2 => n4057, C1 => n6335, C2 => 
                           n4089, A => n1330, ZN => n1327);
   U1358 : AOI221_X1 port map( B1 => n6299, B2 => n4057, C1 => n6296, C2 => 
                           n4089, A => n1537, ZN => n1534);
   U1359 : AOI221_X1 port map( B1 => n6338, B2 => n4056, C1 => n6335, C2 => 
                           n4088, A => n1313, ZN => n1310);
   U1360 : AOI221_X1 port map( B1 => n6299, B2 => n4056, C1 => n6296, C2 => 
                           n4088, A => n1554, ZN => n1551);
   U1361 : AOI221_X1 port map( B1 => n6338, B2 => n4055, C1 => n6335, C2 => 
                           n4087, A => n1296, ZN => n1293);
   U1362 : AOI221_X1 port map( B1 => n6299, B2 => n4055, C1 => n6296, C2 => 
                           n4087, A => n1571, ZN => n1568);
   U1363 : AOI221_X1 port map( B1 => n6338, B2 => n4054, C1 => n6335, C2 => 
                           n4086, A => n1279, ZN => n1276);
   U1364 : AOI221_X1 port map( B1 => n6299, B2 => n4054, C1 => n6296, C2 => 
                           n4086, A => n1588, ZN => n1585);
   U1365 : AOI221_X1 port map( B1 => n6337, B2 => n4053, C1 => n6334, C2 => 
                           n4085, A => n1262, ZN => n1259);
   U1366 : AOI221_X1 port map( B1 => n6299, B2 => n4053, C1 => n6296, C2 => 
                           n4085, A => n1605, ZN => n1602);
   U1367 : AOI221_X1 port map( B1 => n6337, B2 => n4052, C1 => n6334, C2 => 
                           n4084, A => n1245, ZN => n1242);
   U1368 : AOI221_X1 port map( B1 => n6299, B2 => n4052, C1 => n6296, C2 => 
                           n4084, A => n1622, ZN => n1619);
   U1369 : AOI221_X1 port map( B1 => n6337, B2 => n4051, C1 => n6334, C2 => 
                           n4083, A => n1228, ZN => n1225);
   U1370 : AOI221_X1 port map( B1 => n6299, B2 => n4051, C1 => n6296, C2 => 
                           n4083, A => n1639, ZN => n1636);
   U1371 : AOI221_X1 port map( B1 => n6337, B2 => n4050, C1 => n6334, C2 => 
                           n4082, A => n1211, ZN => n1208);
   U1372 : AOI221_X1 port map( B1 => n6299, B2 => n4050, C1 => n6296, C2 => 
                           n4082, A => n1656, ZN => n1653);
   U1373 : AOI221_X1 port map( B1 => n6337, B2 => n4049, C1 => n6334, C2 => 
                           n4081, A => n1194, ZN => n1191);
   U1374 : AOI221_X1 port map( B1 => n6300, B2 => n4049, C1 => n6297, C2 => 
                           n4081, A => n1673, ZN => n1670);
   U1375 : AOI221_X1 port map( B1 => n6337, B2 => n4048, C1 => n6334, C2 => 
                           n4080, A => n1177, ZN => n1174);
   U1376 : AOI221_X1 port map( B1 => n6300, B2 => n4048, C1 => n6297, C2 => 
                           n4080, A => n1690, ZN => n1687);
   U1377 : AOI221_X1 port map( B1 => n6337, B2 => n4047, C1 => n6334, C2 => 
                           n4079, A => n1160, ZN => n1157);
   U1378 : AOI221_X1 port map( B1 => n6300, B2 => n4047, C1 => n6297, C2 => 
                           n4079, A => n1707, ZN => n1704);
   U1379 : AOI221_X1 port map( B1 => n6337, B2 => n4046, C1 => n6334, C2 => 
                           n4078, A => n1143, ZN => n1140);
   U1380 : AOI221_X1 port map( B1 => n6300, B2 => n4046, C1 => n6297, C2 => 
                           n4078, A => n1724, ZN => n1721);
   U1381 : AOI221_X1 port map( B1 => n6337, B2 => n4045, C1 => n6334, C2 => 
                           n4077, A => n1126, ZN => n1123);
   U1382 : AOI221_X1 port map( B1 => n6300, B2 => n4045, C1 => n6297, C2 => 
                           n4077, A => n1741, ZN => n1738);
   U1383 : AOI221_X1 port map( B1 => n6337, B2 => n4044, C1 => n6334, C2 => 
                           n4076, A => n1109, ZN => n1106);
   U1384 : AOI221_X1 port map( B1 => n6300, B2 => n4044, C1 => n6297, C2 => 
                           n4076, A => n1758, ZN => n1755);
   U1385 : AOI221_X1 port map( B1 => n6337, B2 => n4043, C1 => n6334, C2 => 
                           n4075, A => n1092, ZN => n1089);
   U1386 : AOI221_X1 port map( B1 => n6300, B2 => n4043, C1 => n6297, C2 => 
                           n4075, A => n1775, ZN => n1772);
   U1387 : AOI221_X1 port map( B1 => n6337, B2 => n4042, C1 => n6334, C2 => 
                           n4074, A => n1075, ZN => n1072);
   U1388 : AOI221_X1 port map( B1 => n6300, B2 => n4042, C1 => n6297, C2 => 
                           n4074, A => n1792, ZN => n1789);
   U1389 : AOI221_X1 port map( B1 => n6336, B2 => n4041, C1 => n6333, C2 => 
                           n4073, A => n1058, ZN => n1055);
   U1390 : AOI221_X1 port map( B1 => n6300, B2 => n4041, C1 => n6297, C2 => 
                           n4073, A => n1809, ZN => n1806);
   U1391 : AOI221_X1 port map( B1 => n6336, B2 => n4040, C1 => n6333, C2 => 
                           n4072, A => n1041, ZN => n1038);
   U1392 : AOI221_X1 port map( B1 => n6300, B2 => n4040, C1 => n6297, C2 => 
                           n4072, A => n1826, ZN => n1823);
   U1393 : AOI221_X1 port map( B1 => n6336, B2 => n4039, C1 => n6333, C2 => 
                           n4071, A => n1024, ZN => n1021);
   U1394 : AOI221_X1 port map( B1 => n6300, B2 => n4039, C1 => n6297, C2 => 
                           n4071, A => n1843, ZN => n1840);
   U1395 : AOI221_X1 port map( B1 => n6336, B2 => n4038, C1 => n6333, C2 => 
                           n4070, A => n1007, ZN => n1004);
   U1396 : AOI221_X1 port map( B1 => n6300, B2 => n4038, C1 => n6297, C2 => 
                           n4070, A => n1860, ZN => n1857);
   U1397 : AOI221_X1 port map( B1 => n6336, B2 => n4037, C1 => n6333, C2 => 
                           n4069, A => n989, ZN => n984);
   U1398 : AOI221_X1 port map( B1 => n6301, B2 => n4037, C1 => n6298, C2 => 
                           n4069, A => n1877, ZN => n1874);
   U1399 : AOI221_X1 port map( B1 => n6336, B2 => n4036, C1 => n6333, C2 => 
                           n4068, A => n967, ZN => n963);
   U1400 : AOI221_X1 port map( B1 => n6301, B2 => n4036, C1 => n6298, C2 => 
                           n4068, A => n1894, ZN => n1891);
   U1401 : AOI221_X1 port map( B1 => n6336, B2 => n4035, C1 => n6333, C2 => 
                           n4067, A => n946, ZN => n943);
   U1402 : AOI221_X1 port map( B1 => n6301, B2 => n4035, C1 => n6298, C2 => 
                           n4067, A => n1911, ZN => n1908);
   U1403 : AOI221_X1 port map( B1 => n6336, B2 => n4034, C1 => n6333, C2 => 
                           n4066, A => n927, ZN => n924);
   U1404 : AOI221_X1 port map( B1 => n6301, B2 => n4034, C1 => n6298, C2 => 
                           n4066, A => n1928, ZN => n1925);
   U1405 : AOI221_X1 port map( B1 => n6336, B2 => n4033, C1 => n6333, C2 => 
                           n4065, A => n910, ZN => n907);
   U1406 : AOI221_X1 port map( B1 => n6301, B2 => n4033, C1 => n6298, C2 => 
                           n4065, A => n1945, ZN => n1942);
   U1407 : AOI221_X1 port map( B1 => n6336, B2 => n4032, C1 => n6333, C2 => 
                           n4064, A => n893, ZN => n890);
   U1408 : AOI221_X1 port map( B1 => n6301, B2 => n4032, C1 => n6298, C2 => 
                           n4064, A => n1962, ZN => n1959);
   U1409 : AOI221_X1 port map( B1 => n6336, B2 => n4031, C1 => n6333, C2 => 
                           n4063, A => n876, ZN => n873);
   U1410 : AOI221_X1 port map( B1 => n6301, B2 => n4031, C1 => n6298, C2 => 
                           n4063, A => n1979, ZN => n1976);
   U1411 : INV_X1 port map( A => n6084, ZN => n6083);
   U1412 : INV_X1 port map( A => n6093, ZN => n6092);
   U1413 : INV_X1 port map( A => DATAIN(0), ZN => n6339);
   U1414 : INV_X1 port map( A => DATAIN(0), ZN => n6340);
   U1415 : INV_X1 port map( A => DATAIN(1), ZN => n6341);
   U1416 : INV_X1 port map( A => DATAIN(1), ZN => n6342);
   U1417 : INV_X1 port map( A => DATAIN(2), ZN => n6343);
   U1418 : INV_X1 port map( A => DATAIN(2), ZN => n6344);
   U1419 : INV_X1 port map( A => DATAIN(3), ZN => n6345);
   U1420 : INV_X1 port map( A => DATAIN(3), ZN => n6346);
   U1421 : CLKBUF_X1 port map( A => n6478, Z => n6382);
   U1422 : CLKBUF_X1 port map( A => n6478, Z => n6383);
   U1423 : CLKBUF_X1 port map( A => n6478, Z => n6384);
   U1424 : CLKBUF_X1 port map( A => n6478, Z => n6385);
   U1425 : CLKBUF_X1 port map( A => n6478, Z => n6386);
   U1426 : CLKBUF_X1 port map( A => n6477, Z => n6387);
   U1427 : CLKBUF_X1 port map( A => n6477, Z => n6388);
   U1428 : CLKBUF_X1 port map( A => n6477, Z => n6389);
   U1429 : CLKBUF_X1 port map( A => n6477, Z => n6390);
   U1430 : CLKBUF_X1 port map( A => n6477, Z => n6391);
   U1431 : CLKBUF_X1 port map( A => n6477, Z => n6392);
   U1432 : CLKBUF_X1 port map( A => n6476, Z => n6393);
   U1433 : CLKBUF_X1 port map( A => n6476, Z => n6394);
   U1434 : CLKBUF_X1 port map( A => n6476, Z => n6395);
   U1435 : CLKBUF_X1 port map( A => n6476, Z => n6396);
   U1436 : CLKBUF_X1 port map( A => n6476, Z => n6397);
   U1437 : CLKBUF_X1 port map( A => n6476, Z => n6398);
   U1438 : CLKBUF_X1 port map( A => n6475, Z => n6399);
   U1439 : CLKBUF_X1 port map( A => n6475, Z => n6400);
   U1440 : CLKBUF_X1 port map( A => n6475, Z => n6401);
   U1441 : CLKBUF_X1 port map( A => n6475, Z => n6402);
   U1442 : CLKBUF_X1 port map( A => n6475, Z => n6403);
   U1443 : CLKBUF_X1 port map( A => n6475, Z => n6404);
   U1444 : CLKBUF_X1 port map( A => n6474, Z => n6405);
   U1445 : CLKBUF_X1 port map( A => n6474, Z => n6406);
   U1446 : CLKBUF_X1 port map( A => n6474, Z => n6407);
   U1447 : CLKBUF_X1 port map( A => n6474, Z => n6408);
   U1448 : CLKBUF_X1 port map( A => n6474, Z => n6409);
   U1449 : CLKBUF_X1 port map( A => n6474, Z => n6410);
   U1450 : CLKBUF_X1 port map( A => n6473, Z => n6411);
   U1451 : CLKBUF_X1 port map( A => n6473, Z => n6412);
   U1452 : CLKBUF_X1 port map( A => n6473, Z => n6413);
   U1453 : CLKBUF_X1 port map( A => n6473, Z => n6414);
   U1454 : CLKBUF_X1 port map( A => n6473, Z => n6415);
   U1455 : CLKBUF_X1 port map( A => n6473, Z => n6416);
   U1456 : CLKBUF_X1 port map( A => n6472, Z => n6417);
   U1457 : CLKBUF_X1 port map( A => n6472, Z => n6418);
   U1458 : CLKBUF_X1 port map( A => n6472, Z => n6419);
   U1459 : CLKBUF_X1 port map( A => n6472, Z => n6420);
   U1460 : CLKBUF_X1 port map( A => n6472, Z => n6421);
   U1461 : CLKBUF_X1 port map( A => n6472, Z => n6422);
   U1462 : CLKBUF_X1 port map( A => n6471, Z => n6423);
   U1463 : CLKBUF_X1 port map( A => n6471, Z => n6424);
   U1464 : CLKBUF_X1 port map( A => n6471, Z => n6425);
   U1465 : CLKBUF_X1 port map( A => n6471, Z => n6426);
   U1466 : CLKBUF_X1 port map( A => n6471, Z => n6427);
   U1467 : CLKBUF_X1 port map( A => n6471, Z => n6428);
   U1468 : CLKBUF_X1 port map( A => n6470, Z => n6429);
   U1469 : CLKBUF_X1 port map( A => n6470, Z => n6430);
   U1470 : CLKBUF_X1 port map( A => n6470, Z => n6431);
   U1471 : CLKBUF_X1 port map( A => n6470, Z => n6432);
   U1472 : CLKBUF_X1 port map( A => n6470, Z => n6433);
   U1473 : CLKBUF_X1 port map( A => n6470, Z => n6434);
   U1474 : CLKBUF_X1 port map( A => n6469, Z => n6435);
   U1475 : CLKBUF_X1 port map( A => n6469, Z => n6436);
   U1476 : CLKBUF_X1 port map( A => n6469, Z => n6437);
   U1477 : CLKBUF_X1 port map( A => n6469, Z => n6438);
   U1478 : CLKBUF_X1 port map( A => n6469, Z => n6439);
   U1479 : CLKBUF_X1 port map( A => n6469, Z => n6440);
   U1480 : CLKBUF_X1 port map( A => n6468, Z => n6441);
   U1481 : CLKBUF_X1 port map( A => n6468, Z => n6442);
   U1482 : CLKBUF_X1 port map( A => n6468, Z => n6443);
   U1483 : CLKBUF_X1 port map( A => n6468, Z => n6444);
   U1484 : CLKBUF_X1 port map( A => n6468, Z => n6445);
   U1485 : CLKBUF_X1 port map( A => n6468, Z => n6446);
   U1486 : CLKBUF_X1 port map( A => n6467, Z => n6447);
   U1487 : CLKBUF_X1 port map( A => n6467, Z => n6448);
   U1488 : CLKBUF_X1 port map( A => n6467, Z => n6449);
   U1489 : CLKBUF_X1 port map( A => n6467, Z => n6450);
   U1490 : CLKBUF_X1 port map( A => n6467, Z => n6451);
   U1491 : CLKBUF_X1 port map( A => n6467, Z => n6452);
   U1492 : CLKBUF_X1 port map( A => n6466, Z => n6453);
   U1493 : CLKBUF_X1 port map( A => n6466, Z => n6454);
   U1494 : CLKBUF_X1 port map( A => n6466, Z => n6455);
   U1495 : CLKBUF_X1 port map( A => n6466, Z => n6456);
   U1496 : CLKBUF_X1 port map( A => n6466, Z => n6457);
   U1497 : CLKBUF_X1 port map( A => n6466, Z => n6458);
   U1498 : CLKBUF_X1 port map( A => n6465, Z => n6459);
   U1499 : CLKBUF_X1 port map( A => n6465, Z => n6460);
   U1500 : CLKBUF_X1 port map( A => n6465, Z => n6461);
   U1501 : CLKBUF_X1 port map( A => n6465, Z => n6462);
   U1502 : CLKBUF_X1 port map( A => n6465, Z => n6463);
   U1503 : INV_X1 port map( A => ADD_WR(2), ZN => n7591);
   U1504 : INV_X1 port map( A => ADD_WR(3), ZN => n7590);
   U1505 : INV_X1 port map( A => ADD_WR(4), ZN => n7589);
   U1506 : INV_X1 port map( A => ADD_RS1(3), ZN => n7592);
   U1507 : INV_X1 port map( A => ADD_RS1(0), ZN => n7593);
   U1508 : INV_X1 port map( A => ADD_RS1(4), ZN => n7901);
   U1509 : INV_X1 port map( A => ADD_RS1(1), ZN => n6479);
   U1510 : INV_X1 port map( A => n2059, ZN => n7587);
   U1511 : INV_X1 port map( A => n2316, ZN => n7585);
   U1512 : INV_X1 port map( A => ADD_RS2(3), ZN => n7594);
   U1513 : INV_X1 port map( A => ADD_RS2(0), ZN => n7595);
   U1514 : INV_X1 port map( A => ADD_RS2(4), ZN => n7899);
   U1515 : INV_X1 port map( A => ADD_RS2(1), ZN => n6480);
   U1516 : INV_X1 port map( A => n2028, ZN => n7588);
   U1517 : INV_X1 port map( A => n2440, ZN => n7586);
   U1518 : INV_X1 port map( A => n4125, ZN => n6938);
   U1519 : NAND3_X1 port map( A1 => n749, A2 => n7589, A3 => n7590, ZN => n6481
                           );
   U1520 : INV_X1 port map( A => n6481, ZN => n6489);
   U1521 : INV_X1 port map( A => ADD_WR(1), ZN => n6482);
   U1522 : INV_X1 port map( A => n4124, ZN => n6957);
   U1523 : INV_X1 port map( A => n4123, ZN => n6975);
   U1524 : INV_X1 port map( A => n4122, ZN => n6993);
   U1525 : INV_X1 port map( A => n4121, ZN => n7012);
   U1526 : INV_X1 port map( A => n4120, ZN => n7031);
   U1527 : INV_X1 port map( A => n4119, ZN => n7050);
   U1528 : INV_X1 port map( A => n4118, ZN => n7069);
   U1529 : INV_X1 port map( A => n4117, ZN => n7088);
   U1530 : INV_X1 port map( A => n4116, ZN => n7107);
   U1531 : INV_X1 port map( A => n4115, ZN => n7126);
   U1532 : INV_X1 port map( A => n4114, ZN => n7145);
   U1533 : INV_X1 port map( A => n4113, ZN => n7164);
   U1534 : INV_X1 port map( A => n4112, ZN => n7183);
   U1535 : INV_X1 port map( A => n4111, ZN => n7202);
   U1536 : INV_X1 port map( A => n4110, ZN => n7221);
   U1537 : INV_X1 port map( A => n4109, ZN => n7240);
   U1538 : INV_X1 port map( A => n4108, ZN => n7259);
   U1539 : INV_X1 port map( A => n4107, ZN => n7278);
   U1540 : INV_X1 port map( A => n4106, ZN => n7297);
   U1541 : INV_X1 port map( A => n4105, ZN => n7316);
   U1542 : INV_X1 port map( A => n4104, ZN => n7335);
   U1543 : INV_X1 port map( A => n4103, ZN => n7354);
   U1544 : INV_X1 port map( A => n4102, ZN => n7373);
   U1545 : MUX2_X1 port map( A => n5210, B => DATAIN(23), S => n6006, Z => 
                           n4277);
   U1546 : INV_X1 port map( A => n4101, ZN => n7392);
   U1547 : INV_X1 port map( A => n4100, ZN => n7411);
   U1548 : INV_X1 port map( A => n4099, ZN => n7430);
   U1549 : INV_X1 port map( A => n4098, ZN => n7449);
   U1550 : INV_X1 port map( A => n4097, ZN => n7468);
   U1551 : INV_X1 port map( A => n4096, ZN => n7487);
   U1552 : MUX2_X1 port map( A => n5204, B => DATAIN(29), S => n6007, Z => 
                           n4283);
   U1553 : INV_X1 port map( A => n4095, ZN => n7506);
   U1554 : MUX2_X1 port map( A => n5203, B => DATAIN(30), S => n6007, Z => 
                           n4284);
   U1555 : INV_X1 port map( A => n4094, ZN => n7531);
   U1556 : MUX2_X1 port map( A => n5169, B => DATAIN(31), S => n6007, Z => 
                           n4285);
   U1557 : MUX2_X1 port map( A => n5872, B => DATAIN(0), S => n6008, Z => n4158
                           );
   U1558 : MUX2_X1 port map( A => n5871, B => DATAIN(1), S => n6008, Z => n4159
                           );
   U1559 : MUX2_X1 port map( A => n5870, B => DATAIN(2), S => n6008, Z => n4160
                           );
   U1560 : MUX2_X1 port map( A => n5869, B => DATAIN(3), S => n6008, Z => n4161
                           );
   U1561 : MUX2_X1 port map( A => n5868, B => DATAIN(4), S => n6008, Z => n4162
                           );
   U1562 : MUX2_X1 port map( A => n5867, B => DATAIN(5), S => n6008, Z => n4163
                           );
   U1563 : MUX2_X1 port map( A => n5866, B => DATAIN(6), S => n6008, Z => n4164
                           );
   U1564 : MUX2_X1 port map( A => n5865, B => DATAIN(7), S => n6008, Z => n4165
                           );
   U1565 : MUX2_X1 port map( A => n5864, B => DATAIN(8), S => n6008, Z => n4166
                           );
   U1566 : MUX2_X1 port map( A => n5863, B => DATAIN(9), S => n6008, Z => n4167
                           );
   U1567 : MUX2_X1 port map( A => n5862, B => DATAIN(10), S => n6008, Z => 
                           n4168);
   U1568 : MUX2_X1 port map( A => n5861, B => DATAIN(11), S => n6008, Z => 
                           n4169);
   U1569 : MUX2_X1 port map( A => n5860, B => DATAIN(12), S => n6009, Z => 
                           n4170);
   U1570 : MUX2_X1 port map( A => n5859, B => DATAIN(13), S => n6009, Z => 
                           n4171);
   U1571 : MUX2_X1 port map( A => n5858, B => DATAIN(14), S => n6009, Z => 
                           n4172);
   U1572 : MUX2_X1 port map( A => n5857, B => DATAIN(15), S => n6009, Z => 
                           n4173);
   U1573 : MUX2_X1 port map( A => n5856, B => DATAIN(16), S => n6009, Z => 
                           n4174);
   U1574 : MUX2_X1 port map( A => n5855, B => DATAIN(17), S => n6009, Z => 
                           n4175);
   U1575 : MUX2_X1 port map( A => n5854, B => DATAIN(18), S => n6009, Z => 
                           n4176);
   U1576 : MUX2_X1 port map( A => n5853, B => DATAIN(19), S => n6009, Z => 
                           n4177);
   U1577 : MUX2_X1 port map( A => n5852, B => DATAIN(20), S => n6009, Z => 
                           n4178);
   U1578 : MUX2_X1 port map( A => n5851, B => DATAIN(21), S => n6009, Z => 
                           n4179);
   U1579 : MUX2_X1 port map( A => n5850, B => DATAIN(22), S => n6009, Z => 
                           n4180);
   U1580 : MUX2_X1 port map( A => n5849, B => DATAIN(23), S => n6009, Z => 
                           n4181);
   U1581 : MUX2_X1 port map( A => n5848, B => DATAIN(24), S => n6010, Z => 
                           n4182);
   U1582 : MUX2_X1 port map( A => n5847, B => DATAIN(25), S => n6010, Z => 
                           n4183);
   U1583 : MUX2_X1 port map( A => n5846, B => DATAIN(26), S => n6010, Z => 
                           n4184);
   U1584 : MUX2_X1 port map( A => n5845, B => DATAIN(27), S => n6010, Z => 
                           n4185);
   U1585 : MUX2_X1 port map( A => n5844, B => DATAIN(28), S => n6010, Z => 
                           n4186);
   U1586 : MUX2_X1 port map( A => n5843, B => DATAIN(29), S => n6010, Z => 
                           n4187);
   U1587 : MUX2_X1 port map( A => n5842, B => DATAIN(30), S => n6010, Z => 
                           n4188);
   U1588 : MUX2_X1 port map( A => n5841, B => DATAIN(31), S => n6010, Z => 
                           n4189);
   U1589 : MUX2_X1 port map( A => n5874, B => DATAIN(0), S => n6011, Z => n4222
                           );
   U1590 : MUX2_X1 port map( A => n5357, B => DATAIN(1), S => n6011, Z => n4223
                           );
   U1591 : MUX2_X1 port map( A => n5356, B => DATAIN(2), S => n6011, Z => n4224
                           );
   U1592 : MUX2_X1 port map( A => n5355, B => DATAIN(3), S => n6011, Z => n4225
                           );
   U1593 : MUX2_X1 port map( A => n5354, B => DATAIN(4), S => n6011, Z => n4226
                           );
   U1594 : MUX2_X1 port map( A => n5353, B => DATAIN(5), S => n6011, Z => n4227
                           );
   U1595 : MUX2_X1 port map( A => n5352, B => DATAIN(6), S => n6011, Z => n4228
                           );
   U1596 : MUX2_X1 port map( A => n5351, B => DATAIN(7), S => n6011, Z => n4229
                           );
   U1597 : MUX2_X1 port map( A => n5350, B => DATAIN(8), S => n6011, Z => n4230
                           );
   U1598 : MUX2_X1 port map( A => n5349, B => DATAIN(9), S => n6011, Z => n4231
                           );
   U1599 : MUX2_X1 port map( A => n5348, B => DATAIN(10), S => n6011, Z => 
                           n4232);
   U1600 : MUX2_X1 port map( A => n5347, B => DATAIN(11), S => n6011, Z => 
                           n4233);
   U1601 : MUX2_X1 port map( A => n5346, B => DATAIN(12), S => n6012, Z => 
                           n4234);
   U1602 : MUX2_X1 port map( A => n5345, B => DATAIN(13), S => n6012, Z => 
                           n4235);
   U1603 : MUX2_X1 port map( A => n5344, B => DATAIN(14), S => n6012, Z => 
                           n4236);
   U1604 : MUX2_X1 port map( A => n5343, B => DATAIN(15), S => n6012, Z => 
                           n4237);
   U1605 : MUX2_X1 port map( A => n5342, B => DATAIN(16), S => n6012, Z => 
                           n4238);
   U1606 : MUX2_X1 port map( A => n5341, B => DATAIN(17), S => n6012, Z => 
                           n4239);
   U1607 : MUX2_X1 port map( A => n5340, B => DATAIN(18), S => n6012, Z => 
                           n4240);
   U1608 : MUX2_X1 port map( A => n5339, B => DATAIN(19), S => n6012, Z => 
                           n4241);
   U1609 : MUX2_X1 port map( A => n5338, B => DATAIN(20), S => n6012, Z => 
                           n4242);
   U1610 : MUX2_X1 port map( A => n5337, B => DATAIN(21), S => n6012, Z => 
                           n4243);
   U1611 : MUX2_X1 port map( A => n5336, B => DATAIN(22), S => n6012, Z => 
                           n4244);
   U1612 : MUX2_X1 port map( A => n5335, B => DATAIN(23), S => n6012, Z => 
                           n4245);
   U1613 : MUX2_X1 port map( A => n5334, B => DATAIN(24), S => n6013, Z => 
                           n4246);
   U1614 : MUX2_X1 port map( A => n5333, B => DATAIN(25), S => n6013, Z => 
                           n4247);
   U1615 : MUX2_X1 port map( A => n5332, B => DATAIN(26), S => n6013, Z => 
                           n4248);
   U1616 : MUX2_X1 port map( A => n5331, B => DATAIN(27), S => n6013, Z => 
                           n4249);
   U1617 : MUX2_X1 port map( A => n5330, B => DATAIN(28), S => n6013, Z => 
                           n4250);
   U1618 : MUX2_X1 port map( A => n5329, B => DATAIN(29), S => n6013, Z => 
                           n4251);
   U1619 : MUX2_X1 port map( A => n5328, B => DATAIN(30), S => n6013, Z => 
                           n4252);
   U1620 : MUX2_X1 port map( A => n5873, B => DATAIN(31), S => n6013, Z => 
                           n4253);
   U1621 : INV_X1 port map( A => ADD_WR(0), ZN => n6485);
   U1622 : MUX2_X1 port map( A => n5547, B => DATAIN(0), S => n6014, Z => n4350
                           );
   U1623 : MUX2_X1 port map( A => n5452, B => DATAIN(1), S => n6014, Z => n4351
                           );
   U1624 : MUX2_X1 port map( A => n5451, B => DATAIN(2), S => n6014, Z => n4352
                           );
   U1625 : MUX2_X1 port map( A => n5450, B => DATAIN(3), S => n6014, Z => n4353
                           );
   U1626 : MUX2_X1 port map( A => n5449, B => DATAIN(4), S => n6014, Z => n4354
                           );
   U1627 : MUX2_X1 port map( A => n5448, B => DATAIN(5), S => n6014, Z => n4355
                           );
   U1628 : MUX2_X1 port map( A => n5447, B => DATAIN(6), S => n6014, Z => n4356
                           );
   U1629 : MUX2_X1 port map( A => n5446, B => DATAIN(7), S => n6014, Z => n4357
                           );
   U1630 : MUX2_X1 port map( A => n5445, B => DATAIN(8), S => n6014, Z => n4358
                           );
   U1631 : MUX2_X1 port map( A => n5444, B => DATAIN(9), S => n6014, Z => n4359
                           );
   U1632 : MUX2_X1 port map( A => n5443, B => DATAIN(10), S => n6014, Z => 
                           n4360);
   U1633 : MUX2_X1 port map( A => n5442, B => DATAIN(11), S => n6014, Z => 
                           n4361);
   U1634 : MUX2_X1 port map( A => n5441, B => DATAIN(12), S => n6015, Z => 
                           n4362);
   U1635 : MUX2_X1 port map( A => n5440, B => DATAIN(13), S => n6015, Z => 
                           n4363);
   U1636 : MUX2_X1 port map( A => n5439, B => DATAIN(14), S => n6015, Z => 
                           n4364);
   U1637 : MUX2_X1 port map( A => n5438, B => DATAIN(15), S => n6015, Z => 
                           n4365);
   U1638 : MUX2_X1 port map( A => n5437, B => DATAIN(16), S => n6015, Z => 
                           n4366);
   U1639 : MUX2_X1 port map( A => n5436, B => DATAIN(17), S => n6015, Z => 
                           n4367);
   U1640 : MUX2_X1 port map( A => n5435, B => DATAIN(18), S => n6015, Z => 
                           n4368);
   U1641 : MUX2_X1 port map( A => n5434, B => DATAIN(19), S => n6015, Z => 
                           n4369);
   U1642 : MUX2_X1 port map( A => n5433, B => DATAIN(20), S => n6015, Z => 
                           n4370);
   U1643 : MUX2_X1 port map( A => n5432, B => DATAIN(21), S => n6015, Z => 
                           n4371);
   U1644 : MUX2_X1 port map( A => n5431, B => DATAIN(22), S => n6015, Z => 
                           n4372);
   U1645 : MUX2_X1 port map( A => n5430, B => DATAIN(23), S => n6015, Z => 
                           n4373);
   U1646 : MUX2_X1 port map( A => n5429, B => DATAIN(24), S => n6016, Z => 
                           n4374);
   U1647 : MUX2_X1 port map( A => n5428, B => DATAIN(25), S => n6016, Z => 
                           n4375);
   U1648 : MUX2_X1 port map( A => n5427, B => DATAIN(26), S => n6016, Z => 
                           n4376);
   U1649 : MUX2_X1 port map( A => n5426, B => DATAIN(27), S => n6016, Z => 
                           n4377);
   U1650 : MUX2_X1 port map( A => n5425, B => DATAIN(28), S => n6016, Z => 
                           n4378);
   U1651 : MUX2_X1 port map( A => n5424, B => DATAIN(29), S => n6016, Z => 
                           n4379);
   U1652 : MUX2_X1 port map( A => n5423, B => DATAIN(30), S => n6016, Z => 
                           n4380);
   U1653 : MUX2_X1 port map( A => n5422, B => DATAIN(31), S => n6016, Z => 
                           n4381);
   U1654 : INV_X1 port map( A => n2974, ZN => n6934);
   U1655 : MUX2_X1 port map( A => n5136, B => DATAIN(0), S => n6017, Z => n4414
                           );
   U1656 : INV_X1 port map( A => n2975, ZN => n6953);
   U1657 : MUX2_X1 port map( A => n5135, B => DATAIN(1), S => n6017, Z => n4415
                           );
   U1658 : INV_X1 port map( A => n2976, ZN => n6971);
   U1659 : MUX2_X1 port map( A => n5134, B => DATAIN(2), S => n6017, Z => n4416
                           );
   U1660 : INV_X1 port map( A => n2977, ZN => n6989);
   U1661 : MUX2_X1 port map( A => n5133, B => DATAIN(3), S => n6017, Z => n4417
                           );
   U1662 : INV_X1 port map( A => n2978, ZN => n7008);
   U1663 : MUX2_X1 port map( A => n5132, B => DATAIN(4), S => n6017, Z => n4418
                           );
   U1664 : INV_X1 port map( A => n2979, ZN => n7027);
   U1665 : MUX2_X1 port map( A => n5131, B => DATAIN(5), S => n6017, Z => n4419
                           );
   U1666 : INV_X1 port map( A => n2980, ZN => n7046);
   U1667 : MUX2_X1 port map( A => n5130, B => DATAIN(6), S => n6017, Z => n4420
                           );
   U1668 : INV_X1 port map( A => n2981, ZN => n7065);
   U1669 : MUX2_X1 port map( A => n5129, B => DATAIN(7), S => n6017, Z => n4421
                           );
   U1670 : INV_X1 port map( A => n2982, ZN => n7084);
   U1671 : MUX2_X1 port map( A => n5128, B => DATAIN(8), S => n6017, Z => n4422
                           );
   U1672 : INV_X1 port map( A => n3559, ZN => n7103);
   U1673 : MUX2_X1 port map( A => n5127, B => DATAIN(9), S => n6017, Z => n4423
                           );
   U1674 : INV_X1 port map( A => n3560, ZN => n7122);
   U1675 : MUX2_X1 port map( A => n5126, B => DATAIN(10), S => n6017, Z => 
                           n4424);
   U1676 : INV_X1 port map( A => n3561, ZN => n7141);
   U1677 : MUX2_X1 port map( A => n5125, B => DATAIN(11), S => n6017, Z => 
                           n4425);
   U1678 : INV_X1 port map( A => n3562, ZN => n7160);
   U1679 : MUX2_X1 port map( A => n5124, B => DATAIN(12), S => n6018, Z => 
                           n4426);
   U1680 : INV_X1 port map( A => n3563, ZN => n7179);
   U1681 : MUX2_X1 port map( A => n5123, B => DATAIN(13), S => n6018, Z => 
                           n4427);
   U1682 : INV_X1 port map( A => n3564, ZN => n7198);
   U1683 : MUX2_X1 port map( A => n5122, B => DATAIN(14), S => n6018, Z => 
                           n4428);
   U1684 : INV_X1 port map( A => n3565, ZN => n7217);
   U1685 : MUX2_X1 port map( A => n5121, B => DATAIN(15), S => n6018, Z => 
                           n4429);
   U1686 : INV_X1 port map( A => n3566, ZN => n7236);
   U1687 : MUX2_X1 port map( A => n5120, B => DATAIN(16), S => n6018, Z => 
                           n4430);
   U1688 : INV_X1 port map( A => n3567, ZN => n7255);
   U1689 : MUX2_X1 port map( A => n5119, B => DATAIN(17), S => n6018, Z => 
                           n4431);
   U1690 : INV_X1 port map( A => n3568, ZN => n7274);
   U1691 : MUX2_X1 port map( A => n5118, B => DATAIN(18), S => n6018, Z => 
                           n4432);
   U1692 : INV_X1 port map( A => n3569, ZN => n7293);
   U1693 : MUX2_X1 port map( A => n5117, B => DATAIN(19), S => n6018, Z => 
                           n4433);
   U1694 : INV_X1 port map( A => n3570, ZN => n7312);
   U1695 : MUX2_X1 port map( A => n5116, B => DATAIN(20), S => n6018, Z => 
                           n4434);
   U1696 : INV_X1 port map( A => n3571, ZN => n7331);
   U1697 : MUX2_X1 port map( A => n5115, B => DATAIN(21), S => n6018, Z => 
                           n4435);
   U1698 : INV_X1 port map( A => n3572, ZN => n7350);
   U1699 : MUX2_X1 port map( A => n5114, B => DATAIN(22), S => n6018, Z => 
                           n4436);
   U1700 : INV_X1 port map( A => n3573, ZN => n7369);
   U1701 : MUX2_X1 port map( A => n5113, B => DATAIN(23), S => n6018, Z => 
                           n4437);
   U1702 : INV_X1 port map( A => n3574, ZN => n7388);
   U1703 : MUX2_X1 port map( A => n5112, B => DATAIN(24), S => n6019, Z => 
                           n4438);
   U1704 : INV_X1 port map( A => n3575, ZN => n7407);
   U1705 : MUX2_X1 port map( A => n5111, B => DATAIN(25), S => n6019, Z => 
                           n4439);
   U1706 : INV_X1 port map( A => n3576, ZN => n7426);
   U1707 : MUX2_X1 port map( A => n5110, B => DATAIN(26), S => n6019, Z => 
                           n4440);
   U1708 : INV_X1 port map( A => n3577, ZN => n7445);
   U1709 : MUX2_X1 port map( A => n5109, B => DATAIN(27), S => n6019, Z => 
                           n4441);
   U1710 : INV_X1 port map( A => n3578, ZN => n7464);
   U1711 : MUX2_X1 port map( A => n5108, B => DATAIN(28), S => n6019, Z => 
                           n4442);
   U1712 : INV_X1 port map( A => n3579, ZN => n7483);
   U1713 : MUX2_X1 port map( A => n5107, B => DATAIN(29), S => n6019, Z => 
                           n4443);
   U1714 : INV_X1 port map( A => n3580, ZN => n7502);
   U1715 : MUX2_X1 port map( A => n5106, B => DATAIN(30), S => n6019, Z => 
                           n4444);
   U1716 : INV_X1 port map( A => n3581, ZN => n7532);
   U1717 : MUX2_X1 port map( A => n5105, B => DATAIN(31), S => n6019, Z => 
                           n4445);
   U1718 : MUX2_X1 port map( A => n5360, B => DATAIN(0), S => n6020, Z => n4542
                           );
   U1719 : MUX2_X1 port map( A => n5614, B => DATAIN(1), S => n6020, Z => n4543
                           );
   U1720 : MUX2_X1 port map( A => n5613, B => DATAIN(2), S => n6020, Z => n4544
                           );
   U1721 : MUX2_X1 port map( A => n5612, B => DATAIN(3), S => n6020, Z => n4545
                           );
   U1722 : MUX2_X1 port map( A => n5611, B => DATAIN(4), S => n6020, Z => n4546
                           );
   U1723 : MUX2_X1 port map( A => n5610, B => DATAIN(5), S => n6020, Z => n4547
                           );
   U1724 : MUX2_X1 port map( A => n5609, B => DATAIN(6), S => n6020, Z => n4548
                           );
   U1725 : MUX2_X1 port map( A => n5608, B => DATAIN(7), S => n6020, Z => n4549
                           );
   U1726 : MUX2_X1 port map( A => n5607, B => DATAIN(8), S => n6020, Z => n4550
                           );
   U1727 : MUX2_X1 port map( A => n5606, B => DATAIN(9), S => n6020, Z => n4551
                           );
   U1728 : MUX2_X1 port map( A => n5605, B => DATAIN(10), S => n6020, Z => 
                           n4552);
   U1729 : MUX2_X1 port map( A => n5604, B => DATAIN(11), S => n6020, Z => 
                           n4553);
   U1730 : MUX2_X1 port map( A => n5603, B => DATAIN(12), S => n6021, Z => 
                           n4554);
   U1731 : MUX2_X1 port map( A => n5602, B => DATAIN(13), S => n6021, Z => 
                           n4555);
   U1732 : MUX2_X1 port map( A => n5601, B => DATAIN(14), S => n6021, Z => 
                           n4556);
   U1733 : MUX2_X1 port map( A => n5600, B => DATAIN(15), S => n6021, Z => 
                           n4557);
   U1734 : MUX2_X1 port map( A => n5599, B => DATAIN(16), S => n6021, Z => 
                           n4558);
   U1735 : MUX2_X1 port map( A => n5598, B => DATAIN(17), S => n6021, Z => 
                           n4559);
   U1736 : MUX2_X1 port map( A => n5597, B => DATAIN(18), S => n6021, Z => 
                           n4560);
   U1737 : MUX2_X1 port map( A => n5596, B => DATAIN(19), S => n6021, Z => 
                           n4561);
   U1738 : MUX2_X1 port map( A => n5595, B => DATAIN(20), S => n6021, Z => 
                           n4562);
   U1739 : MUX2_X1 port map( A => n5594, B => DATAIN(21), S => n6021, Z => 
                           n4563);
   U1740 : MUX2_X1 port map( A => n5593, B => DATAIN(22), S => n6021, Z => 
                           n4564);
   U1741 : MUX2_X1 port map( A => n5592, B => DATAIN(23), S => n6021, Z => 
                           n4565);
   U1742 : MUX2_X1 port map( A => n5591, B => DATAIN(24), S => n6022, Z => 
                           n4566);
   U1743 : MUX2_X1 port map( A => n5590, B => DATAIN(25), S => n6022, Z => 
                           n4567);
   U1744 : MUX2_X1 port map( A => n5589, B => DATAIN(26), S => n6022, Z => 
                           n4568);
   U1745 : MUX2_X1 port map( A => n5588, B => DATAIN(27), S => n6022, Z => 
                           n4569);
   U1746 : MUX2_X1 port map( A => n5587, B => DATAIN(28), S => n6022, Z => 
                           n4570);
   U1747 : MUX2_X1 port map( A => n5586, B => DATAIN(29), S => n6022, Z => 
                           n4571);
   U1748 : MUX2_X1 port map( A => n5585, B => DATAIN(30), S => n6022, Z => 
                           n4572);
   U1749 : MUX2_X1 port map( A => n5584, B => DATAIN(31), S => n6022, Z => 
                           n4573);
   U1750 : MUX2_X1 port map( A => n5808, B => DATAIN(0), S => n6023, Z => n4126
                           );
   U1751 : MUX2_X1 port map( A => n5807, B => DATAIN(1), S => n6023, Z => n4127
                           );
   U1752 : MUX2_X1 port map( A => n5806, B => DATAIN(2), S => n6023, Z => n4128
                           );
   U1753 : MUX2_X1 port map( A => n5805, B => DATAIN(3), S => n6023, Z => n4129
                           );
   U1754 : MUX2_X1 port map( A => n5804, B => DATAIN(4), S => n6023, Z => n4130
                           );
   U1755 : MUX2_X1 port map( A => n5803, B => DATAIN(5), S => n6023, Z => n4131
                           );
   U1756 : MUX2_X1 port map( A => n5802, B => DATAIN(6), S => n6023, Z => n4132
                           );
   U1757 : MUX2_X1 port map( A => n5801, B => DATAIN(7), S => n6023, Z => n4133
                           );
   U1758 : MUX2_X1 port map( A => n5800, B => DATAIN(8), S => n6023, Z => n4134
                           );
   U1759 : MUX2_X1 port map( A => n5799, B => DATAIN(9), S => n6023, Z => n4135
                           );
   U1760 : MUX2_X1 port map( A => n5798, B => DATAIN(10), S => n6023, Z => 
                           n4136);
   U1761 : MUX2_X1 port map( A => n5797, B => DATAIN(11), S => n6023, Z => 
                           n4137);
   U1762 : MUX2_X1 port map( A => n5796, B => DATAIN(12), S => n6024, Z => 
                           n4138);
   U1763 : MUX2_X1 port map( A => n5795, B => DATAIN(13), S => n6024, Z => 
                           n4139);
   U1764 : MUX2_X1 port map( A => n5794, B => DATAIN(14), S => n6024, Z => 
                           n4140);
   U1765 : MUX2_X1 port map( A => n5793, B => DATAIN(15), S => n6024, Z => 
                           n4141);
   U1766 : MUX2_X1 port map( A => n5792, B => DATAIN(16), S => n6024, Z => 
                           n4142);
   U1767 : MUX2_X1 port map( A => n5791, B => DATAIN(17), S => n6024, Z => 
                           n4143);
   U1768 : MUX2_X1 port map( A => n5790, B => DATAIN(18), S => n6024, Z => 
                           n4144);
   U1769 : MUX2_X1 port map( A => n5789, B => DATAIN(19), S => n6024, Z => 
                           n4145);
   U1770 : MUX2_X1 port map( A => n5788, B => DATAIN(20), S => n6024, Z => 
                           n4146);
   U1771 : MUX2_X1 port map( A => n5787, B => DATAIN(21), S => n6024, Z => 
                           n4147);
   U1772 : MUX2_X1 port map( A => n5786, B => DATAIN(22), S => n6024, Z => 
                           n4148);
   U1773 : MUX2_X1 port map( A => n5785, B => DATAIN(23), S => n6024, Z => 
                           n4149);
   U1774 : MUX2_X1 port map( A => n5784, B => DATAIN(24), S => n6025, Z => 
                           n4150);
   U1775 : MUX2_X1 port map( A => n5783, B => DATAIN(25), S => n6025, Z => 
                           n4151);
   U1776 : MUX2_X1 port map( A => n5782, B => DATAIN(26), S => n6025, Z => 
                           n4152);
   U1777 : MUX2_X1 port map( A => n5781, B => DATAIN(27), S => n6025, Z => 
                           n4153);
   U1778 : MUX2_X1 port map( A => n5780, B => DATAIN(28), S => n6025, Z => 
                           n4154);
   U1779 : MUX2_X1 port map( A => n5779, B => DATAIN(29), S => n6025, Z => 
                           n4155);
   U1780 : MUX2_X1 port map( A => n5778, B => DATAIN(30), S => n6025, Z => 
                           n4156);
   U1781 : MUX2_X1 port map( A => n5777, B => DATAIN(31), S => n6025, Z => 
                           n4157);
   U1782 : MUX2_X1 port map( A => n5646, B => DATAIN(0), S => n6026, Z => n4190
                           );
   U1783 : MUX2_X1 port map( A => n5645, B => DATAIN(1), S => n6026, Z => n4191
                           );
   U1784 : MUX2_X1 port map( A => n5644, B => DATAIN(2), S => n6026, Z => n4192
                           );
   U1785 : MUX2_X1 port map( A => n5643, B => DATAIN(3), S => n6026, Z => n4193
                           );
   U1786 : MUX2_X1 port map( A => n5642, B => DATAIN(4), S => n6026, Z => n4194
                           );
   U1787 : MUX2_X1 port map( A => n5641, B => DATAIN(5), S => n6026, Z => n4195
                           );
   U1788 : MUX2_X1 port map( A => n5640, B => DATAIN(6), S => n6026, Z => n4196
                           );
   U1789 : MUX2_X1 port map( A => n5639, B => DATAIN(7), S => n6026, Z => n4197
                           );
   U1790 : MUX2_X1 port map( A => n5638, B => DATAIN(8), S => n6026, Z => n4198
                           );
   U1791 : MUX2_X1 port map( A => n5637, B => DATAIN(9), S => n6026, Z => n4199
                           );
   U1792 : MUX2_X1 port map( A => n5636, B => DATAIN(10), S => n6026, Z => 
                           n4200);
   U1793 : MUX2_X1 port map( A => n5635, B => DATAIN(11), S => n6026, Z => 
                           n4201);
   U1794 : MUX2_X1 port map( A => n5634, B => DATAIN(12), S => n6027, Z => 
                           n4202);
   U1795 : MUX2_X1 port map( A => n5633, B => DATAIN(13), S => n6027, Z => 
                           n4203);
   U1796 : MUX2_X1 port map( A => n5632, B => DATAIN(14), S => n6027, Z => 
                           n4204);
   U1797 : MUX2_X1 port map( A => n5631, B => DATAIN(15), S => n6027, Z => 
                           n4205);
   U1798 : MUX2_X1 port map( A => n5630, B => DATAIN(16), S => n6027, Z => 
                           n4206);
   U1799 : MUX2_X1 port map( A => n5629, B => DATAIN(17), S => n6027, Z => 
                           n4207);
   U1800 : MUX2_X1 port map( A => n5628, B => DATAIN(18), S => n6027, Z => 
                           n4208);
   U1801 : MUX2_X1 port map( A => n5627, B => DATAIN(19), S => n6027, Z => 
                           n4209);
   U1802 : MUX2_X1 port map( A => n5626, B => DATAIN(20), S => n6027, Z => 
                           n4210);
   U1803 : MUX2_X1 port map( A => n5625, B => DATAIN(21), S => n6027, Z => 
                           n4211);
   U1804 : MUX2_X1 port map( A => n5624, B => DATAIN(22), S => n6027, Z => 
                           n4212);
   U1805 : MUX2_X1 port map( A => n5623, B => DATAIN(23), S => n6027, Z => 
                           n4213);
   U1806 : MUX2_X1 port map( A => n5622, B => DATAIN(24), S => n6028, Z => 
                           n4214);
   U1807 : MUX2_X1 port map( A => n5621, B => DATAIN(25), S => n6028, Z => 
                           n4215);
   U1808 : MUX2_X1 port map( A => n5620, B => DATAIN(26), S => n6028, Z => 
                           n4216);
   U1809 : MUX2_X1 port map( A => n5619, B => DATAIN(27), S => n6028, Z => 
                           n4217);
   U1810 : MUX2_X1 port map( A => n5618, B => DATAIN(28), S => n6028, Z => 
                           n4218);
   U1811 : MUX2_X1 port map( A => n5617, B => DATAIN(29), S => n6028, Z => 
                           n4219);
   U1812 : MUX2_X1 port map( A => n5616, B => DATAIN(30), S => n6028, Z => 
                           n4220);
   U1813 : MUX2_X1 port map( A => n5615, B => DATAIN(31), S => n6028, Z => 
                           n4221);
   U1814 : MUX2_X1 port map( A => n5359, B => DATAIN(0), S => n6029, Z => n4446
                           );
   U1815 : INV_X1 port map( A => n2943, ZN => n6951);
   U1816 : MUX2_X1 port map( A => n5202, B => DATAIN(1), S => n6029, Z => n4447
                           );
   U1817 : INV_X1 port map( A => n2944, ZN => n6969);
   U1818 : MUX2_X1 port map( A => n5201, B => DATAIN(2), S => n6029, Z => n4448
                           );
   U1819 : INV_X1 port map( A => n2945, ZN => n6987);
   U1820 : MUX2_X1 port map( A => n5200, B => DATAIN(3), S => n6029, Z => n4449
                           );
   U1821 : INV_X1 port map( A => n2946, ZN => n7006);
   U1822 : MUX2_X1 port map( A => n5199, B => DATAIN(4), S => n6029, Z => n4450
                           );
   U1823 : INV_X1 port map( A => n2947, ZN => n7025);
   U1824 : MUX2_X1 port map( A => n5198, B => DATAIN(5), S => n6029, Z => n4451
                           );
   U1825 : INV_X1 port map( A => n2948, ZN => n7044);
   U1826 : MUX2_X1 port map( A => n5197, B => DATAIN(6), S => n6029, Z => n4452
                           );
   U1827 : INV_X1 port map( A => n2949, ZN => n7063);
   U1828 : MUX2_X1 port map( A => n5196, B => DATAIN(7), S => n6029, Z => n4453
                           );
   U1829 : INV_X1 port map( A => n2950, ZN => n7082);
   U1830 : MUX2_X1 port map( A => n5195, B => DATAIN(8), S => n6029, Z => n4454
                           );
   U1831 : INV_X1 port map( A => n2951, ZN => n7101);
   U1832 : MUX2_X1 port map( A => n5194, B => DATAIN(9), S => n6029, Z => n4455
                           );
   U1833 : INV_X1 port map( A => n2952, ZN => n7120);
   U1834 : MUX2_X1 port map( A => n5193, B => DATAIN(10), S => n6029, Z => 
                           n4456);
   U1835 : INV_X1 port map( A => n2953, ZN => n7139);
   U1836 : MUX2_X1 port map( A => n5192, B => DATAIN(11), S => n6029, Z => 
                           n4457);
   U1837 : INV_X1 port map( A => n2954, ZN => n7158);
   U1838 : MUX2_X1 port map( A => n5191, B => DATAIN(12), S => n6030, Z => 
                           n4458);
   U1839 : INV_X1 port map( A => n2955, ZN => n7177);
   U1840 : MUX2_X1 port map( A => n5190, B => DATAIN(13), S => n6030, Z => 
                           n4459);
   U1841 : INV_X1 port map( A => n2956, ZN => n7196);
   U1842 : MUX2_X1 port map( A => n5189, B => DATAIN(14), S => n6030, Z => 
                           n4460);
   U1843 : INV_X1 port map( A => n2957, ZN => n7215);
   U1844 : MUX2_X1 port map( A => n5188, B => DATAIN(15), S => n6030, Z => 
                           n4461);
   U1845 : INV_X1 port map( A => n2958, ZN => n7234);
   U1846 : MUX2_X1 port map( A => n5187, B => DATAIN(16), S => n6030, Z => 
                           n4462);
   U1847 : INV_X1 port map( A => n2959, ZN => n7253);
   U1848 : MUX2_X1 port map( A => n5186, B => DATAIN(17), S => n6030, Z => 
                           n4463);
   U1849 : INV_X1 port map( A => n2960, ZN => n7272);
   U1850 : MUX2_X1 port map( A => n5185, B => DATAIN(18), S => n6030, Z => 
                           n4464);
   U1851 : INV_X1 port map( A => n2961, ZN => n7291);
   U1852 : MUX2_X1 port map( A => n5184, B => DATAIN(19), S => n6030, Z => 
                           n4465);
   U1853 : INV_X1 port map( A => n2962, ZN => n7310);
   U1854 : MUX2_X1 port map( A => n5183, B => DATAIN(20), S => n6030, Z => 
                           n4466);
   U1855 : INV_X1 port map( A => n2963, ZN => n7329);
   U1856 : MUX2_X1 port map( A => n5182, B => DATAIN(21), S => n6030, Z => 
                           n4467);
   U1857 : INV_X1 port map( A => n2964, ZN => n7348);
   U1858 : MUX2_X1 port map( A => n5181, B => DATAIN(22), S => n6030, Z => 
                           n4468);
   U1859 : INV_X1 port map( A => n2965, ZN => n7367);
   U1860 : MUX2_X1 port map( A => n5180, B => DATAIN(23), S => n6030, Z => 
                           n4469);
   U1861 : INV_X1 port map( A => n2966, ZN => n7386);
   U1862 : MUX2_X1 port map( A => n5179, B => DATAIN(24), S => n6031, Z => 
                           n4470);
   U1863 : INV_X1 port map( A => n2967, ZN => n7405);
   U1864 : MUX2_X1 port map( A => n5178, B => DATAIN(25), S => n6031, Z => 
                           n4471);
   U1865 : INV_X1 port map( A => n2968, ZN => n7424);
   U1866 : MUX2_X1 port map( A => n5177, B => DATAIN(26), S => n6031, Z => 
                           n4472);
   U1867 : INV_X1 port map( A => n2969, ZN => n7443);
   U1868 : MUX2_X1 port map( A => n5176, B => DATAIN(27), S => n6031, Z => 
                           n4473);
   U1869 : INV_X1 port map( A => n2970, ZN => n7462);
   U1870 : MUX2_X1 port map( A => n5175, B => DATAIN(28), S => n6031, Z => 
                           n4474);
   U1871 : INV_X1 port map( A => n2971, ZN => n7481);
   U1872 : MUX2_X1 port map( A => n5174, B => DATAIN(29), S => n6031, Z => 
                           n4475);
   U1873 : INV_X1 port map( A => n2972, ZN => n7500);
   U1874 : MUX2_X1 port map( A => n5173, B => DATAIN(30), S => n6031, Z => 
                           n4476);
   U1875 : INV_X1 port map( A => n2973, ZN => n7526);
   U1876 : MUX2_X1 port map( A => n5172, B => DATAIN(31), S => n6031, Z => 
                           n4477);
   U1877 : NAND2_X1 port map( A1 => n4606, A2 => n4611, ZN => n6483);
   U1878 : INV_X1 port map( A => n6483, ZN => n6484);
   U1879 : OAI22_X1 port map( A1 => n6034, A2 => n5908, B1 => n6339, B2 => 
                           n6483, ZN => n4574);
   U1880 : OAI22_X1 port map( A1 => n6034, A2 => n5879, B1 => n6341, B2 => 
                           n6483, ZN => n4575);
   U1881 : OAI22_X1 port map( A1 => n6034, A2 => n5878, B1 => n6343, B2 => 
                           n6483, ZN => n4576);
   U1882 : OAI22_X1 port map( A1 => n6034, A2 => n5877, B1 => n6345, B2 => 
                           n6483, ZN => n4577);
   U1883 : MUX2_X1 port map( A => n5514, B => DATAIN(4), S => n6034, Z => n4578
                           );
   U1884 : MUX2_X1 port map( A => n5513, B => DATAIN(5), S => n6034, Z => n4579
                           );
   U1885 : MUX2_X1 port map( A => n5512, B => DATAIN(6), S => n6034, Z => n4580
                           );
   U1886 : MUX2_X1 port map( A => n5511, B => DATAIN(7), S => n6034, Z => n4581
                           );
   U1887 : MUX2_X1 port map( A => n5510, B => DATAIN(8), S => n6033, Z => n4582
                           );
   U1888 : MUX2_X1 port map( A => n5509, B => DATAIN(9), S => n6033, Z => n4583
                           );
   U1889 : MUX2_X1 port map( A => n5508, B => DATAIN(10), S => n6033, Z => 
                           n4584);
   U1890 : MUX2_X1 port map( A => n5507, B => DATAIN(11), S => n6033, Z => 
                           n4585);
   U1891 : MUX2_X1 port map( A => n5506, B => DATAIN(12), S => n6033, Z => 
                           n4586);
   U1892 : MUX2_X1 port map( A => n5505, B => DATAIN(13), S => n6033, Z => 
                           n4587);
   U1893 : MUX2_X1 port map( A => n5504, B => DATAIN(14), S => n6033, Z => 
                           n4588);
   U1894 : MUX2_X1 port map( A => n5503, B => DATAIN(15), S => n6033, Z => 
                           n4589);
   U1895 : MUX2_X1 port map( A => n5502, B => DATAIN(16), S => n6033, Z => 
                           n4590);
   U1896 : MUX2_X1 port map( A => n5501, B => DATAIN(17), S => n6033, Z => 
                           n4591);
   U1897 : MUX2_X1 port map( A => n5500, B => DATAIN(18), S => n6033, Z => 
                           n4592);
   U1898 : MUX2_X1 port map( A => n5499, B => DATAIN(19), S => n6033, Z => 
                           n4593);
   U1899 : MUX2_X1 port map( A => n5498, B => DATAIN(20), S => n6032, Z => 
                           n4594);
   U1900 : MUX2_X1 port map( A => n5497, B => DATAIN(21), S => n6032, Z => 
                           n4595);
   U1901 : MUX2_X1 port map( A => n5496, B => DATAIN(22), S => n6032, Z => 
                           n4596);
   U1902 : MUX2_X1 port map( A => n5495, B => DATAIN(23), S => n6032, Z => 
                           n4597);
   U1903 : MUX2_X1 port map( A => n5494, B => DATAIN(24), S => n6032, Z => 
                           n4598);
   U1904 : MUX2_X1 port map( A => n5493, B => DATAIN(25), S => n6032, Z => 
                           n4599);
   U1905 : MUX2_X1 port map( A => n5492, B => DATAIN(26), S => n6032, Z => 
                           n4600);
   U1906 : MUX2_X1 port map( A => n5491, B => DATAIN(27), S => n6032, Z => 
                           n4601);
   U1907 : MUX2_X1 port map( A => n5490, B => DATAIN(28), S => n6032, Z => 
                           n4602);
   U1908 : MUX2_X1 port map( A => n5489, B => DATAIN(29), S => n6032, Z => 
                           n4603);
   U1909 : MUX2_X1 port map( A => n5488, B => DATAIN(30), S => n6032, Z => 
                           n4604);
   U1910 : MUX2_X1 port map( A => n5487, B => DATAIN(31), S => n6032, Z => 
                           n4605);
   U1911 : MUX2_X1 port map( A => n5840, B => DATAIN(0), S => n6035, Z => n4318
                           );
   U1912 : MUX2_X1 port map( A => n5839, B => DATAIN(1), S => n6035, Z => n4319
                           );
   U1913 : MUX2_X1 port map( A => n5838, B => DATAIN(2), S => n6035, Z => n4320
                           );
   U1914 : MUX2_X1 port map( A => n5837, B => DATAIN(3), S => n6035, Z => n4321
                           );
   U1915 : MUX2_X1 port map( A => n5836, B => DATAIN(4), S => n6035, Z => n4322
                           );
   U1916 : MUX2_X1 port map( A => n5835, B => DATAIN(5), S => n6035, Z => n4323
                           );
   U1917 : MUX2_X1 port map( A => n5834, B => DATAIN(6), S => n6035, Z => n4324
                           );
   U1918 : MUX2_X1 port map( A => n5833, B => DATAIN(7), S => n6035, Z => n4325
                           );
   U1919 : MUX2_X1 port map( A => n5832, B => DATAIN(8), S => n6035, Z => n4326
                           );
   U1920 : MUX2_X1 port map( A => n5831, B => DATAIN(9), S => n6035, Z => n4327
                           );
   U1921 : MUX2_X1 port map( A => n5830, B => DATAIN(10), S => n6035, Z => 
                           n4328);
   U1922 : MUX2_X1 port map( A => n5829, B => DATAIN(11), S => n6035, Z => 
                           n4329);
   U1923 : MUX2_X1 port map( A => n5828, B => DATAIN(12), S => n6036, Z => 
                           n4330);
   U1924 : MUX2_X1 port map( A => n5827, B => DATAIN(13), S => n6036, Z => 
                           n4331);
   U1925 : MUX2_X1 port map( A => n5826, B => DATAIN(14), S => n6036, Z => 
                           n4332);
   U1926 : MUX2_X1 port map( A => n5825, B => DATAIN(15), S => n6036, Z => 
                           n4333);
   U1927 : MUX2_X1 port map( A => n5824, B => DATAIN(16), S => n6036, Z => 
                           n4334);
   U1928 : MUX2_X1 port map( A => n5823, B => DATAIN(17), S => n6036, Z => 
                           n4335);
   U1929 : MUX2_X1 port map( A => n5822, B => DATAIN(18), S => n6036, Z => 
                           n4336);
   U1930 : MUX2_X1 port map( A => n5821, B => DATAIN(19), S => n6036, Z => 
                           n4337);
   U1931 : MUX2_X1 port map( A => n5820, B => DATAIN(20), S => n6036, Z => 
                           n4338);
   U1932 : MUX2_X1 port map( A => n5819, B => DATAIN(21), S => n6036, Z => 
                           n4339);
   U1933 : MUX2_X1 port map( A => n5818, B => DATAIN(22), S => n6036, Z => 
                           n4340);
   U1934 : MUX2_X1 port map( A => n5817, B => DATAIN(23), S => n6036, Z => 
                           n4341);
   U1935 : MUX2_X1 port map( A => n5816, B => DATAIN(24), S => n6037, Z => 
                           n4342);
   U1936 : MUX2_X1 port map( A => n5815, B => DATAIN(25), S => n6037, Z => 
                           n4343);
   U1937 : MUX2_X1 port map( A => n5814, B => DATAIN(26), S => n6037, Z => 
                           n4344);
   U1938 : MUX2_X1 port map( A => n5813, B => DATAIN(27), S => n6037, Z => 
                           n4345);
   U1939 : MUX2_X1 port map( A => n5812, B => DATAIN(28), S => n6037, Z => 
                           n4346);
   U1940 : MUX2_X1 port map( A => n5811, B => DATAIN(29), S => n6037, Z => 
                           n4347);
   U1941 : MUX2_X1 port map( A => n5810, B => DATAIN(30), S => n6037, Z => 
                           n4348);
   U1942 : MUX2_X1 port map( A => n5809, B => DATAIN(31), S => n6037, Z => 
                           n4349);
   U1943 : INV_X1 port map( A => n2252, ZN => n6942);
   U1944 : MUX2_X1 port map( A => n5233, B => DATAIN(0), S => n6038, Z => n4382
                           );
   U1945 : MUX2_X1 port map( A => n5390, B => DATAIN(1), S => n6038, Z => n4383
                           );
   U1946 : MUX2_X1 port map( A => n5389, B => DATAIN(2), S => n6038, Z => n4384
                           );
   U1947 : MUX2_X1 port map( A => n5388, B => DATAIN(3), S => n6038, Z => n4385
                           );
   U1948 : MUX2_X1 port map( A => n5387, B => DATAIN(4), S => n6038, Z => n4386
                           );
   U1949 : MUX2_X1 port map( A => n5386, B => DATAIN(5), S => n6038, Z => n4387
                           );
   U1950 : MUX2_X1 port map( A => n5385, B => DATAIN(6), S => n6038, Z => n4388
                           );
   U1951 : MUX2_X1 port map( A => n5384, B => DATAIN(7), S => n6038, Z => n4389
                           );
   U1952 : MUX2_X1 port map( A => n5383, B => DATAIN(8), S => n6038, Z => n4390
                           );
   U1953 : MUX2_X1 port map( A => n5382, B => DATAIN(9), S => n6038, Z => n4391
                           );
   U1954 : MUX2_X1 port map( A => n5381, B => DATAIN(10), S => n6038, Z => 
                           n4392);
   U1955 : MUX2_X1 port map( A => n5380, B => DATAIN(11), S => n6038, Z => 
                           n4393);
   U1956 : MUX2_X1 port map( A => n5379, B => DATAIN(12), S => n6039, Z => 
                           n4394);
   U1957 : MUX2_X1 port map( A => n5378, B => DATAIN(13), S => n6039, Z => 
                           n4395);
   U1958 : MUX2_X1 port map( A => n5377, B => DATAIN(14), S => n6039, Z => 
                           n4396);
   U1959 : MUX2_X1 port map( A => n5376, B => DATAIN(15), S => n6039, Z => 
                           n4397);
   U1960 : MUX2_X1 port map( A => n5375, B => DATAIN(16), S => n6039, Z => 
                           n4398);
   U1961 : MUX2_X1 port map( A => n5374, B => DATAIN(17), S => n6039, Z => 
                           n4399);
   U1962 : MUX2_X1 port map( A => n5373, B => DATAIN(18), S => n6039, Z => 
                           n4400);
   U1963 : MUX2_X1 port map( A => n5372, B => DATAIN(19), S => n6039, Z => 
                           n4401);
   U1964 : MUX2_X1 port map( A => n5371, B => DATAIN(20), S => n6039, Z => 
                           n4402);
   U1965 : MUX2_X1 port map( A => n5370, B => DATAIN(21), S => n6039, Z => 
                           n4403);
   U1966 : MUX2_X1 port map( A => n5369, B => DATAIN(22), S => n6039, Z => 
                           n4404);
   U1967 : MUX2_X1 port map( A => n5368, B => DATAIN(23), S => n6039, Z => 
                           n4405);
   U1968 : MUX2_X1 port map( A => n5367, B => DATAIN(24), S => n6040, Z => 
                           n4406);
   U1969 : MUX2_X1 port map( A => n5366, B => DATAIN(25), S => n6040, Z => 
                           n4407);
   U1970 : MUX2_X1 port map( A => n5365, B => DATAIN(26), S => n6040, Z => 
                           n4408);
   U1971 : MUX2_X1 port map( A => n5364, B => DATAIN(27), S => n6040, Z => 
                           n4409);
   U1972 : MUX2_X1 port map( A => n5363, B => DATAIN(28), S => n6040, Z => 
                           n4410);
   U1973 : MUX2_X1 port map( A => n5362, B => DATAIN(29), S => n6040, Z => 
                           n4411);
   U1974 : MUX2_X1 port map( A => n5361, B => DATAIN(30), S => n6040, Z => 
                           n4412);
   U1975 : INV_X1 port map( A => n2283, ZN => n7540);
   U1976 : MUX2_X1 port map( A => n5168, B => DATAIN(31), S => n6040, Z => 
                           n4413);
   U1977 : MUX2_X1 port map( A => n5648, B => DATAIN(0), S => n6041, Z => n4478
                           );
   U1978 : MUX2_X1 port map( A => n5679, B => DATAIN(1), S => n6041, Z => n4479
                           );
   U1979 : MUX2_X1 port map( A => n5678, B => DATAIN(2), S => n6041, Z => n4480
                           );
   U1980 : MUX2_X1 port map( A => n5677, B => DATAIN(3), S => n6041, Z => n4481
                           );
   U1981 : MUX2_X1 port map( A => n5676, B => DATAIN(4), S => n6041, Z => n4482
                           );
   U1982 : MUX2_X1 port map( A => n5675, B => DATAIN(5), S => n6041, Z => n4483
                           );
   U1983 : MUX2_X1 port map( A => n5674, B => DATAIN(6), S => n6041, Z => n4484
                           );
   U1984 : MUX2_X1 port map( A => n5673, B => DATAIN(7), S => n6041, Z => n4485
                           );
   U1985 : MUX2_X1 port map( A => n5672, B => DATAIN(8), S => n6041, Z => n4486
                           );
   U1986 : MUX2_X1 port map( A => n5671, B => DATAIN(9), S => n6041, Z => n4487
                           );
   U1987 : MUX2_X1 port map( A => n5670, B => DATAIN(10), S => n6041, Z => 
                           n4488);
   U1988 : MUX2_X1 port map( A => n5669, B => DATAIN(11), S => n6041, Z => 
                           n4489);
   U1989 : MUX2_X1 port map( A => n5668, B => DATAIN(12), S => n6042, Z => 
                           n4490);
   U1990 : MUX2_X1 port map( A => n5667, B => DATAIN(13), S => n6042, Z => 
                           n4491);
   U1991 : MUX2_X1 port map( A => n5666, B => DATAIN(14), S => n6042, Z => 
                           n4492);
   U1992 : MUX2_X1 port map( A => n5665, B => DATAIN(15), S => n6042, Z => 
                           n4493);
   U1993 : MUX2_X1 port map( A => n5664, B => DATAIN(16), S => n6042, Z => 
                           n4494);
   U1994 : MUX2_X1 port map( A => n5663, B => DATAIN(17), S => n6042, Z => 
                           n4495);
   U1995 : MUX2_X1 port map( A => n5662, B => DATAIN(18), S => n6042, Z => 
                           n4496);
   U1996 : MUX2_X1 port map( A => n5661, B => DATAIN(19), S => n6042, Z => 
                           n4497);
   U1997 : MUX2_X1 port map( A => n5660, B => DATAIN(20), S => n6042, Z => 
                           n4498);
   U1998 : MUX2_X1 port map( A => n5659, B => DATAIN(21), S => n6042, Z => 
                           n4499);
   U1999 : MUX2_X1 port map( A => n5658, B => DATAIN(22), S => n6042, Z => 
                           n4500);
   U2000 : MUX2_X1 port map( A => n5657, B => DATAIN(23), S => n6042, Z => 
                           n4501);
   U2001 : MUX2_X1 port map( A => n5656, B => DATAIN(24), S => n6043, Z => 
                           n4502);
   U2002 : MUX2_X1 port map( A => n5655, B => DATAIN(25), S => n6043, Z => 
                           n4503);
   U2003 : MUX2_X1 port map( A => n5654, B => DATAIN(26), S => n6043, Z => 
                           n4504);
   U2004 : MUX2_X1 port map( A => n5653, B => DATAIN(27), S => n6043, Z => 
                           n4505);
   U2005 : MUX2_X1 port map( A => n5652, B => DATAIN(28), S => n6043, Z => 
                           n4506);
   U2006 : MUX2_X1 port map( A => n5651, B => DATAIN(29), S => n6043, Z => 
                           n4507);
   U2007 : MUX2_X1 port map( A => n5650, B => DATAIN(30), S => n6043, Z => 
                           n4508);
   U2008 : MUX2_X1 port map( A => n5649, B => DATAIN(31), S => n6043, Z => 
                           n4509);
   U2009 : MUX2_X1 port map( A => n5876, B => DATAIN(0), S => n6044, Z => n4286
                           );
   U2010 : MUX2_X1 port map( A => n5327, B => DATAIN(1), S => n6044, Z => n4287
                           );
   U2011 : MUX2_X1 port map( A => n5326, B => DATAIN(2), S => n6044, Z => n4288
                           );
   U2012 : MUX2_X1 port map( A => n5325, B => DATAIN(3), S => n6044, Z => n4289
                           );
   U2013 : MUX2_X1 port map( A => n5324, B => DATAIN(4), S => n6044, Z => n4290
                           );
   U2014 : MUX2_X1 port map( A => n5323, B => DATAIN(5), S => n6044, Z => n4291
                           );
   U2015 : MUX2_X1 port map( A => n5322, B => DATAIN(6), S => n6044, Z => n4292
                           );
   U2016 : MUX2_X1 port map( A => n5321, B => DATAIN(7), S => n6044, Z => n4293
                           );
   U2017 : MUX2_X1 port map( A => n5320, B => DATAIN(8), S => n6044, Z => n4294
                           );
   U2018 : MUX2_X1 port map( A => n5319, B => DATAIN(9), S => n6044, Z => n4295
                           );
   U2019 : MUX2_X1 port map( A => n5318, B => DATAIN(10), S => n6044, Z => 
                           n4296);
   U2020 : MUX2_X1 port map( A => n5317, B => DATAIN(11), S => n6044, Z => 
                           n4297);
   U2021 : MUX2_X1 port map( A => n5316, B => DATAIN(12), S => n6045, Z => 
                           n4298);
   U2022 : MUX2_X1 port map( A => n5315, B => DATAIN(13), S => n6045, Z => 
                           n4299);
   U2023 : MUX2_X1 port map( A => n5314, B => DATAIN(14), S => n6045, Z => 
                           n4300);
   U2024 : MUX2_X1 port map( A => n5313, B => DATAIN(15), S => n6045, Z => 
                           n4301);
   U2025 : MUX2_X1 port map( A => n5312, B => DATAIN(16), S => n6045, Z => 
                           n4302);
   U2026 : MUX2_X1 port map( A => n5311, B => DATAIN(17), S => n6045, Z => 
                           n4303);
   U2027 : MUX2_X1 port map( A => n5310, B => DATAIN(18), S => n6045, Z => 
                           n4304);
   U2028 : MUX2_X1 port map( A => n5309, B => DATAIN(19), S => n6045, Z => 
                           n4305);
   U2029 : MUX2_X1 port map( A => n5308, B => DATAIN(20), S => n6045, Z => 
                           n4306);
   U2030 : MUX2_X1 port map( A => n5307, B => DATAIN(21), S => n6045, Z => 
                           n4307);
   U2031 : MUX2_X1 port map( A => n5306, B => DATAIN(22), S => n6045, Z => 
                           n4308);
   U2032 : MUX2_X1 port map( A => n5305, B => DATAIN(23), S => n6045, Z => 
                           n4309);
   U2033 : MUX2_X1 port map( A => n5304, B => DATAIN(24), S => n6046, Z => 
                           n4310);
   U2034 : MUX2_X1 port map( A => n5303, B => DATAIN(25), S => n6046, Z => 
                           n4311);
   U2035 : MUX2_X1 port map( A => n5302, B => DATAIN(26), S => n6046, Z => 
                           n4312);
   U2036 : MUX2_X1 port map( A => n5301, B => DATAIN(27), S => n6046, Z => 
                           n4313);
   U2037 : MUX2_X1 port map( A => n5300, B => DATAIN(28), S => n6046, Z => 
                           n4314);
   U2038 : MUX2_X1 port map( A => n5299, B => DATAIN(29), S => n6046, Z => 
                           n4315);
   U2039 : MUX2_X1 port map( A => n5298, B => DATAIN(30), S => n6046, Z => 
                           n4316);
   U2040 : MUX2_X1 port map( A => n5875, B => DATAIN(31), S => n6046, Z => 
                           n4317);
   U2041 : MUX2_X1 port map( A => n5546, B => DATAIN(0), S => n6047, Z => n4510
                           );
   U2042 : MUX2_X1 port map( A => n5421, B => DATAIN(1), S => n6047, Z => n4511
                           );
   U2043 : MUX2_X1 port map( A => n5420, B => DATAIN(2), S => n6047, Z => n4512
                           );
   U2044 : MUX2_X1 port map( A => n5419, B => DATAIN(3), S => n6047, Z => n4513
                           );
   U2045 : MUX2_X1 port map( A => n5418, B => DATAIN(4), S => n6047, Z => n4514
                           );
   U2046 : MUX2_X1 port map( A => n5417, B => DATAIN(5), S => n6047, Z => n4515
                           );
   U2047 : MUX2_X1 port map( A => n5416, B => DATAIN(6), S => n6047, Z => n4516
                           );
   U2048 : MUX2_X1 port map( A => n5415, B => DATAIN(7), S => n6047, Z => n4517
                           );
   U2049 : MUX2_X1 port map( A => n5414, B => DATAIN(8), S => n6047, Z => n4518
                           );
   U2050 : MUX2_X1 port map( A => n5413, B => DATAIN(9), S => n6047, Z => n4519
                           );
   U2051 : MUX2_X1 port map( A => n5412, B => DATAIN(10), S => n6047, Z => 
                           n4520);
   U2052 : MUX2_X1 port map( A => n5411, B => DATAIN(11), S => n6047, Z => 
                           n4521);
   U2053 : MUX2_X1 port map( A => n5410, B => DATAIN(12), S => n6048, Z => 
                           n4522);
   U2054 : MUX2_X1 port map( A => n5409, B => DATAIN(13), S => n6048, Z => 
                           n4523);
   U2055 : MUX2_X1 port map( A => n5408, B => DATAIN(14), S => n6048, Z => 
                           n4524);
   U2056 : MUX2_X1 port map( A => n5407, B => DATAIN(15), S => n6048, Z => 
                           n4525);
   U2057 : MUX2_X1 port map( A => n5406, B => DATAIN(16), S => n6048, Z => 
                           n4526);
   U2058 : MUX2_X1 port map( A => n5405, B => DATAIN(17), S => n6048, Z => 
                           n4527);
   U2059 : MUX2_X1 port map( A => n5404, B => DATAIN(18), S => n6048, Z => 
                           n4528);
   U2060 : MUX2_X1 port map( A => n5403, B => DATAIN(19), S => n6048, Z => 
                           n4529);
   U2061 : MUX2_X1 port map( A => n5402, B => DATAIN(20), S => n6048, Z => 
                           n4530);
   U2062 : MUX2_X1 port map( A => n5401, B => DATAIN(21), S => n6048, Z => 
                           n4531);
   U2063 : MUX2_X1 port map( A => n5400, B => DATAIN(22), S => n6048, Z => 
                           n4532);
   U2064 : MUX2_X1 port map( A => n5399, B => DATAIN(23), S => n6048, Z => 
                           n4533);
   U2065 : MUX2_X1 port map( A => n5398, B => DATAIN(24), S => n6049, Z => 
                           n4534);
   U2066 : MUX2_X1 port map( A => n5397, B => DATAIN(25), S => n6049, Z => 
                           n4535);
   U2067 : MUX2_X1 port map( A => n5396, B => DATAIN(26), S => n6049, Z => 
                           n4536);
   U2068 : MUX2_X1 port map( A => n5395, B => DATAIN(27), S => n6049, Z => 
                           n4537);
   U2069 : MUX2_X1 port map( A => n5394, B => DATAIN(28), S => n6049, Z => 
                           n4538);
   U2070 : MUX2_X1 port map( A => n5393, B => DATAIN(29), S => n6049, Z => 
                           n4539);
   U2071 : MUX2_X1 port map( A => n5392, B => DATAIN(30), S => n6049, Z => 
                           n4540);
   U2072 : MUX2_X1 port map( A => n5391, B => DATAIN(31), S => n6049, Z => 
                           n4541);
   U2073 : MUX2_X1 port map( A => n5744, B => DATAIN(31), S => n6250, Z => 
                           n3302);
   U2074 : MUX2_X1 port map( A => n5358, B => DATAIN(0), S => n6050, Z => n3079
                           );
   U2075 : MUX2_X1 port map( A => n5711, B => DATAIN(1), S => n6050, Z => n3080
                           );
   U2076 : MUX2_X1 port map( A => n5710, B => DATAIN(2), S => n6050, Z => n3081
                           );
   U2077 : MUX2_X1 port map( A => n5709, B => DATAIN(3), S => n6050, Z => n3082
                           );
   U2078 : MUX2_X1 port map( A => n5708, B => DATAIN(4), S => n6050, Z => n3083
                           );
   U2079 : MUX2_X1 port map( A => n5707, B => DATAIN(5), S => n6050, Z => n3084
                           );
   U2080 : MUX2_X1 port map( A => n5706, B => DATAIN(6), S => n6050, Z => n3085
                           );
   U2081 : MUX2_X1 port map( A => n5705, B => DATAIN(7), S => n6050, Z => n3086
                           );
   U2082 : MUX2_X1 port map( A => n5704, B => DATAIN(8), S => n6050, Z => n3087
                           );
   U2083 : MUX2_X1 port map( A => n5703, B => DATAIN(9), S => n6050, Z => n3088
                           );
   U2084 : MUX2_X1 port map( A => n5702, B => DATAIN(10), S => n6050, Z => 
                           n3089);
   U2085 : MUX2_X1 port map( A => n5701, B => DATAIN(11), S => n6050, Z => 
                           n3090);
   U2086 : MUX2_X1 port map( A => n5700, B => DATAIN(12), S => n6051, Z => 
                           n3091);
   U2087 : MUX2_X1 port map( A => n5699, B => DATAIN(13), S => n6051, Z => 
                           n3092);
   U2088 : MUX2_X1 port map( A => n5698, B => DATAIN(14), S => n6051, Z => 
                           n3093);
   U2089 : MUX2_X1 port map( A => n5697, B => DATAIN(15), S => n6051, Z => 
                           n3094);
   U2090 : MUX2_X1 port map( A => n5696, B => DATAIN(16), S => n6051, Z => 
                           n3095);
   U2091 : MUX2_X1 port map( A => n5695, B => DATAIN(17), S => n6051, Z => 
                           n3096);
   U2092 : MUX2_X1 port map( A => n5694, B => DATAIN(18), S => n6051, Z => 
                           n3097);
   U2093 : MUX2_X1 port map( A => n5693, B => DATAIN(19), S => n6051, Z => 
                           n3098);
   U2094 : MUX2_X1 port map( A => n5692, B => DATAIN(20), S => n6051, Z => 
                           n3099);
   U2095 : MUX2_X1 port map( A => n5691, B => DATAIN(21), S => n6051, Z => 
                           n3100);
   U2096 : MUX2_X1 port map( A => n5690, B => DATAIN(22), S => n6051, Z => 
                           n3101);
   U2097 : MUX2_X1 port map( A => n5689, B => DATAIN(23), S => n6051, Z => 
                           n3102);
   U2098 : MUX2_X1 port map( A => n5688, B => DATAIN(24), S => n6052, Z => 
                           n3103);
   U2099 : MUX2_X1 port map( A => n5687, B => DATAIN(25), S => n6052, Z => 
                           n3104);
   U2100 : MUX2_X1 port map( A => n5686, B => DATAIN(26), S => n6052, Z => 
                           n3105);
   U2101 : MUX2_X1 port map( A => n5685, B => DATAIN(27), S => n6052, Z => 
                           n3106);
   U2102 : MUX2_X1 port map( A => n5684, B => DATAIN(28), S => n6052, Z => 
                           n3107);
   U2103 : MUX2_X1 port map( A => n5683, B => DATAIN(29), S => n6052, Z => 
                           n3108);
   U2104 : MUX2_X1 port map( A => n5682, B => DATAIN(30), S => n6052, Z => 
                           n3109);
   U2105 : MUX2_X1 port map( A => n5681, B => DATAIN(31), S => n6052, Z => 
                           n3110);
   U2106 : NAND2_X1 port map( A1 => n6489, A2 => n4619, ZN => n6486);
   U2107 : OAI22_X1 port map( A1 => n6056, A2 => n5974, B1 => n6340, B2 => 
                           n6057, ZN => n7837);
   U2108 : OAI22_X1 port map( A1 => n6055, A2 => n6004, B1 => n6342, B2 => 
                           n6057, ZN => n7836);
   U2109 : OAI22_X1 port map( A1 => n6056, A2 => n6003, B1 => n6344, B2 => 
                           n6057, ZN => n7835);
   U2110 : OAI22_X1 port map( A1 => n6055, A2 => n6002, B1 => n6346, B2 => 
                           n6057, ZN => n7834);
   U2111 : OAI22_X1 port map( A1 => n6056, A2 => n6001, B1 => n6347, B2 => 
                           n6058, ZN => n7833);
   U2112 : OAI22_X1 port map( A1 => n6055, A2 => n6000, B1 => n6348, B2 => 
                           n6058, ZN => n7832);
   U2113 : OAI22_X1 port map( A1 => n6056, A2 => n5999, B1 => n6349, B2 => 
                           n6058, ZN => n7831);
   U2114 : OAI22_X1 port map( A1 => n6055, A2 => n5998, B1 => n6350, B2 => 
                           n6058, ZN => n7830);
   U2115 : OAI22_X1 port map( A1 => n6056, A2 => n5997, B1 => n6351, B2 => 
                           n6058, ZN => n7829);
   U2116 : OAI22_X1 port map( A1 => n6056, A2 => n5996, B1 => n6352, B2 => 
                           n6058, ZN => n7828);
   U2117 : OAI22_X1 port map( A1 => n6056, A2 => n5995, B1 => n6353, B2 => 
                           n6058, ZN => n7827);
   U2118 : OAI22_X1 port map( A1 => n6056, A2 => n5994, B1 => n6354, B2 => 
                           n6059, ZN => n7826);
   U2119 : OAI22_X1 port map( A1 => n6056, A2 => n5993, B1 => n6355, B2 => 
                           n6059, ZN => n7825);
   U2120 : OAI22_X1 port map( A1 => n6056, A2 => n5992, B1 => n6356, B2 => 
                           n6059, ZN => n7824);
   U2121 : OAI22_X1 port map( A1 => n6056, A2 => n5991, B1 => n6357, B2 => 
                           n6059, ZN => n7823);
   U2122 : OAI22_X1 port map( A1 => n6056, A2 => n5990, B1 => n6358, B2 => 
                           n6059, ZN => n7822);
   U2123 : OAI22_X1 port map( A1 => n6056, A2 => n5989, B1 => n6359, B2 => 
                           n6059, ZN => n7821);
   U2124 : OAI22_X1 port map( A1 => n6056, A2 => n5988, B1 => n6360, B2 => 
                           n6059, ZN => n7820);
   U2125 : OAI22_X1 port map( A1 => n6056, A2 => n5987, B1 => n6361, B2 => 
                           n6060, ZN => n7819);
   U2126 : OAI22_X1 port map( A1 => n6056, A2 => n5986, B1 => n6362, B2 => 
                           n6060, ZN => n7818);
   U2127 : OAI22_X1 port map( A1 => n6055, A2 => n5985, B1 => n6363, B2 => 
                           n6060, ZN => n7817);
   U2128 : OAI22_X1 port map( A1 => n6055, A2 => n5984, B1 => n6364, B2 => 
                           n6060, ZN => n7816);
   U2129 : OAI22_X1 port map( A1 => n6055, A2 => n5983, B1 => n6365, B2 => 
                           n6060, ZN => n7815);
   U2130 : OAI22_X1 port map( A1 => n6055, A2 => n5982, B1 => n6366, B2 => 
                           n6060, ZN => n7814);
   U2131 : OAI22_X1 port map( A1 => n6055, A2 => n5981, B1 => n6367, B2 => 
                           n6060, ZN => n7813);
   U2132 : OAI22_X1 port map( A1 => n6055, A2 => n5980, B1 => n6368, B2 => 
                           n6061, ZN => n7812);
   U2133 : OAI22_X1 port map( A1 => n6055, A2 => n5979, B1 => n6369, B2 => 
                           n6061, ZN => n7811);
   U2134 : OAI22_X1 port map( A1 => n6055, A2 => n5978, B1 => n6370, B2 => 
                           n6061, ZN => n7810);
   U2135 : OAI22_X1 port map( A1 => n6055, A2 => n5977, B1 => n6371, B2 => 
                           n6061, ZN => n7809);
   U2136 : OAI22_X1 port map( A1 => n6055, A2 => n5976, B1 => n6372, B2 => 
                           n6061, ZN => n7808);
   U2137 : OAI22_X1 port map( A1 => n6055, A2 => n5975, B1 => n6373, B2 => 
                           n6061, ZN => n7807);
   U2138 : OAI22_X1 port map( A1 => n6055, A2 => n5973, B1 => n6374, B2 => 
                           n6061, ZN => n7806);
   U2139 : NAND2_X1 port map( A1 => n6489, A2 => n4620, ZN => n6487);
   U2140 : OAI22_X1 port map( A1 => n6065, A2 => n5910, B1 => n6340, B2 => 
                           n6066, ZN => n7805);
   U2141 : OAI22_X1 port map( A1 => n6064, A2 => n5940, B1 => n6342, B2 => 
                           n6066, ZN => n7804);
   U2142 : OAI22_X1 port map( A1 => n6065, A2 => n5939, B1 => n6344, B2 => 
                           n6066, ZN => n7803);
   U2143 : OAI22_X1 port map( A1 => n6064, A2 => n5938, B1 => n6346, B2 => 
                           n6066, ZN => n7802);
   U2144 : OAI22_X1 port map( A1 => n6065, A2 => n5937, B1 => n6347, B2 => 
                           n6067, ZN => n7801);
   U2145 : OAI22_X1 port map( A1 => n6064, A2 => n5936, B1 => n6348, B2 => 
                           n6067, ZN => n7800);
   U2146 : OAI22_X1 port map( A1 => n6065, A2 => n5935, B1 => n6349, B2 => 
                           n6067, ZN => n7799);
   U2147 : OAI22_X1 port map( A1 => n6064, A2 => n5934, B1 => n6350, B2 => 
                           n6067, ZN => n7798);
   U2148 : OAI22_X1 port map( A1 => n6065, A2 => n5933, B1 => n6351, B2 => 
                           n6067, ZN => n7797);
   U2149 : OAI22_X1 port map( A1 => n6065, A2 => n5932, B1 => n6352, B2 => 
                           n6067, ZN => n7796);
   U2150 : OAI22_X1 port map( A1 => n6065, A2 => n5931, B1 => n6353, B2 => 
                           n6067, ZN => n7795);
   U2151 : OAI22_X1 port map( A1 => n6065, A2 => n5930, B1 => n6354, B2 => 
                           n6068, ZN => n7794);
   U2152 : OAI22_X1 port map( A1 => n6065, A2 => n5929, B1 => n6355, B2 => 
                           n6068, ZN => n7793);
   U2153 : OAI22_X1 port map( A1 => n6065, A2 => n5928, B1 => n6356, B2 => 
                           n6068, ZN => n7792);
   U2154 : OAI22_X1 port map( A1 => n6065, A2 => n5927, B1 => n6357, B2 => 
                           n6068, ZN => n7791);
   U2155 : OAI22_X1 port map( A1 => n6065, A2 => n5926, B1 => n6358, B2 => 
                           n6068, ZN => n7790);
   U2156 : OAI22_X1 port map( A1 => n6065, A2 => n5925, B1 => n6359, B2 => 
                           n6068, ZN => n7789);
   U2157 : OAI22_X1 port map( A1 => n6065, A2 => n5924, B1 => n6360, B2 => 
                           n6068, ZN => n7788);
   U2158 : OAI22_X1 port map( A1 => n6065, A2 => n5923, B1 => n6361, B2 => 
                           n6069, ZN => n7787);
   U2159 : OAI22_X1 port map( A1 => n6065, A2 => n5922, B1 => n6362, B2 => 
                           n6069, ZN => n7786);
   U2160 : OAI22_X1 port map( A1 => n6064, A2 => n5921, B1 => n6363, B2 => 
                           n6069, ZN => n7785);
   U2161 : OAI22_X1 port map( A1 => n6064, A2 => n5920, B1 => n6364, B2 => 
                           n6069, ZN => n7784);
   U2162 : OAI22_X1 port map( A1 => n6064, A2 => n5919, B1 => n6365, B2 => 
                           n6069, ZN => n7783);
   U2163 : OAI22_X1 port map( A1 => n6064, A2 => n5918, B1 => n6366, B2 => 
                           n6069, ZN => n7782);
   U2164 : OAI22_X1 port map( A1 => n6064, A2 => n5917, B1 => n6367, B2 => 
                           n6069, ZN => n7781);
   U2165 : OAI22_X1 port map( A1 => n6064, A2 => n5916, B1 => n6368, B2 => 
                           n6070, ZN => n7780);
   U2166 : OAI22_X1 port map( A1 => n6064, A2 => n5915, B1 => n6369, B2 => 
                           n6070, ZN => n7779);
   U2167 : OAI22_X1 port map( A1 => n6064, A2 => n5914, B1 => n6370, B2 => 
                           n6070, ZN => n7778);
   U2168 : OAI22_X1 port map( A1 => n6064, A2 => n5913, B1 => n6371, B2 => 
                           n6070, ZN => n7777);
   U2169 : OAI22_X1 port map( A1 => n6064, A2 => n5912, B1 => n6372, B2 => 
                           n6070, ZN => n7776);
   U2170 : OAI22_X1 port map( A1 => n6064, A2 => n5911, B1 => n6373, B2 => 
                           n6070, ZN => n7775);
   U2171 : OAI22_X1 port map( A1 => n6064, A2 => n5909, B1 => n6374, B2 => 
                           n6070, ZN => n7774);
   U2172 : NAND2_X1 port map( A1 => n6489, A2 => n4614, ZN => n6488);
   U2173 : OAI22_X1 port map( A1 => n6074, A2 => n6936, B1 => n6340, B2 => 
                           n6075, ZN => n7773);
   U2174 : OAI22_X1 port map( A1 => n6073, A2 => n6955, B1 => n6342, B2 => 
                           n6075, ZN => n7772);
   U2175 : OAI22_X1 port map( A1 => n6074, A2 => n6973, B1 => n6344, B2 => 
                           n6075, ZN => n7771);
   U2176 : OAI22_X1 port map( A1 => n6073, A2 => n6991, B1 => n6346, B2 => 
                           n6075, ZN => n7770);
   U2177 : OAI22_X1 port map( A1 => n6074, A2 => n7010, B1 => n6347, B2 => 
                           n6076, ZN => n7769);
   U2178 : OAI22_X1 port map( A1 => n6073, A2 => n7029, B1 => n6348, B2 => 
                           n6076, ZN => n7768);
   U2179 : OAI22_X1 port map( A1 => n6074, A2 => n7048, B1 => n6349, B2 => 
                           n6076, ZN => n7767);
   U2180 : OAI22_X1 port map( A1 => n6073, A2 => n7067, B1 => n6350, B2 => 
                           n6076, ZN => n7766);
   U2181 : OAI22_X1 port map( A1 => n6074, A2 => n7086, B1 => n6351, B2 => 
                           n6076, ZN => n7765);
   U2182 : OAI22_X1 port map( A1 => n6074, A2 => n7105, B1 => n6352, B2 => 
                           n6076, ZN => n7764);
   U2183 : OAI22_X1 port map( A1 => n6074, A2 => n7124, B1 => n6353, B2 => 
                           n6076, ZN => n7763);
   U2184 : OAI22_X1 port map( A1 => n6074, A2 => n7143, B1 => n6354, B2 => 
                           n6077, ZN => n7762);
   U2185 : OAI22_X1 port map( A1 => n6074, A2 => n7162, B1 => n6355, B2 => 
                           n6077, ZN => n7761);
   U2186 : OAI22_X1 port map( A1 => n6074, A2 => n7181, B1 => n6356, B2 => 
                           n6077, ZN => n7760);
   U2187 : OAI22_X1 port map( A1 => n6074, A2 => n7200, B1 => n6357, B2 => 
                           n6077, ZN => n7759);
   U2188 : OAI22_X1 port map( A1 => n6074, A2 => n7219, B1 => n6358, B2 => 
                           n6077, ZN => n7758);
   U2189 : OAI22_X1 port map( A1 => n6074, A2 => n7238, B1 => n6359, B2 => 
                           n6077, ZN => n7757);
   U2190 : OAI22_X1 port map( A1 => n6074, A2 => n7257, B1 => n6360, B2 => 
                           n6077, ZN => n7756);
   U2191 : OAI22_X1 port map( A1 => n6074, A2 => n7276, B1 => n6361, B2 => 
                           n6078, ZN => n7755);
   U2192 : OAI22_X1 port map( A1 => n6074, A2 => n7295, B1 => n6362, B2 => 
                           n6078, ZN => n7754);
   U2193 : OAI22_X1 port map( A1 => n6073, A2 => n7314, B1 => n6363, B2 => 
                           n6078, ZN => n7753);
   U2194 : OAI22_X1 port map( A1 => n6073, A2 => n7333, B1 => n6364, B2 => 
                           n6078, ZN => n7752);
   U2195 : OAI22_X1 port map( A1 => n6073, A2 => n7352, B1 => n6365, B2 => 
                           n6078, ZN => n7751);
   U2196 : OAI22_X1 port map( A1 => n6073, A2 => n7371, B1 => n6366, B2 => 
                           n6078, ZN => n7750);
   U2197 : OAI22_X1 port map( A1 => n6073, A2 => n7390, B1 => n6367, B2 => 
                           n6078, ZN => n7749);
   U2198 : OAI22_X1 port map( A1 => n6073, A2 => n7409, B1 => n6368, B2 => 
                           n6079, ZN => n7748);
   U2199 : OAI22_X1 port map( A1 => n6073, A2 => n7428, B1 => n6369, B2 => 
                           n6079, ZN => n7747);
   U2200 : OAI22_X1 port map( A1 => n6073, A2 => n7447, B1 => n6370, B2 => 
                           n6079, ZN => n7746);
   U2201 : OAI22_X1 port map( A1 => n6073, A2 => n7466, B1 => n6371, B2 => 
                           n6079, ZN => n7745);
   U2202 : OAI22_X1 port map( A1 => n6073, A2 => n7485, B1 => n6372, B2 => 
                           n6079, ZN => n7744);
   U2203 : OAI22_X1 port map( A1 => n6073, A2 => n7504, B1 => n6373, B2 => 
                           n6079, ZN => n7743);
   U2204 : OAI22_X1 port map( A1 => n6073, A2 => n7534, B1 => n6374, B2 => 
                           n6079, ZN => n7742);
   U2205 : NAND2_X1 port map( A1 => n6489, A2 => n4611, ZN => n6490);
   U2206 : OAI22_X1 port map( A1 => n6083, A2 => n6937, B1 => n6339, B2 => 
                           n6084, ZN => n7741);
   U2207 : OAI22_X1 port map( A1 => n6083, A2 => n6956, B1 => n6341, B2 => 
                           n6084, ZN => n7740);
   U2208 : OAI22_X1 port map( A1 => n6083, A2 => n6974, B1 => n6343, B2 => 
                           n6084, ZN => n7739);
   U2209 : OAI22_X1 port map( A1 => n6083, A2 => n6992, B1 => n6345, B2 => 
                           n6084, ZN => n7738);
   U2210 : OAI22_X1 port map( A1 => n6083, A2 => n7011, B1 => n6347, B2 => 
                           n6085, ZN => n7737);
   U2211 : OAI22_X1 port map( A1 => n6083, A2 => n7030, B1 => n6348, B2 => 
                           n6085, ZN => n7736);
   U2212 : OAI22_X1 port map( A1 => n6083, A2 => n7049, B1 => n6349, B2 => 
                           n6085, ZN => n7735);
   U2213 : OAI22_X1 port map( A1 => n6083, A2 => n7068, B1 => n6350, B2 => 
                           n6085, ZN => n7734);
   U2214 : OAI22_X1 port map( A1 => n6082, A2 => n7087, B1 => n6351, B2 => 
                           n6085, ZN => n7733);
   U2215 : OAI22_X1 port map( A1 => n6082, A2 => n7106, B1 => n6352, B2 => 
                           n6085, ZN => n7732);
   U2216 : OAI22_X1 port map( A1 => n6082, A2 => n7125, B1 => n6353, B2 => 
                           n6085, ZN => n7731);
   U2217 : OAI22_X1 port map( A1 => n6082, A2 => n7144, B1 => n6354, B2 => 
                           n6086, ZN => n7730);
   U2218 : OAI22_X1 port map( A1 => n6082, A2 => n7163, B1 => n6355, B2 => 
                           n6086, ZN => n7729);
   U2219 : OAI22_X1 port map( A1 => n6082, A2 => n7182, B1 => n6356, B2 => 
                           n6086, ZN => n7728);
   U2220 : OAI22_X1 port map( A1 => n6082, A2 => n7201, B1 => n6357, B2 => 
                           n6086, ZN => n7727);
   U2221 : OAI22_X1 port map( A1 => n6082, A2 => n7220, B1 => n6358, B2 => 
                           n6086, ZN => n7726);
   U2222 : OAI22_X1 port map( A1 => n6082, A2 => n7239, B1 => n6359, B2 => 
                           n6086, ZN => n7725);
   U2223 : OAI22_X1 port map( A1 => n6082, A2 => n7258, B1 => n6360, B2 => 
                           n6086, ZN => n7724);
   U2224 : OAI22_X1 port map( A1 => n6082, A2 => n7277, B1 => n6361, B2 => 
                           n6087, ZN => n7723);
   U2225 : OAI22_X1 port map( A1 => n6082, A2 => n7296, B1 => n6362, B2 => 
                           n6087, ZN => n7722);
   U2226 : OAI22_X1 port map( A1 => n6083, A2 => n7315, B1 => n6363, B2 => 
                           n6087, ZN => n7721);
   U2227 : OAI22_X1 port map( A1 => n6083, A2 => n7334, B1 => n6364, B2 => 
                           n6087, ZN => n7720);
   U2228 : OAI22_X1 port map( A1 => n6083, A2 => n7353, B1 => n6365, B2 => 
                           n6087, ZN => n7719);
   U2229 : OAI22_X1 port map( A1 => n6083, A2 => n7372, B1 => n6366, B2 => 
                           n6087, ZN => n7718);
   U2230 : OAI22_X1 port map( A1 => n6082, A2 => n7391, B1 => n6367, B2 => 
                           n6087, ZN => n7717);
   U2231 : OAI22_X1 port map( A1 => n6083, A2 => n7410, B1 => n6368, B2 => 
                           n6088, ZN => n7716);
   U2232 : OAI22_X1 port map( A1 => n6082, A2 => n7429, B1 => n6369, B2 => 
                           n6088, ZN => n7715);
   U2233 : OAI22_X1 port map( A1 => n6083, A2 => n7448, B1 => n6370, B2 => 
                           n6088, ZN => n7714);
   U2234 : OAI22_X1 port map( A1 => n6082, A2 => n7467, B1 => n6371, B2 => 
                           n6088, ZN => n7713);
   U2235 : OAI22_X1 port map( A1 => n6083, A2 => n7486, B1 => n6372, B2 => 
                           n6088, ZN => n7712);
   U2236 : OAI22_X1 port map( A1 => n6082, A2 => n7505, B1 => n6373, B2 => 
                           n6088, ZN => n7711);
   U2237 : OAI22_X1 port map( A1 => n6083, A2 => n7535, B1 => n6374, B2 => 
                           n6088, ZN => n7710);
   U2238 : NAND2_X1 port map( A1 => n4607, A2 => n4614, ZN => n6491);
   U2239 : OAI22_X1 port map( A1 => n6092, A2 => n5972, B1 => n6340, B2 => 
                           n6093, ZN => n3207);
   U2240 : OAI22_X1 port map( A1 => n6092, A2 => n5971, B1 => n6342, B2 => 
                           n6093, ZN => n3208);
   U2241 : OAI22_X1 port map( A1 => n6092, A2 => n5970, B1 => n6344, B2 => 
                           n6093, ZN => n3209);
   U2242 : OAI22_X1 port map( A1 => n6092, A2 => n5969, B1 => n6346, B2 => 
                           n6093, ZN => n3210);
   U2243 : OAI22_X1 port map( A1 => n6092, A2 => n5968, B1 => n6347, B2 => 
                           n6094, ZN => n3211);
   U2244 : OAI22_X1 port map( A1 => n6092, A2 => n5967, B1 => n6348, B2 => 
                           n6094, ZN => n3212);
   U2245 : OAI22_X1 port map( A1 => n6092, A2 => n5966, B1 => n6349, B2 => 
                           n6094, ZN => n3213);
   U2246 : OAI22_X1 port map( A1 => n6092, A2 => n5965, B1 => n6350, B2 => 
                           n6094, ZN => n3214);
   U2247 : OAI22_X1 port map( A1 => n6091, A2 => n5964, B1 => n6351, B2 => 
                           n6094, ZN => n3215);
   U2248 : OAI22_X1 port map( A1 => n6091, A2 => n5963, B1 => n6352, B2 => 
                           n6094, ZN => n3216);
   U2249 : OAI22_X1 port map( A1 => n6091, A2 => n5962, B1 => n6353, B2 => 
                           n6094, ZN => n3217);
   U2250 : OAI22_X1 port map( A1 => n6091, A2 => n5961, B1 => n6354, B2 => 
                           n6095, ZN => n3218);
   U2251 : OAI22_X1 port map( A1 => n6091, A2 => n5960, B1 => n6355, B2 => 
                           n6095, ZN => n3219);
   U2252 : OAI22_X1 port map( A1 => n6091, A2 => n5959, B1 => n6356, B2 => 
                           n6095, ZN => n3220);
   U2253 : OAI22_X1 port map( A1 => n6091, A2 => n5958, B1 => n6357, B2 => 
                           n6095, ZN => n3221);
   U2254 : OAI22_X1 port map( A1 => n6091, A2 => n5957, B1 => n6358, B2 => 
                           n6095, ZN => n3222);
   U2255 : OAI22_X1 port map( A1 => n6091, A2 => n5956, B1 => n6359, B2 => 
                           n6095, ZN => n3223);
   U2256 : OAI22_X1 port map( A1 => n6091, A2 => n5955, B1 => n6360, B2 => 
                           n6095, ZN => n3224);
   U2257 : OAI22_X1 port map( A1 => n6091, A2 => n5954, B1 => n6361, B2 => 
                           n6096, ZN => n3225);
   U2258 : OAI22_X1 port map( A1 => n6091, A2 => n5953, B1 => n6362, B2 => 
                           n6096, ZN => n3226);
   U2259 : OAI22_X1 port map( A1 => n6092, A2 => n5952, B1 => n6363, B2 => 
                           n6096, ZN => n3227);
   U2260 : OAI22_X1 port map( A1 => n6092, A2 => n5951, B1 => n6364, B2 => 
                           n6096, ZN => n3228);
   U2261 : OAI22_X1 port map( A1 => n6092, A2 => n5950, B1 => n6365, B2 => 
                           n6096, ZN => n3229);
   U2262 : OAI22_X1 port map( A1 => n6092, A2 => n5949, B1 => n6366, B2 => 
                           n6096, ZN => n3230);
   U2263 : OAI22_X1 port map( A1 => n6091, A2 => n5948, B1 => n6367, B2 => 
                           n6096, ZN => n3231);
   U2264 : OAI22_X1 port map( A1 => n6092, A2 => n5947, B1 => n6368, B2 => 
                           n6097, ZN => n3232);
   U2265 : OAI22_X1 port map( A1 => n6091, A2 => n5946, B1 => n6369, B2 => 
                           n6097, ZN => n3233);
   U2266 : OAI22_X1 port map( A1 => n6092, A2 => n5945, B1 => n6370, B2 => 
                           n6097, ZN => n3234);
   U2267 : OAI22_X1 port map( A1 => n6091, A2 => n5944, B1 => n6371, B2 => 
                           n6097, ZN => n3235);
   U2268 : OAI22_X1 port map( A1 => n6092, A2 => n5943, B1 => n6372, B2 => 
                           n6097, ZN => n3236);
   U2269 : OAI22_X1 port map( A1 => n6091, A2 => n5942, B1 => n6373, B2 => 
                           n6097, ZN => n3237);
   U2270 : OAI22_X1 port map( A1 => n6092, A2 => n5941, B1 => n6374, B2 => 
                           n6097, ZN => n3238);
   U2271 : NAND2_X1 port map( A1 => n4607, A2 => n4611, ZN => n6492);
   U2272 : MUX2_X1 port map( A => n5647, B => DATAIN(0), S => n6100, Z => n3175
                           );
   U2273 : MUX2_X1 port map( A => n5582, B => DATAIN(1), S => n6100, Z => n3176
                           );
   U2274 : MUX2_X1 port map( A => n5581, B => DATAIN(2), S => n6100, Z => n3177
                           );
   U2275 : MUX2_X1 port map( A => n5580, B => DATAIN(3), S => n6100, Z => n3178
                           );
   U2276 : OAI22_X1 port map( A1 => n6100, A2 => n7004, B1 => n6347, B2 => 
                           n6102, ZN => n7709);
   U2277 : OAI22_X1 port map( A1 => n6100, A2 => n7023, B1 => n6348, B2 => 
                           n6102, ZN => n7708);
   U2278 : OAI22_X1 port map( A1 => n6100, A2 => n7042, B1 => n6349, B2 => 
                           n6102, ZN => n7707);
   U2279 : OAI22_X1 port map( A1 => n6100, A2 => n7061, B1 => n6350, B2 => 
                           n6102, ZN => n7706);
   U2280 : OAI22_X1 port map( A1 => n6100, A2 => n7080, B1 => n6351, B2 => 
                           n6103, ZN => n7705);
   U2281 : OAI22_X1 port map( A1 => n6100, A2 => n7099, B1 => n6352, B2 => 
                           n6103, ZN => n7704);
   U2282 : OAI22_X1 port map( A1 => n6100, A2 => n7118, B1 => n6353, B2 => 
                           n6103, ZN => n7703);
   U2283 : OAI22_X1 port map( A1 => n6100, A2 => n7137, B1 => n6354, B2 => 
                           n6103, ZN => n7702);
   U2284 : OAI22_X1 port map( A1 => n6100, A2 => n7156, B1 => n6355, B2 => 
                           n6103, ZN => n7701);
   U2285 : OAI22_X1 port map( A1 => n6101, A2 => n7175, B1 => n6356, B2 => 
                           n6103, ZN => n7700);
   U2286 : OAI22_X1 port map( A1 => n6101, A2 => n7194, B1 => n6357, B2 => 
                           n6103, ZN => n7699);
   U2287 : OAI22_X1 port map( A1 => n6101, A2 => n7213, B1 => n6358, B2 => 
                           n6104, ZN => n7698);
   U2288 : OAI22_X1 port map( A1 => n6101, A2 => n7232, B1 => n6359, B2 => 
                           n6104, ZN => n7697);
   U2289 : OAI22_X1 port map( A1 => n6101, A2 => n7251, B1 => n6360, B2 => 
                           n6104, ZN => n7696);
   U2290 : OAI22_X1 port map( A1 => n6101, A2 => n7270, B1 => n6361, B2 => 
                           n6104, ZN => n7695);
   U2291 : OAI22_X1 port map( A1 => n6101, A2 => n7289, B1 => n6362, B2 => 
                           n6104, ZN => n7694);
   U2292 : OAI22_X1 port map( A1 => n6101, A2 => n7308, B1 => n6363, B2 => 
                           n6104, ZN => n7693);
   U2293 : OAI22_X1 port map( A1 => n6101, A2 => n7327, B1 => n6364, B2 => 
                           n6104, ZN => n7692);
   U2294 : OAI22_X1 port map( A1 => n6101, A2 => n7346, B1 => n6365, B2 => 
                           n6105, ZN => n7691);
   U2295 : OAI22_X1 port map( A1 => n6101, A2 => n7365, B1 => n6366, B2 => 
                           n6105, ZN => n7690);
   U2296 : OAI22_X1 port map( A1 => n6101, A2 => n7384, B1 => n6367, B2 => 
                           n6105, ZN => n7689);
   U2297 : OAI22_X1 port map( A1 => n6101, A2 => n7403, B1 => n6368, B2 => 
                           n6105, ZN => n7688);
   U2298 : OAI22_X1 port map( A1 => n6100, A2 => n7422, B1 => n6369, B2 => 
                           n6105, ZN => n7687);
   U2299 : OAI22_X1 port map( A1 => n6101, A2 => n7441, B1 => n6370, B2 => 
                           n6105, ZN => n7686);
   U2300 : OAI22_X1 port map( A1 => n6100, A2 => n7460, B1 => n6371, B2 => 
                           n6105, ZN => n7685);
   U2301 : OAI22_X1 port map( A1 => n6101, A2 => n7479, B1 => n6372, B2 => 
                           n6106, ZN => n7684);
   U2302 : OAI22_X1 port map( A1 => n6100, A2 => n7498, B1 => n6373, B2 => 
                           n6106, ZN => n7683);
   U2303 : OAI22_X1 port map( A1 => n6101, A2 => n7521, B1 => n6374, B2 => 
                           n6106, ZN => n3206);
   U2304 : NAND2_X1 port map( A1 => n4625, A2 => n4606, ZN => n6493);
   U2305 : MUX2_X1 port map( A => n5583, B => DATAIN(0), S => n6109, Z => n3143
                           );
   U2306 : MUX2_X1 port map( A => n5485, B => DATAIN(1), S => n6109, Z => n3144
                           );
   U2307 : MUX2_X1 port map( A => n5484, B => DATAIN(2), S => n6109, Z => n3145
                           );
   U2308 : MUX2_X1 port map( A => n5483, B => DATAIN(3), S => n6109, Z => n3146
                           );
   U2309 : OAI22_X1 port map( A1 => n6109, A2 => n5907, B1 => n6347, B2 => 
                           n6111, ZN => n7682);
   U2310 : OAI22_X1 port map( A1 => n6109, A2 => n5906, B1 => n6348, B2 => 
                           n6111, ZN => n7681);
   U2311 : OAI22_X1 port map( A1 => n6109, A2 => n5905, B1 => n6349, B2 => 
                           n6111, ZN => n7680);
   U2312 : OAI22_X1 port map( A1 => n6109, A2 => n5904, B1 => n6350, B2 => 
                           n6111, ZN => n7679);
   U2313 : OAI22_X1 port map( A1 => n6109, A2 => n5903, B1 => n6351, B2 => 
                           n6112, ZN => n7678);
   U2314 : OAI22_X1 port map( A1 => n6109, A2 => n5902, B1 => n6352, B2 => 
                           n6112, ZN => n7677);
   U2315 : OAI22_X1 port map( A1 => n6109, A2 => n5901, B1 => n6353, B2 => 
                           n6112, ZN => n7676);
   U2316 : OAI22_X1 port map( A1 => n6109, A2 => n5900, B1 => n6354, B2 => 
                           n6112, ZN => n7675);
   U2317 : OAI22_X1 port map( A1 => n6109, A2 => n5899, B1 => n6355, B2 => 
                           n6112, ZN => n7674);
   U2318 : OAI22_X1 port map( A1 => n6110, A2 => n5898, B1 => n6356, B2 => 
                           n6112, ZN => n7673);
   U2319 : OAI22_X1 port map( A1 => n6110, A2 => n5897, B1 => n6357, B2 => 
                           n6112, ZN => n7672);
   U2320 : OAI22_X1 port map( A1 => n6110, A2 => n5896, B1 => n6358, B2 => 
                           n6113, ZN => n7671);
   U2321 : OAI22_X1 port map( A1 => n6110, A2 => n5895, B1 => n6359, B2 => 
                           n6113, ZN => n7670);
   U2322 : OAI22_X1 port map( A1 => n6110, A2 => n5894, B1 => n6360, B2 => 
                           n6113, ZN => n7669);
   U2323 : OAI22_X1 port map( A1 => n6110, A2 => n5893, B1 => n6361, B2 => 
                           n6113, ZN => n7668);
   U2324 : OAI22_X1 port map( A1 => n6110, A2 => n5892, B1 => n6362, B2 => 
                           n6113, ZN => n7667);
   U2325 : OAI22_X1 port map( A1 => n6110, A2 => n5891, B1 => n6363, B2 => 
                           n6113, ZN => n7666);
   U2326 : OAI22_X1 port map( A1 => n6110, A2 => n5890, B1 => n6364, B2 => 
                           n6113, ZN => n7665);
   U2327 : OAI22_X1 port map( A1 => n6110, A2 => n5889, B1 => n6365, B2 => 
                           n6114, ZN => n7664);
   U2328 : OAI22_X1 port map( A1 => n6110, A2 => n5888, B1 => n6366, B2 => 
                           n6114, ZN => n7663);
   U2329 : OAI22_X1 port map( A1 => n6110, A2 => n5887, B1 => n6367, B2 => 
                           n6114, ZN => n7662);
   U2330 : OAI22_X1 port map( A1 => n6110, A2 => n5886, B1 => n6368, B2 => 
                           n6114, ZN => n7661);
   U2331 : OAI22_X1 port map( A1 => n6109, A2 => n5885, B1 => n6369, B2 => 
                           n6114, ZN => n7660);
   U2332 : OAI22_X1 port map( A1 => n6110, A2 => n5884, B1 => n6370, B2 => 
                           n6114, ZN => n7659);
   U2333 : OAI22_X1 port map( A1 => n6109, A2 => n5883, B1 => n6371, B2 => 
                           n6114, ZN => n7658);
   U2334 : OAI22_X1 port map( A1 => n6110, A2 => n5882, B1 => n6372, B2 => 
                           n6115, ZN => n7657);
   U2335 : OAI22_X1 port map( A1 => n6109, A2 => n5881, B1 => n6373, B2 => 
                           n6115, ZN => n7656);
   U2336 : OAI22_X1 port map( A1 => n6110, A2 => n5880, B1 => n6374, B2 => 
                           n6115, ZN => n3174);
   U2337 : INV_X1 port map( A => n2002, ZN => n6494);
   U2338 : NAND4_X1 port map( A1 => n1997, A2 => n2027, A3 => n1998, A4 => 
                           n6494, ZN => n6495);
   U2339 : NAND2_X1 port map( A1 => n6173, A2 => n6495, ZN => n6502);
   U2340 : INV_X1 port map( A => n6502, ZN => n6916);
   U2341 : NAND2_X1 port map( A1 => n4612, A2 => n4618, ZN => n6906);
   U2342 : NAND2_X1 port map( A1 => n4626, A2 => n4610, ZN => n6907);
   U2343 : OAI22_X1 port map( A1 => n3742, A2 => n4902, B1 => n2284, B2 => 
                           n4900, ZN => n6496);
   U2344 : AOI221_X1 port map( B1 => n6160, B2 => n6938, C1 => n6275, C2 => 
                           n7588, A => n6496, ZN => n6501);
   U2345 : AOI222_X1 port map( A1 => n6298, A2 => n4062, B1 => n6287, B2 => 
                           n7586, C1 => n6301, C2 => n4030, ZN => n6500);
   U2346 : AOI22_X1 port map( A1 => n2910, A2 => n6149, B1 => n6934, B2 => 
                           n6146, ZN => n6497);
   U2347 : OAI221_X1 port map( B1 => n4813, B2 => n6155, C1 => n6936, C2 => 
                           n6152, A => n6497, ZN => n6498);
   U2348 : NOR4_X1 port map( A1 => n6498, A2 => n2025, A3 => n2024, A4 => n2021
                           , ZN => n6499);
   U2349 : AND3_X1 port map( A1 => n6501, A2 => n6500, A3 => n6499, ZN => n6503
                           );
   U2350 : OAI222_X1 port map( A1 => n2124, A2 => n6116, B1 => n939, B2 => 
                           n6121, C1 => n6503, C2 => n6502, ZN => n6510);
   U2351 : NAND2_X1 port map( A1 => n2006, A2 => n4618, ZN => n6910);
   U2352 : NAND2_X1 port map( A1 => n4612, A2 => n4621, ZN => n6513);
   U2353 : INV_X1 port map( A => n2156, ZN => n7553);
   U2354 : AOI22_X1 port map( A1 => n6124, A2 => n7553, B1 => n4897, B2 => 
                           n4972, ZN => n6504);
   U2355 : OAI221_X1 port map( B1 => n2092, B2 => n6130, C1 => n938, C2 => 
                           n6513, A => n6504, ZN => n6509);
   U2356 : NAND2_X1 port map( A1 => n4621, A2 => n1993, ZN => n6913);
   U2357 : NAND2_X1 port map( A1 => n4610, A2 => n4618, ZN => n6515);
   U2358 : AOI22_X1 port map( A1 => n6135, A2 => n950, B1 => n4898, B2 => n4912
                           , ZN => n6505);
   U2359 : OAI221_X1 port map( B1 => n3646, B2 => n6141, C1 => n2188, C2 => 
                           n6515, A => n6505, ZN => n6508);
   U2360 : NAND2_X1 port map( A1 => n1993, A2 => n4618, ZN => n6922);
   U2361 : NAND2_X1 port map( A1 => n4661, A2 => n4610, ZN => n6521);
   U2362 : AOI22_X1 port map( A1 => n6164, A2 => n6942, B1 => n4616, B2 => 
                           DATAIN(0), ZN => n6506);
   U2363 : OAI221_X1 port map( B1 => n2220, B2 => n6170, C1 => n2942, C2 => 
                           n6521, A => n6506, ZN => n6507);
   U2364 : NOR4_X1 port map( A1 => n6510, A2 => n6509, A3 => n6508, A4 => n6507
                           , ZN => n6511);
   U2365 : OAI21_X1 port map( B1 => n6173, B2 => n6512, A => n6511, ZN => n2983
                           );
   U2366 : OAI222_X1 port map( A1 => n956, A2 => n6121, B1 => n2719, B2 => 
                           n6119, C1 => n2125, C2 => n6116, ZN => n6527);
   U2367 : INV_X1 port map( A => n6513, ZN => n6908);
   U2368 : INV_X1 port map( A => n2157, ZN => n7554);
   U2369 : AOI22_X1 port map( A1 => n6127, A2 => n5036, B1 => n6124, B2 => 
                           n7554, ZN => n6514);
   U2370 : OAI221_X1 port map( B1 => n2061, B2 => n6133, C1 => n2093, C2 => 
                           n6130, A => n6514, ZN => n6526);
   U2371 : INV_X1 port map( A => n6515, ZN => n6911);
   U2372 : AOI22_X1 port map( A1 => n6138, A2 => n5033, B1 => n6135, B2 => n966
                           , ZN => n6516);
   U2373 : OAI221_X1 port map( B1 => n6342, B2 => n6144, C1 => n3647, C2 => 
                           n6141, A => n6516, ZN => n6525);
   U2374 : AOI22_X1 port map( A1 => n2911, A2 => n6149, B1 => n6953, B2 => 
                           n6146, ZN => n6517);
   U2375 : OAI221_X1 port map( B1 => n4811, B2 => n6155, C1 => n6955, C2 => 
                           n6152, A => n6517, ZN => n6520);
   U2376 : NAND2_X1 port map( A1 => n6160, A2 => n6957, ZN => n6518);
   U2377 : NAND4_X1 port map( A1 => n1975, A2 => n1976, A3 => n1974, A4 => 
                           n6518, ZN => n6519);
   U2378 : OAI21_X1 port map( B1 => n6520, B2 => n6519, A => n6163, ZN => n6523
                           );
   U2379 : INV_X1 port map( A => n6521, ZN => n6919);
   U2380 : AOI22_X1 port map( A1 => n6167, A2 => n6951, B1 => n6164, B2 => 
                           n4942, ZN => n6522);
   U2381 : OAI211_X1 port map( C1 => n2221, C2 => n6170, A => n6523, B => n6522
                           , ZN => n6524);
   U2382 : NOR4_X1 port map( A1 => n6527, A2 => n6526, A3 => n6525, A4 => n6524
                           , ZN => n6528);
   U2383 : OAI21_X1 port map( B1 => n2623, B2 => n6173, A => n6528, ZN => n2984
                           );
   U2384 : OAI222_X1 port map( A1 => n972, A2 => n6121, B1 => n2720, B2 => 
                           n6119, C1 => n2126, C2 => n6116, ZN => n6540);
   U2385 : INV_X1 port map( A => n2158, ZN => n7555);
   U2386 : AOI22_X1 port map( A1 => n6127, A2 => n5035, B1 => n6124, B2 => 
                           n7555, ZN => n6529);
   U2387 : OAI221_X1 port map( B1 => n2062, B2 => n6133, C1 => n2094, C2 => 
                           n6130, A => n6529, ZN => n6539);
   U2388 : AOI22_X1 port map( A1 => n6138, A2 => n5032, B1 => n6135, B2 => n982
                           , ZN => n6530);
   U2389 : OAI221_X1 port map( B1 => n6344, B2 => n6144, C1 => n3648, C2 => 
                           n6141, A => n6530, ZN => n6538);
   U2390 : AOI22_X1 port map( A1 => n2912, A2 => n6149, B1 => n6971, B2 => 
                           n6146, ZN => n6531);
   U2391 : OAI221_X1 port map( B1 => n4809, B2 => n6155, C1 => n6973, C2 => 
                           n6152, A => n6531, ZN => n6534);
   U2392 : NAND2_X1 port map( A1 => n6160, A2 => n6975, ZN => n6532);
   U2393 : NAND4_X1 port map( A1 => n1958, A2 => n1959, A3 => n1957, A4 => 
                           n6532, ZN => n6533);
   U2394 : OAI21_X1 port map( B1 => n6534, B2 => n6533, A => n6163, ZN => n6536
                           );
   U2395 : AOI22_X1 port map( A1 => n6167, A2 => n6969, B1 => n6164, B2 => 
                           n4941, ZN => n6535);
   U2396 : OAI211_X1 port map( C1 => n2222, C2 => n6170, A => n6536, B => n6535
                           , ZN => n6537);
   U2397 : NOR4_X1 port map( A1 => n6540, A2 => n6539, A3 => n6538, A4 => n6537
                           , ZN => n6541);
   U2398 : OAI21_X1 port map( B1 => n2624, B2 => n6175, A => n6541, ZN => n2985
                           );
   U2399 : OAI222_X1 port map( A1 => n988, A2 => n6121, B1 => n2721, B2 => 
                           n6119, C1 => n2127, C2 => n6116, ZN => n6553);
   U2400 : INV_X1 port map( A => n2159, ZN => n7556);
   U2401 : AOI22_X1 port map( A1 => n6127, A2 => n5034, B1 => n6124, B2 => 
                           n7556, ZN => n6542);
   U2402 : OAI221_X1 port map( B1 => n2063, B2 => n6133, C1 => n2095, C2 => 
                           n6130, A => n6542, ZN => n6552);
   U2403 : AOI22_X1 port map( A1 => n6138, A2 => n5031, B1 => n6135, B2 => n998
                           , ZN => n6543);
   U2404 : OAI221_X1 port map( B1 => n6346, B2 => n6144, C1 => n3649, C2 => 
                           n6141, A => n6543, ZN => n6551);
   U2405 : AOI22_X1 port map( A1 => n2913, A2 => n6149, B1 => n6989, B2 => 
                           n6146, ZN => n6544);
   U2406 : OAI221_X1 port map( B1 => n4807, B2 => n6155, C1 => n6991, C2 => 
                           n6152, A => n6544, ZN => n6547);
   U2407 : NAND2_X1 port map( A1 => n6160, A2 => n6993, ZN => n6545);
   U2408 : NAND4_X1 port map( A1 => n1941, A2 => n1942, A3 => n1940, A4 => 
                           n6545, ZN => n6546);
   U2409 : OAI21_X1 port map( B1 => n6547, B2 => n6546, A => n6163, ZN => n6549
                           );
   U2410 : AOI22_X1 port map( A1 => n6167, A2 => n6987, B1 => n6164, B2 => 
                           n4940, ZN => n6548);
   U2411 : OAI211_X1 port map( C1 => n2223, C2 => n6170, A => n6549, B => n6548
                           , ZN => n6550);
   U2412 : NOR4_X1 port map( A1 => n6553, A2 => n6552, A3 => n6551, A4 => n6550
                           , ZN => n6554);
   U2413 : OAI21_X1 port map( B1 => n2625, B2 => n6175, A => n6554, ZN => n2986
                           );
   U2414 : OAI222_X1 port map( A1 => n4699, A2 => n6121, B1 => n2722, B2 => 
                           n6119, C1 => n2128, C2 => n6116, ZN => n6566);
   U2415 : INV_X1 port map( A => n2160, ZN => n7557);
   U2416 : AOI22_X1 port map( A1 => n6127, A2 => n2850, B1 => n6124, B2 => 
                           n7557, ZN => n6555);
   U2417 : OAI221_X1 port map( B1 => n2064, B2 => n6133, C1 => n2096, C2 => 
                           n6130, A => n6555, ZN => n6565);
   U2418 : AOI22_X1 port map( A1 => n6138, A2 => n5030, B1 => n6135, B2 => 
                           n4970, ZN => n6556);
   U2419 : OAI221_X1 port map( B1 => n6347, B2 => n6144, C1 => n3650, C2 => 
                           n6141, A => n6556, ZN => n6564);
   U2420 : AOI22_X1 port map( A1 => n2914, A2 => n6149, B1 => n7008, B2 => 
                           n6146, ZN => n6557);
   U2421 : OAI221_X1 port map( B1 => n4805, B2 => n6155, C1 => n7010, C2 => 
                           n6152, A => n6557, ZN => n6560);
   U2422 : NAND2_X1 port map( A1 => n6160, A2 => n7012, ZN => n6558);
   U2423 : NAND4_X1 port map( A1 => n1924, A2 => n1925, A3 => n1923, A4 => 
                           n6558, ZN => n6559);
   U2424 : OAI21_X1 port map( B1 => n6560, B2 => n6559, A => n6163, ZN => n6562
                           );
   U2425 : AOI22_X1 port map( A1 => n6167, A2 => n7006, B1 => n6164, B2 => 
                           n4939, ZN => n6561);
   U2426 : OAI211_X1 port map( C1 => n2224, C2 => n6170, A => n6562, B => n6561
                           , ZN => n6563);
   U2427 : NOR4_X1 port map( A1 => n6566, A2 => n6565, A3 => n6564, A4 => n6563
                           , ZN => n6567);
   U2428 : OAI21_X1 port map( B1 => n2626, B2 => n6175, A => n6567, ZN => n2987
                           );
   U2429 : OAI222_X1 port map( A1 => n4697, A2 => n6121, B1 => n2723, B2 => 
                           n6119, C1 => n2129, C2 => n6116, ZN => n6579);
   U2430 : INV_X1 port map( A => n2161, ZN => n7558);
   U2431 : AOI22_X1 port map( A1 => n6127, A2 => n2851, B1 => n6124, B2 => 
                           n7558, ZN => n6568);
   U2432 : OAI221_X1 port map( B1 => n2065, B2 => n6133, C1 => n2097, C2 => 
                           n6130, A => n6568, ZN => n6578);
   U2433 : AOI22_X1 port map( A1 => n6138, A2 => n5029, B1 => n6135, B2 => 
                           n4969, ZN => n6569);
   U2434 : OAI221_X1 port map( B1 => n6348, B2 => n6144, C1 => n3651, C2 => 
                           n6141, A => n6569, ZN => n6577);
   U2435 : AOI22_X1 port map( A1 => n2915, A2 => n6149, B1 => n7027, B2 => 
                           n6146, ZN => n6570);
   U2436 : OAI221_X1 port map( B1 => n4803, B2 => n6155, C1 => n7029, C2 => 
                           n6152, A => n6570, ZN => n6573);
   U2437 : NAND2_X1 port map( A1 => n6160, A2 => n7031, ZN => n6571);
   U2438 : NAND4_X1 port map( A1 => n1907, A2 => n1908, A3 => n1906, A4 => 
                           n6571, ZN => n6572);
   U2439 : OAI21_X1 port map( B1 => n6573, B2 => n6572, A => n6163, ZN => n6575
                           );
   U2440 : AOI22_X1 port map( A1 => n6167, A2 => n7025, B1 => n6164, B2 => 
                           n4938, ZN => n6574);
   U2441 : OAI211_X1 port map( C1 => n2225, C2 => n6170, A => n6575, B => n6574
                           , ZN => n6576);
   U2442 : NOR4_X1 port map( A1 => n6579, A2 => n6578, A3 => n6577, A4 => n6576
                           , ZN => n6580);
   U2443 : OAI21_X1 port map( B1 => n2627, B2 => n6175, A => n6580, ZN => n2988
                           );
   U2444 : OAI222_X1 port map( A1 => n4705, A2 => n6121, B1 => n2724, B2 => 
                           n6119, C1 => n2130, C2 => n6116, ZN => n6592);
   U2445 : INV_X1 port map( A => n2162, ZN => n7559);
   U2446 : AOI22_X1 port map( A1 => n6127, A2 => n2852, B1 => n6124, B2 => 
                           n7559, ZN => n6581);
   U2447 : OAI221_X1 port map( B1 => n2066, B2 => n6133, C1 => n2098, C2 => 
                           n6130, A => n6581, ZN => n6591);
   U2448 : AOI22_X1 port map( A1 => n6138, A2 => n5028, B1 => n6135, B2 => 
                           n4968, ZN => n6582);
   U2449 : OAI221_X1 port map( B1 => n6349, B2 => n6144, C1 => n3652, C2 => 
                           n6141, A => n6582, ZN => n6590);
   U2450 : AOI22_X1 port map( A1 => n2916, A2 => n6149, B1 => n7046, B2 => 
                           n6146, ZN => n6583);
   U2451 : OAI221_X1 port map( B1 => n4801, B2 => n6155, C1 => n7048, C2 => 
                           n6152, A => n6583, ZN => n6586);
   U2452 : NAND2_X1 port map( A1 => n6160, A2 => n7050, ZN => n6584);
   U2453 : NAND4_X1 port map( A1 => n1890, A2 => n1891, A3 => n1889, A4 => 
                           n6584, ZN => n6585);
   U2454 : OAI21_X1 port map( B1 => n6586, B2 => n6585, A => n6163, ZN => n6588
                           );
   U2455 : AOI22_X1 port map( A1 => n6167, A2 => n7044, B1 => n6164, B2 => 
                           n4937, ZN => n6587);
   U2456 : OAI211_X1 port map( C1 => n2226, C2 => n6170, A => n6588, B => n6587
                           , ZN => n6589);
   U2457 : NOR4_X1 port map( A1 => n6592, A2 => n6591, A3 => n6590, A4 => n6589
                           , ZN => n6593);
   U2458 : OAI21_X1 port map( B1 => n2628, B2 => n6175, A => n6593, ZN => n2989
                           );
   U2459 : OAI222_X1 port map( A1 => n4703, A2 => n6121, B1 => n2725, B2 => 
                           n6119, C1 => n2131, C2 => n6116, ZN => n6605);
   U2460 : INV_X1 port map( A => n2163, ZN => n7560);
   U2461 : AOI22_X1 port map( A1 => n6127, A2 => n2853, B1 => n6124, B2 => 
                           n7560, ZN => n6594);
   U2462 : OAI221_X1 port map( B1 => n2067, B2 => n6133, C1 => n2099, C2 => 
                           n6130, A => n6594, ZN => n6604);
   U2463 : AOI22_X1 port map( A1 => n6138, A2 => n5027, B1 => n6135, B2 => 
                           n4967, ZN => n6595);
   U2464 : OAI221_X1 port map( B1 => n6350, B2 => n6144, C1 => n3653, C2 => 
                           n6141, A => n6595, ZN => n6603);
   U2465 : AOI22_X1 port map( A1 => n2917, A2 => n6149, B1 => n7065, B2 => 
                           n6146, ZN => n6596);
   U2466 : OAI221_X1 port map( B1 => n4799, B2 => n6155, C1 => n7067, C2 => 
                           n6152, A => n6596, ZN => n6599);
   U2467 : NAND2_X1 port map( A1 => n6160, A2 => n7069, ZN => n6597);
   U2468 : NAND4_X1 port map( A1 => n1873, A2 => n1874, A3 => n1872, A4 => 
                           n6597, ZN => n6598);
   U2469 : OAI21_X1 port map( B1 => n6599, B2 => n6598, A => n6163, ZN => n6601
                           );
   U2470 : AOI22_X1 port map( A1 => n6167, A2 => n7063, B1 => n6164, B2 => 
                           n4936, ZN => n6600);
   U2471 : OAI211_X1 port map( C1 => n2227, C2 => n6170, A => n6601, B => n6600
                           , ZN => n6602);
   U2472 : NOR4_X1 port map( A1 => n6605, A2 => n6604, A3 => n6603, A4 => n6602
                           , ZN => n6606);
   U2473 : OAI21_X1 port map( B1 => n2629, B2 => n6175, A => n6606, ZN => n2990
                           );
   U2474 : OAI222_X1 port map( A1 => n4701, A2 => n6121, B1 => n2726, B2 => 
                           n6119, C1 => n2132, C2 => n6116, ZN => n6618);
   U2475 : INV_X1 port map( A => n2164, ZN => n7561);
   U2476 : AOI22_X1 port map( A1 => n6127, A2 => n2854, B1 => n6124, B2 => 
                           n7561, ZN => n6607);
   U2477 : OAI221_X1 port map( B1 => n2068, B2 => n6133, C1 => n2100, C2 => 
                           n6130, A => n6607, ZN => n6617);
   U2478 : AOI22_X1 port map( A1 => n6138, A2 => n5026, B1 => n6135, B2 => 
                           n4966, ZN => n6608);
   U2479 : OAI221_X1 port map( B1 => n6351, B2 => n6144, C1 => n3654, C2 => 
                           n6141, A => n6608, ZN => n6616);
   U2480 : AOI22_X1 port map( A1 => n2918, A2 => n6149, B1 => n7084, B2 => 
                           n6146, ZN => n6609);
   U2481 : OAI221_X1 port map( B1 => n4797, B2 => n6155, C1 => n7086, C2 => 
                           n6152, A => n6609, ZN => n6612);
   U2482 : NAND2_X1 port map( A1 => n6159, A2 => n7088, ZN => n6610);
   U2483 : NAND4_X1 port map( A1 => n1856, A2 => n1857, A3 => n1855, A4 => 
                           n6610, ZN => n6611);
   U2484 : OAI21_X1 port map( B1 => n6612, B2 => n6611, A => n6162, ZN => n6614
                           );
   U2485 : AOI22_X1 port map( A1 => n6167, A2 => n7082, B1 => n6164, B2 => 
                           n4935, ZN => n6613);
   U2486 : OAI211_X1 port map( C1 => n2228, C2 => n6170, A => n6614, B => n6613
                           , ZN => n6615);
   U2487 : NOR4_X1 port map( A1 => n6618, A2 => n6617, A3 => n6616, A4 => n6615
                           , ZN => n6619);
   U2488 : OAI21_X1 port map( B1 => n2630, B2 => n6175, A => n6619, ZN => n2991
                           );
   U2489 : OAI222_X1 port map( A1 => n4711, A2 => n6121, B1 => n2727, B2 => 
                           n6119, C1 => n2133, C2 => n6116, ZN => n6631);
   U2490 : INV_X1 port map( A => n2165, ZN => n7562);
   U2491 : AOI22_X1 port map( A1 => n6127, A2 => n2855, B1 => n6124, B2 => 
                           n7562, ZN => n6620);
   U2492 : OAI221_X1 port map( B1 => n2069, B2 => n6133, C1 => n2101, C2 => 
                           n6130, A => n6620, ZN => n6630);
   U2493 : AOI22_X1 port map( A1 => n6138, A2 => n5025, B1 => n6135, B2 => 
                           n4965, ZN => n6621);
   U2494 : OAI221_X1 port map( B1 => n6352, B2 => n6144, C1 => n3655, C2 => 
                           n6141, A => n6621, ZN => n6629);
   U2495 : AOI22_X1 port map( A1 => n2919, A2 => n6149, B1 => n7103, B2 => 
                           n6146, ZN => n6622);
   U2496 : OAI221_X1 port map( B1 => n4795, B2 => n6155, C1 => n7105, C2 => 
                           n6152, A => n6622, ZN => n6625);
   U2497 : NAND2_X1 port map( A1 => n6159, A2 => n7107, ZN => n6623);
   U2498 : NAND4_X1 port map( A1 => n1839, A2 => n1840, A3 => n1838, A4 => 
                           n6623, ZN => n6624);
   U2499 : OAI21_X1 port map( B1 => n6625, B2 => n6624, A => n6162, ZN => n6627
                           );
   U2500 : AOI22_X1 port map( A1 => n6167, A2 => n7101, B1 => n6164, B2 => 
                           n4934, ZN => n6626);
   U2501 : OAI211_X1 port map( C1 => n2229, C2 => n6170, A => n6627, B => n6626
                           , ZN => n6628);
   U2502 : NOR4_X1 port map( A1 => n6631, A2 => n6630, A3 => n6629, A4 => n6628
                           , ZN => n6632);
   U2503 : OAI21_X1 port map( B1 => n2631, B2 => n6175, A => n6632, ZN => n2992
                           );
   U2504 : OAI222_X1 port map( A1 => n4709, A2 => n6121, B1 => n2728, B2 => 
                           n6119, C1 => n2134, C2 => n6116, ZN => n6644);
   U2505 : INV_X1 port map( A => n2166, ZN => n7563);
   U2506 : AOI22_X1 port map( A1 => n6127, A2 => n2856, B1 => n6124, B2 => 
                           n7563, ZN => n6633);
   U2507 : OAI221_X1 port map( B1 => n2070, B2 => n6133, C1 => n2102, C2 => 
                           n6130, A => n6633, ZN => n6643);
   U2508 : AOI22_X1 port map( A1 => n6138, A2 => n5024, B1 => n6135, B2 => 
                           n4964, ZN => n6634);
   U2509 : OAI221_X1 port map( B1 => n6353, B2 => n6144, C1 => n3656, C2 => 
                           n6141, A => n6634, ZN => n6642);
   U2510 : AOI22_X1 port map( A1 => n2920, A2 => n6149, B1 => n7122, B2 => 
                           n6146, ZN => n6635);
   U2511 : OAI221_X1 port map( B1 => n4793, B2 => n6155, C1 => n7124, C2 => 
                           n6152, A => n6635, ZN => n6638);
   U2512 : NAND2_X1 port map( A1 => n6159, A2 => n7126, ZN => n6636);
   U2513 : NAND4_X1 port map( A1 => n1822, A2 => n1823, A3 => n1821, A4 => 
                           n6636, ZN => n6637);
   U2514 : OAI21_X1 port map( B1 => n6638, B2 => n6637, A => n6162, ZN => n6640
                           );
   U2515 : AOI22_X1 port map( A1 => n6167, A2 => n7120, B1 => n6164, B2 => 
                           n4933, ZN => n6639);
   U2516 : OAI211_X1 port map( C1 => n2230, C2 => n6170, A => n6640, B => n6639
                           , ZN => n6641);
   U2517 : NOR4_X1 port map( A1 => n6644, A2 => n6643, A3 => n6642, A4 => n6641
                           , ZN => n6645);
   U2518 : OAI21_X1 port map( B1 => n2632, B2 => n6175, A => n6645, ZN => n2993
                           );
   U2519 : OAI222_X1 port map( A1 => n4707, A2 => n6121, B1 => n2729, B2 => 
                           n6119, C1 => n2135, C2 => n6116, ZN => n6657);
   U2520 : INV_X1 port map( A => n2167, ZN => n7564);
   U2521 : AOI22_X1 port map( A1 => n6127, A2 => n2857, B1 => n6124, B2 => 
                           n7564, ZN => n6646);
   U2522 : OAI221_X1 port map( B1 => n2071, B2 => n6133, C1 => n2103, C2 => 
                           n6130, A => n6646, ZN => n6656);
   U2523 : AOI22_X1 port map( A1 => n6138, A2 => n5023, B1 => n6135, B2 => 
                           n4963, ZN => n6647);
   U2524 : OAI221_X1 port map( B1 => n6354, B2 => n6144, C1 => n3657, C2 => 
                           n6141, A => n6647, ZN => n6655);
   U2525 : AOI22_X1 port map( A1 => n2921, A2 => n6149, B1 => n7141, B2 => 
                           n6146, ZN => n6648);
   U2526 : OAI221_X1 port map( B1 => n4791, B2 => n6155, C1 => n7143, C2 => 
                           n6152, A => n6648, ZN => n6651);
   U2527 : NAND2_X1 port map( A1 => n6159, A2 => n7145, ZN => n6649);
   U2528 : NAND4_X1 port map( A1 => n1805, A2 => n1806, A3 => n1804, A4 => 
                           n6649, ZN => n6650);
   U2529 : OAI21_X1 port map( B1 => n6651, B2 => n6650, A => n6162, ZN => n6653
                           );
   U2530 : AOI22_X1 port map( A1 => n6167, A2 => n7139, B1 => n6164, B2 => 
                           n4932, ZN => n6652);
   U2531 : OAI211_X1 port map( C1 => n2231, C2 => n6170, A => n6653, B => n6652
                           , ZN => n6654);
   U2532 : NOR4_X1 port map( A1 => n6657, A2 => n6656, A3 => n6655, A4 => n6654
                           , ZN => n6658);
   U2533 : OAI21_X1 port map( B1 => n2633, B2 => n6175, A => n6658, ZN => n2994
                           );
   U2534 : OAI222_X1 port map( A1 => n4717, A2 => n6122, B1 => n2730, B2 => 
                           n6119, C1 => n2136, C2 => n6117, ZN => n6670);
   U2535 : INV_X1 port map( A => n2168, ZN => n7565);
   U2536 : AOI22_X1 port map( A1 => n6127, A2 => n2858, B1 => n6125, B2 => 
                           n7565, ZN => n6659);
   U2537 : OAI221_X1 port map( B1 => n2072, B2 => n6133, C1 => n2104, C2 => 
                           n6131, A => n6659, ZN => n6669);
   U2538 : AOI22_X1 port map( A1 => n6138, A2 => n5022, B1 => n6136, B2 => 
                           n4962, ZN => n6660);
   U2539 : OAI221_X1 port map( B1 => n6355, B2 => n6144, C1 => n3658, C2 => 
                           n6142, A => n6660, ZN => n6668);
   U2540 : AOI22_X1 port map( A1 => n2922, A2 => n6150, B1 => n7160, B2 => 
                           n6147, ZN => n6661);
   U2541 : OAI221_X1 port map( B1 => n4789, B2 => n6156, C1 => n7162, C2 => 
                           n6153, A => n6661, ZN => n6664);
   U2542 : NAND2_X1 port map( A1 => n6159, A2 => n7164, ZN => n6662);
   U2543 : NAND4_X1 port map( A1 => n1788, A2 => n1789, A3 => n1787, A4 => 
                           n6662, ZN => n6663);
   U2544 : OAI21_X1 port map( B1 => n6664, B2 => n6663, A => n6162, ZN => n6666
                           );
   U2545 : AOI22_X1 port map( A1 => n6167, A2 => n7158, B1 => n6165, B2 => 
                           n4931, ZN => n6665);
   U2546 : OAI211_X1 port map( C1 => n2232, C2 => n6171, A => n6666, B => n6665
                           , ZN => n6667);
   U2547 : NOR4_X1 port map( A1 => n6670, A2 => n6669, A3 => n6668, A4 => n6667
                           , ZN => n6671);
   U2548 : OAI21_X1 port map( B1 => n2634, B2 => n6174, A => n6671, ZN => n2995
                           );
   U2549 : OAI222_X1 port map( A1 => n4715, A2 => n6122, B1 => n2731, B2 => 
                           n6120, C1 => n2137, C2 => n6117, ZN => n6683);
   U2550 : INV_X1 port map( A => n2169, ZN => n7566);
   U2551 : AOI22_X1 port map( A1 => n6128, A2 => n2859, B1 => n6125, B2 => 
                           n7566, ZN => n6672);
   U2552 : OAI221_X1 port map( B1 => n2073, B2 => n6134, C1 => n2105, C2 => 
                           n6131, A => n6672, ZN => n6682);
   U2553 : AOI22_X1 port map( A1 => n6139, A2 => n5021, B1 => n6136, B2 => 
                           n4961, ZN => n6673);
   U2554 : OAI221_X1 port map( B1 => n6356, B2 => n6145, C1 => n3659, C2 => 
                           n6142, A => n6673, ZN => n6681);
   U2555 : AOI22_X1 port map( A1 => n2923, A2 => n6150, B1 => n7179, B2 => 
                           n6147, ZN => n6674);
   U2556 : OAI221_X1 port map( B1 => n4787, B2 => n6156, C1 => n7181, C2 => 
                           n6153, A => n6674, ZN => n6677);
   U2557 : NAND2_X1 port map( A1 => n6159, A2 => n7183, ZN => n6675);
   U2558 : NAND4_X1 port map( A1 => n1771, A2 => n1772, A3 => n1770, A4 => 
                           n6675, ZN => n6676);
   U2559 : OAI21_X1 port map( B1 => n6677, B2 => n6676, A => n6162, ZN => n6679
                           );
   U2560 : AOI22_X1 port map( A1 => n6168, A2 => n7177, B1 => n6165, B2 => 
                           n4930, ZN => n6678);
   U2561 : OAI211_X1 port map( C1 => n2233, C2 => n6171, A => n6679, B => n6678
                           , ZN => n6680);
   U2562 : NOR4_X1 port map( A1 => n6683, A2 => n6682, A3 => n6681, A4 => n6680
                           , ZN => n6684);
   U2563 : OAI21_X1 port map( B1 => n2635, B2 => n6174, A => n6684, ZN => n2996
                           );
   U2564 : OAI222_X1 port map( A1 => n4713, A2 => n6122, B1 => n2732, B2 => 
                           n6120, C1 => n2138, C2 => n6117, ZN => n6696);
   U2565 : INV_X1 port map( A => n2170, ZN => n7567);
   U2566 : AOI22_X1 port map( A1 => n6128, A2 => n2860, B1 => n6125, B2 => 
                           n7567, ZN => n6685);
   U2567 : OAI221_X1 port map( B1 => n2074, B2 => n6134, C1 => n2106, C2 => 
                           n6131, A => n6685, ZN => n6695);
   U2568 : AOI22_X1 port map( A1 => n6139, A2 => n5020, B1 => n6136, B2 => 
                           n4960, ZN => n6686);
   U2569 : OAI221_X1 port map( B1 => n6357, B2 => n6145, C1 => n3660, C2 => 
                           n6142, A => n6686, ZN => n6694);
   U2570 : AOI22_X1 port map( A1 => n2924, A2 => n6150, B1 => n7198, B2 => 
                           n6147, ZN => n6687);
   U2571 : OAI221_X1 port map( B1 => n4785, B2 => n6156, C1 => n7200, C2 => 
                           n6153, A => n6687, ZN => n6690);
   U2572 : NAND2_X1 port map( A1 => n6159, A2 => n7202, ZN => n6688);
   U2573 : NAND4_X1 port map( A1 => n1754, A2 => n1755, A3 => n1753, A4 => 
                           n6688, ZN => n6689);
   U2574 : OAI21_X1 port map( B1 => n6690, B2 => n6689, A => n6162, ZN => n6692
                           );
   U2575 : AOI22_X1 port map( A1 => n6168, A2 => n7196, B1 => n6165, B2 => 
                           n4929, ZN => n6691);
   U2576 : OAI211_X1 port map( C1 => n2234, C2 => n6171, A => n6692, B => n6691
                           , ZN => n6693);
   U2577 : NOR4_X1 port map( A1 => n6696, A2 => n6695, A3 => n6694, A4 => n6693
                           , ZN => n6697);
   U2578 : OAI21_X1 port map( B1 => n2636, B2 => n6174, A => n6697, ZN => n2997
                           );
   U2579 : OAI222_X1 port map( A1 => n4723, A2 => n6122, B1 => n2733, B2 => 
                           n6120, C1 => n2139, C2 => n6117, ZN => n6709);
   U2580 : INV_X1 port map( A => n2171, ZN => n7568);
   U2581 : AOI22_X1 port map( A1 => n6128, A2 => n2861, B1 => n6125, B2 => 
                           n7568, ZN => n6698);
   U2582 : OAI221_X1 port map( B1 => n2075, B2 => n6134, C1 => n2107, C2 => 
                           n6131, A => n6698, ZN => n6708);
   U2583 : AOI22_X1 port map( A1 => n6139, A2 => n5019, B1 => n6136, B2 => 
                           n4959, ZN => n6699);
   U2584 : OAI221_X1 port map( B1 => n6358, B2 => n6145, C1 => n3661, C2 => 
                           n6142, A => n6699, ZN => n6707);
   U2585 : AOI22_X1 port map( A1 => n2925, A2 => n6150, B1 => n7217, B2 => 
                           n6147, ZN => n6700);
   U2586 : OAI221_X1 port map( B1 => n4783, B2 => n6156, C1 => n7219, C2 => 
                           n6153, A => n6700, ZN => n6703);
   U2587 : NAND2_X1 port map( A1 => n6159, A2 => n7221, ZN => n6701);
   U2588 : NAND4_X1 port map( A1 => n1737, A2 => n1738, A3 => n1736, A4 => 
                           n6701, ZN => n6702);
   U2589 : OAI21_X1 port map( B1 => n6703, B2 => n6702, A => n6162, ZN => n6705
                           );
   U2590 : AOI22_X1 port map( A1 => n6168, A2 => n7215, B1 => n6165, B2 => 
                           n4928, ZN => n6704);
   U2591 : OAI211_X1 port map( C1 => n2235, C2 => n6171, A => n6705, B => n6704
                           , ZN => n6706);
   U2592 : NOR4_X1 port map( A1 => n6709, A2 => n6708, A3 => n6707, A4 => n6706
                           , ZN => n6710);
   U2593 : OAI21_X1 port map( B1 => n2637, B2 => n6174, A => n6710, ZN => n2998
                           );
   U2594 : OAI222_X1 port map( A1 => n4721, A2 => n6122, B1 => n2734, B2 => 
                           n6120, C1 => n2140, C2 => n6117, ZN => n6722);
   U2595 : INV_X1 port map( A => n2172, ZN => n7569);
   U2596 : AOI22_X1 port map( A1 => n6128, A2 => n2862, B1 => n6125, B2 => 
                           n7569, ZN => n6711);
   U2597 : OAI221_X1 port map( B1 => n2076, B2 => n6134, C1 => n2108, C2 => 
                           n6131, A => n6711, ZN => n6721);
   U2598 : AOI22_X1 port map( A1 => n6139, A2 => n5018, B1 => n6136, B2 => 
                           n4958, ZN => n6712);
   U2599 : OAI221_X1 port map( B1 => n6359, B2 => n6145, C1 => n3662, C2 => 
                           n6142, A => n6712, ZN => n6720);
   U2600 : AOI22_X1 port map( A1 => n2926, A2 => n6150, B1 => n7236, B2 => 
                           n6147, ZN => n6713);
   U2601 : OAI221_X1 port map( B1 => n4753, B2 => n6156, C1 => n7238, C2 => 
                           n6153, A => n6713, ZN => n6716);
   U2602 : NAND2_X1 port map( A1 => n6159, A2 => n7240, ZN => n6714);
   U2603 : NAND4_X1 port map( A1 => n1720, A2 => n1721, A3 => n1719, A4 => 
                           n6714, ZN => n6715);
   U2604 : OAI21_X1 port map( B1 => n6716, B2 => n6715, A => n6162, ZN => n6718
                           );
   U2605 : AOI22_X1 port map( A1 => n6168, A2 => n7234, B1 => n6165, B2 => 
                           n4927, ZN => n6717);
   U2606 : OAI211_X1 port map( C1 => n2236, C2 => n6171, A => n6718, B => n6717
                           , ZN => n6719);
   U2607 : NOR4_X1 port map( A1 => n6722, A2 => n6721, A3 => n6720, A4 => n6719
                           , ZN => n6723);
   U2608 : OAI21_X1 port map( B1 => n2638, B2 => n6174, A => n6723, ZN => n2999
                           );
   U2609 : OAI222_X1 port map( A1 => n4719, A2 => n6122, B1 => n2735, B2 => 
                           n6120, C1 => n2141, C2 => n6117, ZN => n6735);
   U2610 : INV_X1 port map( A => n2173, ZN => n7570);
   U2611 : AOI22_X1 port map( A1 => n6128, A2 => n2863, B1 => n6125, B2 => 
                           n7570, ZN => n6724);
   U2612 : OAI221_X1 port map( B1 => n2077, B2 => n6134, C1 => n2109, C2 => 
                           n6131, A => n6724, ZN => n6734);
   U2613 : AOI22_X1 port map( A1 => n6139, A2 => n5017, B1 => n6136, B2 => 
                           n4957, ZN => n6725);
   U2614 : OAI221_X1 port map( B1 => n6360, B2 => n6145, C1 => n3663, C2 => 
                           n6142, A => n6725, ZN => n6733);
   U2615 : AOI22_X1 port map( A1 => n2927, A2 => n6150, B1 => n7255, B2 => 
                           n6147, ZN => n6726);
   U2616 : OAI221_X1 port map( B1 => n4763, B2 => n6156, C1 => n7257, C2 => 
                           n6153, A => n6726, ZN => n6729);
   U2617 : NAND2_X1 port map( A1 => n6159, A2 => n7259, ZN => n6727);
   U2618 : NAND4_X1 port map( A1 => n1703, A2 => n1704, A3 => n1702, A4 => 
                           n6727, ZN => n6728);
   U2619 : OAI21_X1 port map( B1 => n6729, B2 => n6728, A => n6162, ZN => n6731
                           );
   U2620 : AOI22_X1 port map( A1 => n6168, A2 => n7253, B1 => n6165, B2 => 
                           n4926, ZN => n6730);
   U2621 : OAI211_X1 port map( C1 => n2237, C2 => n6171, A => n6731, B => n6730
                           , ZN => n6732);
   U2622 : NOR4_X1 port map( A1 => n6735, A2 => n6734, A3 => n6733, A4 => n6732
                           , ZN => n6736);
   U2623 : OAI21_X1 port map( B1 => n2639, B2 => n6174, A => n6736, ZN => n3000
                           );
   U2624 : OAI222_X1 port map( A1 => n4729, A2 => n6122, B1 => n2736, B2 => 
                           n6120, C1 => n2142, C2 => n6117, ZN => n6748);
   U2625 : INV_X1 port map( A => n2174, ZN => n7571);
   U2626 : AOI22_X1 port map( A1 => n6128, A2 => n2864, B1 => n6125, B2 => 
                           n7571, ZN => n6737);
   U2627 : OAI221_X1 port map( B1 => n2078, B2 => n6134, C1 => n2110, C2 => 
                           n6131, A => n6737, ZN => n6747);
   U2628 : AOI22_X1 port map( A1 => n6139, A2 => n5016, B1 => n6136, B2 => 
                           n4956, ZN => n6738);
   U2629 : OAI221_X1 port map( B1 => n6361, B2 => n6145, C1 => n3664, C2 => 
                           n6142, A => n6738, ZN => n6746);
   U2630 : AOI22_X1 port map( A1 => n2928, A2 => n6150, B1 => n7274, B2 => 
                           n6147, ZN => n6739);
   U2631 : OAI221_X1 port map( B1 => n4757, B2 => n6156, C1 => n7276, C2 => 
                           n6153, A => n6739, ZN => n6742);
   U2632 : NAND2_X1 port map( A1 => n6159, A2 => n7278, ZN => n6740);
   U2633 : NAND4_X1 port map( A1 => n1686, A2 => n1687, A3 => n1685, A4 => 
                           n6740, ZN => n6741);
   U2634 : OAI21_X1 port map( B1 => n6742, B2 => n6741, A => n6162, ZN => n6744
                           );
   U2635 : AOI22_X1 port map( A1 => n6168, A2 => n7272, B1 => n6165, B2 => 
                           n4925, ZN => n6743);
   U2636 : OAI211_X1 port map( C1 => n2238, C2 => n6171, A => n6744, B => n6743
                           , ZN => n6745);
   U2637 : NOR4_X1 port map( A1 => n6748, A2 => n6747, A3 => n6746, A4 => n6745
                           , ZN => n6749);
   U2638 : OAI21_X1 port map( B1 => n2640, B2 => n6174, A => n6749, ZN => n3001
                           );
   U2639 : OAI222_X1 port map( A1 => n4727, A2 => n6122, B1 => n2737, B2 => 
                           n6120, C1 => n2143, C2 => n6117, ZN => n6761);
   U2640 : INV_X1 port map( A => n2175, ZN => n7572);
   U2641 : AOI22_X1 port map( A1 => n6128, A2 => n2865, B1 => n6125, B2 => 
                           n7572, ZN => n6750);
   U2642 : OAI221_X1 port map( B1 => n2079, B2 => n6134, C1 => n2111, C2 => 
                           n6131, A => n6750, ZN => n6760);
   U2643 : AOI22_X1 port map( A1 => n6139, A2 => n5015, B1 => n6136, B2 => 
                           n4955, ZN => n6751);
   U2644 : OAI221_X1 port map( B1 => n6362, B2 => n6145, C1 => n3665, C2 => 
                           n6142, A => n6751, ZN => n6759);
   U2645 : AOI22_X1 port map( A1 => n2929, A2 => n6150, B1 => n7293, B2 => 
                           n6147, ZN => n6752);
   U2646 : OAI221_X1 port map( B1 => n4759, B2 => n6156, C1 => n7295, C2 => 
                           n6153, A => n6752, ZN => n6755);
   U2647 : NAND2_X1 port map( A1 => n6159, A2 => n7297, ZN => n6753);
   U2648 : NAND4_X1 port map( A1 => n1669, A2 => n1670, A3 => n1668, A4 => 
                           n6753, ZN => n6754);
   U2649 : OAI21_X1 port map( B1 => n6755, B2 => n6754, A => n6161, ZN => n6757
                           );
   U2650 : AOI22_X1 port map( A1 => n6168, A2 => n7291, B1 => n6165, B2 => 
                           n4924, ZN => n6756);
   U2651 : OAI211_X1 port map( C1 => n2239, C2 => n6171, A => n6757, B => n6756
                           , ZN => n6758);
   U2652 : NOR4_X1 port map( A1 => n6761, A2 => n6760, A3 => n6759, A4 => n6758
                           , ZN => n6762);
   U2653 : OAI21_X1 port map( B1 => n2641, B2 => n6174, A => n6762, ZN => n3002
                           );
   U2654 : OAI222_X1 port map( A1 => n4725, A2 => n6122, B1 => n2738, B2 => 
                           n6120, C1 => n2144, C2 => n6117, ZN => n6774);
   U2655 : INV_X1 port map( A => n2176, ZN => n7573);
   U2656 : AOI22_X1 port map( A1 => n6128, A2 => n2866, B1 => n6125, B2 => 
                           n7573, ZN => n6763);
   U2657 : OAI221_X1 port map( B1 => n2080, B2 => n6134, C1 => n2112, C2 => 
                           n6131, A => n6763, ZN => n6773);
   U2658 : AOI22_X1 port map( A1 => n6139, A2 => n5014, B1 => n6136, B2 => 
                           n4954, ZN => n6764);
   U2659 : OAI221_X1 port map( B1 => n6363, B2 => n6145, C1 => n3666, C2 => 
                           n6142, A => n6764, ZN => n6772);
   U2660 : AOI22_X1 port map( A1 => n2930, A2 => n6150, B1 => n7312, B2 => 
                           n6147, ZN => n6765);
   U2661 : OAI221_X1 port map( B1 => n4769, B2 => n6156, C1 => n7314, C2 => 
                           n6153, A => n6765, ZN => n6768);
   U2662 : NAND2_X1 port map( A1 => n6158, A2 => n7316, ZN => n6766);
   U2663 : NAND4_X1 port map( A1 => n1652, A2 => n1653, A3 => n1651, A4 => 
                           n6766, ZN => n6767);
   U2664 : OAI21_X1 port map( B1 => n6768, B2 => n6767, A => n6161, ZN => n6770
                           );
   U2665 : AOI22_X1 port map( A1 => n6168, A2 => n7310, B1 => n6165, B2 => 
                           n4923, ZN => n6769);
   U2666 : OAI211_X1 port map( C1 => n2240, C2 => n6171, A => n6770, B => n6769
                           , ZN => n6771);
   U2667 : NOR4_X1 port map( A1 => n6774, A2 => n6773, A3 => n6772, A4 => n6771
                           , ZN => n6775);
   U2668 : OAI21_X1 port map( B1 => n2642, B2 => n6174, A => n6775, ZN => n3003
                           );
   U2669 : OAI222_X1 port map( A1 => n4735, A2 => n6122, B1 => n2739, B2 => 
                           n6120, C1 => n2145, C2 => n6117, ZN => n6787);
   U2670 : INV_X1 port map( A => n2177, ZN => n7574);
   U2671 : AOI22_X1 port map( A1 => n6128, A2 => n2867, B1 => n6125, B2 => 
                           n7574, ZN => n6776);
   U2672 : OAI221_X1 port map( B1 => n2081, B2 => n6134, C1 => n2113, C2 => 
                           n6131, A => n6776, ZN => n6786);
   U2673 : AOI22_X1 port map( A1 => n6139, A2 => n5013, B1 => n6136, B2 => 
                           n4953, ZN => n6777);
   U2674 : OAI221_X1 port map( B1 => n6364, B2 => n6145, C1 => n3667, C2 => 
                           n6142, A => n6777, ZN => n6785);
   U2675 : AOI22_X1 port map( A1 => n2931, A2 => n6150, B1 => n7331, B2 => 
                           n6147, ZN => n6778);
   U2676 : OAI221_X1 port map( B1 => n4761, B2 => n6156, C1 => n7333, C2 => 
                           n6153, A => n6778, ZN => n6781);
   U2677 : NAND2_X1 port map( A1 => n6158, A2 => n7335, ZN => n6779);
   U2678 : NAND4_X1 port map( A1 => n1635, A2 => n1636, A3 => n1634, A4 => 
                           n6779, ZN => n6780);
   U2679 : OAI21_X1 port map( B1 => n6781, B2 => n6780, A => n6161, ZN => n6783
                           );
   U2680 : AOI22_X1 port map( A1 => n6168, A2 => n7329, B1 => n6165, B2 => 
                           n4922, ZN => n6782);
   U2681 : OAI211_X1 port map( C1 => n2241, C2 => n6171, A => n6783, B => n6782
                           , ZN => n6784);
   U2682 : NOR4_X1 port map( A1 => n6787, A2 => n6786, A3 => n6785, A4 => n6784
                           , ZN => n6788);
   U2683 : OAI21_X1 port map( B1 => n2643, B2 => n6174, A => n6788, ZN => n3004
                           );
   U2684 : OAI222_X1 port map( A1 => n4733, A2 => n6122, B1 => n2740, B2 => 
                           n6120, C1 => n2146, C2 => n6117, ZN => n6800);
   U2685 : INV_X1 port map( A => n2178, ZN => n7575);
   U2686 : AOI22_X1 port map( A1 => n6128, A2 => n2868, B1 => n6125, B2 => 
                           n7575, ZN => n6789);
   U2687 : OAI221_X1 port map( B1 => n2082, B2 => n6134, C1 => n2114, C2 => 
                           n6131, A => n6789, ZN => n6799);
   U2688 : AOI22_X1 port map( A1 => n6139, A2 => n5012, B1 => n6136, B2 => 
                           n4952, ZN => n6790);
   U2689 : OAI221_X1 port map( B1 => n6365, B2 => n6145, C1 => n3668, C2 => 
                           n6142, A => n6790, ZN => n6798);
   U2690 : AOI22_X1 port map( A1 => n2932, A2 => n6150, B1 => n7350, B2 => 
                           n6147, ZN => n6791);
   U2691 : OAI221_X1 port map( B1 => n4765, B2 => n6156, C1 => n7352, C2 => 
                           n6153, A => n6791, ZN => n6794);
   U2692 : NAND2_X1 port map( A1 => n6158, A2 => n7354, ZN => n6792);
   U2693 : NAND4_X1 port map( A1 => n1618, A2 => n1619, A3 => n1617, A4 => 
                           n6792, ZN => n6793);
   U2694 : OAI21_X1 port map( B1 => n6794, B2 => n6793, A => n6161, ZN => n6796
                           );
   U2695 : AOI22_X1 port map( A1 => n6168, A2 => n7348, B1 => n6165, B2 => 
                           n4921, ZN => n6795);
   U2696 : OAI211_X1 port map( C1 => n2242, C2 => n6171, A => n6796, B => n6795
                           , ZN => n6797);
   U2697 : NOR4_X1 port map( A1 => n6800, A2 => n6799, A3 => n6798, A4 => n6797
                           , ZN => n6801);
   U2698 : OAI21_X1 port map( B1 => n2644, B2 => n6174, A => n6801, ZN => n3005
                           );
   U2699 : OAI222_X1 port map( A1 => n4731, A2 => n6122, B1 => n2741, B2 => 
                           n6120, C1 => n2147, C2 => n6117, ZN => n6813);
   U2700 : INV_X1 port map( A => n2179, ZN => n7576);
   U2701 : AOI22_X1 port map( A1 => n6128, A2 => n2869, B1 => n6125, B2 => 
                           n7576, ZN => n6802);
   U2702 : OAI221_X1 port map( B1 => n2083, B2 => n6134, C1 => n2115, C2 => 
                           n6131, A => n6802, ZN => n6812);
   U2703 : AOI22_X1 port map( A1 => n6139, A2 => n5011, B1 => n6136, B2 => 
                           n4951, ZN => n6803);
   U2704 : OAI221_X1 port map( B1 => n6366, B2 => n6145, C1 => n3669, C2 => 
                           n6142, A => n6803, ZN => n6811);
   U2705 : AOI22_X1 port map( A1 => n2933, A2 => n6150, B1 => n7369, B2 => 
                           n6147, ZN => n6804);
   U2706 : OAI221_X1 port map( B1 => n4771, B2 => n6156, C1 => n7371, C2 => 
                           n6153, A => n6804, ZN => n6807);
   U2707 : NAND2_X1 port map( A1 => n6158, A2 => n7373, ZN => n6805);
   U2708 : NAND4_X1 port map( A1 => n1601, A2 => n1602, A3 => n1600, A4 => 
                           n6805, ZN => n6806);
   U2709 : OAI21_X1 port map( B1 => n6807, B2 => n6806, A => n6161, ZN => n6809
                           );
   U2710 : AOI22_X1 port map( A1 => n6168, A2 => n7367, B1 => n6165, B2 => 
                           n4920, ZN => n6808);
   U2711 : OAI211_X1 port map( C1 => n2243, C2 => n6171, A => n6809, B => n6808
                           , ZN => n6810);
   U2712 : NOR4_X1 port map( A1 => n6813, A2 => n6812, A3 => n6811, A4 => n6810
                           , ZN => n6814);
   U2713 : OAI21_X1 port map( B1 => n2645, B2 => n6173, A => n6814, ZN => n3006
                           );
   U2714 : OAI222_X1 port map( A1 => n4741, A2 => n6123, B1 => n2742, B2 => 
                           n6120, C1 => n2148, C2 => n6118, ZN => n6826);
   U2715 : INV_X1 port map( A => n2180, ZN => n7577);
   U2716 : AOI22_X1 port map( A1 => n6128, A2 => n2870, B1 => n6126, B2 => 
                           n7577, ZN => n6815);
   U2717 : OAI221_X1 port map( B1 => n2084, B2 => n6134, C1 => n2116, C2 => 
                           n6132, A => n6815, ZN => n6825);
   U2718 : AOI22_X1 port map( A1 => n6139, A2 => n5010, B1 => n6137, B2 => 
                           n4950, ZN => n6816);
   U2719 : OAI221_X1 port map( B1 => n6367, B2 => n6145, C1 => n3670, C2 => 
                           n6143, A => n6816, ZN => n6824);
   U2720 : AOI22_X1 port map( A1 => n2934, A2 => n6151, B1 => n7388, B2 => 
                           n6148, ZN => n6817);
   U2721 : OAI221_X1 port map( B1 => n4767, B2 => n6157, C1 => n7390, C2 => 
                           n6154, A => n6817, ZN => n6820);
   U2722 : NAND2_X1 port map( A1 => n6158, A2 => n7392, ZN => n6818);
   U2723 : NAND4_X1 port map( A1 => n1584, A2 => n1585, A3 => n1583, A4 => 
                           n6818, ZN => n6819);
   U2724 : OAI21_X1 port map( B1 => n6820, B2 => n6819, A => n6161, ZN => n6822
                           );
   U2725 : AOI22_X1 port map( A1 => n6168, A2 => n7386, B1 => n6166, B2 => 
                           n4919, ZN => n6821);
   U2726 : OAI211_X1 port map( C1 => n2244, C2 => n6172, A => n6822, B => n6821
                           , ZN => n6823);
   U2727 : NOR4_X1 port map( A1 => n6826, A2 => n6825, A3 => n6824, A4 => n6823
                           , ZN => n6827);
   U2728 : OAI21_X1 port map( B1 => n2646, B2 => n6173, A => n6827, ZN => n3007
                           );
   U2729 : OAI222_X1 port map( A1 => n4739, A2 => n6123, B1 => n2743, B2 => 
                           n6119, C1 => n2149, C2 => n6118, ZN => n6839);
   U2730 : INV_X1 port map( A => n2181, ZN => n7578);
   U2731 : AOI22_X1 port map( A1 => n6129, A2 => n2871, B1 => n6126, B2 => 
                           n7578, ZN => n6828);
   U2732 : OAI221_X1 port map( B1 => n2085, B2 => n6133, C1 => n2117, C2 => 
                           n6132, A => n6828, ZN => n6838);
   U2733 : AOI22_X1 port map( A1 => n6140, A2 => n5009, B1 => n6137, B2 => 
                           n4949, ZN => n6829);
   U2734 : OAI221_X1 port map( B1 => n6368, B2 => n6144, C1 => n3671, C2 => 
                           n6143, A => n6829, ZN => n6837);
   U2735 : AOI22_X1 port map( A1 => n2935, A2 => n6151, B1 => n7407, B2 => 
                           n6148, ZN => n6830);
   U2736 : OAI221_X1 port map( B1 => n4775, B2 => n6157, C1 => n7409, C2 => 
                           n6154, A => n6830, ZN => n6833);
   U2737 : NAND2_X1 port map( A1 => n6158, A2 => n7411, ZN => n6831);
   U2738 : NAND4_X1 port map( A1 => n1567, A2 => n1568, A3 => n1566, A4 => 
                           n6831, ZN => n6832);
   U2739 : OAI21_X1 port map( B1 => n6833, B2 => n6832, A => n6161, ZN => n6835
                           );
   U2740 : AOI22_X1 port map( A1 => n6169, A2 => n7405, B1 => n6166, B2 => 
                           n4918, ZN => n6834);
   U2741 : OAI211_X1 port map( C1 => n2245, C2 => n6172, A => n6835, B => n6834
                           , ZN => n6836);
   U2742 : NOR4_X1 port map( A1 => n6839, A2 => n6838, A3 => n6837, A4 => n6836
                           , ZN => n6840);
   U2743 : OAI21_X1 port map( B1 => n2647, B2 => n6173, A => n6840, ZN => n3008
                           );
   U2744 : OAI222_X1 port map( A1 => n4737, A2 => n6123, B1 => n2744, B2 => 
                           n6120, C1 => n2150, C2 => n6118, ZN => n6852);
   U2745 : INV_X1 port map( A => n2182, ZN => n7579);
   U2746 : AOI22_X1 port map( A1 => n6129, A2 => n2872, B1 => n6126, B2 => 
                           n7579, ZN => n6841);
   U2747 : OAI221_X1 port map( B1 => n2086, B2 => n6134, C1 => n2118, C2 => 
                           n6132, A => n6841, ZN => n6851);
   U2748 : AOI22_X1 port map( A1 => n6140, A2 => n5008, B1 => n6137, B2 => 
                           n4948, ZN => n6842);
   U2749 : OAI221_X1 port map( B1 => n6369, B2 => n6145, C1 => n3672, C2 => 
                           n6143, A => n6842, ZN => n6850);
   U2750 : AOI22_X1 port map( A1 => n2936, A2 => n6151, B1 => n7426, B2 => 
                           n6148, ZN => n6843);
   U2751 : OAI221_X1 port map( B1 => n4773, B2 => n6157, C1 => n7428, C2 => 
                           n6154, A => n6843, ZN => n6846);
   U2752 : NAND2_X1 port map( A1 => n6158, A2 => n7430, ZN => n6844);
   U2753 : NAND4_X1 port map( A1 => n1550, A2 => n1551, A3 => n1549, A4 => 
                           n6844, ZN => n6845);
   U2754 : OAI21_X1 port map( B1 => n6846, B2 => n6845, A => n6161, ZN => n6848
                           );
   U2755 : AOI22_X1 port map( A1 => n6169, A2 => n7424, B1 => n6166, B2 => 
                           n4917, ZN => n6847);
   U2756 : OAI211_X1 port map( C1 => n2246, C2 => n6172, A => n6848, B => n6847
                           , ZN => n6849);
   U2757 : NOR4_X1 port map( A1 => n6852, A2 => n6851, A3 => n6850, A4 => n6849
                           , ZN => n6853);
   U2758 : OAI21_X1 port map( B1 => n2648, B2 => n6173, A => n6853, ZN => n3009
                           );
   U2759 : OAI222_X1 port map( A1 => n4747, A2 => n6123, B1 => n2745, B2 => 
                           n6119, C1 => n2151, C2 => n6118, ZN => n6865);
   U2760 : INV_X1 port map( A => n2183, ZN => n7580);
   U2761 : AOI22_X1 port map( A1 => n6129, A2 => n2873, B1 => n6126, B2 => 
                           n7580, ZN => n6854);
   U2762 : OAI221_X1 port map( B1 => n2087, B2 => n6133, C1 => n2119, C2 => 
                           n6132, A => n6854, ZN => n6864);
   U2763 : AOI22_X1 port map( A1 => n6140, A2 => n5007, B1 => n6137, B2 => 
                           n4947, ZN => n6855);
   U2764 : OAI221_X1 port map( B1 => n6370, B2 => n6144, C1 => n3673, C2 => 
                           n6143, A => n6855, ZN => n6863);
   U2765 : AOI22_X1 port map( A1 => n2937, A2 => n6151, B1 => n7445, B2 => 
                           n6148, ZN => n6856);
   U2766 : OAI221_X1 port map( B1 => n4755, B2 => n6157, C1 => n7447, C2 => 
                           n6154, A => n6856, ZN => n6859);
   U2767 : NAND2_X1 port map( A1 => n6158, A2 => n7449, ZN => n6857);
   U2768 : NAND4_X1 port map( A1 => n1533, A2 => n1534, A3 => n1532, A4 => 
                           n6857, ZN => n6858);
   U2769 : OAI21_X1 port map( B1 => n6859, B2 => n6858, A => n6161, ZN => n6861
                           );
   U2770 : AOI22_X1 port map( A1 => n6169, A2 => n7443, B1 => n6166, B2 => 
                           n4916, ZN => n6860);
   U2771 : OAI211_X1 port map( C1 => n2247, C2 => n6172, A => n6861, B => n6860
                           , ZN => n6862);
   U2772 : NOR4_X1 port map( A1 => n6865, A2 => n6864, A3 => n6863, A4 => n6862
                           , ZN => n6866);
   U2773 : OAI21_X1 port map( B1 => n2649, B2 => n6173, A => n6866, ZN => n3010
                           );
   U2774 : OAI222_X1 port map( A1 => n4745, A2 => n6123, B1 => n2746, B2 => 
                           n6120, C1 => n2152, C2 => n6118, ZN => n6878);
   U2775 : INV_X1 port map( A => n2184, ZN => n7581);
   U2776 : AOI22_X1 port map( A1 => n6129, A2 => n2874, B1 => n6126, B2 => 
                           n7581, ZN => n6867);
   U2777 : OAI221_X1 port map( B1 => n2088, B2 => n6134, C1 => n2120, C2 => 
                           n6132, A => n6867, ZN => n6877);
   U2778 : AOI22_X1 port map( A1 => n6140, A2 => n5006, B1 => n6137, B2 => 
                           n4946, ZN => n6868);
   U2779 : OAI221_X1 port map( B1 => n6371, B2 => n6145, C1 => n3674, C2 => 
                           n6143, A => n6868, ZN => n6876);
   U2780 : AOI22_X1 port map( A1 => n2938, A2 => n6151, B1 => n7464, B2 => 
                           n6148, ZN => n6869);
   U2781 : OAI221_X1 port map( B1 => n4779, B2 => n6157, C1 => n7466, C2 => 
                           n6154, A => n6869, ZN => n6872);
   U2782 : NAND2_X1 port map( A1 => n6158, A2 => n7468, ZN => n6870);
   U2783 : NAND4_X1 port map( A1 => n1516, A2 => n1517, A3 => n1515, A4 => 
                           n6870, ZN => n6871);
   U2784 : OAI21_X1 port map( B1 => n6872, B2 => n6871, A => n6161, ZN => n6874
                           );
   U2785 : AOI22_X1 port map( A1 => n6169, A2 => n7462, B1 => n6166, B2 => 
                           n4915, ZN => n6873);
   U2786 : OAI211_X1 port map( C1 => n2248, C2 => n6172, A => n6874, B => n6873
                           , ZN => n6875);
   U2787 : NOR4_X1 port map( A1 => n6878, A2 => n6877, A3 => n6876, A4 => n6875
                           , ZN => n6879);
   U2788 : OAI21_X1 port map( B1 => n2650, B2 => n6173, A => n6879, ZN => n3011
                           );
   U2789 : OAI222_X1 port map( A1 => n4743, A2 => n6123, B1 => n2747, B2 => 
                           n6119, C1 => n2153, C2 => n6118, ZN => n6891);
   U2790 : INV_X1 port map( A => n2185, ZN => n7582);
   U2791 : AOI22_X1 port map( A1 => n6129, A2 => n2875, B1 => n6126, B2 => 
                           n7582, ZN => n6880);
   U2792 : OAI221_X1 port map( B1 => n2089, B2 => n6133, C1 => n2121, C2 => 
                           n6132, A => n6880, ZN => n6890);
   U2793 : AOI22_X1 port map( A1 => n6140, A2 => n5005, B1 => n6137, B2 => 
                           n4945, ZN => n6881);
   U2794 : OAI221_X1 port map( B1 => n6372, B2 => n6144, C1 => n3675, C2 => 
                           n6143, A => n6881, ZN => n6889);
   U2795 : AOI22_X1 port map( A1 => n2939, A2 => n6151, B1 => n7483, B2 => 
                           n6148, ZN => n6882);
   U2796 : OAI221_X1 port map( B1 => n4777, B2 => n6157, C1 => n7485, C2 => 
                           n6154, A => n6882, ZN => n6885);
   U2797 : NAND2_X1 port map( A1 => n6158, A2 => n7487, ZN => n6883);
   U2798 : NAND4_X1 port map( A1 => n1499, A2 => n1500, A3 => n1498, A4 => 
                           n6883, ZN => n6884);
   U2799 : OAI21_X1 port map( B1 => n6885, B2 => n6884, A => n6161, ZN => n6887
                           );
   U2800 : AOI22_X1 port map( A1 => n6169, A2 => n7481, B1 => n6166, B2 => 
                           n4914, ZN => n6886);
   U2801 : OAI211_X1 port map( C1 => n2249, C2 => n6172, A => n6887, B => n6886
                           , ZN => n6888);
   U2802 : NOR4_X1 port map( A1 => n6891, A2 => n6890, A3 => n6889, A4 => n6888
                           , ZN => n6892);
   U2803 : OAI21_X1 port map( B1 => n2651, B2 => n6173, A => n6892, ZN => n3012
                           );
   U2804 : OAI222_X1 port map( A1 => n4749, A2 => n6123, B1 => n2748, B2 => 
                           n6120, C1 => n2154, C2 => n6118, ZN => n6904);
   U2805 : INV_X1 port map( A => n2186, ZN => n7583);
   U2806 : AOI22_X1 port map( A1 => n6129, A2 => n2876, B1 => n6126, B2 => 
                           n7583, ZN => n6893);
   U2807 : OAI221_X1 port map( B1 => n2090, B2 => n6134, C1 => n2122, C2 => 
                           n6132, A => n6893, ZN => n6903);
   U2808 : AOI22_X1 port map( A1 => n6140, A2 => n5004, B1 => n6137, B2 => 
                           n4944, ZN => n6894);
   U2809 : OAI221_X1 port map( B1 => n6373, B2 => n6145, C1 => n3676, C2 => 
                           n6143, A => n6894, ZN => n6902);
   U2810 : AOI22_X1 port map( A1 => n2940, A2 => n6151, B1 => n7502, B2 => 
                           n6148, ZN => n6895);
   U2811 : OAI221_X1 port map( B1 => n4781, B2 => n6157, C1 => n7504, C2 => 
                           n6154, A => n6895, ZN => n6898);
   U2812 : NAND2_X1 port map( A1 => n6158, A2 => n7506, ZN => n6896);
   U2813 : NAND4_X1 port map( A1 => n1482, A2 => n1483, A3 => n1481, A4 => 
                           n6896, ZN => n6897);
   U2814 : OAI21_X1 port map( B1 => n6898, B2 => n6897, A => n6161, ZN => n6900
                           );
   U2815 : AOI22_X1 port map( A1 => n6169, A2 => n7500, B1 => n6166, B2 => 
                           n4913, ZN => n6899);
   U2816 : OAI211_X1 port map( C1 => n2250, C2 => n6172, A => n6900, B => n6899
                           , ZN => n6901);
   U2817 : NOR4_X1 port map( A1 => n6904, A2 => n6903, A3 => n6902, A4 => n6901
                           , ZN => n6905);
   U2818 : OAI21_X1 port map( B1 => n2652, B2 => n6173, A => n6905, ZN => n3013
                           );
   U2819 : OAI222_X1 port map( A1 => n4751, A2 => n6123, B1 => n2749, B2 => 
                           n6119, C1 => n2155, C2 => n6118, ZN => n6926);
   U2820 : INV_X1 port map( A => n2187, ZN => n7584);
   U2821 : AOI22_X1 port map( A1 => n6129, A2 => n2877, B1 => n6126, B2 => 
                           n7584, ZN => n6909);
   U2822 : OAI221_X1 port map( B1 => n2091, B2 => n6133, C1 => n2123, C2 => 
                           n6132, A => n6909, ZN => n6925);
   U2823 : AOI22_X1 port map( A1 => n6140, A2 => n5003, B1 => n6137, B2 => 
                           n4943, ZN => n6912);
   U2824 : OAI221_X1 port map( B1 => n6374, B2 => n6144, C1 => n3677, C2 => 
                           n6143, A => n6912, ZN => n6924);
   U2825 : AOI22_X1 port map( A1 => n2941, A2 => n6151, B1 => n7532, B2 => 
                           n6148, ZN => n6914);
   U2826 : OAI221_X1 port map( B1 => n4815, B2 => n6157, C1 => n7534, C2 => 
                           n6154, A => n6914, ZN => n6918);
   U2827 : NAND2_X1 port map( A1 => n6158, A2 => n7531, ZN => n6915);
   U2828 : NAND4_X1 port map( A1 => n1438, A2 => n1439, A3 => n1437, A4 => 
                           n6915, ZN => n6917);
   U2829 : OAI21_X1 port map( B1 => n6918, B2 => n6917, A => n6162, ZN => n6921
                           );
   U2830 : AOI22_X1 port map( A1 => n6169, A2 => n7526, B1 => n6166, B2 => 
                           n7540, ZN => n6920);
   U2831 : OAI211_X1 port map( C1 => n2251, C2 => n6172, A => n6921, B => n6920
                           , ZN => n6923);
   U2832 : NOR4_X1 port map( A1 => n6926, A2 => n6925, A3 => n6924, A4 => n6923
                           , ZN => n6927);
   U2833 : OAI21_X1 port map( B1 => n2653, B2 => n6174, A => n6927, ZN => n3014
                           );
   U2834 : NAND2_X1 port map( A1 => RD2, A2 => n4657, ZN => n6929);
   U2835 : INV_X1 port map( A => n6929, ZN => n7552);
   U2836 : NAND2_X1 port map( A1 => n1412, A2 => n4617, ZN => n7522);
   U2837 : NAND2_X1 port map( A1 => n4615, A2 => n1413, ZN => n7520);
   U2838 : NAND2_X1 port map( A1 => n4615, A2 => n4608, ZN => n7519);
   U2839 : OAI222_X1 port map( A1 => n939, A2 => n6190, B1 => n2124, B2 => 
                           n6187, C1 => n938, C2 => n6186, ZN => n6948);
   U2840 : NAND3_X1 port map( A1 => n1406, A2 => n1412, A3 => n6237, ZN => 
                           n7525);
   U2841 : NAND2_X1 port map( A1 => n1412, A2 => n4615, ZN => n7524);
   U2842 : AOI22_X1 port map( A1 => n6196, A2 => n5068, B1 => n6193, B2 => 
                           n7553, ZN => n6932);
   U2843 : OAI221_X1 port map( B1 => n6202, B2 => n4695, C1 => n2718, C2 => 
                           n6199, A => n6932, ZN => n6947);
   U2844 : NAND2_X1 port map( A1 => n1413, A2 => n4617, ZN => n7529);
   U2845 : NAND2_X1 port map( A1 => n1394, A2 => n4615, ZN => n7528);
   U2846 : AOI22_X1 port map( A1 => n6208, A2 => n5100, B1 => n6205, B2 => 
                           n4971, ZN => n6933);
   U2847 : OAI221_X1 port map( B1 => n2188, B2 => n6214, C1 => n2060, C2 => 
                           n6211, A => n6933, ZN => n6946);
   U2848 : NAND4_X1 port map( A1 => n1399, A2 => n1397, A3 => n6238, A4 => 
                           n1398, ZN => n7544);
   U2849 : AOI22_X1 port map( A1 => n2910, A2 => n6223, B1 => n6934, B2 => 
                           n6220, ZN => n6935);
   U2850 : OAI221_X1 port map( B1 => n6229, B2 => n4813, C1 => n6228, C2 => 
                           n6936, A => n6935, ZN => n6941);
   U2851 : NAND2_X1 port map( A1 => n6217, A2 => n6938, ZN => n6939);
   U2852 : NAND4_X1 port map( A1 => n825, A2 => n826, A3 => n824, A4 => n6939, 
                           ZN => n6940);
   U2853 : OAI21_X1 port map( B1 => n6941, B2 => n6940, A => n6236, ZN => n6944
                           );
   U2854 : NAND3_X1 port map( A1 => n1413, A2 => n1393, A3 => n6236, ZN => 
                           n7545);
   U2855 : INV_X1 port map( A => n7545, ZN => n7511);
   U2856 : AOI22_X1 port map( A1 => n4896, A2 => n6942, B1 => n6181, B2 => 
                           n4911, ZN => n6943);
   U2857 : OAI211_X1 port map( C1 => n7544, C2 => n6340, A => n6944, B => n6943
                           , ZN => n6945);
   U2858 : NOR4_X1 port map( A1 => n6948, A2 => n6947, A3 => n6946, A4 => n6945
                           , ZN => n6949);
   U2859 : OAI21_X1 port map( B1 => n2685, B2 => n6238, A => n6949, ZN => n3046
                           );
   U2860 : OAI222_X1 port map( A1 => n956, A2 => n6190, B1 => n2125, B2 => 
                           n6187, C1 => n955, C2 => n6186, ZN => n6966);
   U2861 : AOI22_X1 port map( A1 => n6196, A2 => n5067, B1 => n6193, B2 => 
                           n7554, ZN => n6950);
   U2862 : OAI221_X1 port map( B1 => n6202, B2 => n4694, C1 => n2719, C2 => 
                           n6199, A => n6950, ZN => n6965);
   U2863 : AOI22_X1 port map( A1 => n6208, A2 => n5099, B1 => n6205, B2 => 
                           n6951, ZN => n6952);
   U2864 : OAI221_X1 port map( B1 => n2189, B2 => n6214, C1 => n2061, C2 => 
                           n6211, A => n6952, ZN => n6964);
   U2865 : AOI22_X1 port map( A1 => n2911, A2 => n6223, B1 => n6953, B2 => 
                           n6220, ZN => n6954);
   U2866 : OAI221_X1 port map( B1 => n6229, B2 => n4811, C1 => n6228, C2 => 
                           n6955, A => n6954, ZN => n6960);
   U2867 : NAND2_X1 port map( A1 => n6217, A2 => n6957, ZN => n6958);
   U2868 : NAND4_X1 port map( A1 => n872, A2 => n873, A3 => n871, A4 => n6958, 
                           ZN => n6959);
   U2869 : OAI21_X1 port map( B1 => n6960, B2 => n6959, A => n6236, ZN => n6962
                           );
   U2870 : INV_X1 port map( A => n7544, ZN => n7510);
   U2871 : AOI22_X1 port map( A1 => n6181, A2 => n5002, B1 => DATAIN(1), B2 => 
                           n6176, ZN => n6961);
   U2872 : OAI211_X1 port map( C1 => n2253, C2 => n6182, A => n6962, B => n6961
                           , ZN => n6963);
   U2873 : NOR4_X1 port map( A1 => n6966, A2 => n6965, A3 => n6964, A4 => n6963
                           , ZN => n6967);
   U2874 : OAI21_X1 port map( B1 => n2684, B2 => n6240, A => n6967, ZN => n3045
                           );
   U2875 : OAI222_X1 port map( A1 => n972, A2 => n6190, B1 => n2126, B2 => 
                           n6187, C1 => n971, C2 => n6186, ZN => n6984);
   U2876 : AOI22_X1 port map( A1 => n6196, A2 => n5066, B1 => n6193, B2 => 
                           n7555, ZN => n6968);
   U2877 : OAI221_X1 port map( B1 => n6202, B2 => n4693, C1 => n2720, C2 => 
                           n6199, A => n6968, ZN => n6983);
   U2878 : AOI22_X1 port map( A1 => n6208, A2 => n5098, B1 => n6205, B2 => 
                           n6969, ZN => n6970);
   U2879 : OAI221_X1 port map( B1 => n2190, B2 => n6214, C1 => n2062, C2 => 
                           n6211, A => n6970, ZN => n6982);
   U2880 : AOI22_X1 port map( A1 => n2912, A2 => n6223, B1 => n6971, B2 => 
                           n6220, ZN => n6972);
   U2881 : OAI221_X1 port map( B1 => n6229, B2 => n4809, C1 => n6228, C2 => 
                           n6973, A => n6972, ZN => n6978);
   U2882 : NAND2_X1 port map( A1 => n6217, A2 => n6975, ZN => n6976);
   U2883 : NAND4_X1 port map( A1 => n889, A2 => n890, A3 => n888, A4 => n6976, 
                           ZN => n6977);
   U2884 : OAI21_X1 port map( B1 => n6978, B2 => n6977, A => n6236, ZN => n6980
                           );
   U2885 : AOI22_X1 port map( A1 => n6181, A2 => n5001, B1 => DATAIN(2), B2 => 
                           n6176, ZN => n6979);
   U2886 : OAI211_X1 port map( C1 => n2254, C2 => n6182, A => n6980, B => n6979
                           , ZN => n6981);
   U2887 : NOR4_X1 port map( A1 => n6984, A2 => n6983, A3 => n6982, A4 => n6981
                           , ZN => n6985);
   U2888 : OAI21_X1 port map( B1 => n2683, B2 => n6240, A => n6985, ZN => n3044
                           );
   U2889 : OAI222_X1 port map( A1 => n988, A2 => n6190, B1 => n2127, B2 => 
                           n6187, C1 => n987, C2 => n6186, ZN => n7002);
   U2890 : AOI22_X1 port map( A1 => n6196, A2 => n5065, B1 => n6193, B2 => 
                           n7556, ZN => n6986);
   U2891 : OAI221_X1 port map( B1 => n6202, B2 => n4692, C1 => n2721, C2 => 
                           n6199, A => n6986, ZN => n7001);
   U2892 : AOI22_X1 port map( A1 => n6208, A2 => n5097, B1 => n6205, B2 => 
                           n6987, ZN => n6988);
   U2893 : OAI221_X1 port map( B1 => n2191, B2 => n6214, C1 => n2063, C2 => 
                           n6211, A => n6988, ZN => n7000);
   U2894 : AOI22_X1 port map( A1 => n2913, A2 => n6223, B1 => n6989, B2 => 
                           n6220, ZN => n6990);
   U2895 : OAI221_X1 port map( B1 => n6229, B2 => n4807, C1 => n6228, C2 => 
                           n6991, A => n6990, ZN => n6996);
   U2896 : NAND2_X1 port map( A1 => n6217, A2 => n6993, ZN => n6994);
   U2897 : NAND4_X1 port map( A1 => n906, A2 => n907, A3 => n905, A4 => n6994, 
                           ZN => n6995);
   U2898 : OAI21_X1 port map( B1 => n6996, B2 => n6995, A => n6236, ZN => n6998
                           );
   U2899 : AOI22_X1 port map( A1 => n6181, A2 => n5000, B1 => DATAIN(3), B2 => 
                           n6176, ZN => n6997);
   U2900 : OAI211_X1 port map( C1 => n2255, C2 => n6182, A => n6998, B => n6997
                           , ZN => n6999);
   U2901 : NOR4_X1 port map( A1 => n7002, A2 => n7001, A3 => n7000, A4 => n6999
                           , ZN => n7003);
   U2902 : OAI21_X1 port map( B1 => n2682, B2 => n6240, A => n7003, ZN => n3043
                           );
   U2903 : OAI222_X1 port map( A1 => n6190, A2 => n4699, B1 => n2128, B2 => 
                           n6187, C1 => n6186, C2 => n4691, ZN => n7021);
   U2904 : AOI22_X1 port map( A1 => n6196, A2 => n5064, B1 => n6193, B2 => 
                           n7557, ZN => n7005);
   U2905 : OAI221_X1 port map( B1 => n2690, B2 => n6202, C1 => n2722, C2 => 
                           n6199, A => n7005, ZN => n7020);
   U2906 : AOI22_X1 port map( A1 => n6208, A2 => n5096, B1 => n6205, B2 => 
                           n7006, ZN => n7007);
   U2907 : OAI221_X1 port map( B1 => n2192, B2 => n6214, C1 => n2064, C2 => 
                           n6211, A => n7007, ZN => n7019);
   U2908 : AOI22_X1 port map( A1 => n2914, A2 => n6223, B1 => n7008, B2 => 
                           n6220, ZN => n7009);
   U2909 : OAI221_X1 port map( B1 => n6229, B2 => n4805, C1 => n6228, C2 => 
                           n7010, A => n7009, ZN => n7015);
   U2910 : NAND2_X1 port map( A1 => n6217, A2 => n7012, ZN => n7013);
   U2911 : NAND4_X1 port map( A1 => n923, A2 => n924, A3 => n922, A4 => n7013, 
                           ZN => n7014);
   U2912 : OAI21_X1 port map( B1 => n7015, B2 => n7014, A => n6236, ZN => n7017
                           );
   U2913 : AOI22_X1 port map( A1 => n6181, A2 => n4999, B1 => DATAIN(4), B2 => 
                           n6176, ZN => n7016);
   U2914 : OAI211_X1 port map( C1 => n2256, C2 => n6182, A => n7017, B => n7016
                           , ZN => n7018);
   U2915 : NOR4_X1 port map( A1 => n7021, A2 => n7020, A3 => n7019, A4 => n7018
                           , ZN => n7022);
   U2916 : OAI21_X1 port map( B1 => n2681, B2 => n6240, A => n7022, ZN => n3042
                           );
   U2917 : OAI222_X1 port map( A1 => n6190, A2 => n4697, B1 => n2129, B2 => 
                           n6187, C1 => n6186, C2 => n4690, ZN => n7040);
   U2918 : AOI22_X1 port map( A1 => n6196, A2 => n5063, B1 => n6193, B2 => 
                           n7558, ZN => n7024);
   U2919 : OAI221_X1 port map( B1 => n2691, B2 => n6202, C1 => n2723, C2 => 
                           n6199, A => n7024, ZN => n7039);
   U2920 : AOI22_X1 port map( A1 => n6208, A2 => n5095, B1 => n6205, B2 => 
                           n7025, ZN => n7026);
   U2921 : OAI221_X1 port map( B1 => n2193, B2 => n6214, C1 => n2065, C2 => 
                           n6211, A => n7026, ZN => n7038);
   U2922 : AOI22_X1 port map( A1 => n2915, A2 => n6223, B1 => n7027, B2 => 
                           n6220, ZN => n7028);
   U2923 : OAI221_X1 port map( B1 => n6229, B2 => n4803, C1 => n6228, C2 => 
                           n7029, A => n7028, ZN => n7034);
   U2924 : NAND2_X1 port map( A1 => n6217, A2 => n7031, ZN => n7032);
   U2925 : NAND4_X1 port map( A1 => n942, A2 => n943, A3 => n941, A4 => n7032, 
                           ZN => n7033);
   U2926 : OAI21_X1 port map( B1 => n7034, B2 => n7033, A => n6236, ZN => n7036
                           );
   U2927 : AOI22_X1 port map( A1 => n6181, A2 => n4998, B1 => DATAIN(5), B2 => 
                           n6176, ZN => n7035);
   U2928 : OAI211_X1 port map( C1 => n2257, C2 => n6182, A => n7036, B => n7035
                           , ZN => n7037);
   U2929 : NOR4_X1 port map( A1 => n7040, A2 => n7039, A3 => n7038, A4 => n7037
                           , ZN => n7041);
   U2930 : OAI21_X1 port map( B1 => n2680, B2 => n6240, A => n7041, ZN => n3041
                           );
   U2931 : OAI222_X1 port map( A1 => n6190, A2 => n4705, B1 => n2130, B2 => 
                           n6187, C1 => n6186, C2 => n4689, ZN => n7059);
   U2932 : AOI22_X1 port map( A1 => n6196, A2 => n5062, B1 => n6193, B2 => 
                           n7559, ZN => n7043);
   U2933 : OAI221_X1 port map( B1 => n2692, B2 => n6202, C1 => n2724, C2 => 
                           n6199, A => n7043, ZN => n7058);
   U2934 : AOI22_X1 port map( A1 => n6208, A2 => n5094, B1 => n6205, B2 => 
                           n7044, ZN => n7045);
   U2935 : OAI221_X1 port map( B1 => n2194, B2 => n6214, C1 => n2066, C2 => 
                           n6211, A => n7045, ZN => n7057);
   U2936 : AOI22_X1 port map( A1 => n2916, A2 => n6223, B1 => n7046, B2 => 
                           n6220, ZN => n7047);
   U2937 : OAI221_X1 port map( B1 => n6229, B2 => n4801, C1 => n6228, C2 => 
                           n7048, A => n7047, ZN => n7053);
   U2938 : NAND2_X1 port map( A1 => n6217, A2 => n7050, ZN => n7051);
   U2939 : NAND4_X1 port map( A1 => n962, A2 => n963, A3 => n961, A4 => n7051, 
                           ZN => n7052);
   U2940 : OAI21_X1 port map( B1 => n7053, B2 => n7052, A => n6236, ZN => n7055
                           );
   U2941 : AOI22_X1 port map( A1 => n6181, A2 => n4997, B1 => DATAIN(6), B2 => 
                           n6176, ZN => n7054);
   U2942 : OAI211_X1 port map( C1 => n2258, C2 => n6182, A => n7055, B => n7054
                           , ZN => n7056);
   U2943 : NOR4_X1 port map( A1 => n7059, A2 => n7058, A3 => n7057, A4 => n7056
                           , ZN => n7060);
   U2944 : OAI21_X1 port map( B1 => n2679, B2 => n6240, A => n7060, ZN => n3040
                           );
   U2945 : OAI222_X1 port map( A1 => n6190, A2 => n4703, B1 => n2131, B2 => 
                           n6187, C1 => n6186, C2 => n4688, ZN => n7078);
   U2946 : AOI22_X1 port map( A1 => n6196, A2 => n5061, B1 => n6193, B2 => 
                           n7560, ZN => n7062);
   U2947 : OAI221_X1 port map( B1 => n2693, B2 => n6202, C1 => n2725, C2 => 
                           n6199, A => n7062, ZN => n7077);
   U2948 : AOI22_X1 port map( A1 => n6208, A2 => n5093, B1 => n6205, B2 => 
                           n7063, ZN => n7064);
   U2949 : OAI221_X1 port map( B1 => n2195, B2 => n6214, C1 => n2067, C2 => 
                           n6211, A => n7064, ZN => n7076);
   U2950 : AOI22_X1 port map( A1 => n2917, A2 => n6223, B1 => n7065, B2 => 
                           n6220, ZN => n7066);
   U2951 : OAI221_X1 port map( B1 => n6229, B2 => n4799, C1 => n6228, C2 => 
                           n7067, A => n7066, ZN => n7072);
   U2952 : NAND2_X1 port map( A1 => n6217, A2 => n7069, ZN => n7070);
   U2953 : NAND4_X1 port map( A1 => n983, A2 => n984, A3 => n981, A4 => n7070, 
                           ZN => n7071);
   U2954 : OAI21_X1 port map( B1 => n7072, B2 => n7071, A => n6236, ZN => n7074
                           );
   U2955 : AOI22_X1 port map( A1 => n6180, A2 => n4996, B1 => DATAIN(7), B2 => 
                           n6176, ZN => n7073);
   U2956 : OAI211_X1 port map( C1 => n2259, C2 => n6182, A => n7074, B => n7073
                           , ZN => n7075);
   U2957 : NOR4_X1 port map( A1 => n7078, A2 => n7077, A3 => n7076, A4 => n7075
                           , ZN => n7079);
   U2958 : OAI21_X1 port map( B1 => n2678, B2 => n6240, A => n7079, ZN => n3039
                           );
   U2959 : OAI222_X1 port map( A1 => n6190, A2 => n4701, B1 => n2132, B2 => 
                           n6187, C1 => n6185, C2 => n4687, ZN => n7097);
   U2960 : AOI22_X1 port map( A1 => n6196, A2 => n5060, B1 => n6193, B2 => 
                           n7561, ZN => n7081);
   U2961 : OAI221_X1 port map( B1 => n2694, B2 => n6202, C1 => n2726, C2 => 
                           n6199, A => n7081, ZN => n7096);
   U2962 : AOI22_X1 port map( A1 => n6208, A2 => n5092, B1 => n6205, B2 => 
                           n7082, ZN => n7083);
   U2963 : OAI221_X1 port map( B1 => n2196, B2 => n6214, C1 => n2068, C2 => 
                           n6211, A => n7083, ZN => n7095);
   U2964 : AOI22_X1 port map( A1 => n2918, A2 => n6223, B1 => n7084, B2 => 
                           n6220, ZN => n7085);
   U2965 : OAI221_X1 port map( B1 => n6229, B2 => n4797, C1 => n6227, C2 => 
                           n7086, A => n7085, ZN => n7091);
   U2966 : NAND2_X1 port map( A1 => n6217, A2 => n7088, ZN => n7089);
   U2967 : NAND4_X1 port map( A1 => n1003, A2 => n1004, A3 => n1002, A4 => 
                           n7089, ZN => n7090);
   U2968 : OAI21_X1 port map( B1 => n7091, B2 => n7090, A => n6235, ZN => n7093
                           );
   U2969 : AOI22_X1 port map( A1 => n6180, A2 => n4995, B1 => DATAIN(8), B2 => 
                           n6176, ZN => n7092);
   U2970 : OAI211_X1 port map( C1 => n2260, C2 => n6182, A => n7093, B => n7092
                           , ZN => n7094);
   U2971 : NOR4_X1 port map( A1 => n7097, A2 => n7096, A3 => n7095, A4 => n7094
                           , ZN => n7098);
   U2972 : OAI21_X1 port map( B1 => n2677, B2 => n6240, A => n7098, ZN => n3038
                           );
   U2973 : OAI222_X1 port map( A1 => n6190, A2 => n4711, B1 => n2133, B2 => 
                           n6187, C1 => n6185, C2 => n4686, ZN => n7116);
   U2974 : AOI22_X1 port map( A1 => n6196, A2 => n5059, B1 => n6193, B2 => 
                           n7562, ZN => n7100);
   U2975 : OAI221_X1 port map( B1 => n2695, B2 => n6202, C1 => n2727, C2 => 
                           n6199, A => n7100, ZN => n7115);
   U2976 : AOI22_X1 port map( A1 => n6208, A2 => n5091, B1 => n6205, B2 => 
                           n7101, ZN => n7102);
   U2977 : OAI221_X1 port map( B1 => n2197, B2 => n6214, C1 => n2069, C2 => 
                           n6211, A => n7102, ZN => n7114);
   U2978 : AOI22_X1 port map( A1 => n2919, A2 => n6223, B1 => n7103, B2 => 
                           n6220, ZN => n7104);
   U2979 : OAI221_X1 port map( B1 => n6229, B2 => n4795, C1 => n6227, C2 => 
                           n7105, A => n7104, ZN => n7110);
   U2980 : NAND2_X1 port map( A1 => n6217, A2 => n7107, ZN => n7108);
   U2981 : NAND4_X1 port map( A1 => n1020, A2 => n1021, A3 => n1019, A4 => 
                           n7108, ZN => n7109);
   U2982 : OAI21_X1 port map( B1 => n7110, B2 => n7109, A => n6235, ZN => n7112
                           );
   U2983 : AOI22_X1 port map( A1 => n6180, A2 => n4994, B1 => DATAIN(9), B2 => 
                           n6176, ZN => n7111);
   U2984 : OAI211_X1 port map( C1 => n2261, C2 => n6182, A => n7112, B => n7111
                           , ZN => n7113);
   U2985 : NOR4_X1 port map( A1 => n7116, A2 => n7115, A3 => n7114, A4 => n7113
                           , ZN => n7117);
   U2986 : OAI21_X1 port map( B1 => n2676, B2 => n6240, A => n7117, ZN => n3037
                           );
   U2987 : OAI222_X1 port map( A1 => n6190, A2 => n4709, B1 => n2134, B2 => 
                           n6187, C1 => n6185, C2 => n4685, ZN => n7135);
   U2988 : AOI22_X1 port map( A1 => n6196, A2 => n5058, B1 => n6193, B2 => 
                           n7563, ZN => n7119);
   U2989 : OAI221_X1 port map( B1 => n2696, B2 => n6202, C1 => n2728, C2 => 
                           n6199, A => n7119, ZN => n7134);
   U2990 : AOI22_X1 port map( A1 => n6208, A2 => n5090, B1 => n6205, B2 => 
                           n7120, ZN => n7121);
   U2991 : OAI221_X1 port map( B1 => n2198, B2 => n6214, C1 => n2070, C2 => 
                           n6211, A => n7121, ZN => n7133);
   U2992 : AOI22_X1 port map( A1 => n2920, A2 => n6223, B1 => n7122, B2 => 
                           n6220, ZN => n7123);
   U2993 : OAI221_X1 port map( B1 => n6229, B2 => n4793, C1 => n6227, C2 => 
                           n7124, A => n7123, ZN => n7129);
   U2994 : NAND2_X1 port map( A1 => n6217, A2 => n7126, ZN => n7127);
   U2995 : NAND4_X1 port map( A1 => n1037, A2 => n1038, A3 => n1036, A4 => 
                           n7127, ZN => n7128);
   U2996 : OAI21_X1 port map( B1 => n7129, B2 => n7128, A => n6235, ZN => n7131
                           );
   U2997 : AOI22_X1 port map( A1 => n6180, A2 => n4993, B1 => DATAIN(10), B2 =>
                           n6176, ZN => n7130);
   U2998 : OAI211_X1 port map( C1 => n2262, C2 => n6182, A => n7131, B => n7130
                           , ZN => n7132);
   U2999 : NOR4_X1 port map( A1 => n7135, A2 => n7134, A3 => n7133, A4 => n7132
                           , ZN => n7136);
   U3000 : OAI21_X1 port map( B1 => n2675, B2 => n6239, A => n7136, ZN => n3036
                           );
   U3001 : OAI222_X1 port map( A1 => n6190, A2 => n4707, B1 => n2135, B2 => 
                           n6187, C1 => n6185, C2 => n4684, ZN => n7154);
   U3002 : AOI22_X1 port map( A1 => n6196, A2 => n5057, B1 => n6193, B2 => 
                           n7564, ZN => n7138);
   U3003 : OAI221_X1 port map( B1 => n2697, B2 => n6202, C1 => n2729, C2 => 
                           n6199, A => n7138, ZN => n7153);
   U3004 : AOI22_X1 port map( A1 => n6208, A2 => n5089, B1 => n6205, B2 => 
                           n7139, ZN => n7140);
   U3005 : OAI221_X1 port map( B1 => n2199, B2 => n6214, C1 => n2071, C2 => 
                           n6211, A => n7140, ZN => n7152);
   U3006 : AOI22_X1 port map( A1 => n2921, A2 => n6223, B1 => n7141, B2 => 
                           n6220, ZN => n7142);
   U3007 : OAI221_X1 port map( B1 => n6229, B2 => n4791, C1 => n6227, C2 => 
                           n7143, A => n7142, ZN => n7148);
   U3008 : NAND2_X1 port map( A1 => n6217, A2 => n7145, ZN => n7146);
   U3009 : NAND4_X1 port map( A1 => n1054, A2 => n1055, A3 => n1053, A4 => 
                           n7146, ZN => n7147);
   U3010 : OAI21_X1 port map( B1 => n7148, B2 => n7147, A => n6235, ZN => n7150
                           );
   U3011 : AOI22_X1 port map( A1 => n6180, A2 => n4992, B1 => DATAIN(11), B2 =>
                           n6176, ZN => n7149);
   U3012 : OAI211_X1 port map( C1 => n2263, C2 => n6182, A => n7150, B => n7149
                           , ZN => n7151);
   U3013 : NOR4_X1 port map( A1 => n7154, A2 => n7153, A3 => n7152, A4 => n7151
                           , ZN => n7155);
   U3014 : OAI21_X1 port map( B1 => n2674, B2 => n6239, A => n7155, ZN => n3035
                           );
   U3015 : OAI222_X1 port map( A1 => n6191, A2 => n4717, B1 => n2136, B2 => 
                           n6188, C1 => n6185, C2 => n4683, ZN => n7173);
   U3016 : AOI22_X1 port map( A1 => n6197, A2 => n5056, B1 => n6194, B2 => 
                           n7565, ZN => n7157);
   U3017 : OAI221_X1 port map( B1 => n2698, B2 => n6203, C1 => n2730, C2 => 
                           n6200, A => n7157, ZN => n7172);
   U3018 : AOI22_X1 port map( A1 => n6209, A2 => n5088, B1 => n6206, B2 => 
                           n7158, ZN => n7159);
   U3019 : OAI221_X1 port map( B1 => n2200, B2 => n6215, C1 => n2072, C2 => 
                           n6212, A => n7159, ZN => n7171);
   U3020 : AOI22_X1 port map( A1 => n2922, A2 => n6224, B1 => n7160, B2 => 
                           n6221, ZN => n7161);
   U3021 : OAI221_X1 port map( B1 => n6230, B2 => n4789, C1 => n6227, C2 => 
                           n7162, A => n7161, ZN => n7167);
   U3022 : NAND2_X1 port map( A1 => n6218, A2 => n7164, ZN => n7165);
   U3023 : NAND4_X1 port map( A1 => n1071, A2 => n1072, A3 => n1070, A4 => 
                           n7165, ZN => n7166);
   U3024 : OAI21_X1 port map( B1 => n7167, B2 => n7166, A => n6235, ZN => n7169
                           );
   U3025 : AOI22_X1 port map( A1 => n6180, A2 => n4991, B1 => DATAIN(12), B2 =>
                           n6176, ZN => n7168);
   U3026 : OAI211_X1 port map( C1 => n2264, C2 => n6182, A => n7169, B => n7168
                           , ZN => n7170);
   U3027 : NOR4_X1 port map( A1 => n7173, A2 => n7172, A3 => n7171, A4 => n7170
                           , ZN => n7174);
   U3028 : OAI21_X1 port map( B1 => n2673, B2 => n6239, A => n7174, ZN => n3034
                           );
   U3029 : OAI222_X1 port map( A1 => n6191, A2 => n4715, B1 => n2137, B2 => 
                           n6188, C1 => n6185, C2 => n4682, ZN => n7192);
   U3030 : AOI22_X1 port map( A1 => n6197, A2 => n5055, B1 => n6194, B2 => 
                           n7566, ZN => n7176);
   U3031 : OAI221_X1 port map( B1 => n2699, B2 => n6203, C1 => n2731, C2 => 
                           n6200, A => n7176, ZN => n7191);
   U3032 : AOI22_X1 port map( A1 => n6209, A2 => n5087, B1 => n6206, B2 => 
                           n7177, ZN => n7178);
   U3033 : OAI221_X1 port map( B1 => n2201, B2 => n6215, C1 => n2073, C2 => 
                           n6212, A => n7178, ZN => n7190);
   U3034 : AOI22_X1 port map( A1 => n2923, A2 => n6224, B1 => n7179, B2 => 
                           n6221, ZN => n7180);
   U3035 : OAI221_X1 port map( B1 => n6230, B2 => n4787, C1 => n6227, C2 => 
                           n7181, A => n7180, ZN => n7186);
   U3036 : NAND2_X1 port map( A1 => n6218, A2 => n7183, ZN => n7184);
   U3037 : NAND4_X1 port map( A1 => n1088, A2 => n1089, A3 => n1087, A4 => 
                           n7184, ZN => n7185);
   U3038 : OAI21_X1 port map( B1 => n7186, B2 => n7185, A => n6235, ZN => n7188
                           );
   U3039 : AOI22_X1 port map( A1 => n6180, A2 => n4990, B1 => DATAIN(13), B2 =>
                           n6177, ZN => n7187);
   U3040 : OAI211_X1 port map( C1 => n2265, C2 => n6183, A => n7188, B => n7187
                           , ZN => n7189);
   U3041 : NOR4_X1 port map( A1 => n7192, A2 => n7191, A3 => n7190, A4 => n7189
                           , ZN => n7193);
   U3042 : OAI21_X1 port map( B1 => n2672, B2 => n6239, A => n7193, ZN => n3033
                           );
   U3043 : OAI222_X1 port map( A1 => n6191, A2 => n4713, B1 => n2138, B2 => 
                           n6188, C1 => n6185, C2 => n4681, ZN => n7211);
   U3044 : AOI22_X1 port map( A1 => n6197, A2 => n5054, B1 => n6194, B2 => 
                           n7567, ZN => n7195);
   U3045 : OAI221_X1 port map( B1 => n2700, B2 => n6203, C1 => n2732, C2 => 
                           n6200, A => n7195, ZN => n7210);
   U3046 : AOI22_X1 port map( A1 => n6209, A2 => n5086, B1 => n6206, B2 => 
                           n7196, ZN => n7197);
   U3047 : OAI221_X1 port map( B1 => n2202, B2 => n6215, C1 => n2074, C2 => 
                           n6212, A => n7197, ZN => n7209);
   U3048 : AOI22_X1 port map( A1 => n2924, A2 => n6224, B1 => n7198, B2 => 
                           n6221, ZN => n7199);
   U3049 : OAI221_X1 port map( B1 => n6230, B2 => n4785, C1 => n6227, C2 => 
                           n7200, A => n7199, ZN => n7205);
   U3050 : NAND2_X1 port map( A1 => n6218, A2 => n7202, ZN => n7203);
   U3051 : NAND4_X1 port map( A1 => n1105, A2 => n1106, A3 => n1104, A4 => 
                           n7203, ZN => n7204);
   U3052 : OAI21_X1 port map( B1 => n7205, B2 => n7204, A => n6235, ZN => n7207
                           );
   U3053 : AOI22_X1 port map( A1 => n6180, A2 => n4989, B1 => DATAIN(14), B2 =>
                           n6177, ZN => n7206);
   U3054 : OAI211_X1 port map( C1 => n2266, C2 => n6183, A => n7207, B => n7206
                           , ZN => n7208);
   U3055 : NOR4_X1 port map( A1 => n7211, A2 => n7210, A3 => n7209, A4 => n7208
                           , ZN => n7212);
   U3056 : OAI21_X1 port map( B1 => n2671, B2 => n6239, A => n7212, ZN => n3032
                           );
   U3057 : OAI222_X1 port map( A1 => n6191, A2 => n4723, B1 => n2139, B2 => 
                           n6188, C1 => n6185, C2 => n4680, ZN => n7230);
   U3058 : AOI22_X1 port map( A1 => n6197, A2 => n5053, B1 => n6194, B2 => 
                           n7568, ZN => n7214);
   U3059 : OAI221_X1 port map( B1 => n2701, B2 => n6203, C1 => n2733, C2 => 
                           n6200, A => n7214, ZN => n7229);
   U3060 : AOI22_X1 port map( A1 => n6209, A2 => n5085, B1 => n6206, B2 => 
                           n7215, ZN => n7216);
   U3061 : OAI221_X1 port map( B1 => n2203, B2 => n6215, C1 => n2075, C2 => 
                           n6212, A => n7216, ZN => n7228);
   U3062 : AOI22_X1 port map( A1 => n2925, A2 => n6224, B1 => n7217, B2 => 
                           n6221, ZN => n7218);
   U3063 : OAI221_X1 port map( B1 => n6230, B2 => n4783, C1 => n6227, C2 => 
                           n7219, A => n7218, ZN => n7224);
   U3064 : NAND2_X1 port map( A1 => n6218, A2 => n7221, ZN => n7222);
   U3065 : NAND4_X1 port map( A1 => n1122, A2 => n1123, A3 => n1121, A4 => 
                           n7222, ZN => n7223);
   U3066 : OAI21_X1 port map( B1 => n7224, B2 => n7223, A => n6235, ZN => n7226
                           );
   U3067 : AOI22_X1 port map( A1 => n6180, A2 => n4988, B1 => DATAIN(15), B2 =>
                           n6177, ZN => n7225);
   U3068 : OAI211_X1 port map( C1 => n2267, C2 => n6183, A => n7226, B => n7225
                           , ZN => n7227);
   U3069 : NOR4_X1 port map( A1 => n7230, A2 => n7229, A3 => n7228, A4 => n7227
                           , ZN => n7231);
   U3070 : OAI21_X1 port map( B1 => n2670, B2 => n6239, A => n7231, ZN => n3031
                           );
   U3071 : OAI222_X1 port map( A1 => n6191, A2 => n4721, B1 => n2140, B2 => 
                           n6188, C1 => n6185, C2 => n4679, ZN => n7249);
   U3072 : AOI22_X1 port map( A1 => n6197, A2 => n5052, B1 => n6194, B2 => 
                           n7569, ZN => n7233);
   U3073 : OAI221_X1 port map( B1 => n2702, B2 => n6203, C1 => n2734, C2 => 
                           n6200, A => n7233, ZN => n7248);
   U3074 : AOI22_X1 port map( A1 => n6209, A2 => n5084, B1 => n6206, B2 => 
                           n7234, ZN => n7235);
   U3075 : OAI221_X1 port map( B1 => n2204, B2 => n6215, C1 => n2076, C2 => 
                           n6212, A => n7235, ZN => n7247);
   U3076 : AOI22_X1 port map( A1 => n2926, A2 => n6224, B1 => n7236, B2 => 
                           n6221, ZN => n7237);
   U3077 : OAI221_X1 port map( B1 => n6230, B2 => n4753, C1 => n6227, C2 => 
                           n7238, A => n7237, ZN => n7243);
   U3078 : NAND2_X1 port map( A1 => n6218, A2 => n7240, ZN => n7241);
   U3079 : NAND4_X1 port map( A1 => n1139, A2 => n1140, A3 => n1138, A4 => 
                           n7241, ZN => n7242);
   U3080 : OAI21_X1 port map( B1 => n7243, B2 => n7242, A => n6235, ZN => n7245
                           );
   U3081 : AOI22_X1 port map( A1 => n6180, A2 => n4987, B1 => DATAIN(16), B2 =>
                           n6177, ZN => n7244);
   U3082 : OAI211_X1 port map( C1 => n2268, C2 => n6183, A => n7245, B => n7244
                           , ZN => n7246);
   U3083 : NOR4_X1 port map( A1 => n7249, A2 => n7248, A3 => n7247, A4 => n7246
                           , ZN => n7250);
   U3084 : OAI21_X1 port map( B1 => n2669, B2 => n6239, A => n7250, ZN => n3030
                           );
   U3085 : OAI222_X1 port map( A1 => n6191, A2 => n4719, B1 => n2141, B2 => 
                           n6188, C1 => n6185, C2 => n4678, ZN => n7268);
   U3086 : AOI22_X1 port map( A1 => n6197, A2 => n5051, B1 => n6194, B2 => 
                           n7570, ZN => n7252);
   U3087 : OAI221_X1 port map( B1 => n2703, B2 => n6203, C1 => n2735, C2 => 
                           n6200, A => n7252, ZN => n7267);
   U3088 : AOI22_X1 port map( A1 => n6209, A2 => n5083, B1 => n6206, B2 => 
                           n7253, ZN => n7254);
   U3089 : OAI221_X1 port map( B1 => n2205, B2 => n6215, C1 => n2077, C2 => 
                           n6212, A => n7254, ZN => n7266);
   U3090 : AOI22_X1 port map( A1 => n2927, A2 => n6224, B1 => n7255, B2 => 
                           n6221, ZN => n7256);
   U3091 : OAI221_X1 port map( B1 => n6230, B2 => n4763, C1 => n6227, C2 => 
                           n7257, A => n7256, ZN => n7262);
   U3092 : NAND2_X1 port map( A1 => n6218, A2 => n7259, ZN => n7260);
   U3093 : NAND4_X1 port map( A1 => n1156, A2 => n1157, A3 => n1155, A4 => 
                           n7260, ZN => n7261);
   U3094 : OAI21_X1 port map( B1 => n7262, B2 => n7261, A => n6235, ZN => n7264
                           );
   U3095 : AOI22_X1 port map( A1 => n6180, A2 => n4986, B1 => DATAIN(17), B2 =>
                           n6177, ZN => n7263);
   U3096 : OAI211_X1 port map( C1 => n2269, C2 => n6183, A => n7264, B => n7263
                           , ZN => n7265);
   U3097 : NOR4_X1 port map( A1 => n7268, A2 => n7267, A3 => n7266, A4 => n7265
                           , ZN => n7269);
   U3098 : OAI21_X1 port map( B1 => n2668, B2 => n6239, A => n7269, ZN => n3029
                           );
   U3099 : OAI222_X1 port map( A1 => n6191, A2 => n4729, B1 => n2142, B2 => 
                           n6188, C1 => n6185, C2 => n4677, ZN => n7287);
   U3100 : AOI22_X1 port map( A1 => n6197, A2 => n5050, B1 => n6194, B2 => 
                           n7571, ZN => n7271);
   U3101 : OAI221_X1 port map( B1 => n2704, B2 => n6203, C1 => n2736, C2 => 
                           n6200, A => n7271, ZN => n7286);
   U3102 : AOI22_X1 port map( A1 => n6209, A2 => n5082, B1 => n6206, B2 => 
                           n7272, ZN => n7273);
   U3103 : OAI221_X1 port map( B1 => n2206, B2 => n6215, C1 => n2078, C2 => 
                           n6212, A => n7273, ZN => n7285);
   U3104 : AOI22_X1 port map( A1 => n2928, A2 => n6224, B1 => n7274, B2 => 
                           n6221, ZN => n7275);
   U3105 : OAI221_X1 port map( B1 => n6230, B2 => n4757, C1 => n6227, C2 => 
                           n7276, A => n7275, ZN => n7281);
   U3106 : NAND2_X1 port map( A1 => n6218, A2 => n7278, ZN => n7279);
   U3107 : NAND4_X1 port map( A1 => n1173, A2 => n1174, A3 => n1172, A4 => 
                           n7279, ZN => n7280);
   U3108 : OAI21_X1 port map( B1 => n7281, B2 => n7280, A => n6235, ZN => n7283
                           );
   U3109 : AOI22_X1 port map( A1 => n6180, A2 => n4985, B1 => DATAIN(18), B2 =>
                           n6177, ZN => n7282);
   U3110 : OAI211_X1 port map( C1 => n2270, C2 => n6183, A => n7283, B => n7282
                           , ZN => n7284);
   U3111 : NOR4_X1 port map( A1 => n7287, A2 => n7286, A3 => n7285, A4 => n7284
                           , ZN => n7288);
   U3112 : OAI21_X1 port map( B1 => n2667, B2 => n6239, A => n7288, ZN => n3028
                           );
   U3113 : OAI222_X1 port map( A1 => n6191, A2 => n4727, B1 => n2143, B2 => 
                           n6188, C1 => n6185, C2 => n4676, ZN => n7306);
   U3114 : AOI22_X1 port map( A1 => n6197, A2 => n5049, B1 => n6194, B2 => 
                           n7572, ZN => n7290);
   U3115 : OAI221_X1 port map( B1 => n2705, B2 => n6203, C1 => n2737, C2 => 
                           n6200, A => n7290, ZN => n7305);
   U3116 : AOI22_X1 port map( A1 => n6209, A2 => n5081, B1 => n6206, B2 => 
                           n7291, ZN => n7292);
   U3117 : OAI221_X1 port map( B1 => n2207, B2 => n6215, C1 => n2079, C2 => 
                           n6212, A => n7292, ZN => n7304);
   U3118 : AOI22_X1 port map( A1 => n2929, A2 => n6224, B1 => n7293, B2 => 
                           n6221, ZN => n7294);
   U3119 : OAI221_X1 port map( B1 => n6230, B2 => n4759, C1 => n6227, C2 => 
                           n7295, A => n7294, ZN => n7300);
   U3120 : NAND2_X1 port map( A1 => n6218, A2 => n7297, ZN => n7298);
   U3121 : NAND4_X1 port map( A1 => n1190, A2 => n1191, A3 => n1189, A4 => 
                           n7298, ZN => n7299);
   U3122 : OAI21_X1 port map( B1 => n7300, B2 => n7299, A => n6234, ZN => n7302
                           );
   U3123 : AOI22_X1 port map( A1 => n6179, A2 => n4984, B1 => DATAIN(19), B2 =>
                           n6177, ZN => n7301);
   U3124 : OAI211_X1 port map( C1 => n2271, C2 => n6183, A => n7302, B => n7301
                           , ZN => n7303);
   U3125 : NOR4_X1 port map( A1 => n7306, A2 => n7305, A3 => n7304, A4 => n7303
                           , ZN => n7307);
   U3126 : OAI21_X1 port map( B1 => n2666, B2 => n6239, A => n7307, ZN => n3027
                           );
   U3127 : OAI222_X1 port map( A1 => n6191, A2 => n4725, B1 => n2144, B2 => 
                           n6188, C1 => n6184, C2 => n4675, ZN => n7325);
   U3128 : AOI22_X1 port map( A1 => n6197, A2 => n5048, B1 => n6194, B2 => 
                           n7573, ZN => n7309);
   U3129 : OAI221_X1 port map( B1 => n2706, B2 => n6203, C1 => n2738, C2 => 
                           n6200, A => n7309, ZN => n7324);
   U3130 : AOI22_X1 port map( A1 => n6209, A2 => n5080, B1 => n6206, B2 => 
                           n7310, ZN => n7311);
   U3131 : OAI221_X1 port map( B1 => n2208, B2 => n6215, C1 => n2080, C2 => 
                           n6212, A => n7311, ZN => n7323);
   U3132 : AOI22_X1 port map( A1 => n2930, A2 => n6224, B1 => n7312, B2 => 
                           n6221, ZN => n7313);
   U3133 : OAI221_X1 port map( B1 => n6230, B2 => n4769, C1 => n6226, C2 => 
                           n7314, A => n7313, ZN => n7319);
   U3134 : NAND2_X1 port map( A1 => n6218, A2 => n7316, ZN => n7317);
   U3135 : NAND4_X1 port map( A1 => n1207, A2 => n1208, A3 => n1206, A4 => 
                           n7317, ZN => n7318);
   U3136 : OAI21_X1 port map( B1 => n7319, B2 => n7318, A => n6235, ZN => n7321
                           );
   U3137 : AOI22_X1 port map( A1 => n6179, A2 => n4983, B1 => DATAIN(20), B2 =>
                           n6177, ZN => n7320);
   U3138 : OAI211_X1 port map( C1 => n2272, C2 => n6183, A => n7321, B => n7320
                           , ZN => n7322);
   U3139 : NOR4_X1 port map( A1 => n7325, A2 => n7324, A3 => n7323, A4 => n7322
                           , ZN => n7326);
   U3140 : OAI21_X1 port map( B1 => n2665, B2 => n6239, A => n7326, ZN => n3026
                           );
   U3141 : OAI222_X1 port map( A1 => n6191, A2 => n4735, B1 => n2145, B2 => 
                           n6188, C1 => n6184, C2 => n4674, ZN => n7344);
   U3142 : AOI22_X1 port map( A1 => n6197, A2 => n5047, B1 => n6194, B2 => 
                           n7574, ZN => n7328);
   U3143 : OAI221_X1 port map( B1 => n2707, B2 => n6203, C1 => n2739, C2 => 
                           n6200, A => n7328, ZN => n7343);
   U3144 : AOI22_X1 port map( A1 => n6209, A2 => n5079, B1 => n6206, B2 => 
                           n7329, ZN => n7330);
   U3145 : OAI221_X1 port map( B1 => n2209, B2 => n6215, C1 => n2081, C2 => 
                           n6212, A => n7330, ZN => n7342);
   U3146 : AOI22_X1 port map( A1 => n2931, A2 => n6224, B1 => n7331, B2 => 
                           n6221, ZN => n7332);
   U3147 : OAI221_X1 port map( B1 => n6230, B2 => n4761, C1 => n6226, C2 => 
                           n7333, A => n7332, ZN => n7338);
   U3148 : NAND2_X1 port map( A1 => n6218, A2 => n7335, ZN => n7336);
   U3149 : NAND4_X1 port map( A1 => n1224, A2 => n1225, A3 => n1223, A4 => 
                           n7336, ZN => n7337);
   U3150 : OAI21_X1 port map( B1 => n7338, B2 => n7337, A => n6234, ZN => n7340
                           );
   U3151 : AOI22_X1 port map( A1 => n6179, A2 => n4982, B1 => DATAIN(21), B2 =>
                           n6177, ZN => n7339);
   U3152 : OAI211_X1 port map( C1 => n2273, C2 => n6183, A => n7340, B => n7339
                           , ZN => n7341);
   U3153 : NOR4_X1 port map( A1 => n7344, A2 => n7343, A3 => n7342, A4 => n7341
                           , ZN => n7345);
   U3154 : OAI21_X1 port map( B1 => n2664, B2 => n6238, A => n7345, ZN => n3025
                           );
   U3155 : OAI222_X1 port map( A1 => n6191, A2 => n4733, B1 => n2146, B2 => 
                           n6188, C1 => n6184, C2 => n4673, ZN => n7363);
   U3156 : AOI22_X1 port map( A1 => n6197, A2 => n5046, B1 => n6194, B2 => 
                           n7575, ZN => n7347);
   U3157 : OAI221_X1 port map( B1 => n2708, B2 => n6203, C1 => n2740, C2 => 
                           n6200, A => n7347, ZN => n7362);
   U3158 : AOI22_X1 port map( A1 => n6209, A2 => n5078, B1 => n6206, B2 => 
                           n7348, ZN => n7349);
   U3159 : OAI221_X1 port map( B1 => n2210, B2 => n6215, C1 => n2082, C2 => 
                           n6212, A => n7349, ZN => n7361);
   U3160 : AOI22_X1 port map( A1 => n2932, A2 => n6224, B1 => n7350, B2 => 
                           n6221, ZN => n7351);
   U3161 : OAI221_X1 port map( B1 => n6230, B2 => n4765, C1 => n6226, C2 => 
                           n7352, A => n7351, ZN => n7357);
   U3162 : NAND2_X1 port map( A1 => n6218, A2 => n7354, ZN => n7355);
   U3163 : NAND4_X1 port map( A1 => n1241, A2 => n1242, A3 => n1240, A4 => 
                           n7355, ZN => n7356);
   U3164 : OAI21_X1 port map( B1 => n7357, B2 => n7356, A => n6234, ZN => n7359
                           );
   U3165 : AOI22_X1 port map( A1 => n6179, A2 => n4981, B1 => DATAIN(22), B2 =>
                           n6177, ZN => n7358);
   U3166 : OAI211_X1 port map( C1 => n2274, C2 => n6183, A => n7359, B => n7358
                           , ZN => n7360);
   U3167 : NOR4_X1 port map( A1 => n7363, A2 => n7362, A3 => n7361, A4 => n7360
                           , ZN => n7364);
   U3168 : OAI21_X1 port map( B1 => n2663, B2 => n6238, A => n7364, ZN => n3024
                           );
   U3169 : OAI222_X1 port map( A1 => n6191, A2 => n4731, B1 => n2147, B2 => 
                           n6188, C1 => n6184, C2 => n4672, ZN => n7382);
   U3170 : AOI22_X1 port map( A1 => n6197, A2 => n5045, B1 => n6194, B2 => 
                           n7576, ZN => n7366);
   U3171 : OAI221_X1 port map( B1 => n2709, B2 => n6203, C1 => n2741, C2 => 
                           n6200, A => n7366, ZN => n7381);
   U3172 : AOI22_X1 port map( A1 => n6209, A2 => n5077, B1 => n6206, B2 => 
                           n7367, ZN => n7368);
   U3173 : OAI221_X1 port map( B1 => n2211, B2 => n6215, C1 => n2083, C2 => 
                           n6212, A => n7368, ZN => n7380);
   U3174 : AOI22_X1 port map( A1 => n2933, A2 => n6224, B1 => n7369, B2 => 
                           n6221, ZN => n7370);
   U3175 : OAI221_X1 port map( B1 => n6230, B2 => n4771, C1 => n6226, C2 => 
                           n7371, A => n7370, ZN => n7376);
   U3176 : NAND2_X1 port map( A1 => n6218, A2 => n7373, ZN => n7374);
   U3177 : NAND4_X1 port map( A1 => n1258, A2 => n1259, A3 => n1257, A4 => 
                           n7374, ZN => n7375);
   U3178 : OAI21_X1 port map( B1 => n7376, B2 => n7375, A => n6234, ZN => n7378
                           );
   U3179 : AOI22_X1 port map( A1 => n6179, A2 => n4980, B1 => DATAIN(23), B2 =>
                           n6177, ZN => n7377);
   U3180 : OAI211_X1 port map( C1 => n2275, C2 => n6183, A => n7378, B => n7377
                           , ZN => n7379);
   U3181 : NOR4_X1 port map( A1 => n7382, A2 => n7381, A3 => n7380, A4 => n7379
                           , ZN => n7383);
   U3182 : OAI21_X1 port map( B1 => n2662, B2 => n6239, A => n7383, ZN => n3023
                           );
   U3183 : OAI222_X1 port map( A1 => n6192, A2 => n4741, B1 => n2148, B2 => 
                           n6189, C1 => n6184, C2 => n4671, ZN => n7401);
   U3184 : AOI22_X1 port map( A1 => n6198, A2 => n5044, B1 => n6195, B2 => 
                           n7577, ZN => n7385);
   U3185 : OAI221_X1 port map( B1 => n2710, B2 => n6204, C1 => n2742, C2 => 
                           n6201, A => n7385, ZN => n7400);
   U3186 : AOI22_X1 port map( A1 => n6210, A2 => n5076, B1 => n6207, B2 => 
                           n7386, ZN => n7387);
   U3187 : OAI221_X1 port map( B1 => n2212, B2 => n6216, C1 => n2084, C2 => 
                           n6213, A => n7387, ZN => n7399);
   U3188 : AOI22_X1 port map( A1 => n2934, A2 => n6225, B1 => n7388, B2 => 
                           n6222, ZN => n7389);
   U3189 : OAI221_X1 port map( B1 => n6231, B2 => n4767, C1 => n6226, C2 => 
                           n7390, A => n7389, ZN => n7395);
   U3190 : NAND2_X1 port map( A1 => n6219, A2 => n7392, ZN => n7393);
   U3191 : NAND4_X1 port map( A1 => n1275, A2 => n1276, A3 => n1274, A4 => 
                           n7393, ZN => n7394);
   U3192 : OAI21_X1 port map( B1 => n7395, B2 => n7394, A => n6234, ZN => n7397
                           );
   U3193 : AOI22_X1 port map( A1 => n6179, A2 => n4979, B1 => DATAIN(24), B2 =>
                           n6177, ZN => n7396);
   U3194 : OAI211_X1 port map( C1 => n2276, C2 => n6183, A => n7397, B => n7396
                           , ZN => n7398);
   U3195 : NOR4_X1 port map( A1 => n7401, A2 => n7400, A3 => n7399, A4 => n7398
                           , ZN => n7402);
   U3196 : OAI21_X1 port map( B1 => n2661, B2 => n6238, A => n7402, ZN => n3022
                           );
   U3197 : OAI222_X1 port map( A1 => n6192, A2 => n4739, B1 => n2149, B2 => 
                           n6189, C1 => n6184, C2 => n4670, ZN => n7420);
   U3198 : AOI22_X1 port map( A1 => n6198, A2 => n5043, B1 => n6195, B2 => 
                           n7578, ZN => n7404);
   U3199 : OAI221_X1 port map( B1 => n2711, B2 => n6204, C1 => n2743, C2 => 
                           n6201, A => n7404, ZN => n7419);
   U3200 : AOI22_X1 port map( A1 => n6210, A2 => n5075, B1 => n6207, B2 => 
                           n7405, ZN => n7406);
   U3201 : OAI221_X1 port map( B1 => n2213, B2 => n6216, C1 => n2085, C2 => 
                           n6213, A => n7406, ZN => n7418);
   U3202 : AOI22_X1 port map( A1 => n2935, A2 => n6225, B1 => n7407, B2 => 
                           n6222, ZN => n7408);
   U3203 : OAI221_X1 port map( B1 => n6231, B2 => n4775, C1 => n6226, C2 => 
                           n7409, A => n7408, ZN => n7414);
   U3204 : NAND2_X1 port map( A1 => n6219, A2 => n7411, ZN => n7412);
   U3205 : NAND4_X1 port map( A1 => n1292, A2 => n1293, A3 => n1291, A4 => 
                           n7412, ZN => n7413);
   U3206 : OAI21_X1 port map( B1 => n7414, B2 => n7413, A => n6234, ZN => n7416
                           );
   U3207 : AOI22_X1 port map( A1 => n6179, A2 => n4978, B1 => DATAIN(25), B2 =>
                           n6178, ZN => n7415);
   U3208 : OAI211_X1 port map( C1 => n2277, C2 => n6183, A => n7416, B => n7415
                           , ZN => n7417);
   U3209 : NOR4_X1 port map( A1 => n7420, A2 => n7419, A3 => n7418, A4 => n7417
                           , ZN => n7421);
   U3210 : OAI21_X1 port map( B1 => n2660, B2 => n6238, A => n7421, ZN => n3021
                           );
   U3211 : OAI222_X1 port map( A1 => n6192, A2 => n4737, B1 => n2150, B2 => 
                           n6189, C1 => n6184, C2 => n4669, ZN => n7439);
   U3212 : AOI22_X1 port map( A1 => n6198, A2 => n5042, B1 => n6195, B2 => 
                           n7579, ZN => n7423);
   U3213 : OAI221_X1 port map( B1 => n2712, B2 => n6204, C1 => n2744, C2 => 
                           n6201, A => n7423, ZN => n7438);
   U3214 : AOI22_X1 port map( A1 => n6210, A2 => n5074, B1 => n6207, B2 => 
                           n7424, ZN => n7425);
   U3215 : OAI221_X1 port map( B1 => n2214, B2 => n6216, C1 => n2086, C2 => 
                           n6213, A => n7425, ZN => n7437);
   U3216 : AOI22_X1 port map( A1 => n2936, A2 => n6225, B1 => n7426, B2 => 
                           n6222, ZN => n7427);
   U3217 : OAI221_X1 port map( B1 => n6231, B2 => n4773, C1 => n6226, C2 => 
                           n7428, A => n7427, ZN => n7433);
   U3218 : NAND2_X1 port map( A1 => n6219, A2 => n7430, ZN => n7431);
   U3219 : NAND4_X1 port map( A1 => n1309, A2 => n1310, A3 => n1308, A4 => 
                           n7431, ZN => n7432);
   U3220 : OAI21_X1 port map( B1 => n7433, B2 => n7432, A => n6234, ZN => n7435
                           );
   U3221 : AOI22_X1 port map( A1 => n6179, A2 => n4977, B1 => DATAIN(26), B2 =>
                           n6178, ZN => n7434);
   U3222 : OAI211_X1 port map( C1 => n2278, C2 => n6182, A => n7435, B => n7434
                           , ZN => n7436);
   U3223 : NOR4_X1 port map( A1 => n7439, A2 => n7438, A3 => n7437, A4 => n7436
                           , ZN => n7440);
   U3224 : OAI21_X1 port map( B1 => n2659, B2 => n6238, A => n7440, ZN => n3020
                           );
   U3225 : OAI222_X1 port map( A1 => n6192, A2 => n4747, B1 => n2151, B2 => 
                           n6189, C1 => n6184, C2 => n4668, ZN => n7458);
   U3226 : AOI22_X1 port map( A1 => n6198, A2 => n5041, B1 => n6195, B2 => 
                           n7580, ZN => n7442);
   U3227 : OAI221_X1 port map( B1 => n2713, B2 => n6204, C1 => n2745, C2 => 
                           n6201, A => n7442, ZN => n7457);
   U3228 : AOI22_X1 port map( A1 => n6210, A2 => n5073, B1 => n6207, B2 => 
                           n7443, ZN => n7444);
   U3229 : OAI221_X1 port map( B1 => n2215, B2 => n6216, C1 => n2087, C2 => 
                           n6213, A => n7444, ZN => n7456);
   U3230 : AOI22_X1 port map( A1 => n2937, A2 => n6225, B1 => n7445, B2 => 
                           n6222, ZN => n7446);
   U3231 : OAI221_X1 port map( B1 => n6231, B2 => n4755, C1 => n6226, C2 => 
                           n7447, A => n7446, ZN => n7452);
   U3232 : NAND2_X1 port map( A1 => n6219, A2 => n7449, ZN => n7450);
   U3233 : NAND4_X1 port map( A1 => n1326, A2 => n1327, A3 => n1325, A4 => 
                           n7450, ZN => n7451);
   U3234 : OAI21_X1 port map( B1 => n7452, B2 => n7451, A => n6234, ZN => n7454
                           );
   U3235 : AOI22_X1 port map( A1 => n6179, A2 => n4976, B1 => DATAIN(27), B2 =>
                           n6178, ZN => n7453);
   U3236 : OAI211_X1 port map( C1 => n2279, C2 => n6183, A => n7454, B => n7453
                           , ZN => n7455);
   U3237 : NOR4_X1 port map( A1 => n7458, A2 => n7457, A3 => n7456, A4 => n7455
                           , ZN => n7459);
   U3238 : OAI21_X1 port map( B1 => n2658, B2 => n6238, A => n7459, ZN => n3019
                           );
   U3239 : OAI222_X1 port map( A1 => n6192, A2 => n4745, B1 => n2152, B2 => 
                           n6189, C1 => n6184, C2 => n4667, ZN => n7477);
   U3240 : AOI22_X1 port map( A1 => n6198, A2 => n5040, B1 => n6195, B2 => 
                           n7581, ZN => n7461);
   U3241 : OAI221_X1 port map( B1 => n2714, B2 => n6204, C1 => n2746, C2 => 
                           n6201, A => n7461, ZN => n7476);
   U3242 : AOI22_X1 port map( A1 => n6210, A2 => n5072, B1 => n6207, B2 => 
                           n7462, ZN => n7463);
   U3243 : OAI221_X1 port map( B1 => n2216, B2 => n6216, C1 => n2088, C2 => 
                           n6213, A => n7463, ZN => n7475);
   U3244 : AOI22_X1 port map( A1 => n2938, A2 => n6225, B1 => n7464, B2 => 
                           n6222, ZN => n7465);
   U3245 : OAI221_X1 port map( B1 => n6231, B2 => n4779, C1 => n6226, C2 => 
                           n7466, A => n7465, ZN => n7471);
   U3246 : NAND2_X1 port map( A1 => n6219, A2 => n7468, ZN => n7469);
   U3247 : NAND4_X1 port map( A1 => n1343, A2 => n1344, A3 => n1342, A4 => 
                           n7469, ZN => n7470);
   U3248 : OAI21_X1 port map( B1 => n7471, B2 => n7470, A => n6234, ZN => n7473
                           );
   U3249 : AOI22_X1 port map( A1 => n6179, A2 => n4975, B1 => DATAIN(28), B2 =>
                           n6178, ZN => n7472);
   U3250 : OAI211_X1 port map( C1 => n2280, C2 => n6182, A => n7473, B => n7472
                           , ZN => n7474);
   U3251 : NOR4_X1 port map( A1 => n7477, A2 => n7476, A3 => n7475, A4 => n7474
                           , ZN => n7478);
   U3252 : OAI21_X1 port map( B1 => n2657, B2 => n6238, A => n7478, ZN => n3018
                           );
   U3253 : OAI222_X1 port map( A1 => n6192, A2 => n4743, B1 => n2153, B2 => 
                           n6189, C1 => n6184, C2 => n4666, ZN => n7496);
   U3254 : AOI22_X1 port map( A1 => n6198, A2 => n5039, B1 => n6195, B2 => 
                           n7582, ZN => n7480);
   U3255 : OAI221_X1 port map( B1 => n2715, B2 => n6204, C1 => n2747, C2 => 
                           n6201, A => n7480, ZN => n7495);
   U3256 : AOI22_X1 port map( A1 => n6210, A2 => n5071, B1 => n6207, B2 => 
                           n7481, ZN => n7482);
   U3257 : OAI221_X1 port map( B1 => n2217, B2 => n6216, C1 => n2089, C2 => 
                           n6213, A => n7482, ZN => n7494);
   U3258 : AOI22_X1 port map( A1 => n2939, A2 => n6225, B1 => n7483, B2 => 
                           n6222, ZN => n7484);
   U3259 : OAI221_X1 port map( B1 => n6231, B2 => n4777, C1 => n6226, C2 => 
                           n7485, A => n7484, ZN => n7490);
   U3260 : NAND2_X1 port map( A1 => n6219, A2 => n7487, ZN => n7488);
   U3261 : NAND4_X1 port map( A1 => n1360, A2 => n1361, A3 => n1359, A4 => 
                           n7488, ZN => n7489);
   U3262 : OAI21_X1 port map( B1 => n7490, B2 => n7489, A => n6234, ZN => n7492
                           );
   U3263 : AOI22_X1 port map( A1 => n6179, A2 => n4974, B1 => DATAIN(29), B2 =>
                           n6178, ZN => n7491);
   U3264 : OAI211_X1 port map( C1 => n2281, C2 => n6183, A => n7492, B => n7491
                           , ZN => n7493);
   U3265 : NOR4_X1 port map( A1 => n7496, A2 => n7495, A3 => n7494, A4 => n7493
                           , ZN => n7497);
   U3266 : OAI21_X1 port map( B1 => n2656, B2 => n6238, A => n7497, ZN => n3017
                           );
   U3267 : OAI222_X1 port map( A1 => n6192, A2 => n4749, B1 => n2154, B2 => 
                           n6189, C1 => n6184, C2 => n4665, ZN => n7517);
   U3268 : AOI22_X1 port map( A1 => n6198, A2 => n5038, B1 => n6195, B2 => 
                           n7583, ZN => n7499);
   U3269 : OAI221_X1 port map( B1 => n2716, B2 => n6204, C1 => n2748, C2 => 
                           n6201, A => n7499, ZN => n7516);
   U3270 : AOI22_X1 port map( A1 => n6210, A2 => n5070, B1 => n6207, B2 => 
                           n7500, ZN => n7501);
   U3271 : OAI221_X1 port map( B1 => n2218, B2 => n6216, C1 => n2090, C2 => 
                           n6213, A => n7501, ZN => n7515);
   U3272 : AOI22_X1 port map( A1 => n2940, A2 => n6225, B1 => n7502, B2 => 
                           n6222, ZN => n7503);
   U3273 : OAI221_X1 port map( B1 => n6231, B2 => n4781, C1 => n6226, C2 => 
                           n7504, A => n7503, ZN => n7509);
   U3274 : NAND2_X1 port map( A1 => n6219, A2 => n7506, ZN => n7507);
   U3275 : NAND4_X1 port map( A1 => n1377, A2 => n1378, A3 => n1376, A4 => 
                           n7507, ZN => n7508);
   U3276 : OAI21_X1 port map( B1 => n7509, B2 => n7508, A => n6234, ZN => n7513
                           );
   U3277 : AOI22_X1 port map( A1 => n6179, A2 => n4973, B1 => DATAIN(30), B2 =>
                           n6178, ZN => n7512);
   U3278 : OAI211_X1 port map( C1 => n2282, C2 => n6182, A => n7513, B => n7512
                           , ZN => n7514);
   U3279 : NOR4_X1 port map( A1 => n7517, A2 => n7516, A3 => n7515, A4 => n7514
                           , ZN => n7518);
   U3280 : OAI21_X1 port map( B1 => n2655, B2 => n6238, A => n7518, ZN => n3016
                           );
   U3281 : OAI222_X1 port map( A1 => n6192, A2 => n4751, B1 => n2155, B2 => 
                           n6189, C1 => n6184, C2 => n4664, ZN => n7549);
   U3282 : AOI22_X1 port map( A1 => n6198, A2 => n5037, B1 => n6195, B2 => 
                           n7584, ZN => n7523);
   U3283 : OAI221_X1 port map( B1 => n2717, B2 => n6204, C1 => n2749, C2 => 
                           n6201, A => n7523, ZN => n7548);
   U3284 : AOI22_X1 port map( A1 => n6210, A2 => n5069, B1 => n6207, B2 => 
                           n7526, ZN => n7527);
   U3285 : OAI221_X1 port map( B1 => n2219, B2 => n6216, C1 => n2091, C2 => 
                           n6213, A => n7527, ZN => n7547);
   U3286 : OAI22_X1 port map( A1 => n3773, A2 => n4901, B1 => n2315, B2 => 
                           n4899, ZN => n7530);
   U3287 : AOI221_X1 port map( B1 => n6219, B2 => n7531, C1 => n6312, C2 => 
                           n7587, A => n7530, ZN => n7539);
   U3288 : AOI222_X1 port map( A1 => n6335, A2 => n4093, B1 => n6324, B2 => 
                           n7585, C1 => n6338, C2 => n4061, ZN => n7538);
   U3289 : AOI22_X1 port map( A1 => n2941, A2 => n6225, B1 => n7532, B2 => 
                           n6222, ZN => n7533);
   U3290 : OAI221_X1 port map( B1 => n4815, B2 => n6231, C1 => n7534, C2 => 
                           n6226, A => n7533, ZN => n7536);
   U3291 : NOR4_X1 port map( A1 => n7536, A2 => n1425, A3 => n1424, A4 => n1421
                           , ZN => n7537);
   U3292 : NAND3_X1 port map( A1 => n7539, A2 => n7538, A3 => n7537, ZN => 
                           n7541);
   U3293 : AOI22_X1 port map( A1 => n6234, A2 => n7541, B1 => n4896, B2 => 
                           n7540, ZN => n7543);
   U3294 : OAI221_X1 port map( B1 => n2251, B2 => n7545, C1 => n7544, C2 => 
                           n6374, A => n7543, ZN => n7546);
   U3295 : NOR4_X1 port map( A1 => n7549, A2 => n7548, A3 => n7547, A4 => n7546
                           , ZN => n7550);
   U3296 : OAI21_X1 port map( B1 => n6238, B2 => n7551, A => n7550, ZN => n3015
                           );
   U3297 : MUX2_X1 port map( A => n5235, B => DATAIN(0), S => n6241, Z => n3047
                           );
   U3298 : MUX2_X1 port map( A => n5297, B => DATAIN(1), S => n6241, Z => n3048
                           );
   U3299 : MUX2_X1 port map( A => n5296, B => DATAIN(2), S => n6241, Z => n3049
                           );
   U3300 : MUX2_X1 port map( A => n5295, B => DATAIN(3), S => n6241, Z => n3050
                           );
   U3301 : MUX2_X1 port map( A => n5294, B => DATAIN(4), S => n6241, Z => n3051
                           );
   U3302 : MUX2_X1 port map( A => n5293, B => DATAIN(5), S => n6241, Z => n3052
                           );
   U3303 : MUX2_X1 port map( A => n5292, B => DATAIN(6), S => n6241, Z => n3053
                           );
   U3304 : MUX2_X1 port map( A => n5291, B => DATAIN(7), S => n6241, Z => n3054
                           );
   U3305 : MUX2_X1 port map( A => n5290, B => DATAIN(8), S => n6241, Z => n3055
                           );
   U3306 : MUX2_X1 port map( A => n5289, B => DATAIN(9), S => n6241, Z => n3056
                           );
   U3307 : MUX2_X1 port map( A => n5288, B => DATAIN(10), S => n6241, Z => 
                           n3057);
   U3308 : MUX2_X1 port map( A => n5287, B => DATAIN(11), S => n6241, Z => 
                           n3058);
   U3309 : MUX2_X1 port map( A => n5286, B => DATAIN(12), S => n6242, Z => 
                           n3059);
   U3310 : MUX2_X1 port map( A => n5285, B => DATAIN(13), S => n6242, Z => 
                           n3060);
   U3311 : MUX2_X1 port map( A => n5284, B => DATAIN(14), S => n6242, Z => 
                           n3061);
   U3312 : MUX2_X1 port map( A => n5283, B => DATAIN(15), S => n6242, Z => 
                           n3062);
   U3313 : MUX2_X1 port map( A => n5282, B => DATAIN(16), S => n6242, Z => 
                           n3063);
   U3314 : MUX2_X1 port map( A => n5281, B => DATAIN(17), S => n6242, Z => 
                           n3064);
   U3315 : MUX2_X1 port map( A => n5280, B => DATAIN(18), S => n6242, Z => 
                           n3065);
   U3316 : MUX2_X1 port map( A => n5279, B => DATAIN(19), S => n6242, Z => 
                           n3066);
   U3317 : MUX2_X1 port map( A => n5278, B => DATAIN(20), S => n6242, Z => 
                           n3067);
   U3318 : MUX2_X1 port map( A => n5277, B => DATAIN(21), S => n6242, Z => 
                           n3068);
   U3319 : MUX2_X1 port map( A => n5276, B => DATAIN(22), S => n6242, Z => 
                           n3069);
   U3320 : MUX2_X1 port map( A => n5275, B => DATAIN(23), S => n6242, Z => 
                           n3070);
   U3321 : MUX2_X1 port map( A => n5274, B => DATAIN(24), S => n6243, Z => 
                           n3071);
   U3322 : MUX2_X1 port map( A => n5273, B => DATAIN(25), S => n6243, Z => 
                           n3072);
   U3323 : MUX2_X1 port map( A => n5272, B => DATAIN(26), S => n6243, Z => 
                           n3073);
   U3324 : MUX2_X1 port map( A => n5271, B => DATAIN(27), S => n6243, Z => 
                           n3074);
   U3325 : MUX2_X1 port map( A => n5270, B => DATAIN(28), S => n6243, Z => 
                           n3075);
   U3326 : MUX2_X1 port map( A => n5269, B => DATAIN(29), S => n6243, Z => 
                           n3076);
   U3327 : MUX2_X1 port map( A => n5268, B => DATAIN(30), S => n6243, Z => 
                           n3077);
   U3328 : MUX2_X1 port map( A => n5234, B => DATAIN(31), S => n6243, Z => 
                           n3078);
   U3329 : MUX2_X1 port map( A => n5171, B => DATAIN(0), S => n6244, Z => n3111
                           );
   U3330 : MUX2_X1 port map( A => n5167, B => DATAIN(1), S => n6244, Z => n3112
                           );
   U3331 : MUX2_X1 port map( A => n5166, B => DATAIN(2), S => n6244, Z => n3113
                           );
   U3332 : MUX2_X1 port map( A => n5165, B => DATAIN(3), S => n6244, Z => n3114
                           );
   U3333 : MUX2_X1 port map( A => n5164, B => DATAIN(4), S => n6244, Z => n3115
                           );
   U3334 : MUX2_X1 port map( A => n5163, B => DATAIN(5), S => n6244, Z => n3116
                           );
   U3335 : MUX2_X1 port map( A => n5162, B => DATAIN(6), S => n6244, Z => n3117
                           );
   U3336 : MUX2_X1 port map( A => n5161, B => DATAIN(7), S => n6244, Z => n3118
                           );
   U3337 : MUX2_X1 port map( A => n5160, B => DATAIN(8), S => n6244, Z => n3119
                           );
   U3338 : MUX2_X1 port map( A => n5159, B => DATAIN(9), S => n6244, Z => n3120
                           );
   U3339 : MUX2_X1 port map( A => n5158, B => DATAIN(10), S => n6244, Z => 
                           n3121);
   U3340 : MUX2_X1 port map( A => n5157, B => DATAIN(11), S => n6244, Z => 
                           n3122);
   U3341 : MUX2_X1 port map( A => n5156, B => DATAIN(12), S => n6245, Z => 
                           n3123);
   U3342 : MUX2_X1 port map( A => n5155, B => DATAIN(13), S => n6245, Z => 
                           n3124);
   U3343 : MUX2_X1 port map( A => n5154, B => DATAIN(14), S => n6245, Z => 
                           n3125);
   U3344 : MUX2_X1 port map( A => n5153, B => DATAIN(15), S => n6245, Z => 
                           n3126);
   U3345 : MUX2_X1 port map( A => n5152, B => DATAIN(16), S => n6245, Z => 
                           n3127);
   U3346 : MUX2_X1 port map( A => n5151, B => DATAIN(17), S => n6245, Z => 
                           n3128);
   U3347 : MUX2_X1 port map( A => n5150, B => DATAIN(18), S => n6245, Z => 
                           n3129);
   U3348 : MUX2_X1 port map( A => n5149, B => DATAIN(19), S => n6245, Z => 
                           n3130);
   U3349 : MUX2_X1 port map( A => n5148, B => DATAIN(20), S => n6245, Z => 
                           n3131);
   U3350 : MUX2_X1 port map( A => n5147, B => DATAIN(21), S => n6245, Z => 
                           n3132);
   U3351 : MUX2_X1 port map( A => n5146, B => DATAIN(22), S => n6245, Z => 
                           n3133);
   U3352 : MUX2_X1 port map( A => n5145, B => DATAIN(23), S => n6245, Z => 
                           n3134);
   U3353 : MUX2_X1 port map( A => n5144, B => DATAIN(24), S => n6246, Z => 
                           n3135);
   U3354 : MUX2_X1 port map( A => n5143, B => DATAIN(25), S => n6246, Z => 
                           n3136);
   U3355 : MUX2_X1 port map( A => n5142, B => DATAIN(26), S => n6246, Z => 
                           n3137);
   U3356 : MUX2_X1 port map( A => n5141, B => DATAIN(27), S => n6246, Z => 
                           n3138);
   U3357 : MUX2_X1 port map( A => n5140, B => DATAIN(28), S => n6246, Z => 
                           n3139);
   U3358 : MUX2_X1 port map( A => n5139, B => DATAIN(29), S => n6246, Z => 
                           n3140);
   U3359 : MUX2_X1 port map( A => n5138, B => DATAIN(30), S => n6246, Z => 
                           n3141);
   U3360 : MUX2_X1 port map( A => n5137, B => DATAIN(31), S => n6246, Z => 
                           n3142);
   U3361 : MUX2_X1 port map( A => n5680, B => DATAIN(0), S => n6247, Z => n3239
                           );
   U3362 : MUX2_X1 port map( A => n5545, B => DATAIN(1), S => n6247, Z => n3240
                           );
   U3363 : MUX2_X1 port map( A => n5544, B => DATAIN(2), S => n6247, Z => n3241
                           );
   U3364 : MUX2_X1 port map( A => n5543, B => DATAIN(3), S => n6247, Z => n3242
                           );
   U3365 : MUX2_X1 port map( A => n5542, B => DATAIN(4), S => n6247, Z => n3243
                           );
   U3366 : MUX2_X1 port map( A => n5541, B => DATAIN(5), S => n6247, Z => n3244
                           );
   U3367 : MUX2_X1 port map( A => n5540, B => DATAIN(6), S => n6247, Z => n3245
                           );
   U3368 : MUX2_X1 port map( A => n5539, B => DATAIN(7), S => n6247, Z => n3246
                           );
   U3369 : MUX2_X1 port map( A => n5538, B => DATAIN(8), S => n6247, Z => n3247
                           );
   U3370 : MUX2_X1 port map( A => n5537, B => DATAIN(9), S => n6247, Z => n3248
                           );
   U3371 : MUX2_X1 port map( A => n5536, B => DATAIN(10), S => n6247, Z => 
                           n3249);
   U3372 : MUX2_X1 port map( A => n5535, B => DATAIN(11), S => n6247, Z => 
                           n3250);
   U3373 : MUX2_X1 port map( A => n5534, B => DATAIN(12), S => n6248, Z => 
                           n3251);
   U3374 : MUX2_X1 port map( A => n5533, B => DATAIN(13), S => n6248, Z => 
                           n3252);
   U3375 : MUX2_X1 port map( A => n5532, B => DATAIN(14), S => n6248, Z => 
                           n3253);
   U3376 : MUX2_X1 port map( A => n5531, B => DATAIN(15), S => n6248, Z => 
                           n3254);
   U3377 : MUX2_X1 port map( A => n5530, B => DATAIN(16), S => n6248, Z => 
                           n3255);
   U3378 : MUX2_X1 port map( A => n5529, B => DATAIN(17), S => n6248, Z => 
                           n3256);
   U3379 : MUX2_X1 port map( A => n5528, B => DATAIN(18), S => n6248, Z => 
                           n3257);
   U3380 : MUX2_X1 port map( A => n5527, B => DATAIN(19), S => n6248, Z => 
                           n3258);
   U3381 : MUX2_X1 port map( A => n5526, B => DATAIN(20), S => n6248, Z => 
                           n3259);
   U3382 : MUX2_X1 port map( A => n5525, B => DATAIN(21), S => n6248, Z => 
                           n3260);
   U3383 : MUX2_X1 port map( A => n5524, B => DATAIN(22), S => n6248, Z => 
                           n3261);
   U3384 : MUX2_X1 port map( A => n5523, B => DATAIN(23), S => n6248, Z => 
                           n3262);
   U3385 : MUX2_X1 port map( A => n5522, B => DATAIN(24), S => n6249, Z => 
                           n3263);
   U3386 : MUX2_X1 port map( A => n5521, B => DATAIN(25), S => n6249, Z => 
                           n3264);
   U3387 : MUX2_X1 port map( A => n5520, B => DATAIN(26), S => n6249, Z => 
                           n3265);
   U3388 : MUX2_X1 port map( A => n5519, B => DATAIN(27), S => n6249, Z => 
                           n3266);
   U3389 : MUX2_X1 port map( A => n5518, B => DATAIN(28), S => n6249, Z => 
                           n3267);
   U3390 : MUX2_X1 port map( A => n5517, B => DATAIN(29), S => n6249, Z => 
                           n3268);
   U3391 : MUX2_X1 port map( A => n5516, B => DATAIN(30), S => n6249, Z => 
                           n3269);
   U3392 : MUX2_X1 port map( A => n5515, B => DATAIN(31), S => n6249, Z => 
                           n3270);
   U3393 : MUX2_X1 port map( A => n5486, B => DATAIN(0), S => n6250, Z => n3271
                           );
   U3394 : MUX2_X1 port map( A => n5482, B => DATAIN(1), S => n6250, Z => n3272
                           );
   U3395 : MUX2_X1 port map( A => n5481, B => DATAIN(2), S => n6250, Z => n3273
                           );
   U3396 : MUX2_X1 port map( A => n5480, B => DATAIN(3), S => n6250, Z => n3274
                           );
   U3397 : MUX2_X1 port map( A => n5479, B => DATAIN(4), S => n6250, Z => n3275
                           );
   U3398 : MUX2_X1 port map( A => n5478, B => DATAIN(5), S => n6250, Z => n3276
                           );
   U3399 : MUX2_X1 port map( A => n5477, B => DATAIN(6), S => n6250, Z => n3277
                           );
   U3400 : MUX2_X1 port map( A => n5476, B => DATAIN(7), S => n6250, Z => n3278
                           );
   U3401 : MUX2_X1 port map( A => n5475, B => DATAIN(8), S => n6250, Z => n3279
                           );
   U3402 : MUX2_X1 port map( A => n5474, B => DATAIN(9), S => n6250, Z => n3280
                           );
   U3403 : MUX2_X1 port map( A => n5473, B => DATAIN(10), S => n6250, Z => 
                           n3281);
   U3404 : MUX2_X1 port map( A => n5472, B => DATAIN(11), S => n6251, Z => 
                           n3282);
   U3405 : MUX2_X1 port map( A => n5471, B => DATAIN(12), S => n6251, Z => 
                           n3283);
   U3406 : MUX2_X1 port map( A => n5470, B => DATAIN(13), S => n6251, Z => 
                           n3284);
   U3407 : MUX2_X1 port map( A => n5469, B => DATAIN(14), S => n6251, Z => 
                           n3285);
   U3408 : MUX2_X1 port map( A => n5468, B => DATAIN(15), S => n6251, Z => 
                           n3286);
   U3409 : MUX2_X1 port map( A => n5467, B => DATAIN(16), S => n6251, Z => 
                           n3287);
   U3410 : MUX2_X1 port map( A => n5466, B => DATAIN(17), S => n6251, Z => 
                           n3288);
   U3411 : MUX2_X1 port map( A => n5465, B => DATAIN(18), S => n6251, Z => 
                           n3289);
   U3412 : MUX2_X1 port map( A => n5464, B => DATAIN(19), S => n6251, Z => 
                           n3290);
   U3413 : MUX2_X1 port map( A => n5463, B => DATAIN(20), S => n6251, Z => 
                           n3291);
   U3414 : MUX2_X1 port map( A => n5462, B => DATAIN(21), S => n6251, Z => 
                           n3292);
   U3415 : MUX2_X1 port map( A => n5461, B => DATAIN(22), S => n6251, Z => 
                           n3293);
   U3416 : MUX2_X1 port map( A => n5460, B => DATAIN(23), S => n6252, Z => 
                           n3294);
   U3417 : MUX2_X1 port map( A => n5459, B => DATAIN(24), S => n6252, Z => 
                           n3295);
   U3418 : MUX2_X1 port map( A => n5458, B => DATAIN(25), S => n6252, Z => 
                           n3296);
   U3419 : MUX2_X1 port map( A => n5457, B => DATAIN(26), S => n6252, Z => 
                           n3297);
   U3420 : MUX2_X1 port map( A => n5456, B => DATAIN(27), S => n6252, Z => 
                           n3298);
   U3421 : MUX2_X1 port map( A => n5455, B => DATAIN(28), S => n6252, Z => 
                           n3299);
   U3422 : MUX2_X1 port map( A => n5454, B => DATAIN(29), S => n6252, Z => 
                           n3300);
   U3423 : MUX2_X1 port map( A => n5453, B => DATAIN(30), S => n6252, Z => 
                           n3301);
   U3424 : MUX2_X1 port map( A => n5776, B => DATAIN(0), S => n6253, Z => n3303
                           );
   U3425 : MUX2_X1 port map( A => n5775, B => DATAIN(1), S => n6253, Z => n3304
                           );
   U3426 : MUX2_X1 port map( A => n5774, B => DATAIN(2), S => n6253, Z => n3305
                           );
   U3427 : MUX2_X1 port map( A => n5773, B => DATAIN(3), S => n6253, Z => n3306
                           );
   U3428 : MUX2_X1 port map( A => n5772, B => DATAIN(4), S => n6253, Z => n3307
                           );
   U3429 : MUX2_X1 port map( A => n5771, B => DATAIN(5), S => n6253, Z => n3308
                           );
   U3430 : MUX2_X1 port map( A => n5770, B => DATAIN(6), S => n6253, Z => n3309
                           );
   U3431 : MUX2_X1 port map( A => n5769, B => DATAIN(7), S => n6253, Z => n3310
                           );
   U3432 : MUX2_X1 port map( A => n5768, B => DATAIN(8), S => n6253, Z => n3311
                           );
   U3433 : MUX2_X1 port map( A => n5767, B => DATAIN(9), S => n6253, Z => n3312
                           );
   U3434 : MUX2_X1 port map( A => n5766, B => DATAIN(10), S => n6253, Z => 
                           n3313);
   U3435 : MUX2_X1 port map( A => n5765, B => DATAIN(11), S => n6253, Z => 
                           n3314);
   U3436 : MUX2_X1 port map( A => n5764, B => DATAIN(12), S => n6254, Z => 
                           n3315);
   U3437 : MUX2_X1 port map( A => n5763, B => DATAIN(13), S => n6254, Z => 
                           n3316);
   U3438 : MUX2_X1 port map( A => n5762, B => DATAIN(14), S => n6254, Z => 
                           n3317);
   U3439 : MUX2_X1 port map( A => n5761, B => DATAIN(15), S => n6254, Z => 
                           n3318);
   U3440 : MUX2_X1 port map( A => n5760, B => DATAIN(16), S => n6254, Z => 
                           n3319);
   U3441 : MUX2_X1 port map( A => n5759, B => DATAIN(17), S => n6254, Z => 
                           n3320);
   U3442 : MUX2_X1 port map( A => n5758, B => DATAIN(18), S => n6254, Z => 
                           n3321);
   U3443 : MUX2_X1 port map( A => n5757, B => DATAIN(19), S => n6254, Z => 
                           n3322);
   U3444 : MUX2_X1 port map( A => n5756, B => DATAIN(20), S => n6254, Z => 
                           n3323);
   U3445 : MUX2_X1 port map( A => n5755, B => DATAIN(21), S => n6254, Z => 
                           n3324);
   U3446 : MUX2_X1 port map( A => n5754, B => DATAIN(22), S => n6254, Z => 
                           n3325);
   U3447 : MUX2_X1 port map( A => n5753, B => DATAIN(23), S => n6254, Z => 
                           n3326);
   U3448 : MUX2_X1 port map( A => n5752, B => DATAIN(24), S => n6255, Z => 
                           n3327);
   U3449 : MUX2_X1 port map( A => n5751, B => DATAIN(25), S => n6255, Z => 
                           n3328);
   U3450 : MUX2_X1 port map( A => n5750, B => DATAIN(26), S => n6255, Z => 
                           n3329);
   U3451 : MUX2_X1 port map( A => n5749, B => DATAIN(27), S => n6255, Z => 
                           n3330);
   U3452 : MUX2_X1 port map( A => n5748, B => DATAIN(28), S => n6255, Z => 
                           n3331);
   U3453 : MUX2_X1 port map( A => n5747, B => DATAIN(29), S => n6255, Z => 
                           n3332);
   U3454 : MUX2_X1 port map( A => n5746, B => DATAIN(30), S => n6255, Z => 
                           n3333);
   U3455 : MUX2_X1 port map( A => n5745, B => DATAIN(31), S => n6255, Z => 
                           n3334);
   U3456 : MUX2_X1 port map( A => n5237, B => DATAIN(0), S => n6256, Z => n3335
                           );
   U3457 : MUX2_X1 port map( A => n5267, B => DATAIN(1), S => n6256, Z => n3336
                           );
   U3458 : MUX2_X1 port map( A => n5266, B => DATAIN(2), S => n6256, Z => n3337
                           );
   U3459 : MUX2_X1 port map( A => n5265, B => DATAIN(3), S => n6256, Z => n3338
                           );
   U3460 : MUX2_X1 port map( A => n5264, B => DATAIN(4), S => n6256, Z => n3339
                           );
   U3461 : MUX2_X1 port map( A => n5263, B => DATAIN(5), S => n6256, Z => n3340
                           );
   U3462 : MUX2_X1 port map( A => n5262, B => DATAIN(6), S => n6256, Z => n3341
                           );
   U3463 : MUX2_X1 port map( A => n5261, B => DATAIN(7), S => n6256, Z => n3342
                           );
   U3464 : MUX2_X1 port map( A => n5260, B => DATAIN(8), S => n6256, Z => n3343
                           );
   U3465 : MUX2_X1 port map( A => n5259, B => DATAIN(9), S => n6256, Z => n3344
                           );
   U3466 : MUX2_X1 port map( A => n5258, B => DATAIN(10), S => n6256, Z => 
                           n3345);
   U3467 : MUX2_X1 port map( A => n5257, B => DATAIN(11), S => n6256, Z => 
                           n3346);
   U3468 : MUX2_X1 port map( A => n5256, B => DATAIN(12), S => n6257, Z => 
                           n3347);
   U3469 : MUX2_X1 port map( A => n5255, B => DATAIN(13), S => n6257, Z => 
                           n3348);
   U3470 : MUX2_X1 port map( A => n5254, B => DATAIN(14), S => n6257, Z => 
                           n3349);
   U3471 : MUX2_X1 port map( A => n5253, B => DATAIN(15), S => n6257, Z => 
                           n3350);
   U3472 : MUX2_X1 port map( A => n5252, B => DATAIN(16), S => n6257, Z => 
                           n3351);
   U3473 : MUX2_X1 port map( A => n5251, B => DATAIN(17), S => n6257, Z => 
                           n3352);
   U3474 : MUX2_X1 port map( A => n5250, B => DATAIN(18), S => n6257, Z => 
                           n3353);
   U3475 : MUX2_X1 port map( A => n5249, B => DATAIN(19), S => n6257, Z => 
                           n3354);
   U3476 : MUX2_X1 port map( A => n5248, B => DATAIN(20), S => n6257, Z => 
                           n3355);
   U3477 : MUX2_X1 port map( A => n5247, B => DATAIN(21), S => n6257, Z => 
                           n3356);
   U3478 : MUX2_X1 port map( A => n5246, B => DATAIN(22), S => n6257, Z => 
                           n3357);
   U3479 : MUX2_X1 port map( A => n5245, B => DATAIN(23), S => n6257, Z => 
                           n3358);
   U3480 : MUX2_X1 port map( A => n5244, B => DATAIN(24), S => n6258, Z => 
                           n3359);
   U3481 : MUX2_X1 port map( A => n5243, B => DATAIN(25), S => n6258, Z => 
                           n3360);
   U3482 : MUX2_X1 port map( A => n5242, B => DATAIN(26), S => n6258, Z => 
                           n3361);
   U3483 : MUX2_X1 port map( A => n5241, B => DATAIN(27), S => n6258, Z => 
                           n3362);
   U3484 : MUX2_X1 port map( A => n5240, B => DATAIN(28), S => n6258, Z => 
                           n3363);
   U3485 : MUX2_X1 port map( A => n5239, B => DATAIN(29), S => n6258, Z => 
                           n3364);
   U3486 : MUX2_X1 port map( A => n5238, B => DATAIN(30), S => n6258, Z => 
                           n3365);
   U3487 : MUX2_X1 port map( A => n5236, B => DATAIN(31), S => n6258, Z => 
                           n3366);
   U3488 : MUX2_X1 port map( A => n5579, B => DATAIN(0), S => n6259, Z => n3367
                           );
   U3489 : MUX2_X1 port map( A => n5578, B => DATAIN(1), S => n6259, Z => n3368
                           );
   U3490 : MUX2_X1 port map( A => n5577, B => DATAIN(2), S => n6259, Z => n3369
                           );
   U3491 : MUX2_X1 port map( A => n5576, B => DATAIN(3), S => n6259, Z => n3370
                           );
   U3492 : MUX2_X1 port map( A => n5575, B => DATAIN(4), S => n6259, Z => n3371
                           );
   U3493 : MUX2_X1 port map( A => n5574, B => DATAIN(5), S => n6259, Z => n3372
                           );
   U3494 : MUX2_X1 port map( A => n5573, B => DATAIN(6), S => n6259, Z => n3373
                           );
   U3495 : MUX2_X1 port map( A => n5572, B => DATAIN(7), S => n6259, Z => n3374
                           );
   U3496 : MUX2_X1 port map( A => n5571, B => DATAIN(8), S => n6259, Z => n3375
                           );
   U3497 : MUX2_X1 port map( A => n5570, B => DATAIN(9), S => n6259, Z => n3376
                           );
   U3498 : MUX2_X1 port map( A => n5569, B => DATAIN(10), S => n6259, Z => 
                           n3377);
   U3499 : MUX2_X1 port map( A => n5568, B => DATAIN(11), S => n6259, Z => 
                           n3378);
   U3500 : MUX2_X1 port map( A => n5567, B => DATAIN(12), S => n6260, Z => 
                           n3379);
   U3501 : MUX2_X1 port map( A => n5566, B => DATAIN(13), S => n6260, Z => 
                           n3380);
   U3502 : MUX2_X1 port map( A => n5565, B => DATAIN(14), S => n6260, Z => 
                           n3381);
   U3503 : MUX2_X1 port map( A => n5564, B => DATAIN(15), S => n6260, Z => 
                           n3382);
   U3504 : MUX2_X1 port map( A => n5563, B => DATAIN(16), S => n6260, Z => 
                           n3383);
   U3505 : MUX2_X1 port map( A => n5562, B => DATAIN(17), S => n6260, Z => 
                           n3384);
   U3506 : MUX2_X1 port map( A => n5561, B => DATAIN(18), S => n6260, Z => 
                           n3385);
   U3507 : MUX2_X1 port map( A => n5560, B => DATAIN(19), S => n6260, Z => 
                           n3386);
   U3508 : MUX2_X1 port map( A => n5559, B => DATAIN(20), S => n6260, Z => 
                           n3387);
   U3509 : MUX2_X1 port map( A => n5558, B => DATAIN(21), S => n6260, Z => 
                           n3388);
   U3510 : MUX2_X1 port map( A => n5557, B => DATAIN(22), S => n6260, Z => 
                           n3389);
   U3511 : MUX2_X1 port map( A => n5556, B => DATAIN(23), S => n6260, Z => 
                           n3390);
   U3512 : MUX2_X1 port map( A => n5555, B => DATAIN(24), S => n6261, Z => 
                           n3391);
   U3513 : MUX2_X1 port map( A => n5554, B => DATAIN(25), S => n6261, Z => 
                           n3392);
   U3514 : MUX2_X1 port map( A => n5553, B => DATAIN(26), S => n6261, Z => 
                           n3393);
   U3515 : MUX2_X1 port map( A => n5552, B => DATAIN(27), S => n6261, Z => 
                           n3394);
   U3516 : MUX2_X1 port map( A => n5551, B => DATAIN(28), S => n6261, Z => 
                           n3395);
   U3517 : MUX2_X1 port map( A => n5550, B => DATAIN(29), S => n6261, Z => 
                           n3396);
   U3518 : MUX2_X1 port map( A => n5549, B => DATAIN(30), S => n6261, Z => 
                           n3397);
   U3519 : MUX2_X1 port map( A => n5548, B => DATAIN(31), S => n6261, Z => 
                           n3398);
   U3520 : MUX2_X1 port map( A => n5743, B => DATAIN(0), S => n6262, Z => n3399
                           );
   U3521 : MUX2_X1 port map( A => n5742, B => DATAIN(1), S => n6262, Z => n3400
                           );
   U3522 : MUX2_X1 port map( A => n5741, B => DATAIN(2), S => n6262, Z => n3401
                           );
   U3523 : MUX2_X1 port map( A => n5740, B => DATAIN(3), S => n6262, Z => n3402
                           );
   U3524 : MUX2_X1 port map( A => n5739, B => DATAIN(4), S => n6262, Z => n3403
                           );
   U3525 : MUX2_X1 port map( A => n5738, B => DATAIN(5), S => n6262, Z => n3404
                           );
   U3526 : MUX2_X1 port map( A => n5737, B => DATAIN(6), S => n6262, Z => n3405
                           );
   U3527 : MUX2_X1 port map( A => n5736, B => DATAIN(7), S => n6262, Z => n3406
                           );
   U3528 : MUX2_X1 port map( A => n5735, B => DATAIN(8), S => n6262, Z => n3407
                           );
   U3529 : MUX2_X1 port map( A => n5734, B => DATAIN(9), S => n6262, Z => n3408
                           );
   U3530 : MUX2_X1 port map( A => n5733, B => DATAIN(10), S => n6262, Z => 
                           n3409);
   U3531 : MUX2_X1 port map( A => n5732, B => DATAIN(11), S => n6262, Z => 
                           n3410);
   U3532 : MUX2_X1 port map( A => n5731, B => DATAIN(12), S => n6263, Z => 
                           n3411);
   U3533 : MUX2_X1 port map( A => n5730, B => DATAIN(13), S => n6263, Z => 
                           n3412);
   U3534 : MUX2_X1 port map( A => n5729, B => DATAIN(14), S => n6263, Z => 
                           n3413);
   U3535 : MUX2_X1 port map( A => n5728, B => DATAIN(15), S => n6263, Z => 
                           n3414);
   U3536 : MUX2_X1 port map( A => n5727, B => DATAIN(16), S => n6263, Z => 
                           n3415);
   U3537 : MUX2_X1 port map( A => n5726, B => DATAIN(17), S => n6263, Z => 
                           n3416);
   U3538 : MUX2_X1 port map( A => n5725, B => DATAIN(18), S => n6263, Z => 
                           n3417);
   U3539 : MUX2_X1 port map( A => n5724, B => DATAIN(19), S => n6263, Z => 
                           n3418);
   U3540 : MUX2_X1 port map( A => n5723, B => DATAIN(20), S => n6263, Z => 
                           n3419);
   U3541 : MUX2_X1 port map( A => n5722, B => DATAIN(21), S => n6263, Z => 
                           n3420);
   U3542 : MUX2_X1 port map( A => n5721, B => DATAIN(22), S => n6263, Z => 
                           n3421);
   U3543 : MUX2_X1 port map( A => n5720, B => DATAIN(23), S => n6263, Z => 
                           n3422);
   U3544 : MUX2_X1 port map( A => n5719, B => DATAIN(24), S => n6264, Z => 
                           n3423);
   U3545 : MUX2_X1 port map( A => n5718, B => DATAIN(25), S => n6264, Z => 
                           n3424);
   U3546 : MUX2_X1 port map( A => n5717, B => DATAIN(26), S => n6264, Z => 
                           n3425);
   U3547 : MUX2_X1 port map( A => n5716, B => DATAIN(27), S => n6264, Z => 
                           n3426);
   U3548 : MUX2_X1 port map( A => n5715, B => DATAIN(28), S => n6264, Z => 
                           n3427);
   U3549 : MUX2_X1 port map( A => n5714, B => DATAIN(29), S => n6264, Z => 
                           n3428);
   U3550 : MUX2_X1 port map( A => n5713, B => DATAIN(30), S => n6264, Z => 
                           n3429);
   U3551 : MUX2_X1 port map( A => n5712, B => DATAIN(31), S => n6264, Z => 
                           n3430);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity instruction_decomposition is

   port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype : in
         std_logic;  ADD_RS1, ADD_RS2, ADD_WR : out std_logic_vector (4 downto 
         0);  IMM : out std_logic_vector (31 downto 0));

end instruction_decomposition;

architecture SYN_bhv of instruction_decomposition is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal IMM_24_port, IMM_23_port, IMM_22_port, IMM_21_port, IMM_20_port, 
      IMM_19_port, IMM_18_port, IMM_17_port, IMM_16_port, IMM_15_port, 
      IMM_14_port, IMM_13_port, IMM_12_port, IMM_11_port, IMM_10_port, 
      IMM_9_port, IMM_8_port, IMM_7_port, IMM_6_port, IMM_5_port, IMM_4_port, 
      IMM_3_port, IMM_2_port, IMM_1_port, IMM_0_port, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, IMM_31_port, n28, n29, n30, n31, n32, n33, n34, n35, 
      n36, n37, n38, n39, n40, n41, n42, n43, n44, n45 : std_logic;

begin
   IMM <= ( IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, 
      IMM_31_port, IMM_31_port, IMM_24_port, IMM_23_port, IMM_22_port, 
      IMM_21_port, IMM_20_port, IMM_19_port, IMM_18_port, IMM_17_port, 
      IMM_16_port, IMM_15_port, IMM_14_port, IMM_13_port, IMM_12_port, 
      IMM_11_port, IMM_10_port, IMM_9_port, IMM_8_port, IMM_7_port, IMM_6_port,
      IMM_5_port, IMM_4_port, IMM_3_port, IMM_2_port, IMM_1_port, IMM_0_port );
   
   U68 : NAND3_X1 port map( A1 => INST_IN(29), A2 => INST_IN(27), A3 => 
                           INST_IN(31), ZN => n26);
   U69 : NAND3_X1 port map( A1 => INST_IN(26), A2 => Itype, A3 => n27, ZN => 
                           n25);
   U2 : NOR2_X1 port map( A1 => n43, A2 => n37, ZN => ADD_RS2(4));
   U3 : NOR2_X1 port map( A1 => n23, A2 => n42, ZN => ADD_RS1(4));
   U4 : NAND2_X1 port map( A1 => Jtype, A2 => n23, ZN => n19);
   U5 : INV_X1 port map( A => n22, ZN => n44);
   U6 : NOR2_X1 port map( A1 => n23, A2 => n41, ZN => ADD_RS1(3));
   U7 : NOR2_X1 port map( A1 => n43, A2 => n36, ZN => ADD_RS2(3));
   U8 : NOR2_X1 port map( A1 => n23, A2 => n38, ZN => ADD_RS1(0));
   U9 : NOR2_X1 port map( A1 => n43, A2 => n33, ZN => ADD_RS2(0));
   U10 : OAI21_X1 port map( B1 => Jtype, B2 => Itype, A => n45, ZN => n22);
   U11 : NOR2_X1 port map( A1 => Itype, A2 => Rtype, ZN => n23);
   U12 : NOR2_X1 port map( A1 => n23, A2 => n39, ZN => ADD_RS1(1));
   U13 : NOR2_X1 port map( A1 => n43, A2 => n34, ZN => ADD_RS2(1));
   U14 : NOR2_X1 port map( A1 => n23, A2 => n40, ZN => ADD_RS1(2));
   U15 : NOR2_X1 port map( A1 => n43, A2 => n35, ZN => ADD_RS2(2));
   U16 : OR2_X1 port map( A1 => n32, A2 => n21, ZN => n20);
   U17 : INV_X1 port map( A => Rtype, ZN => n45);
   U18 : NAND2_X1 port map( A1 => Itype, A2 => n45, ZN => n21);
   U19 : OAI221_X1 port map( B1 => n21, B2 => n33, C1 => n28, C2 => n45, A => 
                           n19, ZN => ADD_WR(0));
   U20 : OAI221_X1 port map( B1 => n21, B2 => n34, C1 => n29, C2 => n45, A => 
                           n19, ZN => ADD_WR(1));
   U21 : OAI221_X1 port map( B1 => n21, B2 => n35, C1 => n30, C2 => n45, A => 
                           n19, ZN => ADD_WR(2));
   U22 : OAI221_X1 port map( B1 => n21, B2 => n36, C1 => n31, C2 => n45, A => 
                           n19, ZN => ADD_WR(3));
   U23 : OAI221_X1 port map( B1 => n21, B2 => n37, C1 => n32, C2 => n45, A => 
                           n19, ZN => ADD_WR(4));
   U24 : OAI21_X1 port map( B1 => n19, B2 => n42, A => n20, ZN => IMM_31_port);
   U25 : OAI21_X1 port map( B1 => n19, B2 => n33, A => n20, ZN => IMM_16_port);
   U26 : OAI21_X1 port map( B1 => n19, B2 => n34, A => n20, ZN => IMM_17_port);
   U27 : OAI21_X1 port map( B1 => n19, B2 => n35, A => n20, ZN => IMM_18_port);
   U28 : OAI21_X1 port map( B1 => n19, B2 => n36, A => n20, ZN => IMM_19_port);
   U29 : OAI21_X1 port map( B1 => n19, B2 => n37, A => n20, ZN => IMM_20_port);
   U30 : OAI21_X1 port map( B1 => n19, B2 => n38, A => n20, ZN => IMM_21_port);
   U31 : OAI21_X1 port map( B1 => n19, B2 => n39, A => n20, ZN => IMM_22_port);
   U32 : OAI21_X1 port map( B1 => n19, B2 => n40, A => n20, ZN => IMM_23_port);
   U33 : OAI21_X1 port map( B1 => n19, B2 => n41, A => n20, ZN => IMM_24_port);
   U34 : NOR2_X1 port map( A1 => n32, A2 => n22, ZN => IMM_15_port);
   U35 : NOR2_X1 port map( A1 => n22, A2 => n28, ZN => IMM_11_port);
   U36 : NOR2_X1 port map( A1 => n22, A2 => n29, ZN => IMM_12_port);
   U37 : NOR2_X1 port map( A1 => n22, A2 => n30, ZN => IMM_13_port);
   U38 : NOR2_X1 port map( A1 => n22, A2 => n31, ZN => IMM_14_port);
   U39 : INV_X1 port map( A => n24, ZN => n43);
   U40 : OAI21_X1 port map( B1 => n25, B2 => n26, A => n45, ZN => n24);
   U41 : INV_X1 port map( A => INST_IN(16), ZN => n33);
   U42 : INV_X1 port map( A => INST_IN(17), ZN => n34);
   U43 : INV_X1 port map( A => INST_IN(18), ZN => n35);
   U44 : INV_X1 port map( A => INST_IN(19), ZN => n36);
   U45 : INV_X1 port map( A => INST_IN(20), ZN => n37);
   U46 : INV_X1 port map( A => INST_IN(15), ZN => n32);
   U47 : NOR2_X1 port map( A1 => INST_IN(30), A2 => INST_IN(28), ZN => n27);
   U48 : INV_X1 port map( A => INST_IN(21), ZN => n38);
   U49 : INV_X1 port map( A => INST_IN(22), ZN => n39);
   U50 : INV_X1 port map( A => INST_IN(23), ZN => n40);
   U51 : INV_X1 port map( A => INST_IN(24), ZN => n41);
   U52 : INV_X1 port map( A => INST_IN(25), ZN => n42);
   U53 : INV_X1 port map( A => INST_IN(11), ZN => n28);
   U54 : INV_X1 port map( A => INST_IN(12), ZN => n29);
   U55 : INV_X1 port map( A => INST_IN(13), ZN => n30);
   U56 : INV_X1 port map( A => INST_IN(14), ZN => n31);
   U57 : AND2_X1 port map( A1 => INST_IN(0), A2 => n44, ZN => IMM_0_port);
   U58 : AND2_X1 port map( A1 => INST_IN(1), A2 => n44, ZN => IMM_1_port);
   U59 : AND2_X1 port map( A1 => INST_IN(2), A2 => n44, ZN => IMM_2_port);
   U60 : AND2_X1 port map( A1 => INST_IN(3), A2 => n44, ZN => IMM_3_port);
   U61 : AND2_X1 port map( A1 => INST_IN(4), A2 => n44, ZN => IMM_4_port);
   U62 : AND2_X1 port map( A1 => INST_IN(5), A2 => n44, ZN => IMM_5_port);
   U63 : AND2_X1 port map( A1 => INST_IN(6), A2 => n44, ZN => IMM_6_port);
   U64 : AND2_X1 port map( A1 => INST_IN(7), A2 => n44, ZN => IMM_7_port);
   U65 : AND2_X1 port map( A1 => INST_IN(8), A2 => n44, ZN => IMM_8_port);
   U66 : AND2_X1 port map( A1 => INST_IN(9), A2 => n44, ZN => IMM_9_port);
   U67 : AND2_X1 port map( A1 => INST_IN(10), A2 => n44, ZN => IMM_10_port);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity instruction_type is

   port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype : 
         out std_logic);

end instruction_type;

architecture SYN_bhv of instruction_type is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15 : std_logic;

begin
   
   U15 : NAND3_X1 port map( A1 => INST_IN(26), A2 => n14, A3 => INST_IN(30), ZN
                           => n12);
   U1 : NOR2_X1 port map( A1 => n4, A2 => n14, ZN => Jtype);
   U2 : NOR3_X1 port map( A1 => n4, A2 => INST_IN(27), A3 => INST_IN(26), ZN =>
                           Rtype);
   U3 : OAI21_X1 port map( B1 => INST_IN(31), B2 => n5, A => n6, ZN => Itype);
   U4 : NAND4_X1 port map( A1 => INST_IN(31), A2 => INST_IN(26), A3 => n7, A4 
                           => INST_IN(27), ZN => n6);
   U5 : AOI21_X1 port map( B1 => INST_IN(29), B2 => n8, A => n13, ZN => n5);
   U6 : NOR2_X1 port map( A1 => INST_IN(30), A2 => INST_IN(28), ZN => n7);
   U7 : OAI21_X1 port map( B1 => INST_IN(30), B2 => INST_IN(26), A => n12, ZN 
                           => n8);
   U8 : OR4_X1 port map( A1 => INST_IN(28), A2 => INST_IN(29), A3 => 
                           INST_IN(30), A4 => INST_IN(31), ZN => n4);
   U9 : INV_X1 port map( A => INST_IN(27), ZN => n14);
   U10 : INV_X1 port map( A => n9, ZN => n13);
   U11 : OAI21_X1 port map( B1 => n10, B2 => n11, A => INST_IN(28), ZN => n9);
   U12 : AOI21_X1 port map( B1 => INST_IN(26), B2 => INST_IN(30), A => 
                           INST_IN(27), ZN => n10);
   U13 : NOR3_X1 port map( A1 => INST_IN(26), A2 => INST_IN(29), A3 => n15, ZN 
                           => n11);
   U14 : INV_X1 port map( A => INST_IN(30), ZN => n15);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Fetch_DW01_add_3 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Fetch_DW01_add_3;

architecture SYN_cla of Fetch_DW01_add_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, n2, n4, n7, n9, n11, n12, n13, n14, 
      n17, n18, n19, n22, n23, n24, n30, n38, n39, n42, n45, n47, n49, n50, n54
      , n55, n56, n57, n58, n59, n61, n62, n63, n64, n65, n69, n70, n71, n73, 
      n76, n77, n79, n82, n85, n86, n87, n89, n94, n95, n96, n97, n101, n102, 
      n103, n104, n109, n110, n114, n115, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, SUM_2_port, n132, n133, 
      n134, n135, n136, n137, n138, n139 : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U13 : XOR2_X1 port map( A => n7, B => A(9), Z => SUM_9_port);
   U20 : XOR2_X1 port map( A => n12, B => A(8), Z => SUM_8_port);
   U23 : XOR2_X1 port map( A => n13, B => A(7), Z => SUM_7_port);
   U24 : XOR2_X1 port map( A => A(12), B => n14, Z => SUM_12_port);
   U40 : XOR2_X1 port map( A => n54, B => A(31), Z => SUM_31_port);
   U86 : NAND3_X1 port map( A1 => A(4), A2 => A(2), A3 => A(9), ZN => n56);
   U105 : XOR2_X1 port map( A => n64, B => A(18), Z => SUM_18_port);
   U106 : XOR2_X1 port map( A => n58, B => A(16), Z => SUM_16_port);
   U107 : XOR2_X1 port map( A => n77, B => A(6), Z => SUM_6_port);
   U108 : XOR2_X1 port map( A => A(2), B => A(3), Z => SUM_3_port);
   U109 : XOR2_X1 port map( A => n18, B => A(4), Z => SUM_4_port);
   U110 : XOR2_X1 port map( A => n70, B => A(10), Z => SUM_10_port);
   U111 : XOR2_X1 port map( A => n89, B => A(24), Z => SUM_24_port);
   U143 : NAND3_X1 port map( A1 => n49, A2 => n42, A3 => A(29), ZN => n82);
   U144 : NAND3_X1 port map( A1 => A(8), A2 => A(11), A3 => A(12), ZN => n104);
   U2 : NOR2_X1 port map( A1 => n19, A2 => n137, ZN => n23);
   U3 : AND2_X1 port map( A1 => n59, A2 => A(14), ZN => n2);
   U4 : AND2_X1 port map( A1 => n4, A2 => A(26), ZN => n39);
   U5 : OR2_X1 port map( A1 => n87, A2 => n138, ZN => n86);
   U6 : NOR2_X1 port map( A1 => n76, A2 => n132, ZN => n12);
   U7 : NAND2_X1 port map( A1 => n58, A2 => n85, ZN => n71);
   U8 : INV_X1 port map( A => n58, ZN => n134);
   U9 : AND2_X1 port map( A1 => n45, A2 => n85, ZN => n89);
   U10 : AND2_X1 port map( A1 => n45, A2 => n85, ZN => n61);
   U11 : AND2_X1 port map( A1 => n101, A2 => n102, ZN => n58);
   U12 : NAND2_X1 port map( A1 => n114, A2 => n115, ZN => n76);
   U14 : AND2_X1 port map( A1 => n101, A2 => n102, ZN => n45);
   U15 : INV_X1 port map( A => n79, ZN => n132);
   U16 : AND2_X1 port map( A1 => n63, A2 => n94, ZN => n85);
   U17 : NAND2_X1 port map( A1 => n114, A2 => n115, ZN => n30);
   U18 : XNOR2_X1 port map( A => n38, B => n138, ZN => SUM_28_port);
   U19 : NOR2_X1 port map( A1 => n71, A2 => n87, ZN => n38);
   U21 : XNOR2_X1 port map( A => n135, B => n69, ZN => SUM_5_port);
   U22 : NAND4_X1 port map( A1 => A(24), A2 => A(25), A3 => A(26), A4 => A(27),
                           ZN => n87);
   U25 : NAND4_X1 port map( A1 => A(8), A2 => A(11), A3 => A(10), A4 => A(9), 
                           ZN => n19);
   U26 : AND2_X1 port map( A1 => n63, A2 => n94, ZN => n49);
   U27 : NOR2_X1 port map( A1 => n87, A2 => n138, ZN => n42);
   U28 : NOR2_X1 port map( A1 => n55, A2 => n56, ZN => n102);
   U29 : NAND4_X1 port map( A1 => A(3), A2 => A(5), A3 => A(6), A4 => A(7), ZN 
                           => n55);
   U30 : NOR2_X1 port map( A1 => n24, A2 => n96, ZN => n94);
   U31 : NAND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n24);
   U32 : NOR2_X1 port map( A1 => n110, A2 => n137, ZN => n109);
   U33 : NAND4_X1 port map( A1 => A(8), A2 => A(11), A3 => A(10), A4 => A(9), 
                           ZN => n110);
   U34 : NOR2_X1 port map( A1 => n76, A2 => n17, ZN => n59);
   U35 : NAND2_X1 port map( A1 => n18, A2 => A(13), ZN => n17);
   U36 : NOR2_X1 port map( A1 => n103, A2 => n104, ZN => n101);
   U37 : NAND4_X1 port map( A1 => A(14), A2 => A(15), A3 => A(13), A4 => A(10),
                           ZN => n103);
   U38 : NOR2_X1 port map( A1 => n96, A2 => n97, ZN => n57);
   U39 : NAND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n97);
   U41 : AND2_X1 port map( A1 => n79, A2 => A(4), ZN => n69);
   U42 : INV_X1 port map( A => A(5), ZN => n135);
   U43 : INV_X1 port map( A => A(28), ZN => n138);
   U44 : NOR2_X1 port map( A1 => n76, A2 => n22, ZN => n7);
   U45 : NAND2_X1 port map( A1 => n18, A2 => A(8), ZN => n22);
   U46 : NOR2_X1 port map( A1 => n133, A2 => n135, ZN => n77);
   U47 : INV_X1 port map( A => n69, ZN => n133);
   U48 : XNOR2_X1 port map( A => n117, B => A(22), ZN => SUM_22_port);
   U49 : NAND3_X1 port map( A1 => n45, A2 => n9, A3 => A(21), ZN => n117);
   U50 : XNOR2_X1 port map( A => n118, B => A(20), ZN => SUM_20_port);
   U51 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => n118);
   U52 : XNOR2_X1 port map( A => n119, B => A(21), ZN => SUM_21_port);
   U53 : NAND2_X1 port map( A1 => n58, A2 => n9, ZN => n119);
   U54 : AND2_X1 port map( A1 => n69, A2 => n11, ZN => n13);
   U55 : NOR2_X1 port map( A1 => n135, A2 => n136, ZN => n11);
   U56 : INV_X1 port map( A => A(6), ZN => n136);
   U57 : XNOR2_X1 port map( A => n120, B => A(14), ZN => SUM_14_port);
   U58 : NAND2_X1 port map( A1 => n109, A2 => n59, ZN => n120);
   U59 : XNOR2_X1 port map( A => n121, B => A(25), ZN => SUM_25_port);
   U60 : NAND2_X1 port map( A1 => A(24), A2 => n89, ZN => n121);
   U61 : NOR2_X1 port map( A1 => n62, A2 => n19, ZN => n14);
   U62 : OR2_X1 port map( A1 => n30, A2 => n132, ZN => n62);
   U63 : XNOR2_X1 port map( A => A(17), B => n122, ZN => SUM_17_port);
   U64 : NAND2_X1 port map( A1 => n58, A2 => A(16), ZN => n122);
   U65 : NOR3_X1 port map( A1 => n134, A2 => n82, A3 => n139, ZN => n54);
   U66 : INV_X1 port map( A => A(30), ZN => n139);
   U67 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n18);
   U68 : NAND2_X1 port map( A1 => A(19), A2 => A(18), ZN => n96);
   U69 : AND2_X1 port map( A1 => A(7), A2 => A(6), ZN => n115);
   U70 : AND2_X1 port map( A1 => A(5), A2 => A(4), ZN => n114);
   U71 : XOR2_X1 port map( A => n123, B => A(30), Z => SUM_30_port);
   U72 : NOR2_X1 port map( A1 => n134, A2 => n82, ZN => n123);
   U73 : XNOR2_X1 port map( A => n95, B => A(23), ZN => SUM_23_port);
   U74 : NAND2_X1 port map( A1 => n65, A2 => A(22), ZN => n95);
   U75 : AND3_X1 port map( A1 => n9, A2 => n45, A3 => A(21), ZN => n65);
   U76 : XNOR2_X1 port map( A => n124, B => A(13), ZN => SUM_13_port);
   U77 : NAND2_X1 port map( A1 => n23, A2 => n12, ZN => n124);
   U78 : XNOR2_X1 port map( A => n125, B => A(15), ZN => SUM_15_port);
   U79 : NAND2_X1 port map( A1 => n2, A2 => n109, ZN => n125);
   U80 : XNOR2_X1 port map( A => n126, B => A(26), ZN => SUM_26_port);
   U81 : NAND2_X1 port map( A1 => n61, A2 => n4, ZN => n126);
   U82 : XNOR2_X1 port map( A => n127, B => A(11), ZN => SUM_11_port);
   U83 : NAND2_X1 port map( A1 => n70, A2 => A(10), ZN => n127);
   U84 : XNOR2_X1 port map( A => n128, B => A(19), ZN => SUM_19_port);
   U85 : NAND2_X1 port map( A1 => n64, A2 => A(18), ZN => n128);
   U87 : XNOR2_X1 port map( A => n129, B => A(27), ZN => SUM_27_port);
   U88 : NAND2_X1 port map( A1 => n61, A2 => n39, ZN => n129);
   U89 : AND3_X1 port map( A1 => n73, A2 => A(9), A3 => A(8), ZN => n70);
   U90 : NOR2_X1 port map( A1 => n30, A2 => n132, ZN => n73);
   U91 : XNOR2_X1 port map( A => n130, B => A(29), ZN => SUM_29_port);
   U92 : OR2_X1 port map( A1 => n71, A2 => n86, ZN => n130);
   U93 : AND2_X1 port map( A1 => n57, A2 => A(20), ZN => n9);
   U94 : INV_X1 port map( A => A(12), ZN => n137);
   U95 : AND2_X1 port map( A1 => A(2), A2 => A(3), ZN => n79);
   U96 : AND2_X1 port map( A1 => n45, A2 => n50, ZN => n64);
   U97 : AND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n50);
   U98 : AND2_X1 port map( A1 => A(24), A2 => A(25), ZN => n4);
   U99 : AND2_X1 port map( A1 => n47, A2 => A(20), ZN => n63);
   U100 : AND3_X1 port map( A1 => A(22), A2 => A(21), A3 => A(23), ZN => n47);
   U101 : INV_X1 port map( A => A(2), ZN => SUM_2_port);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HazardDetection is

   port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : in std_logic_vector (4
         downto 0);  DRAM_R : in std_logic;  INS_IN, PC_IN : in 
         std_logic_vector (31 downto 0);  Bubble : out std_logic;  HDU_INS_OUT,
         HDU_PC_OUT, HDU_NPC_OUT : out std_logic_vector (31 downto 0));

end HazardDetection;

architecture SYN_arch of HazardDetection is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component HazardDetection_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n9, n10, n12, n13, n14, n15, n16, n17, n18, 
      n19, n_1170 : std_logic;

begin
   HDU_INS_OUT <= ( INS_IN(31), INS_IN(30), INS_IN(29), INS_IN(28), INS_IN(27),
      INS_IN(26), INS_IN(25), INS_IN(24), INS_IN(23), INS_IN(22), INS_IN(21), 
      INS_IN(20), INS_IN(19), INS_IN(18), INS_IN(17), INS_IN(16), INS_IN(15), 
      INS_IN(14), INS_IN(13), INS_IN(12), INS_IN(11), INS_IN(10), INS_IN(9), 
      INS_IN(8), INS_IN(7), INS_IN(6), INS_IN(5), INS_IN(4), INS_IN(3), 
      INS_IN(2), INS_IN(1), INS_IN(0) );
   HDU_NPC_OUT <= ( PC_IN(31), PC_IN(30), PC_IN(29), PC_IN(28), PC_IN(27), 
      PC_IN(26), PC_IN(25), PC_IN(24), PC_IN(23), PC_IN(22), PC_IN(21), 
      PC_IN(20), PC_IN(19), PC_IN(18), PC_IN(17), PC_IN(16), PC_IN(15), 
      PC_IN(14), PC_IN(13), PC_IN(12), PC_IN(11), PC_IN(10), PC_IN(9), PC_IN(8)
      , PC_IN(7), PC_IN(6), PC_IN(5), PC_IN(4), PC_IN(3), PC_IN(2), PC_IN(1), 
      PC_IN(0) );
   
   n1 <= '0';
   n2 <= '0';
   n3 <= '1';
   U16 : OAI33_X1 port map( A1 => n5, A2 => n6, A3 => n9, B1 => n10, B2 => n12,
                           B3 => n13, ZN => n4);
   U17 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RS2(4), Z => n13);
   U18 : XOR2_X1 port map( A => ADD_WR(2), B => ADD_RS2(2), Z => n12);
   U19 : NAND3_X1 port map( A1 => n14, A2 => n15, A3 => n16, ZN => n10);
   U20 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RS1(4), Z => n9);
   U21 : XOR2_X1 port map( A => ADD_WR(2), B => ADD_RS1(2), Z => n6);
   U22 : NAND3_X1 port map( A1 => n17, A2 => n18, A3 => n19, ZN => n5);
   sub_25 : HazardDetection_DW01_sub_0 port map( A(31) => PC_IN(31), A(30) => 
                           PC_IN(30), A(29) => PC_IN(29), A(28) => PC_IN(28), 
                           A(27) => PC_IN(27), A(26) => PC_IN(26), A(25) => 
                           PC_IN(25), A(24) => PC_IN(24), A(23) => PC_IN(23), 
                           A(22) => PC_IN(22), A(21) => PC_IN(21), A(20) => 
                           PC_IN(20), A(19) => PC_IN(19), A(18) => PC_IN(18), 
                           A(17) => PC_IN(17), A(16) => PC_IN(16), A(15) => 
                           PC_IN(15), A(14) => PC_IN(14), A(13) => PC_IN(13), 
                           A(12) => PC_IN(12), A(11) => PC_IN(11), A(10) => 
                           PC_IN(10), A(9) => PC_IN(9), A(8) => PC_IN(8), A(7) 
                           => PC_IN(7), A(6) => PC_IN(6), A(5) => PC_IN(5), 
                           A(4) => PC_IN(4), A(3) => PC_IN(3), A(2) => PC_IN(2)
                           , A(1) => PC_IN(1), A(0) => PC_IN(0), B(31) => n2, 
                           B(30) => n2, B(29) => n2, B(28) => n2, B(27) => n2, 
                           B(26) => n2, B(25) => n2, B(24) => n2, B(23) => n2, 
                           B(22) => n2, B(21) => n2, B(20) => n2, B(19) => n2, 
                           B(18) => n2, B(17) => n2, B(16) => n2, B(15) => n2, 
                           B(14) => n2, B(13) => n2, B(12) => n2, B(11) => n2, 
                           B(10) => n2, B(9) => n2, B(8) => n2, B(7) => n2, 
                           B(6) => n2, B(5) => n2, B(4) => n2, B(3) => n2, B(2)
                           => n3, B(1) => n2, B(0) => n2, CI => n1, DIFF(31) =>
                           HDU_PC_OUT(31), DIFF(30) => HDU_PC_OUT(30), DIFF(29)
                           => HDU_PC_OUT(29), DIFF(28) => HDU_PC_OUT(28), 
                           DIFF(27) => HDU_PC_OUT(27), DIFF(26) => 
                           HDU_PC_OUT(26), DIFF(25) => HDU_PC_OUT(25), DIFF(24)
                           => HDU_PC_OUT(24), DIFF(23) => HDU_PC_OUT(23), 
                           DIFF(22) => HDU_PC_OUT(22), DIFF(21) => 
                           HDU_PC_OUT(21), DIFF(20) => HDU_PC_OUT(20), DIFF(19)
                           => HDU_PC_OUT(19), DIFF(18) => HDU_PC_OUT(18), 
                           DIFF(17) => HDU_PC_OUT(17), DIFF(16) => 
                           HDU_PC_OUT(16), DIFF(15) => HDU_PC_OUT(15), DIFF(14)
                           => HDU_PC_OUT(14), DIFF(13) => HDU_PC_OUT(13), 
                           DIFF(12) => HDU_PC_OUT(12), DIFF(11) => 
                           HDU_PC_OUT(11), DIFF(10) => HDU_PC_OUT(10), DIFF(9) 
                           => HDU_PC_OUT(9), DIFF(8) => HDU_PC_OUT(8), DIFF(7) 
                           => HDU_PC_OUT(7), DIFF(6) => HDU_PC_OUT(6), DIFF(5) 
                           => HDU_PC_OUT(5), DIFF(4) => HDU_PC_OUT(4), DIFF(3) 
                           => HDU_PC_OUT(3), DIFF(2) => HDU_PC_OUT(2), DIFF(1) 
                           => HDU_PC_OUT(1), DIFF(0) => HDU_PC_OUT(0), CO => 
                           n_1170);
   U3 : AND3_X1 port map( A1 => DRAM_R, A2 => n4, A3 => RST, ZN => Bubble);
   U7 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS1(3), ZN => n17);
   U8 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS2(3), ZN => n14);
   U9 : XNOR2_X1 port map( A => ADD_WR(0), B => ADD_RS1(0), ZN => n18);
   U10 : XNOR2_X1 port map( A => ADD_WR(0), B => ADD_RS2(0), ZN => n15);
   U11 : XNOR2_X1 port map( A => ADD_WR(1), B => ADD_RS1(1), ZN => n19);
   U12 : XNOR2_X1 port map( A => ADD_WR(1), B => ADD_RS2(1), ZN => n16);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Writeback is

   port( WB_MUX_SEL : in std_logic;  DATA_IN, ALU_RES_IN : in std_logic_vector 
         (31 downto 0);  ADD_WR_IN : in std_logic_vector (4 downto 0);  
         DATA_OUT : out std_logic_vector (31 downto 0);  ADD_WR_OUT : out 
         std_logic_vector (4 downto 0));

end Writeback;

architecture SYN_struct of Writeback is

   component mux21_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;

begin
   ADD_WR_OUT <= ( ADD_WR_IN(4), ADD_WR_IN(3), ADD_WR_IN(2), ADD_WR_IN(1), 
      ADD_WR_IN(0) );
   
   WBmux : mux21_NBIT32_2 port map( A(31) => DATA_IN(31), A(30) => DATA_IN(30),
                           A(29) => DATA_IN(29), A(28) => DATA_IN(28), A(27) =>
                           DATA_IN(27), A(26) => DATA_IN(26), A(25) => 
                           DATA_IN(25), A(24) => DATA_IN(24), A(23) => 
                           DATA_IN(23), A(22) => DATA_IN(22), A(21) => 
                           DATA_IN(21), A(20) => DATA_IN(20), A(19) => 
                           DATA_IN(19), A(18) => DATA_IN(18), A(17) => 
                           DATA_IN(17), A(16) => DATA_IN(16), A(15) => 
                           DATA_IN(15), A(14) => DATA_IN(14), A(13) => 
                           DATA_IN(13), A(12) => DATA_IN(12), A(11) => 
                           DATA_IN(11), A(10) => DATA_IN(10), A(9) => 
                           DATA_IN(9), A(8) => DATA_IN(8), A(7) => DATA_IN(7), 
                           A(6) => DATA_IN(6), A(5) => DATA_IN(5), A(4) => 
                           DATA_IN(4), A(3) => DATA_IN(3), A(2) => DATA_IN(2), 
                           A(1) => DATA_IN(1), A(0) => DATA_IN(0), B(31) => 
                           ALU_RES_IN(31), B(30) => ALU_RES_IN(30), B(29) => 
                           ALU_RES_IN(29), B(28) => ALU_RES_IN(28), B(27) => 
                           ALU_RES_IN(27), B(26) => ALU_RES_IN(26), B(25) => 
                           ALU_RES_IN(25), B(24) => ALU_RES_IN(24), B(23) => 
                           ALU_RES_IN(23), B(22) => ALU_RES_IN(22), B(21) => 
                           ALU_RES_IN(21), B(20) => ALU_RES_IN(20), B(19) => 
                           ALU_RES_IN(19), B(18) => ALU_RES_IN(18), B(17) => 
                           ALU_RES_IN(17), B(16) => ALU_RES_IN(16), B(15) => 
                           ALU_RES_IN(15), B(14) => ALU_RES_IN(14), B(13) => 
                           ALU_RES_IN(13), B(12) => ALU_RES_IN(12), B(11) => 
                           ALU_RES_IN(11), B(10) => ALU_RES_IN(10), B(9) => 
                           ALU_RES_IN(9), B(8) => ALU_RES_IN(8), B(7) => 
                           ALU_RES_IN(7), B(6) => ALU_RES_IN(6), B(5) => 
                           ALU_RES_IN(5), B(4) => ALU_RES_IN(4), B(3) => 
                           ALU_RES_IN(3), B(2) => ALU_RES_IN(2), B(1) => 
                           ALU_RES_IN(1), B(0) => ALU_RES_IN(0), S => 
                           WB_MUX_SEL, Z(31) => DATA_OUT(31), Z(30) => 
                           DATA_OUT(30), Z(29) => DATA_OUT(29), Z(28) => 
                           DATA_OUT(28), Z(27) => DATA_OUT(27), Z(26) => 
                           DATA_OUT(26), Z(25) => DATA_OUT(25), Z(24) => 
                           DATA_OUT(24), Z(23) => DATA_OUT(23), Z(22) => 
                           DATA_OUT(22), Z(21) => DATA_OUT(21), Z(20) => 
                           DATA_OUT(20), Z(19) => DATA_OUT(19), Z(18) => 
                           DATA_OUT(18), Z(17) => DATA_OUT(17), Z(16) => 
                           DATA_OUT(16), Z(15) => DATA_OUT(15), Z(14) => 
                           DATA_OUT(14), Z(13) => DATA_OUT(13), Z(12) => 
                           DATA_OUT(12), Z(11) => DATA_OUT(11), Z(10) => 
                           DATA_OUT(10), Z(9) => DATA_OUT(9), Z(8) => 
                           DATA_OUT(8), Z(7) => DATA_OUT(7), Z(6) => 
                           DATA_OUT(6), Z(5) => DATA_OUT(5), Z(4) => 
                           DATA_OUT(4), Z(3) => DATA_OUT(3), Z(2) => 
                           DATA_OUT(2), Z(1) => DATA_OUT(1), Z(0) => 
                           DATA_OUT(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Memory is

   port( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, DRAM_EN_IN : in std_logic; 
         PC_SEL : in std_logic_vector (1 downto 0);  NPC_IN, NPC_ABS, NPC_REL, 
         ALU_RES_IN, B_IN : in std_logic_vector (31 downto 0);  ADD_WR_IN : in 
         std_logic_vector (4 downto 0);  DRAM_DATA_IN : in std_logic_vector (31
         downto 0);  PC_OUT : out std_logic_vector (31 downto 0);  DRAM_EN_OUT,
         DRAM_R_OUT, DRAM_W_OUT : out std_logic;  DRAM_ADDR_OUT, DRAM_DATA_OUT,
         DATA_OUT, ALU_RES_OUT, OP_MEM : out std_logic_vector (31 downto 0);  
         ADD_WR_MEM, ADD_WR_OUT : out std_logic_vector (4 downto 0));

end Memory;

architecture SYN_struct of Memory is

   component mux41_NBIT32_2
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component regn_N32_1
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N5_1
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N32_2
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   signal n1 : std_logic;

begin
   DRAM_EN_OUT <= DRAM_EN_IN;
   DRAM_R_OUT <= DRAM_R_IN;
   DRAM_W_OUT <= DRAM_W_IN;
   DRAM_ADDR_OUT <= ( ALU_RES_IN(31), ALU_RES_IN(30), ALU_RES_IN(29), 
      ALU_RES_IN(28), ALU_RES_IN(27), ALU_RES_IN(26), ALU_RES_IN(25), 
      ALU_RES_IN(24), ALU_RES_IN(23), ALU_RES_IN(22), ALU_RES_IN(21), 
      ALU_RES_IN(20), ALU_RES_IN(19), ALU_RES_IN(18), ALU_RES_IN(17), 
      ALU_RES_IN(16), ALU_RES_IN(15), ALU_RES_IN(14), ALU_RES_IN(13), 
      ALU_RES_IN(12), ALU_RES_IN(11), ALU_RES_IN(10), ALU_RES_IN(9), 
      ALU_RES_IN(8), ALU_RES_IN(7), ALU_RES_IN(6), ALU_RES_IN(5), ALU_RES_IN(4)
      , ALU_RES_IN(3), ALU_RES_IN(2), ALU_RES_IN(1), ALU_RES_IN(0) );
   DRAM_DATA_OUT <= ( B_IN(31), B_IN(30), B_IN(29), B_IN(28), B_IN(27), 
      B_IN(26), B_IN(25), B_IN(24), B_IN(23), B_IN(22), B_IN(21), B_IN(20), 
      B_IN(19), B_IN(18), B_IN(17), B_IN(16), B_IN(15), B_IN(14), B_IN(13), 
      B_IN(12), B_IN(11), B_IN(10), B_IN(9), B_IN(8), B_IN(7), B_IN(6), B_IN(5)
      , B_IN(4), B_IN(3), B_IN(2), B_IN(1), B_IN(0) );
   OP_MEM <= ( ALU_RES_IN(31), ALU_RES_IN(30), ALU_RES_IN(29), ALU_RES_IN(28), 
      ALU_RES_IN(27), ALU_RES_IN(26), ALU_RES_IN(25), ALU_RES_IN(24), 
      ALU_RES_IN(23), ALU_RES_IN(22), ALU_RES_IN(21), ALU_RES_IN(20), 
      ALU_RES_IN(19), ALU_RES_IN(18), ALU_RES_IN(17), ALU_RES_IN(16), 
      ALU_RES_IN(15), ALU_RES_IN(14), ALU_RES_IN(13), ALU_RES_IN(12), 
      ALU_RES_IN(11), ALU_RES_IN(10), ALU_RES_IN(9), ALU_RES_IN(8), 
      ALU_RES_IN(7), ALU_RES_IN(6), ALU_RES_IN(5), ALU_RES_IN(4), ALU_RES_IN(3)
      , ALU_RES_IN(2), ALU_RES_IN(1), ALU_RES_IN(0) );
   ADD_WR_MEM <= ( ADD_WR_IN(4), ADD_WR_IN(3), ADD_WR_IN(2), ADD_WR_IN(1), 
      ADD_WR_IN(0) );
   
   LMD : regn_N32_2 port map( DIN(31) => DRAM_DATA_IN(31), DIN(30) => 
                           DRAM_DATA_IN(30), DIN(29) => DRAM_DATA_IN(29), 
                           DIN(28) => DRAM_DATA_IN(28), DIN(27) => 
                           DRAM_DATA_IN(27), DIN(26) => DRAM_DATA_IN(26), 
                           DIN(25) => DRAM_DATA_IN(25), DIN(24) => 
                           DRAM_DATA_IN(24), DIN(23) => DRAM_DATA_IN(23), 
                           DIN(22) => DRAM_DATA_IN(22), DIN(21) => 
                           DRAM_DATA_IN(21), DIN(20) => DRAM_DATA_IN(20), 
                           DIN(19) => DRAM_DATA_IN(19), DIN(18) => 
                           DRAM_DATA_IN(18), DIN(17) => DRAM_DATA_IN(17), 
                           DIN(16) => DRAM_DATA_IN(16), DIN(15) => 
                           DRAM_DATA_IN(15), DIN(14) => DRAM_DATA_IN(14), 
                           DIN(13) => DRAM_DATA_IN(13), DIN(12) => 
                           DRAM_DATA_IN(12), DIN(11) => DRAM_DATA_IN(11), 
                           DIN(10) => DRAM_DATA_IN(10), DIN(9) => 
                           DRAM_DATA_IN(9), DIN(8) => DRAM_DATA_IN(8), DIN(7) 
                           => DRAM_DATA_IN(7), DIN(6) => DRAM_DATA_IN(6), 
                           DIN(5) => DRAM_DATA_IN(5), DIN(4) => DRAM_DATA_IN(4)
                           , DIN(3) => DRAM_DATA_IN(3), DIN(2) => 
                           DRAM_DATA_IN(2), DIN(1) => DRAM_DATA_IN(1), DIN(0) 
                           => DRAM_DATA_IN(0), CLK => CLK, EN => MEM_EN_IN, RST
                           => RST, DOUT(31) => DATA_OUT(31), DOUT(30) => 
                           DATA_OUT(30), DOUT(29) => DATA_OUT(29), DOUT(28) => 
                           DATA_OUT(28), DOUT(27) => DATA_OUT(27), DOUT(26) => 
                           DATA_OUT(26), DOUT(25) => DATA_OUT(25), DOUT(24) => 
                           DATA_OUT(24), DOUT(23) => DATA_OUT(23), DOUT(22) => 
                           DATA_OUT(22), DOUT(21) => DATA_OUT(21), DOUT(20) => 
                           DATA_OUT(20), DOUT(19) => DATA_OUT(19), DOUT(18) => 
                           DATA_OUT(18), DOUT(17) => DATA_OUT(17), DOUT(16) => 
                           DATA_OUT(16), DOUT(15) => DATA_OUT(15), DOUT(14) => 
                           DATA_OUT(14), DOUT(13) => DATA_OUT(13), DOUT(12) => 
                           DATA_OUT(12), DOUT(11) => DATA_OUT(11), DOUT(10) => 
                           DATA_OUT(10), DOUT(9) => DATA_OUT(9), DOUT(8) => 
                           DATA_OUT(8), DOUT(7) => DATA_OUT(7), DOUT(6) => 
                           DATA_OUT(6), DOUT(5) => DATA_OUT(5), DOUT(4) => 
                           DATA_OUT(4), DOUT(3) => DATA_OUT(3), DOUT(2) => 
                           DATA_OUT(2), DOUT(1) => DATA_OUT(1), DOUT(0) => 
                           DATA_OUT(0));
   reg0 : regn_N5_1 port map( DIN(4) => ADD_WR_IN(4), DIN(3) => ADD_WR_IN(3), 
                           DIN(2) => ADD_WR_IN(2), DIN(1) => ADD_WR_IN(1), 
                           DIN(0) => ADD_WR_IN(0), CLK => CLK, EN => MEM_EN_IN,
                           RST => RST, DOUT(4) => ADD_WR_OUT(4), DOUT(3) => 
                           ADD_WR_OUT(3), DOUT(2) => ADD_WR_OUT(2), DOUT(1) => 
                           ADD_WR_OUT(1), DOUT(0) => ADD_WR_OUT(0));
   reg1 : regn_N32_1 port map( DIN(31) => ALU_RES_IN(31), DIN(30) => 
                           ALU_RES_IN(30), DIN(29) => ALU_RES_IN(29), DIN(28) 
                           => ALU_RES_IN(28), DIN(27) => ALU_RES_IN(27), 
                           DIN(26) => ALU_RES_IN(26), DIN(25) => ALU_RES_IN(25)
                           , DIN(24) => ALU_RES_IN(24), DIN(23) => 
                           ALU_RES_IN(23), DIN(22) => ALU_RES_IN(22), DIN(21) 
                           => ALU_RES_IN(21), DIN(20) => ALU_RES_IN(20), 
                           DIN(19) => ALU_RES_IN(19), DIN(18) => ALU_RES_IN(18)
                           , DIN(17) => ALU_RES_IN(17), DIN(16) => 
                           ALU_RES_IN(16), DIN(15) => ALU_RES_IN(15), DIN(14) 
                           => ALU_RES_IN(14), DIN(13) => ALU_RES_IN(13), 
                           DIN(12) => ALU_RES_IN(12), DIN(11) => ALU_RES_IN(11)
                           , DIN(10) => ALU_RES_IN(10), DIN(9) => ALU_RES_IN(9)
                           , DIN(8) => ALU_RES_IN(8), DIN(7) => ALU_RES_IN(7), 
                           DIN(6) => ALU_RES_IN(6), DIN(5) => ALU_RES_IN(5), 
                           DIN(4) => ALU_RES_IN(4), DIN(3) => ALU_RES_IN(3), 
                           DIN(2) => ALU_RES_IN(2), DIN(1) => ALU_RES_IN(1), 
                           DIN(0) => ALU_RES_IN(0), CLK => CLK, EN => MEM_EN_IN
                           , RST => RST, DOUT(31) => ALU_RES_OUT(31), DOUT(30) 
                           => ALU_RES_OUT(30), DOUT(29) => ALU_RES_OUT(29), 
                           DOUT(28) => ALU_RES_OUT(28), DOUT(27) => 
                           ALU_RES_OUT(27), DOUT(26) => ALU_RES_OUT(26), 
                           DOUT(25) => ALU_RES_OUT(25), DOUT(24) => 
                           ALU_RES_OUT(24), DOUT(23) => ALU_RES_OUT(23), 
                           DOUT(22) => ALU_RES_OUT(22), DOUT(21) => 
                           ALU_RES_OUT(21), DOUT(20) => ALU_RES_OUT(20), 
                           DOUT(19) => ALU_RES_OUT(19), DOUT(18) => 
                           ALU_RES_OUT(18), DOUT(17) => ALU_RES_OUT(17), 
                           DOUT(16) => ALU_RES_OUT(16), DOUT(15) => 
                           ALU_RES_OUT(15), DOUT(14) => ALU_RES_OUT(14), 
                           DOUT(13) => ALU_RES_OUT(13), DOUT(12) => 
                           ALU_RES_OUT(12), DOUT(11) => ALU_RES_OUT(11), 
                           DOUT(10) => ALU_RES_OUT(10), DOUT(9) => 
                           ALU_RES_OUT(9), DOUT(8) => ALU_RES_OUT(8), DOUT(7) 
                           => ALU_RES_OUT(7), DOUT(6) => ALU_RES_OUT(6), 
                           DOUT(5) => ALU_RES_OUT(5), DOUT(4) => ALU_RES_OUT(4)
                           , DOUT(3) => ALU_RES_OUT(3), DOUT(2) => 
                           ALU_RES_OUT(2), DOUT(1) => ALU_RES_OUT(1), DOUT(0) 
                           => ALU_RES_OUT(0));
   PCsel : mux41_NBIT32_2 port map( A(31) => NPC_IN(31), A(30) => NPC_IN(30), 
                           A(29) => NPC_IN(29), A(28) => NPC_IN(28), A(27) => 
                           NPC_IN(27), A(26) => NPC_IN(26), A(25) => NPC_IN(25)
                           , A(24) => NPC_IN(24), A(23) => NPC_IN(23), A(22) =>
                           NPC_IN(22), A(21) => NPC_IN(21), A(20) => NPC_IN(20)
                           , A(19) => NPC_IN(19), A(18) => NPC_IN(18), A(17) =>
                           NPC_IN(17), A(16) => NPC_IN(16), A(15) => NPC_IN(15)
                           , A(14) => NPC_IN(14), A(13) => NPC_IN(13), A(12) =>
                           NPC_IN(12), A(11) => NPC_IN(11), A(10) => NPC_IN(10)
                           , A(9) => NPC_IN(9), A(8) => NPC_IN(8), A(7) => 
                           NPC_IN(7), A(6) => NPC_IN(6), A(5) => NPC_IN(5), 
                           A(4) => NPC_IN(4), A(3) => NPC_IN(3), A(2) => 
                           NPC_IN(2), A(1) => NPC_IN(1), A(0) => NPC_IN(0), 
                           B(31) => NPC_REL(31), B(30) => NPC_REL(30), B(29) =>
                           NPC_REL(29), B(28) => NPC_REL(28), B(27) => 
                           NPC_REL(27), B(26) => NPC_REL(26), B(25) => 
                           NPC_REL(25), B(24) => NPC_REL(24), B(23) => 
                           NPC_REL(23), B(22) => NPC_REL(22), B(21) => 
                           NPC_REL(21), B(20) => NPC_REL(20), B(19) => 
                           NPC_REL(19), B(18) => NPC_REL(18), B(17) => 
                           NPC_REL(17), B(16) => NPC_REL(16), B(15) => 
                           NPC_REL(15), B(14) => NPC_REL(14), B(13) => 
                           NPC_REL(13), B(12) => NPC_REL(12), B(11) => 
                           NPC_REL(11), B(10) => NPC_REL(10), B(9) => 
                           NPC_REL(9), B(8) => NPC_REL(8), B(7) => NPC_REL(7), 
                           B(6) => NPC_REL(6), B(5) => NPC_REL(5), B(4) => 
                           NPC_REL(4), B(3) => NPC_REL(3), B(2) => NPC_REL(2), 
                           B(1) => NPC_REL(1), B(0) => NPC_REL(0), C(31) => 
                           NPC_ABS(31), C(30) => NPC_ABS(30), C(29) => 
                           NPC_ABS(29), C(28) => NPC_ABS(28), C(27) => 
                           NPC_ABS(27), C(26) => NPC_ABS(26), C(25) => 
                           NPC_ABS(25), C(24) => NPC_ABS(24), C(23) => 
                           NPC_ABS(23), C(22) => NPC_ABS(22), C(21) => 
                           NPC_ABS(21), C(20) => NPC_ABS(20), C(19) => 
                           NPC_ABS(19), C(18) => NPC_ABS(18), C(17) => 
                           NPC_ABS(17), C(16) => NPC_ABS(16), C(15) => 
                           NPC_ABS(15), C(14) => NPC_ABS(14), C(13) => 
                           NPC_ABS(13), C(12) => NPC_ABS(12), C(11) => 
                           NPC_ABS(11), C(10) => NPC_ABS(10), C(9) => 
                           NPC_ABS(9), C(8) => NPC_ABS(8), C(7) => NPC_ABS(7), 
                           C(6) => NPC_ABS(6), C(5) => NPC_ABS(5), C(4) => 
                           NPC_ABS(4), C(3) => NPC_ABS(3), C(2) => NPC_ABS(2), 
                           C(1) => NPC_ABS(1), C(0) => NPC_ABS(0), D(31) => n1,
                           D(30) => n1, D(29) => n1, D(28) => n1, D(27) => n1, 
                           D(26) => n1, D(25) => n1, D(24) => n1, D(23) => n1, 
                           D(22) => n1, D(21) => n1, D(20) => n1, D(19) => n1, 
                           D(18) => n1, D(17) => n1, D(16) => n1, D(15) => n1, 
                           D(14) => n1, D(13) => n1, D(12) => n1, D(11) => n1, 
                           D(10) => n1, D(9) => n1, D(8) => n1, D(7) => n1, 
                           D(6) => n1, D(5) => n1, D(4) => n1, D(3) => n1, D(2)
                           => n1, D(1) => n1, D(0) => n1, S(1) => PC_SEL(1), 
                           S(0) => PC_SEL(0), Z(31) => PC_OUT(31), Z(30) => 
                           PC_OUT(30), Z(29) => PC_OUT(29), Z(28) => PC_OUT(28)
                           , Z(27) => PC_OUT(27), Z(26) => PC_OUT(26), Z(25) =>
                           PC_OUT(25), Z(24) => PC_OUT(24), Z(23) => PC_OUT(23)
                           , Z(22) => PC_OUT(22), Z(21) => PC_OUT(21), Z(20) =>
                           PC_OUT(20), Z(19) => PC_OUT(19), Z(18) => PC_OUT(18)
                           , Z(17) => PC_OUT(17), Z(16) => PC_OUT(16), Z(15) =>
                           PC_OUT(15), Z(14) => PC_OUT(14), Z(13) => PC_OUT(13)
                           , Z(12) => PC_OUT(12), Z(11) => PC_OUT(11), Z(10) =>
                           PC_OUT(10), Z(9) => PC_OUT(9), Z(8) => PC_OUT(8), 
                           Z(7) => PC_OUT(7), Z(6) => PC_OUT(6), Z(5) => 
                           PC_OUT(5), Z(4) => PC_OUT(4), Z(3) => PC_OUT(3), 
                           Z(2) => PC_OUT(2), Z(1) => PC_OUT(1), Z(0) => 
                           PC_OUT(0));
   n1 <= '0';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute is

   port( CLK, RST, MUX_A_SEL : in std_logic;  MUX_B_SEL : in std_logic_vector 
         (1 downto 0);  ALU_OPC : in std_logic_vector (0 to 3);  ALU_OUTREG_EN 
         : in std_logic;  JUMP_TYPE : in std_logic_vector (1 downto 0);  PC_IN,
         A_IN, B_IN, IMM_IN : in std_logic_vector (31 downto 0);  ADD_WR_IN, 
         ADD_RS1_IN, ADD_RS2_IN, ADD_WR_MEM, ADD_WR_WB : in std_logic_vector (4
         downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;  OP_MEM, OP_WB : in 
         std_logic_vector (31 downto 0);  PC_SEL : out std_logic_vector (1 
         downto 0);  ZERO_FLAG : out std_logic;  NPC_ABS, NPC_REL, ALU_RES, 
         B_OUT : out std_logic_vector (31 downto 0);  ADD_WR_OUT : out 
         std_logic_vector (4 downto 0));

end Execute;

architecture SYN_struct of Execute is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component Execute_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component Execute_DW01_add_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component regn_N32_3
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_4
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N5_2
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N32_5
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_6
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component ALU_NBIT32
      port( OP1, OP2 : in std_logic_vector (31 downto 0);  ALU_OPC : in 
            std_logic_vector (0 to 3);  ALU_RES : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux41_NBIT32_3
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux21_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux41_NBIT32_4
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux41_NBIT32_0
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component FWD_Unit
      port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB : in 
            std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;
            FWDA, FWDB : out std_logic_vector (1 downto 0));
   end component;
   
   component regn_N2
      port( DIN : in std_logic_vector (1 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (1 downto 0));
   end component;
   
   component ff_1
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Branch_Cond_Unit_NBIT32
      port( RST : in std_logic;  A : in std_logic_vector (31 downto 0);  
            ALU_OPC : in std_logic_vector (0 to 3);  JUMP_TYPE : in 
            std_logic_vector (1 downto 0);  PC_SEL : out std_logic_vector (1 
            downto 0);  ZERO : out std_logic);
   end component;
   
   signal ZERO_FLAG_port, sig_RST, sig_NPC_ABS_31_port, sig_NPC_ABS_30_port, 
      sig_NPC_ABS_29_port, sig_NPC_ABS_28_port, sig_NPC_ABS_27_port, 
      sig_NPC_ABS_26_port, sig_NPC_ABS_25_port, sig_NPC_ABS_24_port, 
      sig_NPC_ABS_23_port, sig_NPC_ABS_22_port, sig_NPC_ABS_21_port, 
      sig_NPC_ABS_20_port, sig_NPC_ABS_19_port, sig_NPC_ABS_18_port, 
      sig_NPC_ABS_17_port, sig_NPC_ABS_16_port, sig_NPC_ABS_15_port, 
      sig_NPC_ABS_14_port, sig_NPC_ABS_13_port, sig_NPC_ABS_12_port, 
      sig_NPC_ABS_11_port, sig_NPC_ABS_10_port, sig_NPC_ABS_9_port, 
      sig_NPC_ABS_8_port, sig_NPC_ABS_7_port, sig_NPC_ABS_6_port, 
      sig_NPC_ABS_5_port, sig_NPC_ABS_4_port, sig_NPC_ABS_3_port, 
      sig_NPC_ABS_2_port, sig_NPC_ABS_1_port, sig_NPC_ABS_0_port, 
      sig_NPC_REL_31_port, sig_NPC_REL_30_port, sig_NPC_REL_29_port, 
      sig_NPC_REL_28_port, sig_NPC_REL_27_port, sig_NPC_REL_26_port, 
      sig_NPC_REL_25_port, sig_NPC_REL_24_port, sig_NPC_REL_23_port, 
      sig_NPC_REL_22_port, sig_NPC_REL_21_port, sig_NPC_REL_20_port, 
      sig_NPC_REL_19_port, sig_NPC_REL_18_port, sig_NPC_REL_17_port, 
      sig_NPC_REL_16_port, sig_NPC_REL_15_port, sig_NPC_REL_14_port, 
      sig_NPC_REL_13_port, sig_NPC_REL_12_port, sig_NPC_REL_11_port, 
      sig_NPC_REL_10_port, sig_NPC_REL_9_port, sig_NPC_REL_8_port, 
      sig_NPC_REL_7_port, sig_NPC_REL_6_port, sig_NPC_REL_5_port, 
      sig_NPC_REL_4_port, sig_NPC_REL_3_port, sig_NPC_REL_2_port, 
      sig_NPC_REL_1_port, sig_NPC_REL_0_port, sig_PC_SEL_1_port, 
      sig_PC_SEL_0_port, sig_ZERO_FLAG, FWDA_1_port, FWDA_0_port, FWDB_1_port, 
      FWDB_0_port, sig_OP1_31_port, sig_OP1_30_port, sig_OP1_29_port, 
      sig_OP1_28_port, sig_OP1_27_port, sig_OP1_26_port, sig_OP1_25_port, 
      sig_OP1_24_port, sig_OP1_23_port, sig_OP1_22_port, sig_OP1_21_port, 
      sig_OP1_20_port, sig_OP1_19_port, sig_OP1_18_port, sig_OP1_17_port, 
      sig_OP1_16_port, sig_OP1_15_port, sig_OP1_14_port, sig_OP1_13_port, 
      sig_OP1_12_port, sig_OP1_11_port, sig_OP1_10_port, sig_OP1_9_port, 
      sig_OP1_8_port, sig_OP1_7_port, sig_OP1_6_port, sig_OP1_5_port, 
      sig_OP1_4_port, sig_OP1_3_port, sig_OP1_2_port, sig_OP1_1_port, 
      sig_OP1_0_port, sig_OP2_31_port, sig_OP2_30_port, sig_OP2_29_port, 
      sig_OP2_28_port, sig_OP2_27_port, sig_OP2_26_port, sig_OP2_25_port, 
      sig_OP2_24_port, sig_OP2_23_port, sig_OP2_22_port, sig_OP2_21_port, 
      sig_OP2_20_port, sig_OP2_19_port, sig_OP2_18_port, sig_OP2_17_port, 
      sig_OP2_16_port, sig_OP2_15_port, sig_OP2_14_port, sig_OP2_13_port, 
      sig_OP2_12_port, sig_OP2_11_port, sig_OP2_10_port, sig_OP2_9_port, 
      sig_OP2_8_port, sig_OP2_7_port, sig_OP2_6_port, sig_OP2_5_port, 
      sig_OP2_4_port, sig_OP2_3_port, sig_OP2_2_port, sig_OP2_1_port, 
      sig_OP2_0_port, sig_ALU_RES_31_port, sig_ALU_RES_30_port, 
      sig_ALU_RES_29_port, sig_ALU_RES_28_port, sig_ALU_RES_27_port, 
      sig_ALU_RES_26_port, sig_ALU_RES_25_port, sig_ALU_RES_24_port, 
      sig_ALU_RES_23_port, sig_ALU_RES_22_port, sig_ALU_RES_21_port, 
      sig_ALU_RES_20_port, sig_ALU_RES_19_port, sig_ALU_RES_18_port, 
      sig_ALU_RES_17_port, sig_ALU_RES_16_port, sig_ALU_RES_15_port, 
      sig_ALU_RES_14_port, sig_ALU_RES_13_port, sig_ALU_RES_12_port, 
      sig_ALU_RES_11_port, sig_ALU_RES_10_port, sig_ALU_RES_9_port, 
      sig_ALU_RES_8_port, sig_ALU_RES_7_port, sig_ALU_RES_6_port, 
      sig_ALU_RES_5_port, sig_ALU_RES_4_port, sig_ALU_RES_3_port, 
      sig_ALU_RES_2_port, sig_ALU_RES_1_port, sig_ALU_RES_0_port, n7, N9, N8, 
      N7_port, N6, N5, N4, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23, N22
      , N21, N20, N2, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N1, N0,
      n1_port, n8_port, n9_port, n10_port, OP2_FW_9_port, OP2_FW_8_port, 
      OP2_FW_7_port, OP2_FW_6_port, OP2_FW_5_port, OP2_FW_4_port, OP2_FW_3_port
      , OP2_FW_31_port, OP2_FW_30_port, OP2_FW_2_port, OP2_FW_29_port, 
      OP2_FW_28_port, OP2_FW_27_port, OP2_FW_26_port, OP2_FW_25_port, 
      OP2_FW_24_port, OP2_FW_23_port, OP2_FW_22_port, OP2_FW_21_port, 
      OP2_FW_20_port, OP2_FW_1_port, OP2_FW_19_port, OP2_FW_18_port, 
      OP2_FW_17_port, OP2_FW_16_port, OP2_FW_15_port, OP2_FW_14_port, 
      OP2_FW_13_port, OP2_FW_12_port, OP2_FW_11_port, OP2_FW_10_port, 
      OP2_FW_0_port, n11_port, n12_port, n13_port, n_1171, n_1172 : std_logic;

begin
   ZERO_FLAG <= ZERO_FLAG_port;
   
   n7 <= '1';
   n1_port <= '0';
   n8_port <= '1';
   n9_port <= '0';
   n10_port <= '0';
   Branch_Cond : Branch_Cond_Unit_NBIT32 port map( RST => sig_RST, A(31) => 
                           sig_NPC_ABS_31_port, A(30) => sig_NPC_ABS_30_port, 
                           A(29) => sig_NPC_ABS_29_port, A(28) => 
                           sig_NPC_ABS_28_port, A(27) => sig_NPC_ABS_27_port, 
                           A(26) => sig_NPC_ABS_26_port, A(25) => 
                           sig_NPC_ABS_25_port, A(24) => sig_NPC_ABS_24_port, 
                           A(23) => sig_NPC_ABS_23_port, A(22) => 
                           sig_NPC_ABS_22_port, A(21) => sig_NPC_ABS_21_port, 
                           A(20) => sig_NPC_ABS_20_port, A(19) => 
                           sig_NPC_ABS_19_port, A(18) => sig_NPC_ABS_18_port, 
                           A(17) => sig_NPC_ABS_17_port, A(16) => 
                           sig_NPC_ABS_16_port, A(15) => sig_NPC_ABS_15_port, 
                           A(14) => sig_NPC_ABS_14_port, A(13) => 
                           sig_NPC_ABS_13_port, A(12) => sig_NPC_ABS_12_port, 
                           A(11) => sig_NPC_ABS_11_port, A(10) => 
                           sig_NPC_ABS_10_port, A(9) => sig_NPC_ABS_9_port, 
                           A(8) => sig_NPC_ABS_8_port, A(7) => 
                           sig_NPC_ABS_7_port, A(6) => sig_NPC_ABS_6_port, A(5)
                           => sig_NPC_ABS_5_port, A(4) => sig_NPC_ABS_4_port, 
                           A(3) => sig_NPC_ABS_3_port, A(2) => 
                           sig_NPC_ABS_2_port, A(1) => sig_NPC_ABS_1_port, A(0)
                           => sig_NPC_ABS_0_port, ALU_OPC(0) => ALU_OPC(0), 
                           ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => ALU_OPC(2), 
                           ALU_OPC(3) => ALU_OPC(3), JUMP_TYPE(1) => 
                           JUMP_TYPE(1), JUMP_TYPE(0) => JUMP_TYPE(0), 
                           PC_SEL(1) => sig_PC_SEL_1_port, PC_SEL(0) => 
                           sig_PC_SEL_0_port, ZERO => sig_ZERO_FLAG);
   ff0 : ff_1 port map( D => sig_ZERO_FLAG, CLK => CLK, EN => n13_port, RST => 
                           RST, Q => ZERO_FLAG_port);
   reg0 : regn_N2 port map( DIN(1) => sig_PC_SEL_1_port, DIN(0) => 
                           sig_PC_SEL_0_port, CLK => CLK, EN => n7, RST => RST,
                           DOUT(1) => PC_SEL(1), DOUT(0) => PC_SEL(0));
   FWD : FWD_Unit port map( RST => sig_RST, ADD_RS1(4) => ADD_RS1_IN(4), 
                           ADD_RS1(3) => ADD_RS1_IN(3), ADD_RS1(2) => 
                           ADD_RS1_IN(2), ADD_RS1(1) => ADD_RS1_IN(1), 
                           ADD_RS1(0) => ADD_RS1_IN(0), ADD_RS2(4) => 
                           ADD_RS2_IN(4), ADD_RS2(3) => ADD_RS2_IN(3), 
                           ADD_RS2(2) => ADD_RS2_IN(2), ADD_RS2(1) => 
                           ADD_RS2_IN(1), ADD_RS2(0) => ADD_RS2_IN(0), 
                           ADD_WR_MEM(4) => ADD_WR_MEM(4), ADD_WR_MEM(3) => 
                           ADD_WR_MEM(3), ADD_WR_MEM(2) => ADD_WR_MEM(2), 
                           ADD_WR_MEM(1) => ADD_WR_MEM(1), ADD_WR_MEM(0) => 
                           ADD_WR_MEM(0), ADD_WR_WB(4) => ADD_WR_WB(4), 
                           ADD_WR_WB(3) => ADD_WR_WB(3), ADD_WR_WB(2) => 
                           ADD_WR_WB(2), ADD_WR_WB(1) => ADD_WR_WB(1), 
                           ADD_WR_WB(0) => ADD_WR_WB(0), RF_WE_MEM => RF_WE_MEM
                           , RF_WE_WB => RF_WE_WB, FWDA(1) => FWDA_1_port, 
                           FWDA(0) => FWDA_0_port, FWDB(1) => FWDB_1_port, 
                           FWDB(0) => FWDB_0_port);
   FW1 : mux41_NBIT32_0 port map( A(31) => A_IN(31), A(30) => A_IN(30), A(29) 
                           => A_IN(29), A(28) => A_IN(28), A(27) => A_IN(27), 
                           A(26) => A_IN(26), A(25) => A_IN(25), A(24) => 
                           A_IN(24), A(23) => A_IN(23), A(22) => A_IN(22), 
                           A(21) => A_IN(21), A(20) => A_IN(20), A(19) => 
                           A_IN(19), A(18) => A_IN(18), A(17) => A_IN(17), 
                           A(16) => A_IN(16), A(15) => A_IN(15), A(14) => 
                           A_IN(14), A(13) => A_IN(13), A(12) => A_IN(12), 
                           A(11) => A_IN(11), A(10) => A_IN(10), A(9) => 
                           A_IN(9), A(8) => A_IN(8), A(7) => A_IN(7), A(6) => 
                           A_IN(6), A(5) => A_IN(5), A(4) => A_IN(4), A(3) => 
                           A_IN(3), A(2) => A_IN(2), A(1) => A_IN(1), A(0) => 
                           A_IN(0), B(31) => OP_WB(31), B(30) => OP_WB(30), 
                           B(29) => OP_WB(29), B(28) => OP_WB(28), B(27) => 
                           OP_WB(27), B(26) => OP_WB(26), B(25) => OP_WB(25), 
                           B(24) => OP_WB(24), B(23) => OP_WB(23), B(22) => 
                           OP_WB(22), B(21) => OP_WB(21), B(20) => OP_WB(20), 
                           B(19) => OP_WB(19), B(18) => OP_WB(18), B(17) => 
                           OP_WB(17), B(16) => OP_WB(16), B(15) => OP_WB(15), 
                           B(14) => OP_WB(14), B(13) => OP_WB(13), B(12) => 
                           OP_WB(12), B(11) => OP_WB(11), B(10) => OP_WB(10), 
                           B(9) => OP_WB(9), B(8) => OP_WB(8), B(7) => OP_WB(7)
                           , B(6) => OP_WB(6), B(5) => OP_WB(5), B(4) => 
                           OP_WB(4), B(3) => OP_WB(3), B(2) => OP_WB(2), B(1) 
                           => OP_WB(1), B(0) => OP_WB(0), C(31) => OP_MEM(31), 
                           C(30) => OP_MEM(30), C(29) => OP_MEM(29), C(28) => 
                           OP_MEM(28), C(27) => OP_MEM(27), C(26) => OP_MEM(26)
                           , C(25) => OP_MEM(25), C(24) => OP_MEM(24), C(23) =>
                           OP_MEM(23), C(22) => OP_MEM(22), C(21) => OP_MEM(21)
                           , C(20) => OP_MEM(20), C(19) => OP_MEM(19), C(18) =>
                           OP_MEM(18), C(17) => OP_MEM(17), C(16) => OP_MEM(16)
                           , C(15) => OP_MEM(15), C(14) => OP_MEM(14), C(13) =>
                           OP_MEM(13), C(12) => OP_MEM(12), C(11) => OP_MEM(11)
                           , C(10) => OP_MEM(10), C(9) => OP_MEM(9), C(8) => 
                           OP_MEM(8), C(7) => OP_MEM(7), C(6) => OP_MEM(6), 
                           C(5) => OP_MEM(5), C(4) => OP_MEM(4), C(3) => 
                           OP_MEM(3), C(2) => OP_MEM(2), C(1) => OP_MEM(1), 
                           C(0) => OP_MEM(0), D(31) => n12_port, D(30) => 
                           n12_port, D(29) => n12_port, D(28) => n12_port, 
                           D(27) => n12_port, D(26) => n12_port, D(25) => 
                           n12_port, D(24) => n12_port, D(23) => n12_port, 
                           D(22) => n12_port, D(21) => n12_port, D(20) => 
                           n12_port, D(19) => n12_port, D(18) => n12_port, 
                           D(17) => n12_port, D(16) => n12_port, D(15) => 
                           n12_port, D(14) => n12_port, D(13) => n12_port, 
                           D(12) => n12_port, D(11) => n12_port, D(10) => 
                           n12_port, D(9) => n12_port, D(8) => n12_port, D(7) 
                           => n12_port, D(6) => n12_port, D(5) => n12_port, 
                           D(4) => n12_port, D(3) => n12_port, D(2) => n12_port
                           , D(1) => n12_port, D(0) => n12_port, S(1) => 
                           FWDA_1_port, S(0) => FWDA_0_port, Z(31) => 
                           sig_NPC_ABS_31_port, Z(30) => sig_NPC_ABS_30_port, 
                           Z(29) => sig_NPC_ABS_29_port, Z(28) => 
                           sig_NPC_ABS_28_port, Z(27) => sig_NPC_ABS_27_port, 
                           Z(26) => sig_NPC_ABS_26_port, Z(25) => 
                           sig_NPC_ABS_25_port, Z(24) => sig_NPC_ABS_24_port, 
                           Z(23) => sig_NPC_ABS_23_port, Z(22) => 
                           sig_NPC_ABS_22_port, Z(21) => sig_NPC_ABS_21_port, 
                           Z(20) => sig_NPC_ABS_20_port, Z(19) => 
                           sig_NPC_ABS_19_port, Z(18) => sig_NPC_ABS_18_port, 
                           Z(17) => sig_NPC_ABS_17_port, Z(16) => 
                           sig_NPC_ABS_16_port, Z(15) => sig_NPC_ABS_15_port, 
                           Z(14) => sig_NPC_ABS_14_port, Z(13) => 
                           sig_NPC_ABS_13_port, Z(12) => sig_NPC_ABS_12_port, 
                           Z(11) => sig_NPC_ABS_11_port, Z(10) => 
                           sig_NPC_ABS_10_port, Z(9) => sig_NPC_ABS_9_port, 
                           Z(8) => sig_NPC_ABS_8_port, Z(7) => 
                           sig_NPC_ABS_7_port, Z(6) => sig_NPC_ABS_6_port, Z(5)
                           => sig_NPC_ABS_5_port, Z(4) => sig_NPC_ABS_4_port, 
                           Z(3) => sig_NPC_ABS_3_port, Z(2) => 
                           sig_NPC_ABS_2_port, Z(1) => sig_NPC_ABS_1_port, Z(0)
                           => sig_NPC_ABS_0_port);
   FW2 : mux41_NBIT32_4 port map( A(31) => B_IN(31), A(30) => B_IN(30), A(29) 
                           => B_IN(29), A(28) => B_IN(28), A(27) => B_IN(27), 
                           A(26) => B_IN(26), A(25) => B_IN(25), A(24) => 
                           B_IN(24), A(23) => B_IN(23), A(22) => B_IN(22), 
                           A(21) => B_IN(21), A(20) => B_IN(20), A(19) => 
                           B_IN(19), A(18) => B_IN(18), A(17) => B_IN(17), 
                           A(16) => B_IN(16), A(15) => B_IN(15), A(14) => 
                           B_IN(14), A(13) => B_IN(13), A(12) => B_IN(12), 
                           A(11) => B_IN(11), A(10) => B_IN(10), A(9) => 
                           B_IN(9), A(8) => B_IN(8), A(7) => B_IN(7), A(6) => 
                           B_IN(6), A(5) => B_IN(5), A(4) => B_IN(4), A(3) => 
                           B_IN(3), A(2) => B_IN(2), A(1) => B_IN(1), A(0) => 
                           B_IN(0), B(31) => OP_WB(31), B(30) => OP_WB(30), 
                           B(29) => OP_WB(29), B(28) => OP_WB(28), B(27) => 
                           OP_WB(27), B(26) => OP_WB(26), B(25) => OP_WB(25), 
                           B(24) => OP_WB(24), B(23) => OP_WB(23), B(22) => 
                           OP_WB(22), B(21) => OP_WB(21), B(20) => OP_WB(20), 
                           B(19) => OP_WB(19), B(18) => OP_WB(18), B(17) => 
                           OP_WB(17), B(16) => OP_WB(16), B(15) => OP_WB(15), 
                           B(14) => OP_WB(14), B(13) => OP_WB(13), B(12) => 
                           OP_WB(12), B(11) => OP_WB(11), B(10) => OP_WB(10), 
                           B(9) => OP_WB(9), B(8) => OP_WB(8), B(7) => OP_WB(7)
                           , B(6) => OP_WB(6), B(5) => OP_WB(5), B(4) => 
                           OP_WB(4), B(3) => OP_WB(3), B(2) => OP_WB(2), B(1) 
                           => OP_WB(1), B(0) => OP_WB(0), C(31) => OP_MEM(31), 
                           C(30) => OP_MEM(30), C(29) => OP_MEM(29), C(28) => 
                           OP_MEM(28), C(27) => OP_MEM(27), C(26) => OP_MEM(26)
                           , C(25) => OP_MEM(25), C(24) => OP_MEM(24), C(23) =>
                           OP_MEM(23), C(22) => OP_MEM(22), C(21) => OP_MEM(21)
                           , C(20) => OP_MEM(20), C(19) => OP_MEM(19), C(18) =>
                           OP_MEM(18), C(17) => OP_MEM(17), C(16) => OP_MEM(16)
                           , C(15) => OP_MEM(15), C(14) => OP_MEM(14), C(13) =>
                           OP_MEM(13), C(12) => OP_MEM(12), C(11) => OP_MEM(11)
                           , C(10) => OP_MEM(10), C(9) => OP_MEM(9), C(8) => 
                           OP_MEM(8), C(7) => OP_MEM(7), C(6) => OP_MEM(6), 
                           C(5) => OP_MEM(5), C(4) => OP_MEM(4), C(3) => 
                           OP_MEM(3), C(2) => OP_MEM(2), C(1) => OP_MEM(1), 
                           C(0) => OP_MEM(0), D(31) => n12_port, D(30) => 
                           n12_port, D(29) => n12_port, D(28) => n12_port, 
                           D(27) => n12_port, D(26) => n12_port, D(25) => 
                           n12_port, D(24) => n12_port, D(23) => n12_port, 
                           D(22) => n12_port, D(21) => n12_port, D(20) => 
                           n12_port, D(19) => n12_port, D(18) => n12_port, 
                           D(17) => n12_port, D(16) => n12_port, D(15) => 
                           n12_port, D(14) => n12_port, D(13) => n12_port, 
                           D(12) => n12_port, D(11) => n12_port, D(10) => 
                           n12_port, D(9) => n12_port, D(8) => n12_port, D(7) 
                           => n12_port, D(6) => n12_port, D(5) => n12_port, 
                           D(4) => n12_port, D(3) => n12_port, D(2) => n12_port
                           , D(1) => n12_port, D(0) => n12_port, S(1) => 
                           FWDB_1_port, S(0) => FWDB_0_port, Z(31) => 
                           OP2_FW_31_port, Z(30) => OP2_FW_30_port, Z(29) => 
                           OP2_FW_29_port, Z(28) => OP2_FW_28_port, Z(27) => 
                           OP2_FW_27_port, Z(26) => OP2_FW_26_port, Z(25) => 
                           OP2_FW_25_port, Z(24) => OP2_FW_24_port, Z(23) => 
                           OP2_FW_23_port, Z(22) => OP2_FW_22_port, Z(21) => 
                           OP2_FW_21_port, Z(20) => OP2_FW_20_port, Z(19) => 
                           OP2_FW_19_port, Z(18) => OP2_FW_18_port, Z(17) => 
                           OP2_FW_17_port, Z(16) => OP2_FW_16_port, Z(15) => 
                           OP2_FW_15_port, Z(14) => OP2_FW_14_port, Z(13) => 
                           OP2_FW_13_port, Z(12) => OP2_FW_12_port, Z(11) => 
                           OP2_FW_11_port, Z(10) => OP2_FW_10_port, Z(9) => 
                           OP2_FW_9_port, Z(8) => OP2_FW_8_port, Z(7) => 
                           OP2_FW_7_port, Z(6) => OP2_FW_6_port, Z(5) => 
                           OP2_FW_5_port, Z(4) => OP2_FW_4_port, Z(3) => 
                           OP2_FW_3_port, Z(2) => OP2_FW_2_port, Z(1) => 
                           OP2_FW_1_port, Z(0) => OP2_FW_0_port);
   muxA : mux21_NBIT32_3 port map( A(31) => sig_NPC_ABS_31_port, A(30) => 
                           sig_NPC_ABS_30_port, A(29) => sig_NPC_ABS_29_port, 
                           A(28) => sig_NPC_ABS_28_port, A(27) => 
                           sig_NPC_ABS_27_port, A(26) => sig_NPC_ABS_26_port, 
                           A(25) => sig_NPC_ABS_25_port, A(24) => 
                           sig_NPC_ABS_24_port, A(23) => sig_NPC_ABS_23_port, 
                           A(22) => sig_NPC_ABS_22_port, A(21) => 
                           sig_NPC_ABS_21_port, A(20) => sig_NPC_ABS_20_port, 
                           A(19) => sig_NPC_ABS_19_port, A(18) => 
                           sig_NPC_ABS_18_port, A(17) => sig_NPC_ABS_17_port, 
                           A(16) => sig_NPC_ABS_16_port, A(15) => 
                           sig_NPC_ABS_15_port, A(14) => sig_NPC_ABS_14_port, 
                           A(13) => sig_NPC_ABS_13_port, A(12) => 
                           sig_NPC_ABS_12_port, A(11) => sig_NPC_ABS_11_port, 
                           A(10) => sig_NPC_ABS_10_port, A(9) => 
                           sig_NPC_ABS_9_port, A(8) => sig_NPC_ABS_8_port, A(7)
                           => sig_NPC_ABS_7_port, A(6) => sig_NPC_ABS_6_port, 
                           A(5) => sig_NPC_ABS_5_port, A(4) => 
                           sig_NPC_ABS_4_port, A(3) => sig_NPC_ABS_3_port, A(2)
                           => sig_NPC_ABS_2_port, A(1) => sig_NPC_ABS_1_port, 
                           A(0) => sig_NPC_ABS_0_port, B(31) => PC_IN(31), 
                           B(30) => PC_IN(30), B(29) => PC_IN(29), B(28) => 
                           PC_IN(28), B(27) => PC_IN(27), B(26) => PC_IN(26), 
                           B(25) => PC_IN(25), B(24) => PC_IN(24), B(23) => 
                           PC_IN(23), B(22) => PC_IN(22), B(21) => PC_IN(21), 
                           B(20) => PC_IN(20), B(19) => PC_IN(19), B(18) => 
                           PC_IN(18), B(17) => PC_IN(17), B(16) => PC_IN(16), 
                           B(15) => PC_IN(15), B(14) => PC_IN(14), B(13) => 
                           PC_IN(13), B(12) => PC_IN(12), B(11) => PC_IN(11), 
                           B(10) => PC_IN(10), B(9) => PC_IN(9), B(8) => 
                           PC_IN(8), B(7) => PC_IN(7), B(6) => PC_IN(6), B(5) 
                           => PC_IN(5), B(4) => PC_IN(4), B(3) => PC_IN(3), 
                           B(2) => PC_IN(2), B(1) => PC_IN(1), B(0) => PC_IN(0)
                           , S => MUX_A_SEL, Z(31) => sig_OP1_31_port, Z(30) =>
                           sig_OP1_30_port, Z(29) => sig_OP1_29_port, Z(28) => 
                           sig_OP1_28_port, Z(27) => sig_OP1_27_port, Z(26) => 
                           sig_OP1_26_port, Z(25) => sig_OP1_25_port, Z(24) => 
                           sig_OP1_24_port, Z(23) => sig_OP1_23_port, Z(22) => 
                           sig_OP1_22_port, Z(21) => sig_OP1_21_port, Z(20) => 
                           sig_OP1_20_port, Z(19) => sig_OP1_19_port, Z(18) => 
                           sig_OP1_18_port, Z(17) => sig_OP1_17_port, Z(16) => 
                           sig_OP1_16_port, Z(15) => sig_OP1_15_port, Z(14) => 
                           sig_OP1_14_port, Z(13) => sig_OP1_13_port, Z(12) => 
                           sig_OP1_12_port, Z(11) => sig_OP1_11_port, Z(10) => 
                           sig_OP1_10_port, Z(9) => sig_OP1_9_port, Z(8) => 
                           sig_OP1_8_port, Z(7) => sig_OP1_7_port, Z(6) => 
                           sig_OP1_6_port, Z(5) => sig_OP1_5_port, Z(4) => 
                           sig_OP1_4_port, Z(3) => sig_OP1_3_port, Z(2) => 
                           sig_OP1_2_port, Z(1) => sig_OP1_1_port, Z(0) => 
                           sig_OP1_0_port);
   muxB : mux41_NBIT32_3 port map( A(31) => OP2_FW_31_port, A(30) => 
                           OP2_FW_30_port, A(29) => OP2_FW_29_port, A(28) => 
                           OP2_FW_28_port, A(27) => OP2_FW_27_port, A(26) => 
                           OP2_FW_26_port, A(25) => OP2_FW_25_port, A(24) => 
                           OP2_FW_24_port, A(23) => OP2_FW_23_port, A(22) => 
                           OP2_FW_22_port, A(21) => OP2_FW_21_port, A(20) => 
                           OP2_FW_20_port, A(19) => OP2_FW_19_port, A(18) => 
                           OP2_FW_18_port, A(17) => OP2_FW_17_port, A(16) => 
                           OP2_FW_16_port, A(15) => OP2_FW_15_port, A(14) => 
                           OP2_FW_14_port, A(13) => OP2_FW_13_port, A(12) => 
                           OP2_FW_12_port, A(11) => OP2_FW_11_port, A(10) => 
                           OP2_FW_10_port, A(9) => OP2_FW_9_port, A(8) => 
                           OP2_FW_8_port, A(7) => OP2_FW_7_port, A(6) => 
                           OP2_FW_6_port, A(5) => OP2_FW_5_port, A(4) => 
                           OP2_FW_4_port, A(3) => OP2_FW_3_port, A(2) => 
                           OP2_FW_2_port, A(1) => OP2_FW_1_port, A(0) => 
                           OP2_FW_0_port, B(31) => IMM_IN(31), B(30) => 
                           IMM_IN(30), B(29) => IMM_IN(29), B(28) => IMM_IN(28)
                           , B(27) => IMM_IN(27), B(26) => IMM_IN(26), B(25) =>
                           IMM_IN(25), B(24) => IMM_IN(24), B(23) => IMM_IN(23)
                           , B(22) => IMM_IN(22), B(21) => IMM_IN(21), B(20) =>
                           IMM_IN(20), B(19) => IMM_IN(19), B(18) => IMM_IN(18)
                           , B(17) => IMM_IN(17), B(16) => IMM_IN(16), B(15) =>
                           IMM_IN(15), B(14) => IMM_IN(14), B(13) => IMM_IN(13)
                           , B(12) => IMM_IN(12), B(11) => IMM_IN(11), B(10) =>
                           IMM_IN(10), B(9) => IMM_IN(9), B(8) => IMM_IN(8), 
                           B(7) => IMM_IN(7), B(6) => IMM_IN(6), B(5) => 
                           IMM_IN(5), B(4) => IMM_IN(4), B(3) => IMM_IN(3), 
                           B(2) => IMM_IN(2), B(1) => IMM_IN(1), B(0) => 
                           IMM_IN(0), C(31) => n12_port, C(30) => n12_port, 
                           C(29) => n12_port, C(28) => n12_port, C(27) => 
                           n12_port, C(26) => n12_port, C(25) => n12_port, 
                           C(24) => n12_port, C(23) => n12_port, C(22) => 
                           n12_port, C(21) => n12_port, C(20) => n12_port, 
                           C(19) => n12_port, C(18) => n12_port, C(17) => 
                           n12_port, C(16) => n12_port, C(15) => n12_port, 
                           C(14) => n12_port, C(13) => n12_port, C(12) => 
                           n12_port, C(11) => n12_port, C(10) => n12_port, C(9)
                           => n12_port, C(8) => n12_port, C(7) => n12_port, 
                           C(6) => n12_port, C(5) => n12_port, C(4) => n12_port
                           , C(3) => n12_port, C(2) => n13_port, C(1) => 
                           n12_port, C(0) => n12_port, D(31) => n12_port, D(30)
                           => n12_port, D(29) => n12_port, D(28) => n12_port, 
                           D(27) => n12_port, D(26) => n12_port, D(25) => 
                           n12_port, D(24) => n12_port, D(23) => n12_port, 
                           D(22) => n12_port, D(21) => n12_port, D(20) => 
                           n12_port, D(19) => n12_port, D(18) => n12_port, 
                           D(17) => n12_port, D(16) => n12_port, D(15) => 
                           n12_port, D(14) => n12_port, D(13) => n12_port, 
                           D(12) => n12_port, D(11) => n12_port, D(10) => 
                           n12_port, D(9) => n12_port, D(8) => n12_port, D(7) 
                           => n12_port, D(6) => n12_port, D(5) => n12_port, 
                           D(4) => n12_port, D(3) => n12_port, D(2) => n12_port
                           , D(1) => n12_port, D(0) => n12_port, S(1) => 
                           MUX_B_SEL(1), S(0) => MUX_B_SEL(0), Z(31) => 
                           sig_OP2_31_port, Z(30) => sig_OP2_30_port, Z(29) => 
                           sig_OP2_29_port, Z(28) => sig_OP2_28_port, Z(27) => 
                           sig_OP2_27_port, Z(26) => sig_OP2_26_port, Z(25) => 
                           sig_OP2_25_port, Z(24) => sig_OP2_24_port, Z(23) => 
                           sig_OP2_23_port, Z(22) => sig_OP2_22_port, Z(21) => 
                           sig_OP2_21_port, Z(20) => sig_OP2_20_port, Z(19) => 
                           sig_OP2_19_port, Z(18) => sig_OP2_18_port, Z(17) => 
                           sig_OP2_17_port, Z(16) => sig_OP2_16_port, Z(15) => 
                           sig_OP2_15_port, Z(14) => sig_OP2_14_port, Z(13) => 
                           sig_OP2_13_port, Z(12) => sig_OP2_12_port, Z(11) => 
                           sig_OP2_11_port, Z(10) => sig_OP2_10_port, Z(9) => 
                           sig_OP2_9_port, Z(8) => sig_OP2_8_port, Z(7) => 
                           sig_OP2_7_port, Z(6) => sig_OP2_6_port, Z(5) => 
                           sig_OP2_5_port, Z(4) => sig_OP2_4_port, Z(3) => 
                           sig_OP2_3_port, Z(2) => sig_OP2_2_port, Z(1) => 
                           sig_OP2_1_port, Z(0) => sig_OP2_0_port);
   alu0 : ALU_NBIT32 port map( OP1(31) => sig_OP1_31_port, OP1(30) => 
                           sig_OP1_30_port, OP1(29) => sig_OP1_29_port, OP1(28)
                           => sig_OP1_28_port, OP1(27) => sig_OP1_27_port, 
                           OP1(26) => sig_OP1_26_port, OP1(25) => 
                           sig_OP1_25_port, OP1(24) => sig_OP1_24_port, OP1(23)
                           => sig_OP1_23_port, OP1(22) => sig_OP1_22_port, 
                           OP1(21) => sig_OP1_21_port, OP1(20) => 
                           sig_OP1_20_port, OP1(19) => sig_OP1_19_port, OP1(18)
                           => sig_OP1_18_port, OP1(17) => sig_OP1_17_port, 
                           OP1(16) => sig_OP1_16_port, OP1(15) => 
                           sig_OP1_15_port, OP1(14) => sig_OP1_14_port, OP1(13)
                           => sig_OP1_13_port, OP1(12) => sig_OP1_12_port, 
                           OP1(11) => sig_OP1_11_port, OP1(10) => 
                           sig_OP1_10_port, OP1(9) => sig_OP1_9_port, OP1(8) =>
                           sig_OP1_8_port, OP1(7) => sig_OP1_7_port, OP1(6) => 
                           sig_OP1_6_port, OP1(5) => sig_OP1_5_port, OP1(4) => 
                           sig_OP1_4_port, OP1(3) => sig_OP1_3_port, OP1(2) => 
                           sig_OP1_2_port, OP1(1) => sig_OP1_1_port, OP1(0) => 
                           sig_OP1_0_port, OP2(31) => sig_OP2_31_port, OP2(30) 
                           => sig_OP2_30_port, OP2(29) => sig_OP2_29_port, 
                           OP2(28) => sig_OP2_28_port, OP2(27) => 
                           sig_OP2_27_port, OP2(26) => sig_OP2_26_port, OP2(25)
                           => sig_OP2_25_port, OP2(24) => sig_OP2_24_port, 
                           OP2(23) => sig_OP2_23_port, OP2(22) => 
                           sig_OP2_22_port, OP2(21) => sig_OP2_21_port, OP2(20)
                           => sig_OP2_20_port, OP2(19) => sig_OP2_19_port, 
                           OP2(18) => sig_OP2_18_port, OP2(17) => 
                           sig_OP2_17_port, OP2(16) => sig_OP2_16_port, OP2(15)
                           => sig_OP2_15_port, OP2(14) => sig_OP2_14_port, 
                           OP2(13) => sig_OP2_13_port, OP2(12) => 
                           sig_OP2_12_port, OP2(11) => sig_OP2_11_port, OP2(10)
                           => sig_OP2_10_port, OP2(9) => sig_OP2_9_port, OP2(8)
                           => sig_OP2_8_port, OP2(7) => sig_OP2_7_port, OP2(6) 
                           => sig_OP2_6_port, OP2(5) => sig_OP2_5_port, OP2(4) 
                           => sig_OP2_4_port, OP2(3) => sig_OP2_3_port, OP2(2) 
                           => sig_OP2_2_port, OP2(1) => sig_OP2_1_port, OP2(0) 
                           => sig_OP2_0_port, ALU_OPC(0) => ALU_OPC(0), 
                           ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => ALU_OPC(2), 
                           ALU_OPC(3) => ALU_OPC(3), ALU_RES(31) => 
                           sig_ALU_RES_31_port, ALU_RES(30) => 
                           sig_ALU_RES_30_port, ALU_RES(29) => 
                           sig_ALU_RES_29_port, ALU_RES(28) => 
                           sig_ALU_RES_28_port, ALU_RES(27) => 
                           sig_ALU_RES_27_port, ALU_RES(26) => 
                           sig_ALU_RES_26_port, ALU_RES(25) => 
                           sig_ALU_RES_25_port, ALU_RES(24) => 
                           sig_ALU_RES_24_port, ALU_RES(23) => 
                           sig_ALU_RES_23_port, ALU_RES(22) => 
                           sig_ALU_RES_22_port, ALU_RES(21) => 
                           sig_ALU_RES_21_port, ALU_RES(20) => 
                           sig_ALU_RES_20_port, ALU_RES(19) => 
                           sig_ALU_RES_19_port, ALU_RES(18) => 
                           sig_ALU_RES_18_port, ALU_RES(17) => 
                           sig_ALU_RES_17_port, ALU_RES(16) => 
                           sig_ALU_RES_16_port, ALU_RES(15) => 
                           sig_ALU_RES_15_port, ALU_RES(14) => 
                           sig_ALU_RES_14_port, ALU_RES(13) => 
                           sig_ALU_RES_13_port, ALU_RES(12) => 
                           sig_ALU_RES_12_port, ALU_RES(11) => 
                           sig_ALU_RES_11_port, ALU_RES(10) => 
                           sig_ALU_RES_10_port, ALU_RES(9) => 
                           sig_ALU_RES_9_port, ALU_RES(8) => sig_ALU_RES_8_port
                           , ALU_RES(7) => sig_ALU_RES_7_port, ALU_RES(6) => 
                           sig_ALU_RES_6_port, ALU_RES(5) => sig_ALU_RES_5_port
                           , ALU_RES(4) => sig_ALU_RES_4_port, ALU_RES(3) => 
                           sig_ALU_RES_3_port, ALU_RES(2) => sig_ALU_RES_2_port
                           , ALU_RES(1) => sig_ALU_RES_1_port, ALU_RES(0) => 
                           sig_ALU_RES_0_port);
   alureg : regn_N32_6 port map( DIN(31) => sig_ALU_RES_31_port, DIN(30) => 
                           sig_ALU_RES_30_port, DIN(29) => sig_ALU_RES_29_port,
                           DIN(28) => sig_ALU_RES_28_port, DIN(27) => 
                           sig_ALU_RES_27_port, DIN(26) => sig_ALU_RES_26_port,
                           DIN(25) => sig_ALU_RES_25_port, DIN(24) => 
                           sig_ALU_RES_24_port, DIN(23) => sig_ALU_RES_23_port,
                           DIN(22) => sig_ALU_RES_22_port, DIN(21) => 
                           sig_ALU_RES_21_port, DIN(20) => sig_ALU_RES_20_port,
                           DIN(19) => sig_ALU_RES_19_port, DIN(18) => 
                           sig_ALU_RES_18_port, DIN(17) => sig_ALU_RES_17_port,
                           DIN(16) => sig_ALU_RES_16_port, DIN(15) => 
                           sig_ALU_RES_15_port, DIN(14) => sig_ALU_RES_14_port,
                           DIN(13) => sig_ALU_RES_13_port, DIN(12) => 
                           sig_ALU_RES_12_port, DIN(11) => sig_ALU_RES_11_port,
                           DIN(10) => sig_ALU_RES_10_port, DIN(9) => 
                           sig_ALU_RES_9_port, DIN(8) => sig_ALU_RES_8_port, 
                           DIN(7) => sig_ALU_RES_7_port, DIN(6) => 
                           sig_ALU_RES_6_port, DIN(5) => sig_ALU_RES_5_port, 
                           DIN(4) => sig_ALU_RES_4_port, DIN(3) => 
                           sig_ALU_RES_3_port, DIN(2) => sig_ALU_RES_2_port, 
                           DIN(1) => sig_ALU_RES_1_port, DIN(0) => 
                           sig_ALU_RES_0_port, CLK => CLK, EN => ALU_OUTREG_EN,
                           RST => RST, DOUT(31) => ALU_RES(31), DOUT(30) => 
                           ALU_RES(30), DOUT(29) => ALU_RES(29), DOUT(28) => 
                           ALU_RES(28), DOUT(27) => ALU_RES(27), DOUT(26) => 
                           ALU_RES(26), DOUT(25) => ALU_RES(25), DOUT(24) => 
                           ALU_RES(24), DOUT(23) => ALU_RES(23), DOUT(22) => 
                           ALU_RES(22), DOUT(21) => ALU_RES(21), DOUT(20) => 
                           ALU_RES(20), DOUT(19) => ALU_RES(19), DOUT(18) => 
                           ALU_RES(18), DOUT(17) => ALU_RES(17), DOUT(16) => 
                           ALU_RES(16), DOUT(15) => ALU_RES(15), DOUT(14) => 
                           ALU_RES(14), DOUT(13) => ALU_RES(13), DOUT(12) => 
                           ALU_RES(12), DOUT(11) => ALU_RES(11), DOUT(10) => 
                           ALU_RES(10), DOUT(9) => ALU_RES(9), DOUT(8) => 
                           ALU_RES(8), DOUT(7) => ALU_RES(7), DOUT(6) => 
                           ALU_RES(6), DOUT(5) => ALU_RES(5), DOUT(4) => 
                           ALU_RES(4), DOUT(3) => ALU_RES(3), DOUT(2) => 
                           ALU_RES(2), DOUT(1) => ALU_RES(1), DOUT(0) => 
                           ALU_RES(0));
   B_reg : regn_N32_5 port map( DIN(31) => OP2_FW_31_port, DIN(30) => 
                           OP2_FW_30_port, DIN(29) => OP2_FW_29_port, DIN(28) 
                           => OP2_FW_28_port, DIN(27) => OP2_FW_27_port, 
                           DIN(26) => OP2_FW_26_port, DIN(25) => OP2_FW_25_port
                           , DIN(24) => OP2_FW_24_port, DIN(23) => 
                           OP2_FW_23_port, DIN(22) => OP2_FW_22_port, DIN(21) 
                           => OP2_FW_21_port, DIN(20) => OP2_FW_20_port, 
                           DIN(19) => OP2_FW_19_port, DIN(18) => OP2_FW_18_port
                           , DIN(17) => OP2_FW_17_port, DIN(16) => 
                           OP2_FW_16_port, DIN(15) => OP2_FW_15_port, DIN(14) 
                           => OP2_FW_14_port, DIN(13) => OP2_FW_13_port, 
                           DIN(12) => OP2_FW_12_port, DIN(11) => OP2_FW_11_port
                           , DIN(10) => OP2_FW_10_port, DIN(9) => OP2_FW_9_port
                           , DIN(8) => OP2_FW_8_port, DIN(7) => OP2_FW_7_port, 
                           DIN(6) => OP2_FW_6_port, DIN(5) => OP2_FW_5_port, 
                           DIN(4) => OP2_FW_4_port, DIN(3) => OP2_FW_3_port, 
                           DIN(2) => OP2_FW_2_port, DIN(1) => OP2_FW_1_port, 
                           DIN(0) => OP2_FW_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => B_OUT(31), 
                           DOUT(30) => B_OUT(30), DOUT(29) => B_OUT(29), 
                           DOUT(28) => B_OUT(28), DOUT(27) => B_OUT(27), 
                           DOUT(26) => B_OUT(26), DOUT(25) => B_OUT(25), 
                           DOUT(24) => B_OUT(24), DOUT(23) => B_OUT(23), 
                           DOUT(22) => B_OUT(22), DOUT(21) => B_OUT(21), 
                           DOUT(20) => B_OUT(20), DOUT(19) => B_OUT(19), 
                           DOUT(18) => B_OUT(18), DOUT(17) => B_OUT(17), 
                           DOUT(16) => B_OUT(16), DOUT(15) => B_OUT(15), 
                           DOUT(14) => B_OUT(14), DOUT(13) => B_OUT(13), 
                           DOUT(12) => B_OUT(12), DOUT(11) => B_OUT(11), 
                           DOUT(10) => B_OUT(10), DOUT(9) => B_OUT(9), DOUT(8) 
                           => B_OUT(8), DOUT(7) => B_OUT(7), DOUT(6) => 
                           B_OUT(6), DOUT(5) => B_OUT(5), DOUT(4) => B_OUT(4), 
                           DOUT(3) => B_OUT(3), DOUT(2) => B_OUT(2), DOUT(1) =>
                           B_OUT(1), DOUT(0) => B_OUT(0));
   ADD_WR_reg : regn_N5_2 port map( DIN(4) => ADD_WR_IN(4), DIN(3) => 
                           ADD_WR_IN(3), DIN(2) => ADD_WR_IN(2), DIN(1) => 
                           ADD_WR_IN(1), DIN(0) => ADD_WR_IN(0), CLK => CLK, EN
                           => ALU_OUTREG_EN, RST => RST, DOUT(4) => 
                           ADD_WR_OUT(4), DOUT(3) => ADD_WR_OUT(3), DOUT(2) => 
                           ADD_WR_OUT(2), DOUT(1) => ADD_WR_OUT(1), DOUT(0) => 
                           ADD_WR_OUT(0));
   NPC_ABS_reg : regn_N32_4 port map( DIN(31) => sig_NPC_ABS_31_port, DIN(30) 
                           => sig_NPC_ABS_30_port, DIN(29) => 
                           sig_NPC_ABS_29_port, DIN(28) => sig_NPC_ABS_28_port,
                           DIN(27) => sig_NPC_ABS_27_port, DIN(26) => 
                           sig_NPC_ABS_26_port, DIN(25) => sig_NPC_ABS_25_port,
                           DIN(24) => sig_NPC_ABS_24_port, DIN(23) => 
                           sig_NPC_ABS_23_port, DIN(22) => sig_NPC_ABS_22_port,
                           DIN(21) => sig_NPC_ABS_21_port, DIN(20) => 
                           sig_NPC_ABS_20_port, DIN(19) => sig_NPC_ABS_19_port,
                           DIN(18) => sig_NPC_ABS_18_port, DIN(17) => 
                           sig_NPC_ABS_17_port, DIN(16) => sig_NPC_ABS_16_port,
                           DIN(15) => sig_NPC_ABS_15_port, DIN(14) => 
                           sig_NPC_ABS_14_port, DIN(13) => sig_NPC_ABS_13_port,
                           DIN(12) => sig_NPC_ABS_12_port, DIN(11) => 
                           sig_NPC_ABS_11_port, DIN(10) => sig_NPC_ABS_10_port,
                           DIN(9) => sig_NPC_ABS_9_port, DIN(8) => 
                           sig_NPC_ABS_8_port, DIN(7) => sig_NPC_ABS_7_port, 
                           DIN(6) => sig_NPC_ABS_6_port, DIN(5) => 
                           sig_NPC_ABS_5_port, DIN(4) => sig_NPC_ABS_4_port, 
                           DIN(3) => sig_NPC_ABS_3_port, DIN(2) => 
                           sig_NPC_ABS_2_port, DIN(1) => sig_NPC_ABS_1_port, 
                           DIN(0) => sig_NPC_ABS_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => NPC_ABS(31), 
                           DOUT(30) => NPC_ABS(30), DOUT(29) => NPC_ABS(29), 
                           DOUT(28) => NPC_ABS(28), DOUT(27) => NPC_ABS(27), 
                           DOUT(26) => NPC_ABS(26), DOUT(25) => NPC_ABS(25), 
                           DOUT(24) => NPC_ABS(24), DOUT(23) => NPC_ABS(23), 
                           DOUT(22) => NPC_ABS(22), DOUT(21) => NPC_ABS(21), 
                           DOUT(20) => NPC_ABS(20), DOUT(19) => NPC_ABS(19), 
                           DOUT(18) => NPC_ABS(18), DOUT(17) => NPC_ABS(17), 
                           DOUT(16) => NPC_ABS(16), DOUT(15) => NPC_ABS(15), 
                           DOUT(14) => NPC_ABS(14), DOUT(13) => NPC_ABS(13), 
                           DOUT(12) => NPC_ABS(12), DOUT(11) => NPC_ABS(11), 
                           DOUT(10) => NPC_ABS(10), DOUT(9) => NPC_ABS(9), 
                           DOUT(8) => NPC_ABS(8), DOUT(7) => NPC_ABS(7), 
                           DOUT(6) => NPC_ABS(6), DOUT(5) => NPC_ABS(5), 
                           DOUT(4) => NPC_ABS(4), DOUT(3) => NPC_ABS(3), 
                           DOUT(2) => NPC_ABS(2), DOUT(1) => NPC_ABS(1), 
                           DOUT(0) => NPC_ABS(0));
   NPC_REL_reg : regn_N32_3 port map( DIN(31) => sig_NPC_REL_31_port, DIN(30) 
                           => sig_NPC_REL_30_port, DIN(29) => 
                           sig_NPC_REL_29_port, DIN(28) => sig_NPC_REL_28_port,
                           DIN(27) => sig_NPC_REL_27_port, DIN(26) => 
                           sig_NPC_REL_26_port, DIN(25) => sig_NPC_REL_25_port,
                           DIN(24) => sig_NPC_REL_24_port, DIN(23) => 
                           sig_NPC_REL_23_port, DIN(22) => sig_NPC_REL_22_port,
                           DIN(21) => sig_NPC_REL_21_port, DIN(20) => 
                           sig_NPC_REL_20_port, DIN(19) => sig_NPC_REL_19_port,
                           DIN(18) => sig_NPC_REL_18_port, DIN(17) => 
                           sig_NPC_REL_17_port, DIN(16) => sig_NPC_REL_16_port,
                           DIN(15) => sig_NPC_REL_15_port, DIN(14) => 
                           sig_NPC_REL_14_port, DIN(13) => sig_NPC_REL_13_port,
                           DIN(12) => sig_NPC_REL_12_port, DIN(11) => 
                           sig_NPC_REL_11_port, DIN(10) => sig_NPC_REL_10_port,
                           DIN(9) => sig_NPC_REL_9_port, DIN(8) => 
                           sig_NPC_REL_8_port, DIN(7) => sig_NPC_REL_7_port, 
                           DIN(6) => sig_NPC_REL_6_port, DIN(5) => 
                           sig_NPC_REL_5_port, DIN(4) => sig_NPC_REL_4_port, 
                           DIN(3) => sig_NPC_REL_3_port, DIN(2) => 
                           sig_NPC_REL_2_port, DIN(1) => sig_NPC_REL_1_port, 
                           DIN(0) => sig_NPC_REL_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => NPC_REL(31), 
                           DOUT(30) => NPC_REL(30), DOUT(29) => NPC_REL(29), 
                           DOUT(28) => NPC_REL(28), DOUT(27) => NPC_REL(27), 
                           DOUT(26) => NPC_REL(26), DOUT(25) => NPC_REL(25), 
                           DOUT(24) => NPC_REL(24), DOUT(23) => NPC_REL(23), 
                           DOUT(22) => NPC_REL(22), DOUT(21) => NPC_REL(21), 
                           DOUT(20) => NPC_REL(20), DOUT(19) => NPC_REL(19), 
                           DOUT(18) => NPC_REL(18), DOUT(17) => NPC_REL(17), 
                           DOUT(16) => NPC_REL(16), DOUT(15) => NPC_REL(15), 
                           DOUT(14) => NPC_REL(14), DOUT(13) => NPC_REL(13), 
                           DOUT(12) => NPC_REL(12), DOUT(11) => NPC_REL(11), 
                           DOUT(10) => NPC_REL(10), DOUT(9) => NPC_REL(9), 
                           DOUT(8) => NPC_REL(8), DOUT(7) => NPC_REL(7), 
                           DOUT(6) => NPC_REL(6), DOUT(5) => NPC_REL(5), 
                           DOUT(4) => NPC_REL(4), DOUT(3) => NPC_REL(3), 
                           DOUT(2) => NPC_REL(2), DOUT(1) => NPC_REL(1), 
                           DOUT(0) => NPC_REL(0));
   add_1_root_add_0_root_add_118_2 : Execute_DW01_add_1 port map( A(31) => 
                           n1_port, A(30) => n1_port, A(29) => n1_port, A(28) 
                           => n1_port, A(27) => n1_port, A(26) => n1_port, 
                           A(25) => n1_port, A(24) => n1_port, A(23) => n1_port
                           , A(22) => n1_port, A(21) => n1_port, A(20) => 
                           n1_port, A(19) => n1_port, A(18) => n1_port, A(17) 
                           => n1_port, A(16) => n1_port, A(15) => n1_port, 
                           A(14) => n1_port, A(13) => n1_port, A(12) => n1_port
                           , A(11) => n1_port, A(10) => n1_port, A(9) => 
                           n1_port, A(8) => n1_port, A(7) => n1_port, A(6) => 
                           n1_port, A(5) => n1_port, A(4) => n1_port, A(3) => 
                           n1_port, A(2) => n8_port, A(1) => n1_port, A(0) => 
                           n1_port, B(31) => IMM_IN(31), B(30) => IMM_IN(30), 
                           B(29) => IMM_IN(29), B(28) => IMM_IN(28), B(27) => 
                           IMM_IN(27), B(26) => IMM_IN(26), B(25) => IMM_IN(25)
                           , B(24) => IMM_IN(24), B(23) => IMM_IN(23), B(22) =>
                           IMM_IN(22), B(21) => IMM_IN(21), B(20) => IMM_IN(20)
                           , B(19) => IMM_IN(19), B(18) => IMM_IN(18), B(17) =>
                           IMM_IN(17), B(16) => IMM_IN(16), B(15) => IMM_IN(15)
                           , B(14) => IMM_IN(14), B(13) => IMM_IN(13), B(12) =>
                           IMM_IN(12), B(11) => IMM_IN(11), B(10) => IMM_IN(10)
                           , B(9) => IMM_IN(9), B(8) => IMM_IN(8), B(7) => 
                           IMM_IN(7), B(6) => IMM_IN(6), B(5) => IMM_IN(5), 
                           B(4) => IMM_IN(4), B(3) => IMM_IN(3), B(2) => 
                           IMM_IN(2), B(1) => IMM_IN(1), B(0) => IMM_IN(0), CI 
                           => n9_port, SUM(31) => N31, SUM(30) => N30, SUM(29) 
                           => N29, SUM(28) => N28, SUM(27) => N27, SUM(26) => 
                           N26, SUM(25) => N25, SUM(24) => N24, SUM(23) => N23,
                           SUM(22) => N22, SUM(21) => N21, SUM(20) => N20, 
                           SUM(19) => N19, SUM(18) => N18, SUM(17) => N17, 
                           SUM(16) => N16, SUM(15) => N15, SUM(14) => N14, 
                           SUM(13) => N13, SUM(12) => N12, SUM(11) => N11, 
                           SUM(10) => N10, SUM(9) => N9, SUM(8) => N8, SUM(7) 
                           => N7_port, SUM(6) => N6, SUM(5) => N5, SUM(4) => N4
                           , SUM(3) => N3, SUM(2) => N2, SUM(1) => N1, SUM(0) 
                           => N0, CO => n_1171);
   add_0_root_add_0_root_add_118_2 : Execute_DW01_add_0 port map( A(31) => 
                           PC_IN(31), A(30) => PC_IN(30), A(29) => PC_IN(29), 
                           A(28) => PC_IN(28), A(27) => PC_IN(27), A(26) => 
                           PC_IN(26), A(25) => PC_IN(25), A(24) => PC_IN(24), 
                           A(23) => PC_IN(23), A(22) => PC_IN(22), A(21) => 
                           PC_IN(21), A(20) => PC_IN(20), A(19) => PC_IN(19), 
                           A(18) => PC_IN(18), A(17) => PC_IN(17), A(16) => 
                           PC_IN(16), A(15) => PC_IN(15), A(14) => PC_IN(14), 
                           A(13) => PC_IN(13), A(12) => PC_IN(12), A(11) => 
                           PC_IN(11), A(10) => PC_IN(10), A(9) => PC_IN(9), 
                           A(8) => PC_IN(8), A(7) => PC_IN(7), A(6) => PC_IN(6)
                           , A(5) => PC_IN(5), A(4) => PC_IN(4), A(3) => 
                           PC_IN(3), A(2) => PC_IN(2), A(1) => PC_IN(1), A(0) 
                           => PC_IN(0), B(31) => N31, B(30) => N30, B(29) => 
                           N29, B(28) => N28, B(27) => N27, B(26) => N26, B(25)
                           => N25, B(24) => N24, B(23) => N23, B(22) => N22, 
                           B(21) => N21, B(20) => N20, B(19) => N19, B(18) => 
                           N18, B(17) => N17, B(16) => N16, B(15) => N15, B(14)
                           => N14, B(13) => N13, B(12) => N12, B(11) => N11, 
                           B(10) => N10, B(9) => N9, B(8) => N8, B(7) => 
                           N7_port, B(6) => N6, B(5) => N5, B(4) => N4, B(3) =>
                           N3, B(2) => N2, B(1) => N1, B(0) => N0, CI => 
                           n10_port, SUM(31) => sig_NPC_REL_31_port, SUM(30) =>
                           sig_NPC_REL_30_port, SUM(29) => sig_NPC_REL_29_port,
                           SUM(28) => sig_NPC_REL_28_port, SUM(27) => 
                           sig_NPC_REL_27_port, SUM(26) => sig_NPC_REL_26_port,
                           SUM(25) => sig_NPC_REL_25_port, SUM(24) => 
                           sig_NPC_REL_24_port, SUM(23) => sig_NPC_REL_23_port,
                           SUM(22) => sig_NPC_REL_22_port, SUM(21) => 
                           sig_NPC_REL_21_port, SUM(20) => sig_NPC_REL_20_port,
                           SUM(19) => sig_NPC_REL_19_port, SUM(18) => 
                           sig_NPC_REL_18_port, SUM(17) => sig_NPC_REL_17_port,
                           SUM(16) => sig_NPC_REL_16_port, SUM(15) => 
                           sig_NPC_REL_15_port, SUM(14) => sig_NPC_REL_14_port,
                           SUM(13) => sig_NPC_REL_13_port, SUM(12) => 
                           sig_NPC_REL_12_port, SUM(11) => sig_NPC_REL_11_port,
                           SUM(10) => sig_NPC_REL_10_port, SUM(9) => 
                           sig_NPC_REL_9_port, SUM(8) => sig_NPC_REL_8_port, 
                           SUM(7) => sig_NPC_REL_7_port, SUM(6) => 
                           sig_NPC_REL_6_port, SUM(5) => sig_NPC_REL_5_port, 
                           SUM(4) => sig_NPC_REL_4_port, SUM(3) => 
                           sig_NPC_REL_3_port, SUM(2) => sig_NPC_REL_2_port, 
                           SUM(1) => sig_NPC_REL_1_port, SUM(0) => 
                           sig_NPC_REL_0_port, CO => n_1172);
   U5 : NOR2_X1 port map( A1 => ZERO_FLAG_port, A2 => n11_port, ZN => sig_RST);
   U6 : INV_X1 port map( A => RST, ZN => n11_port);
   n12_port <= '0';
   n13_port <= '1';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Decode is

   port( CLK, RST, REG_LATCH_EN, RD1, RD2, RF_WE, ZERO_FLAG : in std_logic;  
         PC_IN, INS_IN : in std_logic_vector (31 downto 0);  ADD_WR : in 
         std_logic_vector (4 downto 0);  DATA_WR_IN : in std_logic_vector (31 
         downto 0);  PC_OUT, A_OUT, B_OUT, IMM_OUT : out std_logic_vector (31 
         downto 0);  ADD_RS1_HDU, ADD_RS2_HDU, ADD_WR_OUT, ADD_RS1_OUT, 
         ADD_RS2_OUT : out std_logic_vector (4 downto 0));

end Decode;

architecture SYN_struct of Decode is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component register_file_NBIT_ADD5_NBIT_DATA32
      port( CLK, RST, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RS1, 
            ADD_RS2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component regn_N5_3
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N5_4
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N5_0
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N32_7
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_8
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component instruction_decomposition
      port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype :
            in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : out std_logic_vector (4 
            downto 0);  IMM : out std_logic_vector (31 downto 0));
   end component;
   
   component instruction_type
      port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype :
            out std_logic);
   end component;
   
   signal ADD_RS1_HDU_4_port, ADD_RS1_HDU_3_port, ADD_RS1_HDU_2_port, 
      ADD_RS1_HDU_1_port, ADD_RS1_HDU_0_port, ADD_RS2_HDU_4_port, 
      ADD_RS2_HDU_3_port, ADD_RS2_HDU_2_port, ADD_RS2_HDU_1_port, 
      ADD_RS2_HDU_0_port, sig_RST, sig_Rtype, sig_Itype, sig_Jtype, 
      sig_ADD_WR_4_port, sig_ADD_WR_3_port, sig_ADD_WR_2_port, 
      sig_ADD_WR_1_port, sig_ADD_WR_0_port, sig_IMM_31_port, sig_IMM_30_port, 
      sig_IMM_29_port, sig_IMM_28_port, sig_IMM_27_port, sig_IMM_26_port, 
      sig_IMM_25_port, sig_IMM_24_port, sig_IMM_23_port, sig_IMM_22_port, 
      sig_IMM_21_port, sig_IMM_20_port, sig_IMM_19_port, sig_IMM_18_port, 
      sig_IMM_17_port, sig_IMM_16_port, sig_IMM_15_port, sig_IMM_14_port, 
      sig_IMM_13_port, sig_IMM_12_port, sig_IMM_11_port, sig_IMM_10_port, 
      sig_IMM_9_port, sig_IMM_8_port, sig_IMM_7_port, sig_IMM_6_port, 
      sig_IMM_5_port, sig_IMM_4_port, sig_IMM_3_port, sig_IMM_2_port, 
      sig_IMM_1_port, sig_IMM_0_port, n2, n3 : std_logic;

begin
   ADD_RS1_HDU <= ( ADD_RS1_HDU_4_port, ADD_RS1_HDU_3_port, ADD_RS1_HDU_2_port,
      ADD_RS1_HDU_1_port, ADD_RS1_HDU_0_port );
   ADD_RS2_HDU <= ( ADD_RS2_HDU_4_port, ADD_RS2_HDU_3_port, ADD_RS2_HDU_2_port,
      ADD_RS2_HDU_1_port, ADD_RS2_HDU_0_port );
   
   ins_type : instruction_type port map( INST_IN(31) => INS_IN(31), INST_IN(30)
                           => INS_IN(30), INST_IN(29) => INS_IN(29), 
                           INST_IN(28) => INS_IN(28), INST_IN(27) => INS_IN(27)
                           , INST_IN(26) => INS_IN(26), INST_IN(25) => 
                           INS_IN(25), INST_IN(24) => INS_IN(24), INST_IN(23) 
                           => INS_IN(23), INST_IN(22) => INS_IN(22), 
                           INST_IN(21) => INS_IN(21), INST_IN(20) => INS_IN(20)
                           , INST_IN(19) => INS_IN(19), INST_IN(18) => 
                           INS_IN(18), INST_IN(17) => INS_IN(17), INST_IN(16) 
                           => INS_IN(16), INST_IN(15) => INS_IN(15), 
                           INST_IN(14) => INS_IN(14), INST_IN(13) => INS_IN(13)
                           , INST_IN(12) => INS_IN(12), INST_IN(11) => 
                           INS_IN(11), INST_IN(10) => INS_IN(10), INST_IN(9) =>
                           INS_IN(9), INST_IN(8) => INS_IN(8), INST_IN(7) => 
                           INS_IN(7), INST_IN(6) => INS_IN(6), INST_IN(5) => 
                           INS_IN(5), INST_IN(4) => INS_IN(4), INST_IN(3) => 
                           INS_IN(3), INST_IN(2) => INS_IN(2), INST_IN(1) => 
                           INS_IN(1), INST_IN(0) => INS_IN(0), Rtype => 
                           sig_Rtype, Itype => sig_Itype, Jtype => sig_Jtype);
   ins_dec : instruction_decomposition port map( INST_IN(31) => INS_IN(31), 
                           INST_IN(30) => INS_IN(30), INST_IN(29) => INS_IN(29)
                           , INST_IN(28) => INS_IN(28), INST_IN(27) => 
                           INS_IN(27), INST_IN(26) => INS_IN(26), INST_IN(25) 
                           => INS_IN(25), INST_IN(24) => INS_IN(24), 
                           INST_IN(23) => INS_IN(23), INST_IN(22) => INS_IN(22)
                           , INST_IN(21) => INS_IN(21), INST_IN(20) => 
                           INS_IN(20), INST_IN(19) => INS_IN(19), INST_IN(18) 
                           => INS_IN(18), INST_IN(17) => INS_IN(17), 
                           INST_IN(16) => INS_IN(16), INST_IN(15) => INS_IN(15)
                           , INST_IN(14) => INS_IN(14), INST_IN(13) => 
                           INS_IN(13), INST_IN(12) => INS_IN(12), INST_IN(11) 
                           => INS_IN(11), INST_IN(10) => INS_IN(10), INST_IN(9)
                           => INS_IN(9), INST_IN(8) => INS_IN(8), INST_IN(7) =>
                           INS_IN(7), INST_IN(6) => INS_IN(6), INST_IN(5) => 
                           INS_IN(5), INST_IN(4) => INS_IN(4), INST_IN(3) => 
                           INS_IN(3), INST_IN(2) => INS_IN(2), INST_IN(1) => 
                           INS_IN(1), INST_IN(0) => INS_IN(0), Rtype => 
                           sig_Rtype, Itype => sig_Itype, Jtype => sig_Jtype, 
                           ADD_RS1(4) => ADD_RS1_HDU_4_port, ADD_RS1(3) => 
                           ADD_RS1_HDU_3_port, ADD_RS1(2) => ADD_RS1_HDU_2_port
                           , ADD_RS1(1) => ADD_RS1_HDU_1_port, ADD_RS1(0) => 
                           ADD_RS1_HDU_0_port, ADD_RS2(4) => ADD_RS2_HDU_4_port
                           , ADD_RS2(3) => ADD_RS2_HDU_3_port, ADD_RS2(2) => 
                           ADD_RS2_HDU_2_port, ADD_RS2(1) => ADD_RS2_HDU_1_port
                           , ADD_RS2(0) => ADD_RS2_HDU_0_port, ADD_WR(4) => 
                           sig_ADD_WR_4_port, ADD_WR(3) => sig_ADD_WR_3_port, 
                           ADD_WR(2) => sig_ADD_WR_2_port, ADD_WR(1) => 
                           sig_ADD_WR_1_port, ADD_WR(0) => sig_ADD_WR_0_port, 
                           IMM(31) => sig_IMM_31_port, IMM(30) => 
                           sig_IMM_30_port, IMM(29) => sig_IMM_29_port, IMM(28)
                           => sig_IMM_28_port, IMM(27) => sig_IMM_27_port, 
                           IMM(26) => sig_IMM_26_port, IMM(25) => 
                           sig_IMM_25_port, IMM(24) => sig_IMM_24_port, IMM(23)
                           => sig_IMM_23_port, IMM(22) => sig_IMM_22_port, 
                           IMM(21) => sig_IMM_21_port, IMM(20) => 
                           sig_IMM_20_port, IMM(19) => sig_IMM_19_port, IMM(18)
                           => sig_IMM_18_port, IMM(17) => sig_IMM_17_port, 
                           IMM(16) => sig_IMM_16_port, IMM(15) => 
                           sig_IMM_15_port, IMM(14) => sig_IMM_14_port, IMM(13)
                           => sig_IMM_13_port, IMM(12) => sig_IMM_12_port, 
                           IMM(11) => sig_IMM_11_port, IMM(10) => 
                           sig_IMM_10_port, IMM(9) => sig_IMM_9_port, IMM(8) =>
                           sig_IMM_8_port, IMM(7) => sig_IMM_7_port, IMM(6) => 
                           sig_IMM_6_port, IMM(5) => sig_IMM_5_port, IMM(4) => 
                           sig_IMM_4_port, IMM(3) => sig_IMM_3_port, IMM(2) => 
                           sig_IMM_2_port, IMM(1) => sig_IMM_1_port, IMM(0) => 
                           sig_IMM_0_port);
   regPC : regn_N32_8 port map( DIN(31) => PC_IN(31), DIN(30) => PC_IN(30), 
                           DIN(29) => PC_IN(29), DIN(28) => PC_IN(28), DIN(27) 
                           => PC_IN(27), DIN(26) => PC_IN(26), DIN(25) => 
                           PC_IN(25), DIN(24) => PC_IN(24), DIN(23) => 
                           PC_IN(23), DIN(22) => PC_IN(22), DIN(21) => 
                           PC_IN(21), DIN(20) => PC_IN(20), DIN(19) => 
                           PC_IN(19), DIN(18) => PC_IN(18), DIN(17) => 
                           PC_IN(17), DIN(16) => PC_IN(16), DIN(15) => 
                           PC_IN(15), DIN(14) => PC_IN(14), DIN(13) => 
                           PC_IN(13), DIN(12) => PC_IN(12), DIN(11) => 
                           PC_IN(11), DIN(10) => PC_IN(10), DIN(9) => PC_IN(9),
                           DIN(8) => PC_IN(8), DIN(7) => PC_IN(7), DIN(6) => 
                           PC_IN(6), DIN(5) => PC_IN(5), DIN(4) => PC_IN(4), 
                           DIN(3) => PC_IN(3), DIN(2) => PC_IN(2), DIN(1) => 
                           PC_IN(1), DIN(0) => PC_IN(0), CLK => CLK, EN => n3, 
                           RST => sig_RST, DOUT(31) => PC_OUT(31), DOUT(30) => 
                           PC_OUT(30), DOUT(29) => PC_OUT(29), DOUT(28) => 
                           PC_OUT(28), DOUT(27) => PC_OUT(27), DOUT(26) => 
                           PC_OUT(26), DOUT(25) => PC_OUT(25), DOUT(24) => 
                           PC_OUT(24), DOUT(23) => PC_OUT(23), DOUT(22) => 
                           PC_OUT(22), DOUT(21) => PC_OUT(21), DOUT(20) => 
                           PC_OUT(20), DOUT(19) => PC_OUT(19), DOUT(18) => 
                           PC_OUT(18), DOUT(17) => PC_OUT(17), DOUT(16) => 
                           PC_OUT(16), DOUT(15) => PC_OUT(15), DOUT(14) => 
                           PC_OUT(14), DOUT(13) => PC_OUT(13), DOUT(12) => 
                           PC_OUT(12), DOUT(11) => PC_OUT(11), DOUT(10) => 
                           PC_OUT(10), DOUT(9) => PC_OUT(9), DOUT(8) => 
                           PC_OUT(8), DOUT(7) => PC_OUT(7), DOUT(6) => 
                           PC_OUT(6), DOUT(5) => PC_OUT(5), DOUT(4) => 
                           PC_OUT(4), DOUT(3) => PC_OUT(3), DOUT(2) => 
                           PC_OUT(2), DOUT(1) => PC_OUT(1), DOUT(0) => 
                           PC_OUT(0));
   regIMM : regn_N32_7 port map( DIN(31) => sig_IMM_31_port, DIN(30) => 
                           sig_IMM_30_port, DIN(29) => sig_IMM_29_port, DIN(28)
                           => sig_IMM_28_port, DIN(27) => sig_IMM_27_port, 
                           DIN(26) => sig_IMM_26_port, DIN(25) => 
                           sig_IMM_25_port, DIN(24) => sig_IMM_24_port, DIN(23)
                           => sig_IMM_23_port, DIN(22) => sig_IMM_22_port, 
                           DIN(21) => sig_IMM_21_port, DIN(20) => 
                           sig_IMM_20_port, DIN(19) => sig_IMM_19_port, DIN(18)
                           => sig_IMM_18_port, DIN(17) => sig_IMM_17_port, 
                           DIN(16) => sig_IMM_16_port, DIN(15) => 
                           sig_IMM_15_port, DIN(14) => sig_IMM_14_port, DIN(13)
                           => sig_IMM_13_port, DIN(12) => sig_IMM_12_port, 
                           DIN(11) => sig_IMM_11_port, DIN(10) => 
                           sig_IMM_10_port, DIN(9) => sig_IMM_9_port, DIN(8) =>
                           sig_IMM_8_port, DIN(7) => sig_IMM_7_port, DIN(6) => 
                           sig_IMM_6_port, DIN(5) => sig_IMM_5_port, DIN(4) => 
                           sig_IMM_4_port, DIN(3) => sig_IMM_3_port, DIN(2) => 
                           sig_IMM_2_port, DIN(1) => sig_IMM_1_port, DIN(0) => 
                           sig_IMM_0_port, CLK => CLK, EN => REG_LATCH_EN, RST 
                           => sig_RST, DOUT(31) => IMM_OUT(31), DOUT(30) => 
                           IMM_OUT(30), DOUT(29) => IMM_OUT(29), DOUT(28) => 
                           IMM_OUT(28), DOUT(27) => IMM_OUT(27), DOUT(26) => 
                           IMM_OUT(26), DOUT(25) => IMM_OUT(25), DOUT(24) => 
                           IMM_OUT(24), DOUT(23) => IMM_OUT(23), DOUT(22) => 
                           IMM_OUT(22), DOUT(21) => IMM_OUT(21), DOUT(20) => 
                           IMM_OUT(20), DOUT(19) => IMM_OUT(19), DOUT(18) => 
                           IMM_OUT(18), DOUT(17) => IMM_OUT(17), DOUT(16) => 
                           IMM_OUT(16), DOUT(15) => IMM_OUT(15), DOUT(14) => 
                           IMM_OUT(14), DOUT(13) => IMM_OUT(13), DOUT(12) => 
                           IMM_OUT(12), DOUT(11) => IMM_OUT(11), DOUT(10) => 
                           IMM_OUT(10), DOUT(9) => IMM_OUT(9), DOUT(8) => 
                           IMM_OUT(8), DOUT(7) => IMM_OUT(7), DOUT(6) => 
                           IMM_OUT(6), DOUT(5) => IMM_OUT(5), DOUT(4) => 
                           IMM_OUT(4), DOUT(3) => IMM_OUT(3), DOUT(2) => 
                           IMM_OUT(2), DOUT(1) => IMM_OUT(1), DOUT(0) => 
                           IMM_OUT(0));
   regWR : regn_N5_0 port map( DIN(4) => sig_ADD_WR_4_port, DIN(3) => 
                           sig_ADD_WR_3_port, DIN(2) => sig_ADD_WR_2_port, 
                           DIN(1) => sig_ADD_WR_1_port, DIN(0) => 
                           sig_ADD_WR_0_port, CLK => CLK, EN => REG_LATCH_EN, 
                           RST => sig_RST, DOUT(4) => ADD_WR_OUT(4), DOUT(3) =>
                           ADD_WR_OUT(3), DOUT(2) => ADD_WR_OUT(2), DOUT(1) => 
                           ADD_WR_OUT(1), DOUT(0) => ADD_WR_OUT(0));
   regRS1 : regn_N5_4 port map( DIN(4) => ADD_RS1_HDU_4_port, DIN(3) => 
                           ADD_RS1_HDU_3_port, DIN(2) => ADD_RS1_HDU_2_port, 
                           DIN(1) => ADD_RS1_HDU_1_port, DIN(0) => 
                           ADD_RS1_HDU_0_port, CLK => CLK, EN => REG_LATCH_EN, 
                           RST => sig_RST, DOUT(4) => ADD_RS1_OUT(4), DOUT(3) 
                           => ADD_RS1_OUT(3), DOUT(2) => ADD_RS1_OUT(2), 
                           DOUT(1) => ADD_RS1_OUT(1), DOUT(0) => ADD_RS1_OUT(0)
                           );
   regRS2 : regn_N5_3 port map( DIN(4) => ADD_RS2_HDU_4_port, DIN(3) => 
                           ADD_RS2_HDU_3_port, DIN(2) => ADD_RS2_HDU_2_port, 
                           DIN(1) => ADD_RS2_HDU_1_port, DIN(0) => 
                           ADD_RS2_HDU_0_port, CLK => CLK, EN => REG_LATCH_EN, 
                           RST => sig_RST, DOUT(4) => ADD_RS2_OUT(4), DOUT(3) 
                           => ADD_RS2_OUT(3), DOUT(2) => ADD_RS2_OUT(2), 
                           DOUT(1) => ADD_RS2_OUT(1), DOUT(0) => ADD_RS2_OUT(0)
                           );
   rf : register_file_NBIT_ADD5_NBIT_DATA32 port map( CLK => CLK, RST => RST, 
                           ENABLE => REG_LATCH_EN, RD1 => RD1, RD2 => RD2, WR 
                           => RF_WE, ADD_WR(4) => ADD_WR(4), ADD_WR(3) => 
                           ADD_WR(3), ADD_WR(2) => ADD_WR(2), ADD_WR(1) => 
                           ADD_WR(1), ADD_WR(0) => ADD_WR(0), ADD_RS1(4) => 
                           ADD_RS1_HDU_4_port, ADD_RS1(3) => ADD_RS1_HDU_3_port
                           , ADD_RS1(2) => ADD_RS1_HDU_2_port, ADD_RS1(1) => 
                           ADD_RS1_HDU_1_port, ADD_RS1(0) => ADD_RS1_HDU_0_port
                           , ADD_RS2(4) => ADD_RS2_HDU_4_port, ADD_RS2(3) => 
                           ADD_RS2_HDU_3_port, ADD_RS2(2) => ADD_RS2_HDU_2_port
                           , ADD_RS2(1) => ADD_RS2_HDU_1_port, ADD_RS2(0) => 
                           ADD_RS2_HDU_0_port, DATAIN(31) => DATA_WR_IN(31), 
                           DATAIN(30) => DATA_WR_IN(30), DATAIN(29) => 
                           DATA_WR_IN(29), DATAIN(28) => DATA_WR_IN(28), 
                           DATAIN(27) => DATA_WR_IN(27), DATAIN(26) => 
                           DATA_WR_IN(26), DATAIN(25) => DATA_WR_IN(25), 
                           DATAIN(24) => DATA_WR_IN(24), DATAIN(23) => 
                           DATA_WR_IN(23), DATAIN(22) => DATA_WR_IN(22), 
                           DATAIN(21) => DATA_WR_IN(21), DATAIN(20) => 
                           DATA_WR_IN(20), DATAIN(19) => DATA_WR_IN(19), 
                           DATAIN(18) => DATA_WR_IN(18), DATAIN(17) => 
                           DATA_WR_IN(17), DATAIN(16) => DATA_WR_IN(16), 
                           DATAIN(15) => DATA_WR_IN(15), DATAIN(14) => 
                           DATA_WR_IN(14), DATAIN(13) => DATA_WR_IN(13), 
                           DATAIN(12) => DATA_WR_IN(12), DATAIN(11) => 
                           DATA_WR_IN(11), DATAIN(10) => DATA_WR_IN(10), 
                           DATAIN(9) => DATA_WR_IN(9), DATAIN(8) => 
                           DATA_WR_IN(8), DATAIN(7) => DATA_WR_IN(7), DATAIN(6)
                           => DATA_WR_IN(6), DATAIN(5) => DATA_WR_IN(5), 
                           DATAIN(4) => DATA_WR_IN(4), DATAIN(3) => 
                           DATA_WR_IN(3), DATAIN(2) => DATA_WR_IN(2), DATAIN(1)
                           => DATA_WR_IN(1), DATAIN(0) => DATA_WR_IN(0), 
                           OUT1(31) => A_OUT(31), OUT1(30) => A_OUT(30), 
                           OUT1(29) => A_OUT(29), OUT1(28) => A_OUT(28), 
                           OUT1(27) => A_OUT(27), OUT1(26) => A_OUT(26), 
                           OUT1(25) => A_OUT(25), OUT1(24) => A_OUT(24), 
                           OUT1(23) => A_OUT(23), OUT1(22) => A_OUT(22), 
                           OUT1(21) => A_OUT(21), OUT1(20) => A_OUT(20), 
                           OUT1(19) => A_OUT(19), OUT1(18) => A_OUT(18), 
                           OUT1(17) => A_OUT(17), OUT1(16) => A_OUT(16), 
                           OUT1(15) => A_OUT(15), OUT1(14) => A_OUT(14), 
                           OUT1(13) => A_OUT(13), OUT1(12) => A_OUT(12), 
                           OUT1(11) => A_OUT(11), OUT1(10) => A_OUT(10), 
                           OUT1(9) => A_OUT(9), OUT1(8) => A_OUT(8), OUT1(7) =>
                           A_OUT(7), OUT1(6) => A_OUT(6), OUT1(5) => A_OUT(5), 
                           OUT1(4) => A_OUT(4), OUT1(3) => A_OUT(3), OUT1(2) =>
                           A_OUT(2), OUT1(1) => A_OUT(1), OUT1(0) => A_OUT(0), 
                           OUT2(31) => B_OUT(31), OUT2(30) => B_OUT(30), 
                           OUT2(29) => B_OUT(29), OUT2(28) => B_OUT(28), 
                           OUT2(27) => B_OUT(27), OUT2(26) => B_OUT(26), 
                           OUT2(25) => B_OUT(25), OUT2(24) => B_OUT(24), 
                           OUT2(23) => B_OUT(23), OUT2(22) => B_OUT(22), 
                           OUT2(21) => B_OUT(21), OUT2(20) => B_OUT(20), 
                           OUT2(19) => B_OUT(19), OUT2(18) => B_OUT(18), 
                           OUT2(17) => B_OUT(17), OUT2(16) => B_OUT(16), 
                           OUT2(15) => B_OUT(15), OUT2(14) => B_OUT(14), 
                           OUT2(13) => B_OUT(13), OUT2(12) => B_OUT(12), 
                           OUT2(11) => B_OUT(11), OUT2(10) => B_OUT(10), 
                           OUT2(9) => B_OUT(9), OUT2(8) => B_OUT(8), OUT2(7) =>
                           B_OUT(7), OUT2(6) => B_OUT(6), OUT2(5) => B_OUT(5), 
                           OUT2(4) => B_OUT(4), OUT2(3) => B_OUT(3), OUT2(2) =>
                           B_OUT(2), OUT2(1) => B_OUT(1), OUT2(0) => B_OUT(0));
   U2 : NOR2_X1 port map( A1 => ZERO_FLAG, A2 => n2, ZN => sig_RST);
   U3 : INV_X1 port map( A => RST, ZN => n2);
   n3 <= '1';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Fetch is

   port( CLK, RST, ZERO_FLAG : in std_logic;  PC_EXT, INS_IN : in 
         std_logic_vector (31 downto 0);  Bubble_in : in std_logic;  HDU_INS_IN
         , HDU_PC_IN, HDU_NPC_IN : in std_logic_vector (31 downto 0);  PC_OUT, 
         ADDR_OUT, NPC_OUT, INS_OUT : out std_logic_vector (31 downto 0));

end Fetch;

architecture SYN_struct of Fetch is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component Fetch_DW01_add_3
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component regn_N32_9
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_10
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_0
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   signal ADDR_OUT_31_port, ADDR_OUT_30_port, ADDR_OUT_29_port, 
      ADDR_OUT_28_port, n27, n28, ADDR_OUT_25_port, ADDR_OUT_24_port, n29, n30,
      n31, ADDR_OUT_20_port, n32, n33, n34, n35, n36, n37, n38, 
      ADDR_OUT_12_port, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      ADDR_OUT_1_port, ADDR_OUT_0_port, sig_RST, n4, n5, n6, sig_NPC_9_port, 
      sig_NPC_8_port, sig_NPC_7_port, sig_NPC_6_port, sig_NPC_5_port, 
      sig_NPC_4_port, sig_NPC_3_port, sig_NPC_31_port, sig_NPC_30_port, 
      sig_NPC_2_port, sig_NPC_29_port, sig_NPC_28_port, sig_NPC_27_port, 
      sig_NPC_26_port, sig_NPC_25_port, sig_NPC_24_port, sig_NPC_23_port, 
      sig_NPC_22_port, sig_NPC_21_port, sig_NPC_20_port, sig_NPC_1_port, 
      sig_NPC_19_port, sig_NPC_18_port, sig_NPC_17_port, sig_NPC_16_port, 
      sig_NPC_15_port, sig_NPC_14_port, sig_NPC_13_port, sig_NPC_12_port, 
      sig_NPC_11_port, sig_NPC_10_port, sig_NPC_0_port, sig_INS_9_port, 
      sig_INS_8_port, sig_INS_7_port, sig_INS_6_port, sig_INS_5_port, 
      sig_INS_4_port, sig_INS_3_port, sig_INS_31_port, sig_INS_30_port, 
      sig_INS_2_port, sig_INS_29_port, sig_INS_28_port, sig_INS_27_port, 
      sig_INS_26_port, sig_INS_25_port, sig_INS_24_port, sig_INS_23_port, 
      sig_INS_22_port, sig_INS_21_port, sig_INS_20_port, sig_INS_1_port, 
      sig_INS_19_port, sig_INS_18_port, sig_INS_17_port, sig_INS_16_port, 
      sig_INS_15_port, sig_INS_14_port, sig_INS_13_port, sig_INS_12_port, 
      sig_INS_11_port, sig_INS_10_port, sig_INS_0_port, PC_MUX_OUT_9_port, 
      PC_MUX_OUT_8_port, PC_MUX_OUT_7_port, PC_MUX_OUT_6_port, 
      PC_MUX_OUT_5_port, PC_MUX_OUT_4_port, PC_MUX_OUT_3_port, 
      PC_MUX_OUT_31_port, PC_MUX_OUT_30_port, PC_MUX_OUT_2_port, 
      PC_MUX_OUT_29_port, PC_MUX_OUT_28_port, PC_MUX_OUT_27_port, 
      PC_MUX_OUT_26_port, PC_MUX_OUT_25_port, PC_MUX_OUT_24_port, 
      PC_MUX_OUT_23_port, PC_MUX_OUT_22_port, PC_MUX_OUT_21_port, 
      PC_MUX_OUT_20_port, PC_MUX_OUT_1_port, PC_MUX_OUT_19_port, 
      PC_MUX_OUT_18_port, PC_MUX_OUT_17_port, PC_MUX_OUT_16_port, 
      PC_MUX_OUT_15_port, PC_MUX_OUT_14_port, PC_MUX_OUT_13_port, 
      PC_MUX_OUT_12_port, PC_MUX_OUT_11_port, PC_MUX_OUT_10_port, 
      PC_MUX_OUT_0_port, n49, n50, n_1173 : std_logic;

begin
   ADDR_OUT <= ( ADDR_OUT_31_port, ADDR_OUT_30_port, ADDR_OUT_29_port, 
      ADDR_OUT_28_port, n27, n28, ADDR_OUT_25_port, ADDR_OUT_24_port, n29, n30,
      n31, ADDR_OUT_20_port, n32, n33, n34, n35, n36, n37, n38, 
      ADDR_OUT_12_port, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      ADDR_OUT_1_port, ADDR_OUT_0_port );
   
   n4 <= '0';
   n5 <= '1';
   n6 <= '0';
   NPC_or_NPC_HDU : mux21_NBIT32_0 port map( A(31) => PC_EXT(31), A(30) => 
                           PC_EXT(30), A(29) => PC_EXT(29), A(28) => PC_EXT(28)
                           , A(27) => PC_EXT(27), A(26) => PC_EXT(26), A(25) =>
                           PC_EXT(25), A(24) => PC_EXT(24), A(23) => PC_EXT(23)
                           , A(22) => PC_EXT(22), A(21) => PC_EXT(21), A(20) =>
                           PC_EXT(20), A(19) => PC_EXT(19), A(18) => PC_EXT(18)
                           , A(17) => PC_EXT(17), A(16) => PC_EXT(16), A(15) =>
                           PC_EXT(15), A(14) => PC_EXT(14), A(13) => PC_EXT(13)
                           , A(12) => PC_EXT(12), A(11) => PC_EXT(11), A(10) =>
                           PC_EXT(10), A(9) => PC_EXT(9), A(8) => PC_EXT(8), 
                           A(7) => PC_EXT(7), A(6) => PC_EXT(6), A(5) => 
                           PC_EXT(5), A(4) => PC_EXT(4), A(3) => PC_EXT(3), 
                           A(2) => PC_EXT(2), A(1) => PC_EXT(1), A(0) => 
                           PC_EXT(0), B(31) => HDU_NPC_IN(31), B(30) => 
                           HDU_NPC_IN(30), B(29) => HDU_NPC_IN(29), B(28) => 
                           HDU_NPC_IN(28), B(27) => HDU_NPC_IN(27), B(26) => 
                           HDU_NPC_IN(26), B(25) => HDU_NPC_IN(25), B(24) => 
                           HDU_NPC_IN(24), B(23) => HDU_NPC_IN(23), B(22) => 
                           HDU_NPC_IN(22), B(21) => HDU_NPC_IN(21), B(20) => 
                           HDU_NPC_IN(20), B(19) => HDU_NPC_IN(19), B(18) => 
                           HDU_NPC_IN(18), B(17) => HDU_NPC_IN(17), B(16) => 
                           HDU_NPC_IN(16), B(15) => HDU_NPC_IN(15), B(14) => 
                           HDU_NPC_IN(14), B(13) => HDU_NPC_IN(13), B(12) => 
                           HDU_NPC_IN(12), B(11) => HDU_NPC_IN(11), B(10) => 
                           HDU_NPC_IN(10), B(9) => HDU_NPC_IN(9), B(8) => 
                           HDU_NPC_IN(8), B(7) => HDU_NPC_IN(7), B(6) => 
                           HDU_NPC_IN(6), B(5) => HDU_NPC_IN(5), B(4) => 
                           HDU_NPC_IN(4), B(3) => HDU_NPC_IN(3), B(2) => 
                           HDU_NPC_IN(2), B(1) => HDU_NPC_IN(1), B(0) => 
                           HDU_NPC_IN(0), S => Bubble_in, Z(31) => 
                           sig_NPC_31_port, Z(30) => sig_NPC_30_port, Z(29) => 
                           sig_NPC_29_port, Z(28) => sig_NPC_28_port, Z(27) => 
                           sig_NPC_27_port, Z(26) => sig_NPC_26_port, Z(25) => 
                           sig_NPC_25_port, Z(24) => sig_NPC_24_port, Z(23) => 
                           sig_NPC_23_port, Z(22) => sig_NPC_22_port, Z(21) => 
                           sig_NPC_21_port, Z(20) => sig_NPC_20_port, Z(19) => 
                           sig_NPC_19_port, Z(18) => sig_NPC_18_port, Z(17) => 
                           sig_NPC_17_port, Z(16) => sig_NPC_16_port, Z(15) => 
                           sig_NPC_15_port, Z(14) => sig_NPC_14_port, Z(13) => 
                           sig_NPC_13_port, Z(12) => sig_NPC_12_port, Z(11) => 
                           sig_NPC_11_port, Z(10) => sig_NPC_10_port, Z(9) => 
                           sig_NPC_9_port, Z(8) => sig_NPC_8_port, Z(7) => 
                           sig_NPC_7_port, Z(6) => sig_NPC_6_port, Z(5) => 
                           sig_NPC_5_port, Z(4) => sig_NPC_4_port, Z(3) => 
                           sig_NPC_3_port, Z(2) => sig_NPC_2_port, Z(1) => 
                           sig_NPC_1_port, Z(0) => sig_NPC_0_port);
   PC_or_PC_HDU : mux21_NBIT32_5 port map( A(31) => ADDR_OUT_31_port, A(30) => 
                           ADDR_OUT_30_port, A(29) => ADDR_OUT_29_port, A(28) 
                           => ADDR_OUT_28_port, A(27) => n27, A(26) => n28, 
                           A(25) => ADDR_OUT_25_port, A(24) => ADDR_OUT_24_port
                           , A(23) => n29, A(22) => n30, A(21) => n31, A(20) =>
                           ADDR_OUT_20_port, A(19) => n32, A(18) => n33, A(17) 
                           => n34, A(16) => n35, A(15) => n36, A(14) => n37, 
                           A(13) => n38, A(12) => ADDR_OUT_12_port, A(11) => 
                           n39, A(10) => n40, A(9) => n41, A(8) => n42, A(7) =>
                           n43, A(6) => n44, A(5) => n45, A(4) => n46, A(3) => 
                           n47, A(2) => n48, A(1) => ADDR_OUT_1_port, A(0) => 
                           ADDR_OUT_0_port, B(31) => HDU_PC_IN(31), B(30) => 
                           HDU_PC_IN(30), B(29) => HDU_PC_IN(29), B(28) => 
                           HDU_PC_IN(28), B(27) => HDU_PC_IN(27), B(26) => 
                           HDU_PC_IN(26), B(25) => HDU_PC_IN(25), B(24) => 
                           HDU_PC_IN(24), B(23) => HDU_PC_IN(23), B(22) => 
                           HDU_PC_IN(22), B(21) => HDU_PC_IN(21), B(20) => 
                           HDU_PC_IN(20), B(19) => HDU_PC_IN(19), B(18) => 
                           HDU_PC_IN(18), B(17) => HDU_PC_IN(17), B(16) => 
                           HDU_PC_IN(16), B(15) => HDU_PC_IN(15), B(14) => 
                           HDU_PC_IN(14), B(13) => HDU_PC_IN(13), B(12) => 
                           HDU_PC_IN(12), B(11) => HDU_PC_IN(11), B(10) => 
                           HDU_PC_IN(10), B(9) => HDU_PC_IN(9), B(8) => 
                           HDU_PC_IN(8), B(7) => HDU_PC_IN(7), B(6) => 
                           HDU_PC_IN(6), B(5) => HDU_PC_IN(5), B(4) => 
                           HDU_PC_IN(4), B(3) => HDU_PC_IN(3), B(2) => 
                           HDU_PC_IN(2), B(1) => HDU_PC_IN(1), B(0) => 
                           HDU_PC_IN(0), S => Bubble_in, Z(31) => 
                           PC_MUX_OUT_31_port, Z(30) => PC_MUX_OUT_30_port, 
                           Z(29) => PC_MUX_OUT_29_port, Z(28) => 
                           PC_MUX_OUT_28_port, Z(27) => PC_MUX_OUT_27_port, 
                           Z(26) => PC_MUX_OUT_26_port, Z(25) => 
                           PC_MUX_OUT_25_port, Z(24) => PC_MUX_OUT_24_port, 
                           Z(23) => PC_MUX_OUT_23_port, Z(22) => 
                           PC_MUX_OUT_22_port, Z(21) => PC_MUX_OUT_21_port, 
                           Z(20) => PC_MUX_OUT_20_port, Z(19) => 
                           PC_MUX_OUT_19_port, Z(18) => PC_MUX_OUT_18_port, 
                           Z(17) => PC_MUX_OUT_17_port, Z(16) => 
                           PC_MUX_OUT_16_port, Z(15) => PC_MUX_OUT_15_port, 
                           Z(14) => PC_MUX_OUT_14_port, Z(13) => 
                           PC_MUX_OUT_13_port, Z(12) => PC_MUX_OUT_12_port, 
                           Z(11) => PC_MUX_OUT_11_port, Z(10) => 
                           PC_MUX_OUT_10_port, Z(9) => PC_MUX_OUT_9_port, Z(8) 
                           => PC_MUX_OUT_8_port, Z(7) => PC_MUX_OUT_7_port, 
                           Z(6) => PC_MUX_OUT_6_port, Z(5) => PC_MUX_OUT_5_port
                           , Z(4) => PC_MUX_OUT_4_port, Z(3) => 
                           PC_MUX_OUT_3_port, Z(2) => PC_MUX_OUT_2_port, Z(1) 
                           => PC_MUX_OUT_1_port, Z(0) => PC_MUX_OUT_0_port);
   INS_or_HDU_INS : mux21_NBIT32_4 port map( A(31) => INS_IN(31), A(30) => 
                           INS_IN(30), A(29) => INS_IN(29), A(28) => INS_IN(28)
                           , A(27) => INS_IN(27), A(26) => INS_IN(26), A(25) =>
                           INS_IN(25), A(24) => INS_IN(24), A(23) => INS_IN(23)
                           , A(22) => INS_IN(22), A(21) => INS_IN(21), A(20) =>
                           INS_IN(20), A(19) => INS_IN(19), A(18) => INS_IN(18)
                           , A(17) => INS_IN(17), A(16) => INS_IN(16), A(15) =>
                           INS_IN(15), A(14) => INS_IN(14), A(13) => INS_IN(13)
                           , A(12) => INS_IN(12), A(11) => INS_IN(11), A(10) =>
                           INS_IN(10), A(9) => INS_IN(9), A(8) => INS_IN(8), 
                           A(7) => INS_IN(7), A(6) => INS_IN(6), A(5) => 
                           INS_IN(5), A(4) => INS_IN(4), A(3) => INS_IN(3), 
                           A(2) => INS_IN(2), A(1) => INS_IN(1), A(0) => 
                           INS_IN(0), B(31) => HDU_INS_IN(31), B(30) => 
                           HDU_INS_IN(30), B(29) => HDU_INS_IN(29), B(28) => 
                           HDU_INS_IN(28), B(27) => HDU_INS_IN(27), B(26) => 
                           HDU_INS_IN(26), B(25) => HDU_INS_IN(25), B(24) => 
                           HDU_INS_IN(24), B(23) => HDU_INS_IN(23), B(22) => 
                           HDU_INS_IN(22), B(21) => HDU_INS_IN(21), B(20) => 
                           HDU_INS_IN(20), B(19) => HDU_INS_IN(19), B(18) => 
                           HDU_INS_IN(18), B(17) => HDU_INS_IN(17), B(16) => 
                           HDU_INS_IN(16), B(15) => HDU_INS_IN(15), B(14) => 
                           HDU_INS_IN(14), B(13) => HDU_INS_IN(13), B(12) => 
                           HDU_INS_IN(12), B(11) => HDU_INS_IN(11), B(10) => 
                           HDU_INS_IN(10), B(9) => HDU_INS_IN(9), B(8) => 
                           HDU_INS_IN(8), B(7) => HDU_INS_IN(7), B(6) => 
                           HDU_INS_IN(6), B(5) => HDU_INS_IN(5), B(4) => 
                           HDU_INS_IN(4), B(3) => HDU_INS_IN(3), B(2) => 
                           HDU_INS_IN(2), B(1) => HDU_INS_IN(1), B(0) => 
                           HDU_INS_IN(0), S => Bubble_in, Z(31) => 
                           sig_INS_31_port, Z(30) => sig_INS_30_port, Z(29) => 
                           sig_INS_29_port, Z(28) => sig_INS_28_port, Z(27) => 
                           sig_INS_27_port, Z(26) => sig_INS_26_port, Z(25) => 
                           sig_INS_25_port, Z(24) => sig_INS_24_port, Z(23) => 
                           sig_INS_23_port, Z(22) => sig_INS_22_port, Z(21) => 
                           sig_INS_21_port, Z(20) => sig_INS_20_port, Z(19) => 
                           sig_INS_19_port, Z(18) => sig_INS_18_port, Z(17) => 
                           sig_INS_17_port, Z(16) => sig_INS_16_port, Z(15) => 
                           sig_INS_15_port, Z(14) => sig_INS_14_port, Z(13) => 
                           sig_INS_13_port, Z(12) => sig_INS_12_port, Z(11) => 
                           sig_INS_11_port, Z(10) => sig_INS_10_port, Z(9) => 
                           sig_INS_9_port, Z(8) => sig_INS_8_port, Z(7) => 
                           sig_INS_7_port, Z(6) => sig_INS_6_port, Z(5) => 
                           sig_INS_5_port, Z(4) => sig_INS_4_port, Z(3) => 
                           sig_INS_3_port, Z(2) => sig_INS_2_port, Z(1) => 
                           sig_INS_1_port, Z(0) => sig_INS_0_port);
   PC : regn_N32_0 port map( DIN(31) => sig_NPC_31_port, DIN(30) => 
                           sig_NPC_30_port, DIN(29) => sig_NPC_29_port, DIN(28)
                           => sig_NPC_28_port, DIN(27) => sig_NPC_27_port, 
                           DIN(26) => sig_NPC_26_port, DIN(25) => 
                           sig_NPC_25_port, DIN(24) => sig_NPC_24_port, DIN(23)
                           => sig_NPC_23_port, DIN(22) => sig_NPC_22_port, 
                           DIN(21) => sig_NPC_21_port, DIN(20) => 
                           sig_NPC_20_port, DIN(19) => sig_NPC_19_port, DIN(18)
                           => sig_NPC_18_port, DIN(17) => sig_NPC_17_port, 
                           DIN(16) => sig_NPC_16_port, DIN(15) => 
                           sig_NPC_15_port, DIN(14) => sig_NPC_14_port, DIN(13)
                           => sig_NPC_13_port, DIN(12) => sig_NPC_12_port, 
                           DIN(11) => sig_NPC_11_port, DIN(10) => 
                           sig_NPC_10_port, DIN(9) => sig_NPC_9_port, DIN(8) =>
                           sig_NPC_8_port, DIN(7) => sig_NPC_7_port, DIN(6) => 
                           sig_NPC_6_port, DIN(5) => sig_NPC_5_port, DIN(4) => 
                           sig_NPC_4_port, DIN(3) => sig_NPC_3_port, DIN(2) => 
                           sig_NPC_2_port, DIN(1) => sig_NPC_1_port, DIN(0) => 
                           sig_NPC_0_port, CLK => CLK, EN => n50, RST => RST, 
                           DOUT(31) => ADDR_OUT_31_port, DOUT(30) => 
                           ADDR_OUT_30_port, DOUT(29) => ADDR_OUT_29_port, 
                           DOUT(28) => ADDR_OUT_28_port, DOUT(27) => n27, 
                           DOUT(26) => n28, DOUT(25) => ADDR_OUT_25_port, 
                           DOUT(24) => ADDR_OUT_24_port, DOUT(23) => n29, 
                           DOUT(22) => n30, DOUT(21) => n31, DOUT(20) => 
                           ADDR_OUT_20_port, DOUT(19) => n32, DOUT(18) => n33, 
                           DOUT(17) => n34, DOUT(16) => n35, DOUT(15) => n36, 
                           DOUT(14) => n37, DOUT(13) => n38, DOUT(12) => 
                           ADDR_OUT_12_port, DOUT(11) => n39, DOUT(10) => n40, 
                           DOUT(9) => n41, DOUT(8) => n42, DOUT(7) => n43, 
                           DOUT(6) => n44, DOUT(5) => n45, DOUT(4) => n46, 
                           DOUT(3) => n47, DOUT(2) => n48, DOUT(1) => 
                           ADDR_OUT_1_port, DOUT(0) => ADDR_OUT_0_port);
   PC_reg : regn_N32_10 port map( DIN(31) => PC_MUX_OUT_31_port, DIN(30) => 
                           PC_MUX_OUT_30_port, DIN(29) => PC_MUX_OUT_29_port, 
                           DIN(28) => PC_MUX_OUT_28_port, DIN(27) => 
                           PC_MUX_OUT_27_port, DIN(26) => PC_MUX_OUT_26_port, 
                           DIN(25) => PC_MUX_OUT_25_port, DIN(24) => 
                           PC_MUX_OUT_24_port, DIN(23) => PC_MUX_OUT_23_port, 
                           DIN(22) => PC_MUX_OUT_22_port, DIN(21) => 
                           PC_MUX_OUT_21_port, DIN(20) => PC_MUX_OUT_20_port, 
                           DIN(19) => PC_MUX_OUT_19_port, DIN(18) => 
                           PC_MUX_OUT_18_port, DIN(17) => PC_MUX_OUT_17_port, 
                           DIN(16) => PC_MUX_OUT_16_port, DIN(15) => 
                           PC_MUX_OUT_15_port, DIN(14) => PC_MUX_OUT_14_port, 
                           DIN(13) => PC_MUX_OUT_13_port, DIN(12) => 
                           PC_MUX_OUT_12_port, DIN(11) => PC_MUX_OUT_11_port, 
                           DIN(10) => PC_MUX_OUT_10_port, DIN(9) => 
                           PC_MUX_OUT_9_port, DIN(8) => PC_MUX_OUT_8_port, 
                           DIN(7) => PC_MUX_OUT_7_port, DIN(6) => 
                           PC_MUX_OUT_6_port, DIN(5) => PC_MUX_OUT_5_port, 
                           DIN(4) => PC_MUX_OUT_4_port, DIN(3) => 
                           PC_MUX_OUT_3_port, DIN(2) => PC_MUX_OUT_2_port, 
                           DIN(1) => PC_MUX_OUT_1_port, DIN(0) => 
                           PC_MUX_OUT_0_port, CLK => CLK, EN => n50, RST => 
                           sig_RST, DOUT(31) => PC_OUT(31), DOUT(30) => 
                           PC_OUT(30), DOUT(29) => PC_OUT(29), DOUT(28) => 
                           PC_OUT(28), DOUT(27) => PC_OUT(27), DOUT(26) => 
                           PC_OUT(26), DOUT(25) => PC_OUT(25), DOUT(24) => 
                           PC_OUT(24), DOUT(23) => PC_OUT(23), DOUT(22) => 
                           PC_OUT(22), DOUT(21) => PC_OUT(21), DOUT(20) => 
                           PC_OUT(20), DOUT(19) => PC_OUT(19), DOUT(18) => 
                           PC_OUT(18), DOUT(17) => PC_OUT(17), DOUT(16) => 
                           PC_OUT(16), DOUT(15) => PC_OUT(15), DOUT(14) => 
                           PC_OUT(14), DOUT(13) => PC_OUT(13), DOUT(12) => 
                           PC_OUT(12), DOUT(11) => PC_OUT(11), DOUT(10) => 
                           PC_OUT(10), DOUT(9) => PC_OUT(9), DOUT(8) => 
                           PC_OUT(8), DOUT(7) => PC_OUT(7), DOUT(6) => 
                           PC_OUT(6), DOUT(5) => PC_OUT(5), DOUT(4) => 
                           PC_OUT(4), DOUT(3) => PC_OUT(3), DOUT(2) => 
                           PC_OUT(2), DOUT(1) => PC_OUT(1), DOUT(0) => 
                           PC_OUT(0));
   IR : regn_N32_9 port map( DIN(31) => sig_INS_31_port, DIN(30) => 
                           sig_INS_30_port, DIN(29) => sig_INS_29_port, DIN(28)
                           => sig_INS_28_port, DIN(27) => sig_INS_27_port, 
                           DIN(26) => sig_INS_26_port, DIN(25) => 
                           sig_INS_25_port, DIN(24) => sig_INS_24_port, DIN(23)
                           => sig_INS_23_port, DIN(22) => sig_INS_22_port, 
                           DIN(21) => sig_INS_21_port, DIN(20) => 
                           sig_INS_20_port, DIN(19) => sig_INS_19_port, DIN(18)
                           => sig_INS_18_port, DIN(17) => sig_INS_17_port, 
                           DIN(16) => sig_INS_16_port, DIN(15) => 
                           sig_INS_15_port, DIN(14) => sig_INS_14_port, DIN(13)
                           => sig_INS_13_port, DIN(12) => sig_INS_12_port, 
                           DIN(11) => sig_INS_11_port, DIN(10) => 
                           sig_INS_10_port, DIN(9) => sig_INS_9_port, DIN(8) =>
                           sig_INS_8_port, DIN(7) => sig_INS_7_port, DIN(6) => 
                           sig_INS_6_port, DIN(5) => sig_INS_5_port, DIN(4) => 
                           sig_INS_4_port, DIN(3) => sig_INS_3_port, DIN(2) => 
                           sig_INS_2_port, DIN(1) => sig_INS_1_port, DIN(0) => 
                           sig_INS_0_port, CLK => CLK, EN => n50, RST => 
                           sig_RST, DOUT(31) => INS_OUT(31), DOUT(30) => 
                           INS_OUT(30), DOUT(29) => INS_OUT(29), DOUT(28) => 
                           INS_OUT(28), DOUT(27) => INS_OUT(27), DOUT(26) => 
                           INS_OUT(26), DOUT(25) => INS_OUT(25), DOUT(24) => 
                           INS_OUT(24), DOUT(23) => INS_OUT(23), DOUT(22) => 
                           INS_OUT(22), DOUT(21) => INS_OUT(21), DOUT(20) => 
                           INS_OUT(20), DOUT(19) => INS_OUT(19), DOUT(18) => 
                           INS_OUT(18), DOUT(17) => INS_OUT(17), DOUT(16) => 
                           INS_OUT(16), DOUT(15) => INS_OUT(15), DOUT(14) => 
                           INS_OUT(14), DOUT(13) => INS_OUT(13), DOUT(12) => 
                           INS_OUT(12), DOUT(11) => INS_OUT(11), DOUT(10) => 
                           INS_OUT(10), DOUT(9) => INS_OUT(9), DOUT(8) => 
                           INS_OUT(8), DOUT(7) => INS_OUT(7), DOUT(6) => 
                           INS_OUT(6), DOUT(5) => INS_OUT(5), DOUT(4) => 
                           INS_OUT(4), DOUT(3) => INS_OUT(3), DOUT(2) => 
                           INS_OUT(2), DOUT(1) => INS_OUT(1), DOUT(0) => 
                           INS_OUT(0));
   add_54 : Fetch_DW01_add_3 port map( A(31) => ADDR_OUT_31_port, A(30) => 
                           ADDR_OUT_30_port, A(29) => ADDR_OUT_29_port, A(28) 
                           => ADDR_OUT_28_port, A(27) => n27, A(26) => n28, 
                           A(25) => ADDR_OUT_25_port, A(24) => ADDR_OUT_24_port
                           , A(23) => n29, A(22) => n30, A(21) => n31, A(20) =>
                           ADDR_OUT_20_port, A(19) => n32, A(18) => n33, A(17) 
                           => n34, A(16) => n35, A(15) => n36, A(14) => n37, 
                           A(13) => n38, A(12) => ADDR_OUT_12_port, A(11) => 
                           n39, A(10) => n40, A(9) => n41, A(8) => n42, A(7) =>
                           n43, A(6) => n44, A(5) => n45, A(4) => n46, A(3) => 
                           n47, A(2) => n48, A(1) => ADDR_OUT_1_port, A(0) => 
                           ADDR_OUT_0_port, B(31) => n4, B(30) => n4, B(29) => 
                           n4, B(28) => n4, B(27) => n4, B(26) => n4, B(25) => 
                           n4, B(24) => n4, B(23) => n4, B(22) => n4, B(21) => 
                           n4, B(20) => n4, B(19) => n4, B(18) => n4, B(17) => 
                           n4, B(16) => n4, B(15) => n4, B(14) => n4, B(13) => 
                           n4, B(12) => n4, B(11) => n4, B(10) => n4, B(9) => 
                           n4, B(8) => n4, B(7) => n4, B(6) => n4, B(5) => n4, 
                           B(4) => n4, B(3) => n4, B(2) => n5, B(1) => n4, B(0)
                           => n4, CI => n6, SUM(31) => NPC_OUT(31), SUM(30) => 
                           NPC_OUT(30), SUM(29) => NPC_OUT(29), SUM(28) => 
                           NPC_OUT(28), SUM(27) => NPC_OUT(27), SUM(26) => 
                           NPC_OUT(26), SUM(25) => NPC_OUT(25), SUM(24) => 
                           NPC_OUT(24), SUM(23) => NPC_OUT(23), SUM(22) => 
                           NPC_OUT(22), SUM(21) => NPC_OUT(21), SUM(20) => 
                           NPC_OUT(20), SUM(19) => NPC_OUT(19), SUM(18) => 
                           NPC_OUT(18), SUM(17) => NPC_OUT(17), SUM(16) => 
                           NPC_OUT(16), SUM(15) => NPC_OUT(15), SUM(14) => 
                           NPC_OUT(14), SUM(13) => NPC_OUT(13), SUM(12) => 
                           NPC_OUT(12), SUM(11) => NPC_OUT(11), SUM(10) => 
                           NPC_OUT(10), SUM(9) => NPC_OUT(9), SUM(8) => 
                           NPC_OUT(8), SUM(7) => NPC_OUT(7), SUM(6) => 
                           NPC_OUT(6), SUM(5) => NPC_OUT(5), SUM(4) => 
                           NPC_OUT(4), SUM(3) => NPC_OUT(3), SUM(2) => 
                           NPC_OUT(2), SUM(1) => NPC_OUT(1), SUM(0) => 
                           NPC_OUT(0), CO => n_1173);
   U3 : NOR2_X1 port map( A1 => ZERO_FLAG, A2 => n49, ZN => sig_RST);
   U4 : INV_X1 port map( A => RST, ZN => n49);
   n50 <= '1';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity hardwired_cu_NBIT32 is

   port( REG_LATCH_EN, RD1, RD2, MUX_A_SEL : out std_logic;  MUX_B_SEL : out 
         std_logic_vector (1 downto 0);  ALU_OPC : out std_logic_vector (0 to 
         3);  ALU_OUTREG_EN, DRAM_R_IN : out std_logic;  JUMP_TYPE : out 
         std_logic_vector (1 downto 0);  MEM_EN_IN, DRAM_W_IN, RF_WE, 
         DRAM_EN_IN, WB_MUX_SEL : out std_logic;  INS_IN : in std_logic_vector 
         (31 downto 0);  Bubble, Clk, Rst : in std_logic);

end hardwired_cu_NBIT32;

architecture SYN_bhv of hardwired_cu_NBIT32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal AluOP_E_3_port, AluOP_E_2_port, AluOP_E_1_port, AluOP_E_0_port, N24, 
      N25, N26, N27, n18, n19, n20, n21, n22, n23, n24_port, n25_port, n26_port
      , n27_port, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181 : std_logic;

begin
   
   AluOP_E_reg_3_inst : DFFR_X1 port map( D => N27, CK => Clk, RN => Rst, Q => 
                           AluOP_E_3_port, QN => n_1174);
   ALU_OPC_reg_3_inst : DFFR_X1 port map( D => AluOP_E_3_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(0), QN => n_1175);
   AluOP_E_reg_2_inst : DFFR_X1 port map( D => N26, CK => Clk, RN => Rst, Q => 
                           AluOP_E_2_port, QN => n_1176);
   ALU_OPC_reg_2_inst : DFFR_X1 port map( D => AluOP_E_2_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(1), QN => n_1177);
   AluOP_E_reg_1_inst : DFFR_X1 port map( D => N25, CK => Clk, RN => Rst, Q => 
                           AluOP_E_1_port, QN => n_1178);
   ALU_OPC_reg_1_inst : DFFR_X1 port map( D => AluOP_E_1_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(2), QN => n_1179);
   AluOP_E_reg_0_inst : DFFR_X1 port map( D => N24, CK => Clk, RN => Rst, Q => 
                           AluOP_E_0_port, QN => n_1180);
   ALU_OPC_reg_0_inst : DFFR_X1 port map( D => AluOP_E_0_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(3), QN => n_1181);
   WB_MUX_SEL <= '0';
   DRAM_EN_IN <= '0';
   RF_WE <= '0';
   DRAM_W_IN <= '0';
   MEM_EN_IN <= '0';
   JUMP_TYPE(0) <= '0';
   JUMP_TYPE(1) <= '0';
   DRAM_R_IN <= '0';
   ALU_OUTREG_EN <= '0';
   MUX_B_SEL(0) <= '0';
   MUX_B_SEL(1) <= '0';
   MUX_A_SEL <= '0';
   RD2 <= '0';
   RD1 <= '0';
   REG_LATCH_EN <= '0';
   U73 : XOR2_X1 port map( A => INS_IN(1), B => INS_IN(0), Z => n25_port);
   U74 : NAND3_X1 port map( A1 => n37, A2 => n38, A3 => n61, ZN => n27_port);
   U75 : NAND3_X1 port map( A1 => n39, A2 => INS_IN(30), A3 => n40, ZN => n37);
   U76 : NAND3_X1 port map( A1 => n43, A2 => n26_port, A3 => INS_IN(30), ZN => 
                           n30);
   U77 : NAND3_X1 port map( A1 => n63, A2 => n66, A3 => n24_port, ZN => n31);
   U78 : OAI33_X1 port map( A1 => n53, A2 => n71, A3 => n73, B1 => n54, B2 => 
                           INS_IN(1), B3 => n55, ZN => n20);
   U79 : NAND3_X1 port map( A1 => n43, A2 => n75, A3 => INS_IN(28), ZN => n52);
   U80 : NAND3_X1 port map( A1 => n73, A2 => n75, A3 => n43, ZN => n42);
   U18 : INV_X1 port map( A => n36, ZN => n62);
   U19 : OAI22_X1 port map( A1 => n73, A2 => n30, B1 => n41, B2 => n42, ZN => 
                           n35);
   U20 : AOI21_X1 port map( B1 => n39, B2 => n74, A => n20, ZN => n36);
   U21 : NOR2_X1 port map( A1 => n41, A2 => n52, ZN => n29);
   U22 : INV_X1 port map( A => n40, ZN => n72);
   U23 : INV_X1 port map( A => n30, ZN => n69);
   U24 : INV_X1 port map( A => n52, ZN => n74);
   U25 : INV_X1 port map( A => n39, ZN => n71);
   U26 : INV_X1 port map( A => n26_port, ZN => n67);
   U27 : INV_X1 port map( A => n56, ZN => n61);
   U28 : OAI21_X1 port map( B1 => n65, B2 => n38, A => n57, ZN => n56);
   U29 : OR3_X1 port map( A1 => n72, A2 => n75, A3 => n41, ZN => n57);
   U30 : INV_X1 port map( A => n28, ZN => n68);
   U31 : AOI21_X1 port map( B1 => n73, B2 => n69, A => n29, ZN => n28);
   U32 : NAND2_X1 port map( A1 => INS_IN(5), A2 => INS_IN(3), ZN => n54);
   U33 : NAND2_X1 port map( A1 => INS_IN(30), A2 => n43, ZN => n53);
   U34 : NOR4_X1 port map( A1 => INS_IN(6), A2 => INS_IN(4), A3 => INS_IN(10), 
                           A4 => n59, ZN => n46);
   U35 : OR3_X1 port map( A1 => INS_IN(9), A2 => INS_IN(8), A3 => INS_IN(7), ZN
                           => n59);
   U36 : NOR3_X1 port map( A1 => INS_IN(29), A2 => INS_IN(31), A3 => n73, ZN =>
                           n40);
   U37 : NOR2_X1 port map( A1 => INS_IN(27), A2 => INS_IN(26), ZN => n39);
   U38 : OAI221_X1 port map( B1 => n64, B2 => n31, C1 => Bubble, C2 => n32, A 
                           => n33, ZN => N25);
   U39 : INV_X1 port map( A => n44, ZN => n64);
   U40 : OAI211_X1 port map( C1 => INS_IN(3), C2 => n63, A => n65, B => n34, ZN
                           => n33);
   U41 : NOR3_X1 port map( A1 => n35, A2 => n27_port, A3 => n62, ZN => n32);
   U42 : OAI221_X1 port map( B1 => INS_IN(2), B2 => n19, C1 => Bubble, C2 => 
                           n22, A => n23, ZN => N26);
   U43 : NAND4_X1 port map( A1 => n24_port, A2 => INS_IN(2), A3 => n25_port, A4
                           => n66, ZN => n23);
   U44 : AOI211_X1 port map( C1 => n74, C2 => n26_port, A => n68, B => n27_port
                           , ZN => n22);
   U45 : OAI22_X1 port map( A1 => INS_IN(29), A2 => INS_IN(31), B1 => n76, B2 
                           => INS_IN(30), ZN => n51);
   U46 : NOR2_X1 port map( A1 => n70, A2 => INS_IN(27), ZN => n26_port);
   U47 : NOR3_X1 port map( A1 => n72, A2 => INS_IN(30), A3 => n67, ZN => n49);
   U48 : INV_X1 port map( A => INS_IN(28), ZN => n73);
   U49 : NAND4_X1 port map( A1 => INS_IN(2), A2 => n46, A3 => n47, A4 => n63, 
                           ZN => n55);
   U50 : OAI22_X1 port map( A1 => Bubble, A2 => n45, B1 => n44, B2 => n31, ZN 
                           => N24);
   U51 : NOR4_X1 port map( A1 => n48, A2 => n49, A3 => n29, A4 => n50, ZN => 
                           n45);
   U52 : AND4_X1 port map( A1 => n73, A2 => n51, A3 => INS_IN(26), A4 => 
                           INS_IN(27), ZN => n50);
   U53 : OAI211_X1 port map( C1 => n71, C2 => n42, A => n61, B => n36, ZN => 
                           n48);
   U54 : NOR2_X1 port map( A1 => n65, A2 => INS_IN(2), ZN => n44);
   U55 : NAND4_X1 port map( A1 => INS_IN(0), A2 => n24_port, A3 => INS_IN(3), 
                           A4 => n65, ZN => n19);
   U56 : INV_X1 port map( A => INS_IN(1), ZN => n65);
   U57 : NAND2_X1 port map( A1 => INS_IN(27), A2 => n70, ZN => n41);
   U58 : AND2_X1 port map( A1 => INS_IN(29), A2 => n76, ZN => n43);
   U59 : AND3_X1 port map( A1 => n39, A2 => n73, A3 => n58, ZN => n47);
   U60 : NOR3_X1 port map( A1 => INS_IN(29), A2 => INS_IN(31), A3 => INS_IN(30)
                           , ZN => n58);
   U61 : AND4_X1 port map( A1 => INS_IN(5), A2 => n46, A3 => n47, A4 => n60, ZN
                           => n24_port);
   U62 : INV_X1 port map( A => Bubble, ZN => n60);
   U63 : OAI21_X1 port map( B1 => Bubble, B2 => n18, A => n19, ZN => N27);
   U64 : NOR3_X1 port map( A1 => n20, A2 => n69, A3 => n21, ZN => n18);
   U65 : AOI211_X1 port map( C1 => n71, C2 => n67, A => n72, B => INS_IN(30), 
                           ZN => n21);
   U66 : INV_X1 port map( A => INS_IN(0), ZN => n63);
   U67 : OR3_X1 port map( A1 => INS_IN(3), A2 => INS_IN(5), A3 => n55, ZN => 
                           n38);
   U68 : INV_X1 port map( A => INS_IN(30), ZN => n75);
   U69 : INV_X1 port map( A => INS_IN(26), ZN => n70);
   U70 : INV_X1 port map( A => INS_IN(3), ZN => n66);
   U71 : INV_X1 port map( A => INS_IN(31), ZN => n76);
   U72 : AND2_X1 port map( A1 => INS_IN(2), A2 => n24_port, ZN => n34);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Datapath is

   port( CLK, RST : in std_logic;  INS_IN, DATA_IN : in std_logic_vector (31 
         downto 0);  REG_LATCH_EN, RD1, RD2, MUX_A_SEL : in std_logic;  
         MUX_B_SEL : in std_logic_vector (1 downto 0);  ALU_OPC : in 
         std_logic_vector (0 to 3);  ALU_OUTREG_EN : in std_logic;  JUMP_TYPE :
         in std_logic_vector (1 downto 0);  DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, 
         RF_WE, DRAM_EN_IN, WB_MUX_SEL : in std_logic;  INS_OUT, IRAM_ADDR_OUT,
         DRAM_ADDR_OUT, DATA_OUT : out std_logic_vector (31 downto 0);  
         DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble_out : out std_logic);

end Datapath;

architecture SYN_struct of Datapath is

   component HazardDetection
      port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : in std_logic_vector
            (4 downto 0);  DRAM_R : in std_logic;  INS_IN, PC_IN : in 
            std_logic_vector (31 downto 0);  Bubble : out std_logic;  
            HDU_INS_OUT, HDU_PC_OUT, HDU_NPC_OUT : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Writeback
      port( WB_MUX_SEL : in std_logic;  DATA_IN, ALU_RES_IN : in 
            std_logic_vector (31 downto 0);  ADD_WR_IN : in std_logic_vector (4
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0);  
            ADD_WR_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component ff_2
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Memory
      port( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, DRAM_EN_IN : in 
            std_logic;  PC_SEL : in std_logic_vector (1 downto 0);  NPC_IN, 
            NPC_ABS, NPC_REL, ALU_RES_IN, B_IN : in std_logic_vector (31 downto
            0);  ADD_WR_IN : in std_logic_vector (4 downto 0);  DRAM_DATA_IN : 
            in std_logic_vector (31 downto 0);  PC_OUT : out std_logic_vector 
            (31 downto 0);  DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT : out std_logic
            ;  DRAM_ADDR_OUT, DRAM_DATA_OUT, DATA_OUT, ALU_RES_OUT, OP_MEM : 
            out std_logic_vector (31 downto 0);  ADD_WR_MEM, ADD_WR_OUT : out 
            std_logic_vector (4 downto 0));
   end component;
   
   component ff_0
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Execute
      port( CLK, RST, MUX_A_SEL : in std_logic;  MUX_B_SEL : in 
            std_logic_vector (1 downto 0);  ALU_OPC : in std_logic_vector (0 to
            3);  ALU_OUTREG_EN : in std_logic;  JUMP_TYPE : in std_logic_vector
            (1 downto 0);  PC_IN, A_IN, B_IN, IMM_IN : in std_logic_vector (31 
            downto 0);  ADD_WR_IN, ADD_RS1_IN, ADD_RS2_IN, ADD_WR_MEM, 
            ADD_WR_WB : in std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB 
            : in std_logic;  OP_MEM, OP_WB : in std_logic_vector (31 downto 0);
            PC_SEL : out std_logic_vector (1 downto 0);  ZERO_FLAG : out 
            std_logic;  NPC_ABS, NPC_REL, ALU_RES, B_OUT : out std_logic_vector
            (31 downto 0);  ADD_WR_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component Decode
      port( CLK, RST, REG_LATCH_EN, RD1, RD2, RF_WE, ZERO_FLAG : in std_logic; 
            PC_IN, INS_IN : in std_logic_vector (31 downto 0);  ADD_WR : in 
            std_logic_vector (4 downto 0);  DATA_WR_IN : in std_logic_vector 
            (31 downto 0);  PC_OUT, A_OUT, B_OUT, IMM_OUT : out 
            std_logic_vector (31 downto 0);  ADD_RS1_HDU, ADD_RS2_HDU, 
            ADD_WR_OUT, ADD_RS1_OUT, ADD_RS2_OUT : out std_logic_vector (4 
            downto 0));
   end component;
   
   component Fetch
      port( CLK, RST, ZERO_FLAG : in std_logic;  PC_EXT, INS_IN : in 
            std_logic_vector (31 downto 0);  Bubble_in : in std_logic;  
            HDU_INS_IN, HDU_PC_IN, HDU_NPC_IN : in std_logic_vector (31 downto 
            0);  PC_OUT, ADDR_OUT, NPC_OUT, INS_OUT : out std_logic_vector (31 
            downto 0));
   end component;
   
   signal INS_OUT_31_port, INS_OUT_30_port, INS_OUT_29_port, INS_OUT_28_port, 
      INS_OUT_27_port, INS_OUT_26_port, INS_OUT_25_port, INS_OUT_24_port, 
      INS_OUT_23_port, INS_OUT_22_port, INS_OUT_21_port, INS_OUT_20_port, 
      INS_OUT_19_port, INS_OUT_18_port, INS_OUT_17_port, INS_OUT_16_port, 
      INS_OUT_15_port, INS_OUT_14_port, INS_OUT_13_port, INS_OUT_12_port, 
      INS_OUT_11_port, INS_OUT_10_port, INS_OUT_9_port, INS_OUT_8_port, 
      INS_OUT_7_port, INS_OUT_6_port, INS_OUT_5_port, INS_OUT_4_port, 
      INS_OUT_3_port, INS_OUT_2_port, INS_OUT_1_port, INS_OUT_0_port, 
      Bubble_out_port, ZERO_FLAG_EX, PC_MEM_OUT_31_port, PC_MEM_OUT_30_port, 
      PC_MEM_OUT_29_port, PC_MEM_OUT_28_port, PC_MEM_OUT_27_port, 
      PC_MEM_OUT_26_port, PC_MEM_OUT_25_port, PC_MEM_OUT_24_port, 
      PC_MEM_OUT_23_port, PC_MEM_OUT_22_port, PC_MEM_OUT_21_port, 
      PC_MEM_OUT_20_port, PC_MEM_OUT_19_port, PC_MEM_OUT_18_port, 
      PC_MEM_OUT_17_port, PC_MEM_OUT_16_port, PC_MEM_OUT_15_port, 
      PC_MEM_OUT_14_port, PC_MEM_OUT_13_port, PC_MEM_OUT_12_port, 
      PC_MEM_OUT_11_port, PC_MEM_OUT_10_port, PC_MEM_OUT_9_port, 
      PC_MEM_OUT_8_port, PC_MEM_OUT_7_port, PC_MEM_OUT_6_port, 
      PC_MEM_OUT_5_port, PC_MEM_OUT_4_port, PC_MEM_OUT_3_port, 
      PC_MEM_OUT_2_port, PC_MEM_OUT_1_port, PC_MEM_OUT_0_port, 
      sig_HDU_INS_OUT_31_port, sig_HDU_INS_OUT_30_port, sig_HDU_INS_OUT_29_port
      , sig_HDU_INS_OUT_28_port, sig_HDU_INS_OUT_27_port, 
      sig_HDU_INS_OUT_26_port, sig_HDU_INS_OUT_25_port, sig_HDU_INS_OUT_24_port
      , sig_HDU_INS_OUT_23_port, sig_HDU_INS_OUT_22_port, 
      sig_HDU_INS_OUT_21_port, sig_HDU_INS_OUT_20_port, sig_HDU_INS_OUT_19_port
      , sig_HDU_INS_OUT_18_port, sig_HDU_INS_OUT_17_port, 
      sig_HDU_INS_OUT_16_port, sig_HDU_INS_OUT_15_port, sig_HDU_INS_OUT_14_port
      , sig_HDU_INS_OUT_13_port, sig_HDU_INS_OUT_12_port, 
      sig_HDU_INS_OUT_11_port, sig_HDU_INS_OUT_10_port, sig_HDU_INS_OUT_9_port,
      sig_HDU_INS_OUT_8_port, sig_HDU_INS_OUT_7_port, sig_HDU_INS_OUT_6_port, 
      sig_HDU_INS_OUT_5_port, sig_HDU_INS_OUT_4_port, sig_HDU_INS_OUT_3_port, 
      sig_HDU_INS_OUT_2_port, sig_HDU_INS_OUT_1_port, sig_HDU_INS_OUT_0_port, 
      sig_HDU_PC_OUT_31_port, sig_HDU_PC_OUT_30_port, sig_HDU_PC_OUT_29_port, 
      sig_HDU_PC_OUT_28_port, sig_HDU_PC_OUT_27_port, sig_HDU_PC_OUT_26_port, 
      sig_HDU_PC_OUT_25_port, sig_HDU_PC_OUT_24_port, sig_HDU_PC_OUT_23_port, 
      sig_HDU_PC_OUT_22_port, sig_HDU_PC_OUT_21_port, sig_HDU_PC_OUT_20_port, 
      sig_HDU_PC_OUT_19_port, sig_HDU_PC_OUT_18_port, sig_HDU_PC_OUT_17_port, 
      sig_HDU_PC_OUT_16_port, sig_HDU_PC_OUT_15_port, sig_HDU_PC_OUT_14_port, 
      sig_HDU_PC_OUT_13_port, sig_HDU_PC_OUT_12_port, sig_HDU_PC_OUT_11_port, 
      sig_HDU_PC_OUT_10_port, sig_HDU_PC_OUT_9_port, sig_HDU_PC_OUT_8_port, 
      sig_HDU_PC_OUT_7_port, sig_HDU_PC_OUT_6_port, sig_HDU_PC_OUT_5_port, 
      sig_HDU_PC_OUT_4_port, sig_HDU_PC_OUT_3_port, sig_HDU_PC_OUT_2_port, 
      sig_HDU_PC_OUT_1_port, sig_HDU_PC_OUT_0_port, sig_HDU_NPC_OUT_31_port, 
      sig_HDU_NPC_OUT_30_port, sig_HDU_NPC_OUT_29_port, sig_HDU_NPC_OUT_28_port
      , sig_HDU_NPC_OUT_27_port, sig_HDU_NPC_OUT_26_port, 
      sig_HDU_NPC_OUT_25_port, sig_HDU_NPC_OUT_24_port, sig_HDU_NPC_OUT_23_port
      , sig_HDU_NPC_OUT_22_port, sig_HDU_NPC_OUT_21_port, 
      sig_HDU_NPC_OUT_20_port, sig_HDU_NPC_OUT_19_port, sig_HDU_NPC_OUT_18_port
      , sig_HDU_NPC_OUT_17_port, sig_HDU_NPC_OUT_16_port, 
      sig_HDU_NPC_OUT_15_port, sig_HDU_NPC_OUT_14_port, sig_HDU_NPC_OUT_13_port
      , sig_HDU_NPC_OUT_12_port, sig_HDU_NPC_OUT_11_port, 
      sig_HDU_NPC_OUT_10_port, sig_HDU_NPC_OUT_9_port, sig_HDU_NPC_OUT_8_port, 
      sig_HDU_NPC_OUT_7_port, sig_HDU_NPC_OUT_6_port, sig_HDU_NPC_OUT_5_port, 
      sig_HDU_NPC_OUT_4_port, sig_HDU_NPC_OUT_3_port, sig_HDU_NPC_OUT_2_port, 
      sig_HDU_NPC_OUT_1_port, sig_HDU_NPC_OUT_0_port, PC_FETCH_OUT_31_port, 
      PC_FETCH_OUT_30_port, PC_FETCH_OUT_29_port, PC_FETCH_OUT_28_port, 
      PC_FETCH_OUT_27_port, PC_FETCH_OUT_26_port, PC_FETCH_OUT_25_port, 
      PC_FETCH_OUT_24_port, PC_FETCH_OUT_23_port, PC_FETCH_OUT_22_port, 
      PC_FETCH_OUT_21_port, PC_FETCH_OUT_20_port, PC_FETCH_OUT_19_port, 
      PC_FETCH_OUT_18_port, PC_FETCH_OUT_17_port, PC_FETCH_OUT_16_port, 
      PC_FETCH_OUT_15_port, PC_FETCH_OUT_14_port, PC_FETCH_OUT_13_port, 
      PC_FETCH_OUT_12_port, PC_FETCH_OUT_11_port, PC_FETCH_OUT_10_port, 
      PC_FETCH_OUT_9_port, PC_FETCH_OUT_8_port, PC_FETCH_OUT_7_port, 
      PC_FETCH_OUT_6_port, PC_FETCH_OUT_5_port, PC_FETCH_OUT_4_port, 
      PC_FETCH_OUT_3_port, PC_FETCH_OUT_2_port, PC_FETCH_OUT_1_port, 
      PC_FETCH_OUT_0_port, NPC_FETCH_OUT_31_port, NPC_FETCH_OUT_30_port, 
      NPC_FETCH_OUT_29_port, NPC_FETCH_OUT_28_port, NPC_FETCH_OUT_27_port, 
      NPC_FETCH_OUT_26_port, NPC_FETCH_OUT_25_port, NPC_FETCH_OUT_24_port, 
      NPC_FETCH_OUT_23_port, NPC_FETCH_OUT_22_port, NPC_FETCH_OUT_21_port, 
      NPC_FETCH_OUT_20_port, NPC_FETCH_OUT_19_port, NPC_FETCH_OUT_18_port, 
      NPC_FETCH_OUT_17_port, NPC_FETCH_OUT_16_port, NPC_FETCH_OUT_15_port, 
      NPC_FETCH_OUT_14_port, NPC_FETCH_OUT_13_port, NPC_FETCH_OUT_12_port, 
      NPC_FETCH_OUT_11_port, NPC_FETCH_OUT_10_port, NPC_FETCH_OUT_9_port, 
      NPC_FETCH_OUT_8_port, NPC_FETCH_OUT_7_port, NPC_FETCH_OUT_6_port, 
      NPC_FETCH_OUT_5_port, NPC_FETCH_OUT_4_port, NPC_FETCH_OUT_3_port, 
      NPC_FETCH_OUT_2_port, NPC_FETCH_OUT_1_port, NPC_FETCH_OUT_0_port, 
      RF_WE_WB, ADD_WR_WB_4_port, ADD_WR_WB_3_port, ADD_WR_WB_2_port, 
      ADD_WR_WB_1_port, ADD_WR_WB_0_port, OP_WB_31_port, OP_WB_30_port, 
      OP_WB_29_port, OP_WB_28_port, OP_WB_27_port, OP_WB_26_port, OP_WB_25_port
      , OP_WB_24_port, OP_WB_23_port, OP_WB_22_port, OP_WB_21_port, 
      OP_WB_20_port, OP_WB_19_port, OP_WB_18_port, OP_WB_17_port, OP_WB_16_port
      , OP_WB_15_port, OP_WB_14_port, OP_WB_13_port, OP_WB_12_port, 
      OP_WB_11_port, OP_WB_10_port, OP_WB_9_port, OP_WB_8_port, OP_WB_7_port, 
      OP_WB_6_port, OP_WB_5_port, OP_WB_4_port, OP_WB_3_port, OP_WB_2_port, 
      OP_WB_1_port, OP_WB_0_port, PC_DECODE_OUT_31_port, PC_DECODE_OUT_30_port,
      PC_DECODE_OUT_29_port, PC_DECODE_OUT_28_port, PC_DECODE_OUT_27_port, 
      PC_DECODE_OUT_26_port, PC_DECODE_OUT_25_port, PC_DECODE_OUT_24_port, 
      PC_DECODE_OUT_23_port, PC_DECODE_OUT_22_port, PC_DECODE_OUT_21_port, 
      PC_DECODE_OUT_20_port, PC_DECODE_OUT_19_port, PC_DECODE_OUT_18_port, 
      PC_DECODE_OUT_17_port, PC_DECODE_OUT_16_port, PC_DECODE_OUT_15_port, 
      PC_DECODE_OUT_14_port, PC_DECODE_OUT_13_port, PC_DECODE_OUT_12_port, 
      PC_DECODE_OUT_11_port, PC_DECODE_OUT_10_port, PC_DECODE_OUT_9_port, 
      PC_DECODE_OUT_8_port, PC_DECODE_OUT_7_port, PC_DECODE_OUT_6_port, 
      PC_DECODE_OUT_5_port, PC_DECODE_OUT_4_port, PC_DECODE_OUT_3_port, 
      PC_DECODE_OUT_2_port, PC_DECODE_OUT_1_port, PC_DECODE_OUT_0_port, 
      A_DECODE_OUT_31_port, A_DECODE_OUT_30_port, A_DECODE_OUT_29_port, 
      A_DECODE_OUT_28_port, A_DECODE_OUT_27_port, A_DECODE_OUT_26_port, 
      A_DECODE_OUT_25_port, A_DECODE_OUT_24_port, A_DECODE_OUT_23_port, 
      A_DECODE_OUT_22_port, A_DECODE_OUT_21_port, A_DECODE_OUT_20_port, 
      A_DECODE_OUT_19_port, A_DECODE_OUT_18_port, A_DECODE_OUT_17_port, 
      A_DECODE_OUT_16_port, A_DECODE_OUT_15_port, A_DECODE_OUT_14_port, 
      A_DECODE_OUT_13_port, A_DECODE_OUT_12_port, A_DECODE_OUT_11_port, 
      A_DECODE_OUT_10_port, A_DECODE_OUT_9_port, A_DECODE_OUT_8_port, 
      A_DECODE_OUT_7_port, A_DECODE_OUT_6_port, A_DECODE_OUT_5_port, 
      A_DECODE_OUT_4_port, A_DECODE_OUT_3_port, A_DECODE_OUT_2_port, 
      A_DECODE_OUT_1_port, A_DECODE_OUT_0_port, B_DECODE_OUT_31_port, 
      B_DECODE_OUT_30_port, B_DECODE_OUT_29_port, B_DECODE_OUT_28_port, 
      B_DECODE_OUT_27_port, B_DECODE_OUT_26_port, B_DECODE_OUT_25_port, 
      B_DECODE_OUT_24_port, B_DECODE_OUT_23_port, B_DECODE_OUT_22_port, 
      B_DECODE_OUT_21_port, B_DECODE_OUT_20_port, B_DECODE_OUT_19_port, 
      B_DECODE_OUT_18_port, B_DECODE_OUT_17_port, B_DECODE_OUT_16_port, 
      B_DECODE_OUT_15_port, B_DECODE_OUT_14_port, B_DECODE_OUT_13_port, 
      B_DECODE_OUT_12_port, B_DECODE_OUT_11_port, B_DECODE_OUT_10_port, 
      B_DECODE_OUT_9_port, B_DECODE_OUT_8_port, B_DECODE_OUT_7_port, 
      B_DECODE_OUT_6_port, B_DECODE_OUT_5_port, B_DECODE_OUT_4_port, 
      B_DECODE_OUT_3_port, B_DECODE_OUT_2_port, B_DECODE_OUT_1_port, 
      B_DECODE_OUT_0_port, IMM_DECODE_OUT_31_port, IMM_DECODE_OUT_30_port, 
      IMM_DECODE_OUT_29_port, IMM_DECODE_OUT_28_port, IMM_DECODE_OUT_27_port, 
      IMM_DECODE_OUT_26_port, IMM_DECODE_OUT_25_port, IMM_DECODE_OUT_24_port, 
      IMM_DECODE_OUT_23_port, IMM_DECODE_OUT_22_port, IMM_DECODE_OUT_21_port, 
      IMM_DECODE_OUT_20_port, IMM_DECODE_OUT_19_port, IMM_DECODE_OUT_18_port, 
      IMM_DECODE_OUT_17_port, IMM_DECODE_OUT_16_port, IMM_DECODE_OUT_15_port, 
      IMM_DECODE_OUT_14_port, IMM_DECODE_OUT_13_port, IMM_DECODE_OUT_12_port, 
      IMM_DECODE_OUT_11_port, IMM_DECODE_OUT_10_port, IMM_DECODE_OUT_9_port, 
      IMM_DECODE_OUT_8_port, IMM_DECODE_OUT_7_port, IMM_DECODE_OUT_6_port, 
      IMM_DECODE_OUT_5_port, IMM_DECODE_OUT_4_port, IMM_DECODE_OUT_3_port, 
      IMM_DECODE_OUT_2_port, IMM_DECODE_OUT_1_port, IMM_DECODE_OUT_0_port, 
      ADD_RS1_HDU_4_port, ADD_RS1_HDU_3_port, ADD_RS1_HDU_2_port, 
      ADD_RS1_HDU_1_port, ADD_RS1_HDU_0_port, ADD_RS2_HDU_4_port, 
      ADD_RS2_HDU_3_port, ADD_RS2_HDU_2_port, ADD_RS2_HDU_1_port, 
      ADD_RS2_HDU_0_port, ADD_WR_DECODE_OUT_4_port, ADD_WR_DECODE_OUT_3_port, 
      ADD_WR_DECODE_OUT_2_port, ADD_WR_DECODE_OUT_1_port, 
      ADD_WR_DECODE_OUT_0_port, ADD_RS1_DECODE_OUT_4_port, 
      ADD_RS1_DECODE_OUT_3_port, ADD_RS1_DECODE_OUT_2_port, 
      ADD_RS1_DECODE_OUT_1_port, ADD_RS1_DECODE_OUT_0_port, 
      ADD_RS2_DECODE_OUT_4_port, ADD_RS2_DECODE_OUT_3_port, 
      ADD_RS2_DECODE_OUT_2_port, ADD_RS2_DECODE_OUT_1_port, 
      ADD_RS2_DECODE_OUT_0_port, ADD_WR_MEM_4_port, ADD_WR_MEM_3_port, 
      ADD_WR_MEM_2_port, ADD_WR_MEM_1_port, ADD_WR_MEM_0_port, OP_MEM_31_port, 
      OP_MEM_30_port, OP_MEM_29_port, OP_MEM_28_port, OP_MEM_27_port, 
      OP_MEM_26_port, OP_MEM_25_port, OP_MEM_24_port, OP_MEM_23_port, 
      OP_MEM_22_port, OP_MEM_21_port, OP_MEM_20_port, OP_MEM_19_port, 
      OP_MEM_18_port, OP_MEM_17_port, OP_MEM_16_port, OP_MEM_15_port, 
      OP_MEM_14_port, OP_MEM_13_port, OP_MEM_12_port, OP_MEM_11_port, 
      OP_MEM_10_port, OP_MEM_9_port, OP_MEM_8_port, OP_MEM_7_port, 
      OP_MEM_6_port, OP_MEM_5_port, OP_MEM_4_port, OP_MEM_3_port, OP_MEM_2_port
      , OP_MEM_1_port, OP_MEM_0_port, PC_SEL_EX_1_port, PC_SEL_EX_0_port, 
      NPC_ABS_EX_31_port, NPC_ABS_EX_30_port, NPC_ABS_EX_29_port, 
      NPC_ABS_EX_28_port, NPC_ABS_EX_27_port, NPC_ABS_EX_26_port, 
      NPC_ABS_EX_25_port, NPC_ABS_EX_24_port, NPC_ABS_EX_23_port, 
      NPC_ABS_EX_22_port, NPC_ABS_EX_21_port, NPC_ABS_EX_20_port, 
      NPC_ABS_EX_19_port, NPC_ABS_EX_18_port, NPC_ABS_EX_17_port, 
      NPC_ABS_EX_16_port, NPC_ABS_EX_15_port, NPC_ABS_EX_14_port, 
      NPC_ABS_EX_13_port, NPC_ABS_EX_12_port, NPC_ABS_EX_11_port, 
      NPC_ABS_EX_10_port, NPC_ABS_EX_9_port, NPC_ABS_EX_8_port, 
      NPC_ABS_EX_7_port, NPC_ABS_EX_6_port, NPC_ABS_EX_5_port, 
      NPC_ABS_EX_4_port, NPC_ABS_EX_3_port, NPC_ABS_EX_2_port, 
      NPC_ABS_EX_1_port, NPC_ABS_EX_0_port, NPC_REL_EX_31_port, 
      NPC_REL_EX_30_port, NPC_REL_EX_29_port, NPC_REL_EX_28_port, 
      NPC_REL_EX_27_port, NPC_REL_EX_26_port, NPC_REL_EX_25_port, 
      NPC_REL_EX_24_port, NPC_REL_EX_23_port, NPC_REL_EX_22_port, 
      NPC_REL_EX_21_port, NPC_REL_EX_20_port, NPC_REL_EX_19_port, 
      NPC_REL_EX_18_port, NPC_REL_EX_17_port, NPC_REL_EX_16_port, 
      NPC_REL_EX_15_port, NPC_REL_EX_14_port, NPC_REL_EX_13_port, 
      NPC_REL_EX_12_port, NPC_REL_EX_11_port, NPC_REL_EX_10_port, 
      NPC_REL_EX_9_port, NPC_REL_EX_8_port, NPC_REL_EX_7_port, 
      NPC_REL_EX_6_port, NPC_REL_EX_5_port, NPC_REL_EX_4_port, 
      NPC_REL_EX_3_port, NPC_REL_EX_2_port, NPC_REL_EX_1_port, 
      NPC_REL_EX_0_port, ALU_RES_EX_31_port, ALU_RES_EX_30_port, 
      ALU_RES_EX_29_port, ALU_RES_EX_28_port, ALU_RES_EX_27_port, 
      ALU_RES_EX_26_port, ALU_RES_EX_25_port, ALU_RES_EX_24_port, 
      ALU_RES_EX_23_port, ALU_RES_EX_22_port, ALU_RES_EX_21_port, 
      ALU_RES_EX_20_port, ALU_RES_EX_19_port, ALU_RES_EX_18_port, 
      ALU_RES_EX_17_port, ALU_RES_EX_16_port, ALU_RES_EX_15_port, 
      ALU_RES_EX_14_port, ALU_RES_EX_13_port, ALU_RES_EX_12_port, 
      ALU_RES_EX_11_port, ALU_RES_EX_10_port, ALU_RES_EX_9_port, 
      ALU_RES_EX_8_port, ALU_RES_EX_7_port, ALU_RES_EX_6_port, 
      ALU_RES_EX_5_port, ALU_RES_EX_4_port, ALU_RES_EX_3_port, 
      ALU_RES_EX_2_port, ALU_RES_EX_1_port, ALU_RES_EX_0_port, B_EX_OUT_31_port
      , B_EX_OUT_30_port, B_EX_OUT_29_port, B_EX_OUT_28_port, B_EX_OUT_27_port,
      B_EX_OUT_26_port, B_EX_OUT_25_port, B_EX_OUT_24_port, B_EX_OUT_23_port, 
      B_EX_OUT_22_port, B_EX_OUT_21_port, B_EX_OUT_20_port, B_EX_OUT_19_port, 
      B_EX_OUT_18_port, B_EX_OUT_17_port, B_EX_OUT_16_port, B_EX_OUT_15_port, 
      B_EX_OUT_14_port, B_EX_OUT_13_port, B_EX_OUT_12_port, B_EX_OUT_11_port, 
      B_EX_OUT_10_port, B_EX_OUT_9_port, B_EX_OUT_8_port, B_EX_OUT_7_port, 
      B_EX_OUT_6_port, B_EX_OUT_5_port, B_EX_OUT_4_port, B_EX_OUT_3_port, 
      B_EX_OUT_2_port, B_EX_OUT_1_port, B_EX_OUT_0_port, ADD_WR_EX_OUT_4_port, 
      ADD_WR_EX_OUT_3_port, ADD_WR_EX_OUT_2_port, ADD_WR_EX_OUT_1_port, 
      ADD_WR_EX_OUT_0_port, DRAM_R_MEM, DATA_MEM_OUT_31_port, 
      DATA_MEM_OUT_30_port, DATA_MEM_OUT_29_port, DATA_MEM_OUT_28_port, 
      DATA_MEM_OUT_27_port, DATA_MEM_OUT_26_port, DATA_MEM_OUT_25_port, 
      DATA_MEM_OUT_24_port, DATA_MEM_OUT_23_port, DATA_MEM_OUT_22_port, 
      DATA_MEM_OUT_21_port, DATA_MEM_OUT_20_port, DATA_MEM_OUT_19_port, 
      DATA_MEM_OUT_18_port, DATA_MEM_OUT_17_port, DATA_MEM_OUT_16_port, 
      DATA_MEM_OUT_15_port, DATA_MEM_OUT_14_port, DATA_MEM_OUT_13_port, 
      DATA_MEM_OUT_12_port, DATA_MEM_OUT_11_port, DATA_MEM_OUT_10_port, 
      DATA_MEM_OUT_9_port, DATA_MEM_OUT_8_port, DATA_MEM_OUT_7_port, 
      DATA_MEM_OUT_6_port, DATA_MEM_OUT_5_port, DATA_MEM_OUT_4_port, 
      DATA_MEM_OUT_3_port, DATA_MEM_OUT_2_port, DATA_MEM_OUT_1_port, 
      DATA_MEM_OUT_0_port, ALU_RES_MEM_31_port, ALU_RES_MEM_30_port, 
      ALU_RES_MEM_29_port, ALU_RES_MEM_28_port, ALU_RES_MEM_27_port, 
      ALU_RES_MEM_26_port, ALU_RES_MEM_25_port, ALU_RES_MEM_24_port, 
      ALU_RES_MEM_23_port, ALU_RES_MEM_22_port, ALU_RES_MEM_21_port, 
      ALU_RES_MEM_20_port, ALU_RES_MEM_19_port, ALU_RES_MEM_18_port, 
      ALU_RES_MEM_17_port, ALU_RES_MEM_16_port, ALU_RES_MEM_15_port, 
      ALU_RES_MEM_14_port, ALU_RES_MEM_13_port, ALU_RES_MEM_12_port, 
      ALU_RES_MEM_11_port, ALU_RES_MEM_10_port, ALU_RES_MEM_9_port, 
      ALU_RES_MEM_8_port, ALU_RES_MEM_7_port, ALU_RES_MEM_6_port, 
      ALU_RES_MEM_5_port, ALU_RES_MEM_4_port, ALU_RES_MEM_3_port, 
      ALU_RES_MEM_2_port, ALU_RES_MEM_1_port, ALU_RES_MEM_0_port, 
      ADD_WR_MEM_OUT_4_port, ADD_WR_MEM_OUT_3_port, ADD_WR_MEM_OUT_2_port, 
      ADD_WR_MEM_OUT_1_port, ADD_WR_MEM_OUT_0_port, n1 : std_logic;

begin
   INS_OUT <= ( INS_OUT_31_port, INS_OUT_30_port, INS_OUT_29_port, 
      INS_OUT_28_port, INS_OUT_27_port, INS_OUT_26_port, INS_OUT_25_port, 
      INS_OUT_24_port, INS_OUT_23_port, INS_OUT_22_port, INS_OUT_21_port, 
      INS_OUT_20_port, INS_OUT_19_port, INS_OUT_18_port, INS_OUT_17_port, 
      INS_OUT_16_port, INS_OUT_15_port, INS_OUT_14_port, INS_OUT_13_port, 
      INS_OUT_12_port, INS_OUT_11_port, INS_OUT_10_port, INS_OUT_9_port, 
      INS_OUT_8_port, INS_OUT_7_port, INS_OUT_6_port, INS_OUT_5_port, 
      INS_OUT_4_port, INS_OUT_3_port, INS_OUT_2_port, INS_OUT_1_port, 
      INS_OUT_0_port );
   Bubble_out <= Bubble_out_port;
   
   FetchStage : Fetch port map( CLK => CLK, RST => RST, ZERO_FLAG => 
                           ZERO_FLAG_EX, PC_EXT(31) => PC_MEM_OUT_31_port, 
                           PC_EXT(30) => PC_MEM_OUT_30_port, PC_EXT(29) => 
                           PC_MEM_OUT_29_port, PC_EXT(28) => PC_MEM_OUT_28_port
                           , PC_EXT(27) => PC_MEM_OUT_27_port, PC_EXT(26) => 
                           PC_MEM_OUT_26_port, PC_EXT(25) => PC_MEM_OUT_25_port
                           , PC_EXT(24) => PC_MEM_OUT_24_port, PC_EXT(23) => 
                           PC_MEM_OUT_23_port, PC_EXT(22) => PC_MEM_OUT_22_port
                           , PC_EXT(21) => PC_MEM_OUT_21_port, PC_EXT(20) => 
                           PC_MEM_OUT_20_port, PC_EXT(19) => PC_MEM_OUT_19_port
                           , PC_EXT(18) => PC_MEM_OUT_18_port, PC_EXT(17) => 
                           PC_MEM_OUT_17_port, PC_EXT(16) => PC_MEM_OUT_16_port
                           , PC_EXT(15) => PC_MEM_OUT_15_port, PC_EXT(14) => 
                           PC_MEM_OUT_14_port, PC_EXT(13) => PC_MEM_OUT_13_port
                           , PC_EXT(12) => PC_MEM_OUT_12_port, PC_EXT(11) => 
                           PC_MEM_OUT_11_port, PC_EXT(10) => PC_MEM_OUT_10_port
                           , PC_EXT(9) => PC_MEM_OUT_9_port, PC_EXT(8) => 
                           PC_MEM_OUT_8_port, PC_EXT(7) => PC_MEM_OUT_7_port, 
                           PC_EXT(6) => PC_MEM_OUT_6_port, PC_EXT(5) => 
                           PC_MEM_OUT_5_port, PC_EXT(4) => PC_MEM_OUT_4_port, 
                           PC_EXT(3) => PC_MEM_OUT_3_port, PC_EXT(2) => 
                           PC_MEM_OUT_2_port, PC_EXT(1) => PC_MEM_OUT_1_port, 
                           PC_EXT(0) => PC_MEM_OUT_0_port, INS_IN(31) => 
                           INS_IN(31), INS_IN(30) => INS_IN(30), INS_IN(29) => 
                           INS_IN(29), INS_IN(28) => INS_IN(28), INS_IN(27) => 
                           INS_IN(27), INS_IN(26) => INS_IN(26), INS_IN(25) => 
                           INS_IN(25), INS_IN(24) => INS_IN(24), INS_IN(23) => 
                           INS_IN(23), INS_IN(22) => INS_IN(22), INS_IN(21) => 
                           INS_IN(21), INS_IN(20) => INS_IN(20), INS_IN(19) => 
                           INS_IN(19), INS_IN(18) => INS_IN(18), INS_IN(17) => 
                           INS_IN(17), INS_IN(16) => INS_IN(16), INS_IN(15) => 
                           INS_IN(15), INS_IN(14) => INS_IN(14), INS_IN(13) => 
                           INS_IN(13), INS_IN(12) => INS_IN(12), INS_IN(11) => 
                           INS_IN(11), INS_IN(10) => INS_IN(10), INS_IN(9) => 
                           INS_IN(9), INS_IN(8) => INS_IN(8), INS_IN(7) => 
                           INS_IN(7), INS_IN(6) => INS_IN(6), INS_IN(5) => 
                           INS_IN(5), INS_IN(4) => INS_IN(4), INS_IN(3) => 
                           INS_IN(3), INS_IN(2) => INS_IN(2), INS_IN(1) => 
                           INS_IN(1), INS_IN(0) => INS_IN(0), Bubble_in => 
                           Bubble_out_port, HDU_INS_IN(31) => 
                           sig_HDU_INS_OUT_31_port, HDU_INS_IN(30) => 
                           sig_HDU_INS_OUT_30_port, HDU_INS_IN(29) => 
                           sig_HDU_INS_OUT_29_port, HDU_INS_IN(28) => 
                           sig_HDU_INS_OUT_28_port, HDU_INS_IN(27) => 
                           sig_HDU_INS_OUT_27_port, HDU_INS_IN(26) => 
                           sig_HDU_INS_OUT_26_port, HDU_INS_IN(25) => 
                           sig_HDU_INS_OUT_25_port, HDU_INS_IN(24) => 
                           sig_HDU_INS_OUT_24_port, HDU_INS_IN(23) => 
                           sig_HDU_INS_OUT_23_port, HDU_INS_IN(22) => 
                           sig_HDU_INS_OUT_22_port, HDU_INS_IN(21) => 
                           sig_HDU_INS_OUT_21_port, HDU_INS_IN(20) => 
                           sig_HDU_INS_OUT_20_port, HDU_INS_IN(19) => 
                           sig_HDU_INS_OUT_19_port, HDU_INS_IN(18) => 
                           sig_HDU_INS_OUT_18_port, HDU_INS_IN(17) => 
                           sig_HDU_INS_OUT_17_port, HDU_INS_IN(16) => 
                           sig_HDU_INS_OUT_16_port, HDU_INS_IN(15) => 
                           sig_HDU_INS_OUT_15_port, HDU_INS_IN(14) => 
                           sig_HDU_INS_OUT_14_port, HDU_INS_IN(13) => 
                           sig_HDU_INS_OUT_13_port, HDU_INS_IN(12) => 
                           sig_HDU_INS_OUT_12_port, HDU_INS_IN(11) => 
                           sig_HDU_INS_OUT_11_port, HDU_INS_IN(10) => 
                           sig_HDU_INS_OUT_10_port, HDU_INS_IN(9) => 
                           sig_HDU_INS_OUT_9_port, HDU_INS_IN(8) => 
                           sig_HDU_INS_OUT_8_port, HDU_INS_IN(7) => 
                           sig_HDU_INS_OUT_7_port, HDU_INS_IN(6) => 
                           sig_HDU_INS_OUT_6_port, HDU_INS_IN(5) => 
                           sig_HDU_INS_OUT_5_port, HDU_INS_IN(4) => 
                           sig_HDU_INS_OUT_4_port, HDU_INS_IN(3) => 
                           sig_HDU_INS_OUT_3_port, HDU_INS_IN(2) => 
                           sig_HDU_INS_OUT_2_port, HDU_INS_IN(1) => 
                           sig_HDU_INS_OUT_1_port, HDU_INS_IN(0) => 
                           sig_HDU_INS_OUT_0_port, HDU_PC_IN(31) => 
                           sig_HDU_PC_OUT_31_port, HDU_PC_IN(30) => 
                           sig_HDU_PC_OUT_30_port, HDU_PC_IN(29) => 
                           sig_HDU_PC_OUT_29_port, HDU_PC_IN(28) => 
                           sig_HDU_PC_OUT_28_port, HDU_PC_IN(27) => 
                           sig_HDU_PC_OUT_27_port, HDU_PC_IN(26) => 
                           sig_HDU_PC_OUT_26_port, HDU_PC_IN(25) => 
                           sig_HDU_PC_OUT_25_port, HDU_PC_IN(24) => 
                           sig_HDU_PC_OUT_24_port, HDU_PC_IN(23) => 
                           sig_HDU_PC_OUT_23_port, HDU_PC_IN(22) => 
                           sig_HDU_PC_OUT_22_port, HDU_PC_IN(21) => 
                           sig_HDU_PC_OUT_21_port, HDU_PC_IN(20) => 
                           sig_HDU_PC_OUT_20_port, HDU_PC_IN(19) => 
                           sig_HDU_PC_OUT_19_port, HDU_PC_IN(18) => 
                           sig_HDU_PC_OUT_18_port, HDU_PC_IN(17) => 
                           sig_HDU_PC_OUT_17_port, HDU_PC_IN(16) => 
                           sig_HDU_PC_OUT_16_port, HDU_PC_IN(15) => 
                           sig_HDU_PC_OUT_15_port, HDU_PC_IN(14) => 
                           sig_HDU_PC_OUT_14_port, HDU_PC_IN(13) => 
                           sig_HDU_PC_OUT_13_port, HDU_PC_IN(12) => 
                           sig_HDU_PC_OUT_12_port, HDU_PC_IN(11) => 
                           sig_HDU_PC_OUT_11_port, HDU_PC_IN(10) => 
                           sig_HDU_PC_OUT_10_port, HDU_PC_IN(9) => 
                           sig_HDU_PC_OUT_9_port, HDU_PC_IN(8) => 
                           sig_HDU_PC_OUT_8_port, HDU_PC_IN(7) => 
                           sig_HDU_PC_OUT_7_port, HDU_PC_IN(6) => 
                           sig_HDU_PC_OUT_6_port, HDU_PC_IN(5) => 
                           sig_HDU_PC_OUT_5_port, HDU_PC_IN(4) => 
                           sig_HDU_PC_OUT_4_port, HDU_PC_IN(3) => 
                           sig_HDU_PC_OUT_3_port, HDU_PC_IN(2) => 
                           sig_HDU_PC_OUT_2_port, HDU_PC_IN(1) => 
                           sig_HDU_PC_OUT_1_port, HDU_PC_IN(0) => 
                           sig_HDU_PC_OUT_0_port, HDU_NPC_IN(31) => 
                           sig_HDU_NPC_OUT_31_port, HDU_NPC_IN(30) => 
                           sig_HDU_NPC_OUT_30_port, HDU_NPC_IN(29) => 
                           sig_HDU_NPC_OUT_29_port, HDU_NPC_IN(28) => 
                           sig_HDU_NPC_OUT_28_port, HDU_NPC_IN(27) => 
                           sig_HDU_NPC_OUT_27_port, HDU_NPC_IN(26) => 
                           sig_HDU_NPC_OUT_26_port, HDU_NPC_IN(25) => 
                           sig_HDU_NPC_OUT_25_port, HDU_NPC_IN(24) => 
                           sig_HDU_NPC_OUT_24_port, HDU_NPC_IN(23) => 
                           sig_HDU_NPC_OUT_23_port, HDU_NPC_IN(22) => 
                           sig_HDU_NPC_OUT_22_port, HDU_NPC_IN(21) => 
                           sig_HDU_NPC_OUT_21_port, HDU_NPC_IN(20) => 
                           sig_HDU_NPC_OUT_20_port, HDU_NPC_IN(19) => 
                           sig_HDU_NPC_OUT_19_port, HDU_NPC_IN(18) => 
                           sig_HDU_NPC_OUT_18_port, HDU_NPC_IN(17) => 
                           sig_HDU_NPC_OUT_17_port, HDU_NPC_IN(16) => 
                           sig_HDU_NPC_OUT_16_port, HDU_NPC_IN(15) => 
                           sig_HDU_NPC_OUT_15_port, HDU_NPC_IN(14) => 
                           sig_HDU_NPC_OUT_14_port, HDU_NPC_IN(13) => 
                           sig_HDU_NPC_OUT_13_port, HDU_NPC_IN(12) => 
                           sig_HDU_NPC_OUT_12_port, HDU_NPC_IN(11) => 
                           sig_HDU_NPC_OUT_11_port, HDU_NPC_IN(10) => 
                           sig_HDU_NPC_OUT_10_port, HDU_NPC_IN(9) => 
                           sig_HDU_NPC_OUT_9_port, HDU_NPC_IN(8) => 
                           sig_HDU_NPC_OUT_8_port, HDU_NPC_IN(7) => 
                           sig_HDU_NPC_OUT_7_port, HDU_NPC_IN(6) => 
                           sig_HDU_NPC_OUT_6_port, HDU_NPC_IN(5) => 
                           sig_HDU_NPC_OUT_5_port, HDU_NPC_IN(4) => 
                           sig_HDU_NPC_OUT_4_port, HDU_NPC_IN(3) => 
                           sig_HDU_NPC_OUT_3_port, HDU_NPC_IN(2) => 
                           sig_HDU_NPC_OUT_2_port, HDU_NPC_IN(1) => 
                           sig_HDU_NPC_OUT_1_port, HDU_NPC_IN(0) => 
                           sig_HDU_NPC_OUT_0_port, PC_OUT(31) => 
                           PC_FETCH_OUT_31_port, PC_OUT(30) => 
                           PC_FETCH_OUT_30_port, PC_OUT(29) => 
                           PC_FETCH_OUT_29_port, PC_OUT(28) => 
                           PC_FETCH_OUT_28_port, PC_OUT(27) => 
                           PC_FETCH_OUT_27_port, PC_OUT(26) => 
                           PC_FETCH_OUT_26_port, PC_OUT(25) => 
                           PC_FETCH_OUT_25_port, PC_OUT(24) => 
                           PC_FETCH_OUT_24_port, PC_OUT(23) => 
                           PC_FETCH_OUT_23_port, PC_OUT(22) => 
                           PC_FETCH_OUT_22_port, PC_OUT(21) => 
                           PC_FETCH_OUT_21_port, PC_OUT(20) => 
                           PC_FETCH_OUT_20_port, PC_OUT(19) => 
                           PC_FETCH_OUT_19_port, PC_OUT(18) => 
                           PC_FETCH_OUT_18_port, PC_OUT(17) => 
                           PC_FETCH_OUT_17_port, PC_OUT(16) => 
                           PC_FETCH_OUT_16_port, PC_OUT(15) => 
                           PC_FETCH_OUT_15_port, PC_OUT(14) => 
                           PC_FETCH_OUT_14_port, PC_OUT(13) => 
                           PC_FETCH_OUT_13_port, PC_OUT(12) => 
                           PC_FETCH_OUT_12_port, PC_OUT(11) => 
                           PC_FETCH_OUT_11_port, PC_OUT(10) => 
                           PC_FETCH_OUT_10_port, PC_OUT(9) => 
                           PC_FETCH_OUT_9_port, PC_OUT(8) => 
                           PC_FETCH_OUT_8_port, PC_OUT(7) => 
                           PC_FETCH_OUT_7_port, PC_OUT(6) => 
                           PC_FETCH_OUT_6_port, PC_OUT(5) => 
                           PC_FETCH_OUT_5_port, PC_OUT(4) => 
                           PC_FETCH_OUT_4_port, PC_OUT(3) => 
                           PC_FETCH_OUT_3_port, PC_OUT(2) => 
                           PC_FETCH_OUT_2_port, PC_OUT(1) => 
                           PC_FETCH_OUT_1_port, PC_OUT(0) => 
                           PC_FETCH_OUT_0_port, ADDR_OUT(31) => 
                           IRAM_ADDR_OUT(31), ADDR_OUT(30) => IRAM_ADDR_OUT(30)
                           , ADDR_OUT(29) => IRAM_ADDR_OUT(29), ADDR_OUT(28) =>
                           IRAM_ADDR_OUT(28), ADDR_OUT(27) => IRAM_ADDR_OUT(27)
                           , ADDR_OUT(26) => IRAM_ADDR_OUT(26), ADDR_OUT(25) =>
                           IRAM_ADDR_OUT(25), ADDR_OUT(24) => IRAM_ADDR_OUT(24)
                           , ADDR_OUT(23) => IRAM_ADDR_OUT(23), ADDR_OUT(22) =>
                           IRAM_ADDR_OUT(22), ADDR_OUT(21) => IRAM_ADDR_OUT(21)
                           , ADDR_OUT(20) => IRAM_ADDR_OUT(20), ADDR_OUT(19) =>
                           IRAM_ADDR_OUT(19), ADDR_OUT(18) => IRAM_ADDR_OUT(18)
                           , ADDR_OUT(17) => IRAM_ADDR_OUT(17), ADDR_OUT(16) =>
                           IRAM_ADDR_OUT(16), ADDR_OUT(15) => IRAM_ADDR_OUT(15)
                           , ADDR_OUT(14) => IRAM_ADDR_OUT(14), ADDR_OUT(13) =>
                           IRAM_ADDR_OUT(13), ADDR_OUT(12) => IRAM_ADDR_OUT(12)
                           , ADDR_OUT(11) => IRAM_ADDR_OUT(11), ADDR_OUT(10) =>
                           IRAM_ADDR_OUT(10), ADDR_OUT(9) => IRAM_ADDR_OUT(9), 
                           ADDR_OUT(8) => IRAM_ADDR_OUT(8), ADDR_OUT(7) => 
                           IRAM_ADDR_OUT(7), ADDR_OUT(6) => IRAM_ADDR_OUT(6), 
                           ADDR_OUT(5) => IRAM_ADDR_OUT(5), ADDR_OUT(4) => 
                           IRAM_ADDR_OUT(4), ADDR_OUT(3) => IRAM_ADDR_OUT(3), 
                           ADDR_OUT(2) => IRAM_ADDR_OUT(2), ADDR_OUT(1) => 
                           IRAM_ADDR_OUT(1), ADDR_OUT(0) => IRAM_ADDR_OUT(0), 
                           NPC_OUT(31) => NPC_FETCH_OUT_31_port, NPC_OUT(30) =>
                           NPC_FETCH_OUT_30_port, NPC_OUT(29) => 
                           NPC_FETCH_OUT_29_port, NPC_OUT(28) => 
                           NPC_FETCH_OUT_28_port, NPC_OUT(27) => 
                           NPC_FETCH_OUT_27_port, NPC_OUT(26) => 
                           NPC_FETCH_OUT_26_port, NPC_OUT(25) => 
                           NPC_FETCH_OUT_25_port, NPC_OUT(24) => 
                           NPC_FETCH_OUT_24_port, NPC_OUT(23) => 
                           NPC_FETCH_OUT_23_port, NPC_OUT(22) => 
                           NPC_FETCH_OUT_22_port, NPC_OUT(21) => 
                           NPC_FETCH_OUT_21_port, NPC_OUT(20) => 
                           NPC_FETCH_OUT_20_port, NPC_OUT(19) => 
                           NPC_FETCH_OUT_19_port, NPC_OUT(18) => 
                           NPC_FETCH_OUT_18_port, NPC_OUT(17) => 
                           NPC_FETCH_OUT_17_port, NPC_OUT(16) => 
                           NPC_FETCH_OUT_16_port, NPC_OUT(15) => 
                           NPC_FETCH_OUT_15_port, NPC_OUT(14) => 
                           NPC_FETCH_OUT_14_port, NPC_OUT(13) => 
                           NPC_FETCH_OUT_13_port, NPC_OUT(12) => 
                           NPC_FETCH_OUT_12_port, NPC_OUT(11) => 
                           NPC_FETCH_OUT_11_port, NPC_OUT(10) => 
                           NPC_FETCH_OUT_10_port, NPC_OUT(9) => 
                           NPC_FETCH_OUT_9_port, NPC_OUT(8) => 
                           NPC_FETCH_OUT_8_port, NPC_OUT(7) => 
                           NPC_FETCH_OUT_7_port, NPC_OUT(6) => 
                           NPC_FETCH_OUT_6_port, NPC_OUT(5) => 
                           NPC_FETCH_OUT_5_port, NPC_OUT(4) => 
                           NPC_FETCH_OUT_4_port, NPC_OUT(3) => 
                           NPC_FETCH_OUT_3_port, NPC_OUT(2) => 
                           NPC_FETCH_OUT_2_port, NPC_OUT(1) => 
                           NPC_FETCH_OUT_1_port, NPC_OUT(0) => 
                           NPC_FETCH_OUT_0_port, INS_OUT(31) => INS_OUT_31_port
                           , INS_OUT(30) => INS_OUT_30_port, INS_OUT(29) => 
                           INS_OUT_29_port, INS_OUT(28) => INS_OUT_28_port, 
                           INS_OUT(27) => INS_OUT_27_port, INS_OUT(26) => 
                           INS_OUT_26_port, INS_OUT(25) => INS_OUT_25_port, 
                           INS_OUT(24) => INS_OUT_24_port, INS_OUT(23) => 
                           INS_OUT_23_port, INS_OUT(22) => INS_OUT_22_port, 
                           INS_OUT(21) => INS_OUT_21_port, INS_OUT(20) => 
                           INS_OUT_20_port, INS_OUT(19) => INS_OUT_19_port, 
                           INS_OUT(18) => INS_OUT_18_port, INS_OUT(17) => 
                           INS_OUT_17_port, INS_OUT(16) => INS_OUT_16_port, 
                           INS_OUT(15) => INS_OUT_15_port, INS_OUT(14) => 
                           INS_OUT_14_port, INS_OUT(13) => INS_OUT_13_port, 
                           INS_OUT(12) => INS_OUT_12_port, INS_OUT(11) => 
                           INS_OUT_11_port, INS_OUT(10) => INS_OUT_10_port, 
                           INS_OUT(9) => INS_OUT_9_port, INS_OUT(8) => 
                           INS_OUT_8_port, INS_OUT(7) => INS_OUT_7_port, 
                           INS_OUT(6) => INS_OUT_6_port, INS_OUT(5) => 
                           INS_OUT_5_port, INS_OUT(4) => INS_OUT_4_port, 
                           INS_OUT(3) => INS_OUT_3_port, INS_OUT(2) => 
                           INS_OUT_2_port, INS_OUT(1) => INS_OUT_1_port, 
                           INS_OUT(0) => INS_OUT_0_port);
   DecodeStage : Decode port map( CLK => CLK, RST => RST, REG_LATCH_EN => 
                           REG_LATCH_EN, RD1 => RD1, RD2 => RD2, RF_WE => 
                           RF_WE_WB, ZERO_FLAG => ZERO_FLAG_EX, PC_IN(31) => 
                           PC_FETCH_OUT_31_port, PC_IN(30) => 
                           PC_FETCH_OUT_30_port, PC_IN(29) => 
                           PC_FETCH_OUT_29_port, PC_IN(28) => 
                           PC_FETCH_OUT_28_port, PC_IN(27) => 
                           PC_FETCH_OUT_27_port, PC_IN(26) => 
                           PC_FETCH_OUT_26_port, PC_IN(25) => 
                           PC_FETCH_OUT_25_port, PC_IN(24) => 
                           PC_FETCH_OUT_24_port, PC_IN(23) => 
                           PC_FETCH_OUT_23_port, PC_IN(22) => 
                           PC_FETCH_OUT_22_port, PC_IN(21) => 
                           PC_FETCH_OUT_21_port, PC_IN(20) => 
                           PC_FETCH_OUT_20_port, PC_IN(19) => 
                           PC_FETCH_OUT_19_port, PC_IN(18) => 
                           PC_FETCH_OUT_18_port, PC_IN(17) => 
                           PC_FETCH_OUT_17_port, PC_IN(16) => 
                           PC_FETCH_OUT_16_port, PC_IN(15) => 
                           PC_FETCH_OUT_15_port, PC_IN(14) => 
                           PC_FETCH_OUT_14_port, PC_IN(13) => 
                           PC_FETCH_OUT_13_port, PC_IN(12) => 
                           PC_FETCH_OUT_12_port, PC_IN(11) => 
                           PC_FETCH_OUT_11_port, PC_IN(10) => 
                           PC_FETCH_OUT_10_port, PC_IN(9) => 
                           PC_FETCH_OUT_9_port, PC_IN(8) => PC_FETCH_OUT_8_port
                           , PC_IN(7) => PC_FETCH_OUT_7_port, PC_IN(6) => 
                           PC_FETCH_OUT_6_port, PC_IN(5) => PC_FETCH_OUT_5_port
                           , PC_IN(4) => PC_FETCH_OUT_4_port, PC_IN(3) => 
                           PC_FETCH_OUT_3_port, PC_IN(2) => PC_FETCH_OUT_2_port
                           , PC_IN(1) => PC_FETCH_OUT_1_port, PC_IN(0) => 
                           PC_FETCH_OUT_0_port, INS_IN(31) => INS_OUT_31_port, 
                           INS_IN(30) => INS_OUT_30_port, INS_IN(29) => 
                           INS_OUT_29_port, INS_IN(28) => INS_OUT_28_port, 
                           INS_IN(27) => INS_OUT_27_port, INS_IN(26) => 
                           INS_OUT_26_port, INS_IN(25) => INS_OUT_25_port, 
                           INS_IN(24) => INS_OUT_24_port, INS_IN(23) => 
                           INS_OUT_23_port, INS_IN(22) => INS_OUT_22_port, 
                           INS_IN(21) => INS_OUT_21_port, INS_IN(20) => 
                           INS_OUT_20_port, INS_IN(19) => INS_OUT_19_port, 
                           INS_IN(18) => INS_OUT_18_port, INS_IN(17) => 
                           INS_OUT_17_port, INS_IN(16) => INS_OUT_16_port, 
                           INS_IN(15) => INS_OUT_15_port, INS_IN(14) => 
                           INS_OUT_14_port, INS_IN(13) => INS_OUT_13_port, 
                           INS_IN(12) => INS_OUT_12_port, INS_IN(11) => 
                           INS_OUT_11_port, INS_IN(10) => INS_OUT_10_port, 
                           INS_IN(9) => INS_OUT_9_port, INS_IN(8) => 
                           INS_OUT_8_port, INS_IN(7) => INS_OUT_7_port, 
                           INS_IN(6) => INS_OUT_6_port, INS_IN(5) => 
                           INS_OUT_5_port, INS_IN(4) => INS_OUT_4_port, 
                           INS_IN(3) => INS_OUT_3_port, INS_IN(2) => 
                           INS_OUT_2_port, INS_IN(1) => INS_OUT_1_port, 
                           INS_IN(0) => INS_OUT_0_port, ADD_WR(4) => 
                           ADD_WR_WB_4_port, ADD_WR(3) => ADD_WR_WB_3_port, 
                           ADD_WR(2) => ADD_WR_WB_2_port, ADD_WR(1) => 
                           ADD_WR_WB_1_port, ADD_WR(0) => ADD_WR_WB_0_port, 
                           DATA_WR_IN(31) => OP_WB_31_port, DATA_WR_IN(30) => 
                           OP_WB_30_port, DATA_WR_IN(29) => OP_WB_29_port, 
                           DATA_WR_IN(28) => OP_WB_28_port, DATA_WR_IN(27) => 
                           OP_WB_27_port, DATA_WR_IN(26) => OP_WB_26_port, 
                           DATA_WR_IN(25) => OP_WB_25_port, DATA_WR_IN(24) => 
                           OP_WB_24_port, DATA_WR_IN(23) => OP_WB_23_port, 
                           DATA_WR_IN(22) => OP_WB_22_port, DATA_WR_IN(21) => 
                           OP_WB_21_port, DATA_WR_IN(20) => OP_WB_20_port, 
                           DATA_WR_IN(19) => OP_WB_19_port, DATA_WR_IN(18) => 
                           OP_WB_18_port, DATA_WR_IN(17) => OP_WB_17_port, 
                           DATA_WR_IN(16) => OP_WB_16_port, DATA_WR_IN(15) => 
                           OP_WB_15_port, DATA_WR_IN(14) => OP_WB_14_port, 
                           DATA_WR_IN(13) => OP_WB_13_port, DATA_WR_IN(12) => 
                           OP_WB_12_port, DATA_WR_IN(11) => OP_WB_11_port, 
                           DATA_WR_IN(10) => OP_WB_10_port, DATA_WR_IN(9) => 
                           OP_WB_9_port, DATA_WR_IN(8) => OP_WB_8_port, 
                           DATA_WR_IN(7) => OP_WB_7_port, DATA_WR_IN(6) => 
                           OP_WB_6_port, DATA_WR_IN(5) => OP_WB_5_port, 
                           DATA_WR_IN(4) => OP_WB_4_port, DATA_WR_IN(3) => 
                           OP_WB_3_port, DATA_WR_IN(2) => OP_WB_2_port, 
                           DATA_WR_IN(1) => OP_WB_1_port, DATA_WR_IN(0) => 
                           OP_WB_0_port, PC_OUT(31) => PC_DECODE_OUT_31_port, 
                           PC_OUT(30) => PC_DECODE_OUT_30_port, PC_OUT(29) => 
                           PC_DECODE_OUT_29_port, PC_OUT(28) => 
                           PC_DECODE_OUT_28_port, PC_OUT(27) => 
                           PC_DECODE_OUT_27_port, PC_OUT(26) => 
                           PC_DECODE_OUT_26_port, PC_OUT(25) => 
                           PC_DECODE_OUT_25_port, PC_OUT(24) => 
                           PC_DECODE_OUT_24_port, PC_OUT(23) => 
                           PC_DECODE_OUT_23_port, PC_OUT(22) => 
                           PC_DECODE_OUT_22_port, PC_OUT(21) => 
                           PC_DECODE_OUT_21_port, PC_OUT(20) => 
                           PC_DECODE_OUT_20_port, PC_OUT(19) => 
                           PC_DECODE_OUT_19_port, PC_OUT(18) => 
                           PC_DECODE_OUT_18_port, PC_OUT(17) => 
                           PC_DECODE_OUT_17_port, PC_OUT(16) => 
                           PC_DECODE_OUT_16_port, PC_OUT(15) => 
                           PC_DECODE_OUT_15_port, PC_OUT(14) => 
                           PC_DECODE_OUT_14_port, PC_OUT(13) => 
                           PC_DECODE_OUT_13_port, PC_OUT(12) => 
                           PC_DECODE_OUT_12_port, PC_OUT(11) => 
                           PC_DECODE_OUT_11_port, PC_OUT(10) => 
                           PC_DECODE_OUT_10_port, PC_OUT(9) => 
                           PC_DECODE_OUT_9_port, PC_OUT(8) => 
                           PC_DECODE_OUT_8_port, PC_OUT(7) => 
                           PC_DECODE_OUT_7_port, PC_OUT(6) => 
                           PC_DECODE_OUT_6_port, PC_OUT(5) => 
                           PC_DECODE_OUT_5_port, PC_OUT(4) => 
                           PC_DECODE_OUT_4_port, PC_OUT(3) => 
                           PC_DECODE_OUT_3_port, PC_OUT(2) => 
                           PC_DECODE_OUT_2_port, PC_OUT(1) => 
                           PC_DECODE_OUT_1_port, PC_OUT(0) => 
                           PC_DECODE_OUT_0_port, A_OUT(31) => 
                           A_DECODE_OUT_31_port, A_OUT(30) => 
                           A_DECODE_OUT_30_port, A_OUT(29) => 
                           A_DECODE_OUT_29_port, A_OUT(28) => 
                           A_DECODE_OUT_28_port, A_OUT(27) => 
                           A_DECODE_OUT_27_port, A_OUT(26) => 
                           A_DECODE_OUT_26_port, A_OUT(25) => 
                           A_DECODE_OUT_25_port, A_OUT(24) => 
                           A_DECODE_OUT_24_port, A_OUT(23) => 
                           A_DECODE_OUT_23_port, A_OUT(22) => 
                           A_DECODE_OUT_22_port, A_OUT(21) => 
                           A_DECODE_OUT_21_port, A_OUT(20) => 
                           A_DECODE_OUT_20_port, A_OUT(19) => 
                           A_DECODE_OUT_19_port, A_OUT(18) => 
                           A_DECODE_OUT_18_port, A_OUT(17) => 
                           A_DECODE_OUT_17_port, A_OUT(16) => 
                           A_DECODE_OUT_16_port, A_OUT(15) => 
                           A_DECODE_OUT_15_port, A_OUT(14) => 
                           A_DECODE_OUT_14_port, A_OUT(13) => 
                           A_DECODE_OUT_13_port, A_OUT(12) => 
                           A_DECODE_OUT_12_port, A_OUT(11) => 
                           A_DECODE_OUT_11_port, A_OUT(10) => 
                           A_DECODE_OUT_10_port, A_OUT(9) => 
                           A_DECODE_OUT_9_port, A_OUT(8) => A_DECODE_OUT_8_port
                           , A_OUT(7) => A_DECODE_OUT_7_port, A_OUT(6) => 
                           A_DECODE_OUT_6_port, A_OUT(5) => A_DECODE_OUT_5_port
                           , A_OUT(4) => A_DECODE_OUT_4_port, A_OUT(3) => 
                           A_DECODE_OUT_3_port, A_OUT(2) => A_DECODE_OUT_2_port
                           , A_OUT(1) => A_DECODE_OUT_1_port, A_OUT(0) => 
                           A_DECODE_OUT_0_port, B_OUT(31) => 
                           B_DECODE_OUT_31_port, B_OUT(30) => 
                           B_DECODE_OUT_30_port, B_OUT(29) => 
                           B_DECODE_OUT_29_port, B_OUT(28) => 
                           B_DECODE_OUT_28_port, B_OUT(27) => 
                           B_DECODE_OUT_27_port, B_OUT(26) => 
                           B_DECODE_OUT_26_port, B_OUT(25) => 
                           B_DECODE_OUT_25_port, B_OUT(24) => 
                           B_DECODE_OUT_24_port, B_OUT(23) => 
                           B_DECODE_OUT_23_port, B_OUT(22) => 
                           B_DECODE_OUT_22_port, B_OUT(21) => 
                           B_DECODE_OUT_21_port, B_OUT(20) => 
                           B_DECODE_OUT_20_port, B_OUT(19) => 
                           B_DECODE_OUT_19_port, B_OUT(18) => 
                           B_DECODE_OUT_18_port, B_OUT(17) => 
                           B_DECODE_OUT_17_port, B_OUT(16) => 
                           B_DECODE_OUT_16_port, B_OUT(15) => 
                           B_DECODE_OUT_15_port, B_OUT(14) => 
                           B_DECODE_OUT_14_port, B_OUT(13) => 
                           B_DECODE_OUT_13_port, B_OUT(12) => 
                           B_DECODE_OUT_12_port, B_OUT(11) => 
                           B_DECODE_OUT_11_port, B_OUT(10) => 
                           B_DECODE_OUT_10_port, B_OUT(9) => 
                           B_DECODE_OUT_9_port, B_OUT(8) => B_DECODE_OUT_8_port
                           , B_OUT(7) => B_DECODE_OUT_7_port, B_OUT(6) => 
                           B_DECODE_OUT_6_port, B_OUT(5) => B_DECODE_OUT_5_port
                           , B_OUT(4) => B_DECODE_OUT_4_port, B_OUT(3) => 
                           B_DECODE_OUT_3_port, B_OUT(2) => B_DECODE_OUT_2_port
                           , B_OUT(1) => B_DECODE_OUT_1_port, B_OUT(0) => 
                           B_DECODE_OUT_0_port, IMM_OUT(31) => 
                           IMM_DECODE_OUT_31_port, IMM_OUT(30) => 
                           IMM_DECODE_OUT_30_port, IMM_OUT(29) => 
                           IMM_DECODE_OUT_29_port, IMM_OUT(28) => 
                           IMM_DECODE_OUT_28_port, IMM_OUT(27) => 
                           IMM_DECODE_OUT_27_port, IMM_OUT(26) => 
                           IMM_DECODE_OUT_26_port, IMM_OUT(25) => 
                           IMM_DECODE_OUT_25_port, IMM_OUT(24) => 
                           IMM_DECODE_OUT_24_port, IMM_OUT(23) => 
                           IMM_DECODE_OUT_23_port, IMM_OUT(22) => 
                           IMM_DECODE_OUT_22_port, IMM_OUT(21) => 
                           IMM_DECODE_OUT_21_port, IMM_OUT(20) => 
                           IMM_DECODE_OUT_20_port, IMM_OUT(19) => 
                           IMM_DECODE_OUT_19_port, IMM_OUT(18) => 
                           IMM_DECODE_OUT_18_port, IMM_OUT(17) => 
                           IMM_DECODE_OUT_17_port, IMM_OUT(16) => 
                           IMM_DECODE_OUT_16_port, IMM_OUT(15) => 
                           IMM_DECODE_OUT_15_port, IMM_OUT(14) => 
                           IMM_DECODE_OUT_14_port, IMM_OUT(13) => 
                           IMM_DECODE_OUT_13_port, IMM_OUT(12) => 
                           IMM_DECODE_OUT_12_port, IMM_OUT(11) => 
                           IMM_DECODE_OUT_11_port, IMM_OUT(10) => 
                           IMM_DECODE_OUT_10_port, IMM_OUT(9) => 
                           IMM_DECODE_OUT_9_port, IMM_OUT(8) => 
                           IMM_DECODE_OUT_8_port, IMM_OUT(7) => 
                           IMM_DECODE_OUT_7_port, IMM_OUT(6) => 
                           IMM_DECODE_OUT_6_port, IMM_OUT(5) => 
                           IMM_DECODE_OUT_5_port, IMM_OUT(4) => 
                           IMM_DECODE_OUT_4_port, IMM_OUT(3) => 
                           IMM_DECODE_OUT_3_port, IMM_OUT(2) => 
                           IMM_DECODE_OUT_2_port, IMM_OUT(1) => 
                           IMM_DECODE_OUT_1_port, IMM_OUT(0) => 
                           IMM_DECODE_OUT_0_port, ADD_RS1_HDU(4) => 
                           ADD_RS1_HDU_4_port, ADD_RS1_HDU(3) => 
                           ADD_RS1_HDU_3_port, ADD_RS1_HDU(2) => 
                           ADD_RS1_HDU_2_port, ADD_RS1_HDU(1) => 
                           ADD_RS1_HDU_1_port, ADD_RS1_HDU(0) => 
                           ADD_RS1_HDU_0_port, ADD_RS2_HDU(4) => 
                           ADD_RS2_HDU_4_port, ADD_RS2_HDU(3) => 
                           ADD_RS2_HDU_3_port, ADD_RS2_HDU(2) => 
                           ADD_RS2_HDU_2_port, ADD_RS2_HDU(1) => 
                           ADD_RS2_HDU_1_port, ADD_RS2_HDU(0) => 
                           ADD_RS2_HDU_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_DECODE_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_DECODE_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_DECODE_OUT_0_port, ADD_RS1_OUT(4) => 
                           ADD_RS1_DECODE_OUT_4_port, ADD_RS1_OUT(3) => 
                           ADD_RS1_DECODE_OUT_3_port, ADD_RS1_OUT(2) => 
                           ADD_RS1_DECODE_OUT_2_port, ADD_RS1_OUT(1) => 
                           ADD_RS1_DECODE_OUT_1_port, ADD_RS1_OUT(0) => 
                           ADD_RS1_DECODE_OUT_0_port, ADD_RS2_OUT(4) => 
                           ADD_RS2_DECODE_OUT_4_port, ADD_RS2_OUT(3) => 
                           ADD_RS2_DECODE_OUT_3_port, ADD_RS2_OUT(2) => 
                           ADD_RS2_DECODE_OUT_2_port, ADD_RS2_OUT(1) => 
                           ADD_RS2_DECODE_OUT_1_port, ADD_RS2_OUT(0) => 
                           ADD_RS2_DECODE_OUT_0_port);
   ExecuteStage : Execute port map( CLK => CLK, RST => RST, MUX_A_SEL => 
                           MUX_A_SEL, MUX_B_SEL(1) => MUX_B_SEL(1), 
                           MUX_B_SEL(0) => MUX_B_SEL(0), ALU_OPC(0) => 
                           ALU_OPC(0), ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => 
                           ALU_OPC(2), ALU_OPC(3) => ALU_OPC(3), ALU_OUTREG_EN 
                           => ALU_OUTREG_EN, JUMP_TYPE(1) => JUMP_TYPE(1), 
                           JUMP_TYPE(0) => JUMP_TYPE(0), PC_IN(31) => 
                           PC_DECODE_OUT_31_port, PC_IN(30) => 
                           PC_DECODE_OUT_30_port, PC_IN(29) => 
                           PC_DECODE_OUT_29_port, PC_IN(28) => 
                           PC_DECODE_OUT_28_port, PC_IN(27) => 
                           PC_DECODE_OUT_27_port, PC_IN(26) => 
                           PC_DECODE_OUT_26_port, PC_IN(25) => 
                           PC_DECODE_OUT_25_port, PC_IN(24) => 
                           PC_DECODE_OUT_24_port, PC_IN(23) => 
                           PC_DECODE_OUT_23_port, PC_IN(22) => 
                           PC_DECODE_OUT_22_port, PC_IN(21) => 
                           PC_DECODE_OUT_21_port, PC_IN(20) => 
                           PC_DECODE_OUT_20_port, PC_IN(19) => 
                           PC_DECODE_OUT_19_port, PC_IN(18) => 
                           PC_DECODE_OUT_18_port, PC_IN(17) => 
                           PC_DECODE_OUT_17_port, PC_IN(16) => 
                           PC_DECODE_OUT_16_port, PC_IN(15) => 
                           PC_DECODE_OUT_15_port, PC_IN(14) => 
                           PC_DECODE_OUT_14_port, PC_IN(13) => 
                           PC_DECODE_OUT_13_port, PC_IN(12) => 
                           PC_DECODE_OUT_12_port, PC_IN(11) => 
                           PC_DECODE_OUT_11_port, PC_IN(10) => 
                           PC_DECODE_OUT_10_port, PC_IN(9) => 
                           PC_DECODE_OUT_9_port, PC_IN(8) => 
                           PC_DECODE_OUT_8_port, PC_IN(7) => 
                           PC_DECODE_OUT_7_port, PC_IN(6) => 
                           PC_DECODE_OUT_6_port, PC_IN(5) => 
                           PC_DECODE_OUT_5_port, PC_IN(4) => 
                           PC_DECODE_OUT_4_port, PC_IN(3) => 
                           PC_DECODE_OUT_3_port, PC_IN(2) => 
                           PC_DECODE_OUT_2_port, PC_IN(1) => 
                           PC_DECODE_OUT_1_port, PC_IN(0) => 
                           PC_DECODE_OUT_0_port, A_IN(31) => 
                           A_DECODE_OUT_31_port, A_IN(30) => 
                           A_DECODE_OUT_30_port, A_IN(29) => 
                           A_DECODE_OUT_29_port, A_IN(28) => 
                           A_DECODE_OUT_28_port, A_IN(27) => 
                           A_DECODE_OUT_27_port, A_IN(26) => 
                           A_DECODE_OUT_26_port, A_IN(25) => 
                           A_DECODE_OUT_25_port, A_IN(24) => 
                           A_DECODE_OUT_24_port, A_IN(23) => 
                           A_DECODE_OUT_23_port, A_IN(22) => 
                           A_DECODE_OUT_22_port, A_IN(21) => 
                           A_DECODE_OUT_21_port, A_IN(20) => 
                           A_DECODE_OUT_20_port, A_IN(19) => 
                           A_DECODE_OUT_19_port, A_IN(18) => 
                           A_DECODE_OUT_18_port, A_IN(17) => 
                           A_DECODE_OUT_17_port, A_IN(16) => 
                           A_DECODE_OUT_16_port, A_IN(15) => 
                           A_DECODE_OUT_15_port, A_IN(14) => 
                           A_DECODE_OUT_14_port, A_IN(13) => 
                           A_DECODE_OUT_13_port, A_IN(12) => 
                           A_DECODE_OUT_12_port, A_IN(11) => 
                           A_DECODE_OUT_11_port, A_IN(10) => 
                           A_DECODE_OUT_10_port, A_IN(9) => A_DECODE_OUT_9_port
                           , A_IN(8) => A_DECODE_OUT_8_port, A_IN(7) => 
                           A_DECODE_OUT_7_port, A_IN(6) => A_DECODE_OUT_6_port,
                           A_IN(5) => A_DECODE_OUT_5_port, A_IN(4) => 
                           A_DECODE_OUT_4_port, A_IN(3) => A_DECODE_OUT_3_port,
                           A_IN(2) => A_DECODE_OUT_2_port, A_IN(1) => 
                           A_DECODE_OUT_1_port, A_IN(0) => A_DECODE_OUT_0_port,
                           B_IN(31) => B_DECODE_OUT_31_port, B_IN(30) => 
                           B_DECODE_OUT_30_port, B_IN(29) => 
                           B_DECODE_OUT_29_port, B_IN(28) => 
                           B_DECODE_OUT_28_port, B_IN(27) => 
                           B_DECODE_OUT_27_port, B_IN(26) => 
                           B_DECODE_OUT_26_port, B_IN(25) => 
                           B_DECODE_OUT_25_port, B_IN(24) => 
                           B_DECODE_OUT_24_port, B_IN(23) => 
                           B_DECODE_OUT_23_port, B_IN(22) => 
                           B_DECODE_OUT_22_port, B_IN(21) => 
                           B_DECODE_OUT_21_port, B_IN(20) => 
                           B_DECODE_OUT_20_port, B_IN(19) => 
                           B_DECODE_OUT_19_port, B_IN(18) => 
                           B_DECODE_OUT_18_port, B_IN(17) => 
                           B_DECODE_OUT_17_port, B_IN(16) => 
                           B_DECODE_OUT_16_port, B_IN(15) => 
                           B_DECODE_OUT_15_port, B_IN(14) => 
                           B_DECODE_OUT_14_port, B_IN(13) => 
                           B_DECODE_OUT_13_port, B_IN(12) => 
                           B_DECODE_OUT_12_port, B_IN(11) => 
                           B_DECODE_OUT_11_port, B_IN(10) => 
                           B_DECODE_OUT_10_port, B_IN(9) => B_DECODE_OUT_9_port
                           , B_IN(8) => B_DECODE_OUT_8_port, B_IN(7) => 
                           B_DECODE_OUT_7_port, B_IN(6) => B_DECODE_OUT_6_port,
                           B_IN(5) => B_DECODE_OUT_5_port, B_IN(4) => 
                           B_DECODE_OUT_4_port, B_IN(3) => B_DECODE_OUT_3_port,
                           B_IN(2) => B_DECODE_OUT_2_port, B_IN(1) => 
                           B_DECODE_OUT_1_port, B_IN(0) => B_DECODE_OUT_0_port,
                           IMM_IN(31) => IMM_DECODE_OUT_31_port, IMM_IN(30) => 
                           IMM_DECODE_OUT_30_port, IMM_IN(29) => 
                           IMM_DECODE_OUT_29_port, IMM_IN(28) => 
                           IMM_DECODE_OUT_28_port, IMM_IN(27) => 
                           IMM_DECODE_OUT_27_port, IMM_IN(26) => 
                           IMM_DECODE_OUT_26_port, IMM_IN(25) => 
                           IMM_DECODE_OUT_25_port, IMM_IN(24) => 
                           IMM_DECODE_OUT_24_port, IMM_IN(23) => 
                           IMM_DECODE_OUT_23_port, IMM_IN(22) => 
                           IMM_DECODE_OUT_22_port, IMM_IN(21) => 
                           IMM_DECODE_OUT_21_port, IMM_IN(20) => 
                           IMM_DECODE_OUT_20_port, IMM_IN(19) => 
                           IMM_DECODE_OUT_19_port, IMM_IN(18) => 
                           IMM_DECODE_OUT_18_port, IMM_IN(17) => 
                           IMM_DECODE_OUT_17_port, IMM_IN(16) => 
                           IMM_DECODE_OUT_16_port, IMM_IN(15) => 
                           IMM_DECODE_OUT_15_port, IMM_IN(14) => 
                           IMM_DECODE_OUT_14_port, IMM_IN(13) => 
                           IMM_DECODE_OUT_13_port, IMM_IN(12) => 
                           IMM_DECODE_OUT_12_port, IMM_IN(11) => 
                           IMM_DECODE_OUT_11_port, IMM_IN(10) => 
                           IMM_DECODE_OUT_10_port, IMM_IN(9) => 
                           IMM_DECODE_OUT_9_port, IMM_IN(8) => 
                           IMM_DECODE_OUT_8_port, IMM_IN(7) => 
                           IMM_DECODE_OUT_7_port, IMM_IN(6) => 
                           IMM_DECODE_OUT_6_port, IMM_IN(5) => 
                           IMM_DECODE_OUT_5_port, IMM_IN(4) => 
                           IMM_DECODE_OUT_4_port, IMM_IN(3) => 
                           IMM_DECODE_OUT_3_port, IMM_IN(2) => 
                           IMM_DECODE_OUT_2_port, IMM_IN(1) => 
                           IMM_DECODE_OUT_1_port, IMM_IN(0) => 
                           IMM_DECODE_OUT_0_port, ADD_WR_IN(4) => 
                           ADD_WR_DECODE_OUT_4_port, ADD_WR_IN(3) => 
                           ADD_WR_DECODE_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_DECODE_OUT_0_port, ADD_RS1_IN(4) => 
                           ADD_RS1_DECODE_OUT_4_port, ADD_RS1_IN(3) => 
                           ADD_RS1_DECODE_OUT_3_port, ADD_RS1_IN(2) => 
                           ADD_RS1_DECODE_OUT_2_port, ADD_RS1_IN(1) => 
                           ADD_RS1_DECODE_OUT_1_port, ADD_RS1_IN(0) => 
                           ADD_RS1_DECODE_OUT_0_port, ADD_RS2_IN(4) => 
                           ADD_RS2_DECODE_OUT_4_port, ADD_RS2_IN(3) => 
                           ADD_RS2_DECODE_OUT_3_port, ADD_RS2_IN(2) => 
                           ADD_RS2_DECODE_OUT_2_port, ADD_RS2_IN(1) => 
                           ADD_RS2_DECODE_OUT_1_port, ADD_RS2_IN(0) => 
                           ADD_RS2_DECODE_OUT_0_port, ADD_WR_MEM(4) => 
                           ADD_WR_MEM_4_port, ADD_WR_MEM(3) => 
                           ADD_WR_MEM_3_port, ADD_WR_MEM(2) => 
                           ADD_WR_MEM_2_port, ADD_WR_MEM(1) => 
                           ADD_WR_MEM_1_port, ADD_WR_MEM(0) => 
                           ADD_WR_MEM_0_port, ADD_WR_WB(4) => ADD_WR_WB_4_port,
                           ADD_WR_WB(3) => ADD_WR_WB_3_port, ADD_WR_WB(2) => 
                           ADD_WR_WB_2_port, ADD_WR_WB(1) => ADD_WR_WB_1_port, 
                           ADD_WR_WB(0) => ADD_WR_WB_0_port, RF_WE_MEM => RF_WE
                           , RF_WE_WB => RF_WE_WB, OP_MEM(31) => OP_MEM_31_port
                           , OP_MEM(30) => OP_MEM_30_port, OP_MEM(29) => 
                           OP_MEM_29_port, OP_MEM(28) => OP_MEM_28_port, 
                           OP_MEM(27) => OP_MEM_27_port, OP_MEM(26) => 
                           OP_MEM_26_port, OP_MEM(25) => OP_MEM_25_port, 
                           OP_MEM(24) => OP_MEM_24_port, OP_MEM(23) => 
                           OP_MEM_23_port, OP_MEM(22) => OP_MEM_22_port, 
                           OP_MEM(21) => OP_MEM_21_port, OP_MEM(20) => 
                           OP_MEM_20_port, OP_MEM(19) => OP_MEM_19_port, 
                           OP_MEM(18) => OP_MEM_18_port, OP_MEM(17) => 
                           OP_MEM_17_port, OP_MEM(16) => OP_MEM_16_port, 
                           OP_MEM(15) => OP_MEM_15_port, OP_MEM(14) => 
                           OP_MEM_14_port, OP_MEM(13) => OP_MEM_13_port, 
                           OP_MEM(12) => OP_MEM_12_port, OP_MEM(11) => 
                           OP_MEM_11_port, OP_MEM(10) => OP_MEM_10_port, 
                           OP_MEM(9) => OP_MEM_9_port, OP_MEM(8) => 
                           OP_MEM_8_port, OP_MEM(7) => OP_MEM_7_port, OP_MEM(6)
                           => OP_MEM_6_port, OP_MEM(5) => OP_MEM_5_port, 
                           OP_MEM(4) => OP_MEM_4_port, OP_MEM(3) => 
                           OP_MEM_3_port, OP_MEM(2) => OP_MEM_2_port, OP_MEM(1)
                           => OP_MEM_1_port, OP_MEM(0) => OP_MEM_0_port, 
                           OP_WB(31) => OP_WB_31_port, OP_WB(30) => 
                           OP_WB_30_port, OP_WB(29) => OP_WB_29_port, OP_WB(28)
                           => OP_WB_28_port, OP_WB(27) => OP_WB_27_port, 
                           OP_WB(26) => OP_WB_26_port, OP_WB(25) => 
                           OP_WB_25_port, OP_WB(24) => OP_WB_24_port, OP_WB(23)
                           => OP_WB_23_port, OP_WB(22) => OP_WB_22_port, 
                           OP_WB(21) => OP_WB_21_port, OP_WB(20) => 
                           OP_WB_20_port, OP_WB(19) => OP_WB_19_port, OP_WB(18)
                           => OP_WB_18_port, OP_WB(17) => OP_WB_17_port, 
                           OP_WB(16) => OP_WB_16_port, OP_WB(15) => 
                           OP_WB_15_port, OP_WB(14) => OP_WB_14_port, OP_WB(13)
                           => OP_WB_13_port, OP_WB(12) => OP_WB_12_port, 
                           OP_WB(11) => OP_WB_11_port, OP_WB(10) => 
                           OP_WB_10_port, OP_WB(9) => OP_WB_9_port, OP_WB(8) =>
                           OP_WB_8_port, OP_WB(7) => OP_WB_7_port, OP_WB(6) => 
                           OP_WB_6_port, OP_WB(5) => OP_WB_5_port, OP_WB(4) => 
                           OP_WB_4_port, OP_WB(3) => OP_WB_3_port, OP_WB(2) => 
                           OP_WB_2_port, OP_WB(1) => OP_WB_1_port, OP_WB(0) => 
                           OP_WB_0_port, PC_SEL(1) => PC_SEL_EX_1_port, 
                           PC_SEL(0) => PC_SEL_EX_0_port, ZERO_FLAG => 
                           ZERO_FLAG_EX, NPC_ABS(31) => NPC_ABS_EX_31_port, 
                           NPC_ABS(30) => NPC_ABS_EX_30_port, NPC_ABS(29) => 
                           NPC_ABS_EX_29_port, NPC_ABS(28) => 
                           NPC_ABS_EX_28_port, NPC_ABS(27) => 
                           NPC_ABS_EX_27_port, NPC_ABS(26) => 
                           NPC_ABS_EX_26_port, NPC_ABS(25) => 
                           NPC_ABS_EX_25_port, NPC_ABS(24) => 
                           NPC_ABS_EX_24_port, NPC_ABS(23) => 
                           NPC_ABS_EX_23_port, NPC_ABS(22) => 
                           NPC_ABS_EX_22_port, NPC_ABS(21) => 
                           NPC_ABS_EX_21_port, NPC_ABS(20) => 
                           NPC_ABS_EX_20_port, NPC_ABS(19) => 
                           NPC_ABS_EX_19_port, NPC_ABS(18) => 
                           NPC_ABS_EX_18_port, NPC_ABS(17) => 
                           NPC_ABS_EX_17_port, NPC_ABS(16) => 
                           NPC_ABS_EX_16_port, NPC_ABS(15) => 
                           NPC_ABS_EX_15_port, NPC_ABS(14) => 
                           NPC_ABS_EX_14_port, NPC_ABS(13) => 
                           NPC_ABS_EX_13_port, NPC_ABS(12) => 
                           NPC_ABS_EX_12_port, NPC_ABS(11) => 
                           NPC_ABS_EX_11_port, NPC_ABS(10) => 
                           NPC_ABS_EX_10_port, NPC_ABS(9) => NPC_ABS_EX_9_port,
                           NPC_ABS(8) => NPC_ABS_EX_8_port, NPC_ABS(7) => 
                           NPC_ABS_EX_7_port, NPC_ABS(6) => NPC_ABS_EX_6_port, 
                           NPC_ABS(5) => NPC_ABS_EX_5_port, NPC_ABS(4) => 
                           NPC_ABS_EX_4_port, NPC_ABS(3) => NPC_ABS_EX_3_port, 
                           NPC_ABS(2) => NPC_ABS_EX_2_port, NPC_ABS(1) => 
                           NPC_ABS_EX_1_port, NPC_ABS(0) => NPC_ABS_EX_0_port, 
                           NPC_REL(31) => NPC_REL_EX_31_port, NPC_REL(30) => 
                           NPC_REL_EX_30_port, NPC_REL(29) => 
                           NPC_REL_EX_29_port, NPC_REL(28) => 
                           NPC_REL_EX_28_port, NPC_REL(27) => 
                           NPC_REL_EX_27_port, NPC_REL(26) => 
                           NPC_REL_EX_26_port, NPC_REL(25) => 
                           NPC_REL_EX_25_port, NPC_REL(24) => 
                           NPC_REL_EX_24_port, NPC_REL(23) => 
                           NPC_REL_EX_23_port, NPC_REL(22) => 
                           NPC_REL_EX_22_port, NPC_REL(21) => 
                           NPC_REL_EX_21_port, NPC_REL(20) => 
                           NPC_REL_EX_20_port, NPC_REL(19) => 
                           NPC_REL_EX_19_port, NPC_REL(18) => 
                           NPC_REL_EX_18_port, NPC_REL(17) => 
                           NPC_REL_EX_17_port, NPC_REL(16) => 
                           NPC_REL_EX_16_port, NPC_REL(15) => 
                           NPC_REL_EX_15_port, NPC_REL(14) => 
                           NPC_REL_EX_14_port, NPC_REL(13) => 
                           NPC_REL_EX_13_port, NPC_REL(12) => 
                           NPC_REL_EX_12_port, NPC_REL(11) => 
                           NPC_REL_EX_11_port, NPC_REL(10) => 
                           NPC_REL_EX_10_port, NPC_REL(9) => NPC_REL_EX_9_port,
                           NPC_REL(8) => NPC_REL_EX_8_port, NPC_REL(7) => 
                           NPC_REL_EX_7_port, NPC_REL(6) => NPC_REL_EX_6_port, 
                           NPC_REL(5) => NPC_REL_EX_5_port, NPC_REL(4) => 
                           NPC_REL_EX_4_port, NPC_REL(3) => NPC_REL_EX_3_port, 
                           NPC_REL(2) => NPC_REL_EX_2_port, NPC_REL(1) => 
                           NPC_REL_EX_1_port, NPC_REL(0) => NPC_REL_EX_0_port, 
                           ALU_RES(31) => ALU_RES_EX_31_port, ALU_RES(30) => 
                           ALU_RES_EX_30_port, ALU_RES(29) => 
                           ALU_RES_EX_29_port, ALU_RES(28) => 
                           ALU_RES_EX_28_port, ALU_RES(27) => 
                           ALU_RES_EX_27_port, ALU_RES(26) => 
                           ALU_RES_EX_26_port, ALU_RES(25) => 
                           ALU_RES_EX_25_port, ALU_RES(24) => 
                           ALU_RES_EX_24_port, ALU_RES(23) => 
                           ALU_RES_EX_23_port, ALU_RES(22) => 
                           ALU_RES_EX_22_port, ALU_RES(21) => 
                           ALU_RES_EX_21_port, ALU_RES(20) => 
                           ALU_RES_EX_20_port, ALU_RES(19) => 
                           ALU_RES_EX_19_port, ALU_RES(18) => 
                           ALU_RES_EX_18_port, ALU_RES(17) => 
                           ALU_RES_EX_17_port, ALU_RES(16) => 
                           ALU_RES_EX_16_port, ALU_RES(15) => 
                           ALU_RES_EX_15_port, ALU_RES(14) => 
                           ALU_RES_EX_14_port, ALU_RES(13) => 
                           ALU_RES_EX_13_port, ALU_RES(12) => 
                           ALU_RES_EX_12_port, ALU_RES(11) => 
                           ALU_RES_EX_11_port, ALU_RES(10) => 
                           ALU_RES_EX_10_port, ALU_RES(9) => ALU_RES_EX_9_port,
                           ALU_RES(8) => ALU_RES_EX_8_port, ALU_RES(7) => 
                           ALU_RES_EX_7_port, ALU_RES(6) => ALU_RES_EX_6_port, 
                           ALU_RES(5) => ALU_RES_EX_5_port, ALU_RES(4) => 
                           ALU_RES_EX_4_port, ALU_RES(3) => ALU_RES_EX_3_port, 
                           ALU_RES(2) => ALU_RES_EX_2_port, ALU_RES(1) => 
                           ALU_RES_EX_1_port, ALU_RES(0) => ALU_RES_EX_0_port, 
                           B_OUT(31) => B_EX_OUT_31_port, B_OUT(30) => 
                           B_EX_OUT_30_port, B_OUT(29) => B_EX_OUT_29_port, 
                           B_OUT(28) => B_EX_OUT_28_port, B_OUT(27) => 
                           B_EX_OUT_27_port, B_OUT(26) => B_EX_OUT_26_port, 
                           B_OUT(25) => B_EX_OUT_25_port, B_OUT(24) => 
                           B_EX_OUT_24_port, B_OUT(23) => B_EX_OUT_23_port, 
                           B_OUT(22) => B_EX_OUT_22_port, B_OUT(21) => 
                           B_EX_OUT_21_port, B_OUT(20) => B_EX_OUT_20_port, 
                           B_OUT(19) => B_EX_OUT_19_port, B_OUT(18) => 
                           B_EX_OUT_18_port, B_OUT(17) => B_EX_OUT_17_port, 
                           B_OUT(16) => B_EX_OUT_16_port, B_OUT(15) => 
                           B_EX_OUT_15_port, B_OUT(14) => B_EX_OUT_14_port, 
                           B_OUT(13) => B_EX_OUT_13_port, B_OUT(12) => 
                           B_EX_OUT_12_port, B_OUT(11) => B_EX_OUT_11_port, 
                           B_OUT(10) => B_EX_OUT_10_port, B_OUT(9) => 
                           B_EX_OUT_9_port, B_OUT(8) => B_EX_OUT_8_port, 
                           B_OUT(7) => B_EX_OUT_7_port, B_OUT(6) => 
                           B_EX_OUT_6_port, B_OUT(5) => B_EX_OUT_5_port, 
                           B_OUT(4) => B_EX_OUT_4_port, B_OUT(3) => 
                           B_EX_OUT_3_port, B_OUT(2) => B_EX_OUT_2_port, 
                           B_OUT(1) => B_EX_OUT_1_port, B_OUT(0) => 
                           B_EX_OUT_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_EX_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_EX_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_EX_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_EX_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_EX_OUT_0_port);
   DRAM_R_ff : ff_0 port map( D => DRAM_R_IN, CLK => CLK, EN => n1, RST => RST,
                           Q => DRAM_R_MEM);
   MemoryStage : Memory port map( CLK => CLK, RST => RST, MEM_EN_IN => 
                           MEM_EN_IN, DRAM_R_IN => DRAM_R_MEM, DRAM_W_IN => 
                           DRAM_W_IN, DRAM_EN_IN => DRAM_EN_IN, PC_SEL(1) => 
                           PC_SEL_EX_1_port, PC_SEL(0) => PC_SEL_EX_0_port, 
                           NPC_IN(31) => NPC_FETCH_OUT_31_port, NPC_IN(30) => 
                           NPC_FETCH_OUT_30_port, NPC_IN(29) => 
                           NPC_FETCH_OUT_29_port, NPC_IN(28) => 
                           NPC_FETCH_OUT_28_port, NPC_IN(27) => 
                           NPC_FETCH_OUT_27_port, NPC_IN(26) => 
                           NPC_FETCH_OUT_26_port, NPC_IN(25) => 
                           NPC_FETCH_OUT_25_port, NPC_IN(24) => 
                           NPC_FETCH_OUT_24_port, NPC_IN(23) => 
                           NPC_FETCH_OUT_23_port, NPC_IN(22) => 
                           NPC_FETCH_OUT_22_port, NPC_IN(21) => 
                           NPC_FETCH_OUT_21_port, NPC_IN(20) => 
                           NPC_FETCH_OUT_20_port, NPC_IN(19) => 
                           NPC_FETCH_OUT_19_port, NPC_IN(18) => 
                           NPC_FETCH_OUT_18_port, NPC_IN(17) => 
                           NPC_FETCH_OUT_17_port, NPC_IN(16) => 
                           NPC_FETCH_OUT_16_port, NPC_IN(15) => 
                           NPC_FETCH_OUT_15_port, NPC_IN(14) => 
                           NPC_FETCH_OUT_14_port, NPC_IN(13) => 
                           NPC_FETCH_OUT_13_port, NPC_IN(12) => 
                           NPC_FETCH_OUT_12_port, NPC_IN(11) => 
                           NPC_FETCH_OUT_11_port, NPC_IN(10) => 
                           NPC_FETCH_OUT_10_port, NPC_IN(9) => 
                           NPC_FETCH_OUT_9_port, NPC_IN(8) => 
                           NPC_FETCH_OUT_8_port, NPC_IN(7) => 
                           NPC_FETCH_OUT_7_port, NPC_IN(6) => 
                           NPC_FETCH_OUT_6_port, NPC_IN(5) => 
                           NPC_FETCH_OUT_5_port, NPC_IN(4) => 
                           NPC_FETCH_OUT_4_port, NPC_IN(3) => 
                           NPC_FETCH_OUT_3_port, NPC_IN(2) => 
                           NPC_FETCH_OUT_2_port, NPC_IN(1) => 
                           NPC_FETCH_OUT_1_port, NPC_IN(0) => 
                           NPC_FETCH_OUT_0_port, NPC_ABS(31) => 
                           NPC_ABS_EX_31_port, NPC_ABS(30) => 
                           NPC_ABS_EX_30_port, NPC_ABS(29) => 
                           NPC_ABS_EX_29_port, NPC_ABS(28) => 
                           NPC_ABS_EX_28_port, NPC_ABS(27) => 
                           NPC_ABS_EX_27_port, NPC_ABS(26) => 
                           NPC_ABS_EX_26_port, NPC_ABS(25) => 
                           NPC_ABS_EX_25_port, NPC_ABS(24) => 
                           NPC_ABS_EX_24_port, NPC_ABS(23) => 
                           NPC_ABS_EX_23_port, NPC_ABS(22) => 
                           NPC_ABS_EX_22_port, NPC_ABS(21) => 
                           NPC_ABS_EX_21_port, NPC_ABS(20) => 
                           NPC_ABS_EX_20_port, NPC_ABS(19) => 
                           NPC_ABS_EX_19_port, NPC_ABS(18) => 
                           NPC_ABS_EX_18_port, NPC_ABS(17) => 
                           NPC_ABS_EX_17_port, NPC_ABS(16) => 
                           NPC_ABS_EX_16_port, NPC_ABS(15) => 
                           NPC_ABS_EX_15_port, NPC_ABS(14) => 
                           NPC_ABS_EX_14_port, NPC_ABS(13) => 
                           NPC_ABS_EX_13_port, NPC_ABS(12) => 
                           NPC_ABS_EX_12_port, NPC_ABS(11) => 
                           NPC_ABS_EX_11_port, NPC_ABS(10) => 
                           NPC_ABS_EX_10_port, NPC_ABS(9) => NPC_ABS_EX_9_port,
                           NPC_ABS(8) => NPC_ABS_EX_8_port, NPC_ABS(7) => 
                           NPC_ABS_EX_7_port, NPC_ABS(6) => NPC_ABS_EX_6_port, 
                           NPC_ABS(5) => NPC_ABS_EX_5_port, NPC_ABS(4) => 
                           NPC_ABS_EX_4_port, NPC_ABS(3) => NPC_ABS_EX_3_port, 
                           NPC_ABS(2) => NPC_ABS_EX_2_port, NPC_ABS(1) => 
                           NPC_ABS_EX_1_port, NPC_ABS(0) => NPC_ABS_EX_0_port, 
                           NPC_REL(31) => NPC_REL_EX_31_port, NPC_REL(30) => 
                           NPC_REL_EX_30_port, NPC_REL(29) => 
                           NPC_REL_EX_29_port, NPC_REL(28) => 
                           NPC_REL_EX_28_port, NPC_REL(27) => 
                           NPC_REL_EX_27_port, NPC_REL(26) => 
                           NPC_REL_EX_26_port, NPC_REL(25) => 
                           NPC_REL_EX_25_port, NPC_REL(24) => 
                           NPC_REL_EX_24_port, NPC_REL(23) => 
                           NPC_REL_EX_23_port, NPC_REL(22) => 
                           NPC_REL_EX_22_port, NPC_REL(21) => 
                           NPC_REL_EX_21_port, NPC_REL(20) => 
                           NPC_REL_EX_20_port, NPC_REL(19) => 
                           NPC_REL_EX_19_port, NPC_REL(18) => 
                           NPC_REL_EX_18_port, NPC_REL(17) => 
                           NPC_REL_EX_17_port, NPC_REL(16) => 
                           NPC_REL_EX_16_port, NPC_REL(15) => 
                           NPC_REL_EX_15_port, NPC_REL(14) => 
                           NPC_REL_EX_14_port, NPC_REL(13) => 
                           NPC_REL_EX_13_port, NPC_REL(12) => 
                           NPC_REL_EX_12_port, NPC_REL(11) => 
                           NPC_REL_EX_11_port, NPC_REL(10) => 
                           NPC_REL_EX_10_port, NPC_REL(9) => NPC_REL_EX_9_port,
                           NPC_REL(8) => NPC_REL_EX_8_port, NPC_REL(7) => 
                           NPC_REL_EX_7_port, NPC_REL(6) => NPC_REL_EX_6_port, 
                           NPC_REL(5) => NPC_REL_EX_5_port, NPC_REL(4) => 
                           NPC_REL_EX_4_port, NPC_REL(3) => NPC_REL_EX_3_port, 
                           NPC_REL(2) => NPC_REL_EX_2_port, NPC_REL(1) => 
                           NPC_REL_EX_1_port, NPC_REL(0) => NPC_REL_EX_0_port, 
                           ALU_RES_IN(31) => ALU_RES_EX_31_port, ALU_RES_IN(30)
                           => ALU_RES_EX_30_port, ALU_RES_IN(29) => 
                           ALU_RES_EX_29_port, ALU_RES_IN(28) => 
                           ALU_RES_EX_28_port, ALU_RES_IN(27) => 
                           ALU_RES_EX_27_port, ALU_RES_IN(26) => 
                           ALU_RES_EX_26_port, ALU_RES_IN(25) => 
                           ALU_RES_EX_25_port, ALU_RES_IN(24) => 
                           ALU_RES_EX_24_port, ALU_RES_IN(23) => 
                           ALU_RES_EX_23_port, ALU_RES_IN(22) => 
                           ALU_RES_EX_22_port, ALU_RES_IN(21) => 
                           ALU_RES_EX_21_port, ALU_RES_IN(20) => 
                           ALU_RES_EX_20_port, ALU_RES_IN(19) => 
                           ALU_RES_EX_19_port, ALU_RES_IN(18) => 
                           ALU_RES_EX_18_port, ALU_RES_IN(17) => 
                           ALU_RES_EX_17_port, ALU_RES_IN(16) => 
                           ALU_RES_EX_16_port, ALU_RES_IN(15) => 
                           ALU_RES_EX_15_port, ALU_RES_IN(14) => 
                           ALU_RES_EX_14_port, ALU_RES_IN(13) => 
                           ALU_RES_EX_13_port, ALU_RES_IN(12) => 
                           ALU_RES_EX_12_port, ALU_RES_IN(11) => 
                           ALU_RES_EX_11_port, ALU_RES_IN(10) => 
                           ALU_RES_EX_10_port, ALU_RES_IN(9) => 
                           ALU_RES_EX_9_port, ALU_RES_IN(8) => 
                           ALU_RES_EX_8_port, ALU_RES_IN(7) => 
                           ALU_RES_EX_7_port, ALU_RES_IN(6) => 
                           ALU_RES_EX_6_port, ALU_RES_IN(5) => 
                           ALU_RES_EX_5_port, ALU_RES_IN(4) => 
                           ALU_RES_EX_4_port, ALU_RES_IN(3) => 
                           ALU_RES_EX_3_port, ALU_RES_IN(2) => 
                           ALU_RES_EX_2_port, ALU_RES_IN(1) => 
                           ALU_RES_EX_1_port, ALU_RES_IN(0) => 
                           ALU_RES_EX_0_port, B_IN(31) => B_EX_OUT_31_port, 
                           B_IN(30) => B_EX_OUT_30_port, B_IN(29) => 
                           B_EX_OUT_29_port, B_IN(28) => B_EX_OUT_28_port, 
                           B_IN(27) => B_EX_OUT_27_port, B_IN(26) => 
                           B_EX_OUT_26_port, B_IN(25) => B_EX_OUT_25_port, 
                           B_IN(24) => B_EX_OUT_24_port, B_IN(23) => 
                           B_EX_OUT_23_port, B_IN(22) => B_EX_OUT_22_port, 
                           B_IN(21) => B_EX_OUT_21_port, B_IN(20) => 
                           B_EX_OUT_20_port, B_IN(19) => B_EX_OUT_19_port, 
                           B_IN(18) => B_EX_OUT_18_port, B_IN(17) => 
                           B_EX_OUT_17_port, B_IN(16) => B_EX_OUT_16_port, 
                           B_IN(15) => B_EX_OUT_15_port, B_IN(14) => 
                           B_EX_OUT_14_port, B_IN(13) => B_EX_OUT_13_port, 
                           B_IN(12) => B_EX_OUT_12_port, B_IN(11) => 
                           B_EX_OUT_11_port, B_IN(10) => B_EX_OUT_10_port, 
                           B_IN(9) => B_EX_OUT_9_port, B_IN(8) => 
                           B_EX_OUT_8_port, B_IN(7) => B_EX_OUT_7_port, B_IN(6)
                           => B_EX_OUT_6_port, B_IN(5) => B_EX_OUT_5_port, 
                           B_IN(4) => B_EX_OUT_4_port, B_IN(3) => 
                           B_EX_OUT_3_port, B_IN(2) => B_EX_OUT_2_port, B_IN(1)
                           => B_EX_OUT_1_port, B_IN(0) => B_EX_OUT_0_port, 
                           ADD_WR_IN(4) => ADD_WR_EX_OUT_4_port, ADD_WR_IN(3) 
                           => ADD_WR_EX_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_EX_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_EX_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_EX_OUT_0_port, DRAM_DATA_IN(31) => 
                           DATA_IN(31), DRAM_DATA_IN(30) => DATA_IN(30), 
                           DRAM_DATA_IN(29) => DATA_IN(29), DRAM_DATA_IN(28) =>
                           DATA_IN(28), DRAM_DATA_IN(27) => DATA_IN(27), 
                           DRAM_DATA_IN(26) => DATA_IN(26), DRAM_DATA_IN(25) =>
                           DATA_IN(25), DRAM_DATA_IN(24) => DATA_IN(24), 
                           DRAM_DATA_IN(23) => DATA_IN(23), DRAM_DATA_IN(22) =>
                           DATA_IN(22), DRAM_DATA_IN(21) => DATA_IN(21), 
                           DRAM_DATA_IN(20) => DATA_IN(20), DRAM_DATA_IN(19) =>
                           DATA_IN(19), DRAM_DATA_IN(18) => DATA_IN(18), 
                           DRAM_DATA_IN(17) => DATA_IN(17), DRAM_DATA_IN(16) =>
                           DATA_IN(16), DRAM_DATA_IN(15) => DATA_IN(15), 
                           DRAM_DATA_IN(14) => DATA_IN(14), DRAM_DATA_IN(13) =>
                           DATA_IN(13), DRAM_DATA_IN(12) => DATA_IN(12), 
                           DRAM_DATA_IN(11) => DATA_IN(11), DRAM_DATA_IN(10) =>
                           DATA_IN(10), DRAM_DATA_IN(9) => DATA_IN(9), 
                           DRAM_DATA_IN(8) => DATA_IN(8), DRAM_DATA_IN(7) => 
                           DATA_IN(7), DRAM_DATA_IN(6) => DATA_IN(6), 
                           DRAM_DATA_IN(5) => DATA_IN(5), DRAM_DATA_IN(4) => 
                           DATA_IN(4), DRAM_DATA_IN(3) => DATA_IN(3), 
                           DRAM_DATA_IN(2) => DATA_IN(2), DRAM_DATA_IN(1) => 
                           DATA_IN(1), DRAM_DATA_IN(0) => DATA_IN(0), 
                           PC_OUT(31) => PC_MEM_OUT_31_port, PC_OUT(30) => 
                           PC_MEM_OUT_30_port, PC_OUT(29) => PC_MEM_OUT_29_port
                           , PC_OUT(28) => PC_MEM_OUT_28_port, PC_OUT(27) => 
                           PC_MEM_OUT_27_port, PC_OUT(26) => PC_MEM_OUT_26_port
                           , PC_OUT(25) => PC_MEM_OUT_25_port, PC_OUT(24) => 
                           PC_MEM_OUT_24_port, PC_OUT(23) => PC_MEM_OUT_23_port
                           , PC_OUT(22) => PC_MEM_OUT_22_port, PC_OUT(21) => 
                           PC_MEM_OUT_21_port, PC_OUT(20) => PC_MEM_OUT_20_port
                           , PC_OUT(19) => PC_MEM_OUT_19_port, PC_OUT(18) => 
                           PC_MEM_OUT_18_port, PC_OUT(17) => PC_MEM_OUT_17_port
                           , PC_OUT(16) => PC_MEM_OUT_16_port, PC_OUT(15) => 
                           PC_MEM_OUT_15_port, PC_OUT(14) => PC_MEM_OUT_14_port
                           , PC_OUT(13) => PC_MEM_OUT_13_port, PC_OUT(12) => 
                           PC_MEM_OUT_12_port, PC_OUT(11) => PC_MEM_OUT_11_port
                           , PC_OUT(10) => PC_MEM_OUT_10_port, PC_OUT(9) => 
                           PC_MEM_OUT_9_port, PC_OUT(8) => PC_MEM_OUT_8_port, 
                           PC_OUT(7) => PC_MEM_OUT_7_port, PC_OUT(6) => 
                           PC_MEM_OUT_6_port, PC_OUT(5) => PC_MEM_OUT_5_port, 
                           PC_OUT(4) => PC_MEM_OUT_4_port, PC_OUT(3) => 
                           PC_MEM_OUT_3_port, PC_OUT(2) => PC_MEM_OUT_2_port, 
                           PC_OUT(1) => PC_MEM_OUT_1_port, PC_OUT(0) => 
                           PC_MEM_OUT_0_port, DRAM_EN_OUT => DRAM_EN_OUT, 
                           DRAM_R_OUT => DRAM_R_OUT, DRAM_W_OUT => DRAM_W_OUT, 
                           DRAM_ADDR_OUT(31) => DRAM_ADDR_OUT(31), 
                           DRAM_ADDR_OUT(30) => DRAM_ADDR_OUT(30), 
                           DRAM_ADDR_OUT(29) => DRAM_ADDR_OUT(29), 
                           DRAM_ADDR_OUT(28) => DRAM_ADDR_OUT(28), 
                           DRAM_ADDR_OUT(27) => DRAM_ADDR_OUT(27), 
                           DRAM_ADDR_OUT(26) => DRAM_ADDR_OUT(26), 
                           DRAM_ADDR_OUT(25) => DRAM_ADDR_OUT(25), 
                           DRAM_ADDR_OUT(24) => DRAM_ADDR_OUT(24), 
                           DRAM_ADDR_OUT(23) => DRAM_ADDR_OUT(23), 
                           DRAM_ADDR_OUT(22) => DRAM_ADDR_OUT(22), 
                           DRAM_ADDR_OUT(21) => DRAM_ADDR_OUT(21), 
                           DRAM_ADDR_OUT(20) => DRAM_ADDR_OUT(20), 
                           DRAM_ADDR_OUT(19) => DRAM_ADDR_OUT(19), 
                           DRAM_ADDR_OUT(18) => DRAM_ADDR_OUT(18), 
                           DRAM_ADDR_OUT(17) => DRAM_ADDR_OUT(17), 
                           DRAM_ADDR_OUT(16) => DRAM_ADDR_OUT(16), 
                           DRAM_ADDR_OUT(15) => DRAM_ADDR_OUT(15), 
                           DRAM_ADDR_OUT(14) => DRAM_ADDR_OUT(14), 
                           DRAM_ADDR_OUT(13) => DRAM_ADDR_OUT(13), 
                           DRAM_ADDR_OUT(12) => DRAM_ADDR_OUT(12), 
                           DRAM_ADDR_OUT(11) => DRAM_ADDR_OUT(11), 
                           DRAM_ADDR_OUT(10) => DRAM_ADDR_OUT(10), 
                           DRAM_ADDR_OUT(9) => DRAM_ADDR_OUT(9), 
                           DRAM_ADDR_OUT(8) => DRAM_ADDR_OUT(8), 
                           DRAM_ADDR_OUT(7) => DRAM_ADDR_OUT(7), 
                           DRAM_ADDR_OUT(6) => DRAM_ADDR_OUT(6), 
                           DRAM_ADDR_OUT(5) => DRAM_ADDR_OUT(5), 
                           DRAM_ADDR_OUT(4) => DRAM_ADDR_OUT(4), 
                           DRAM_ADDR_OUT(3) => DRAM_ADDR_OUT(3), 
                           DRAM_ADDR_OUT(2) => DRAM_ADDR_OUT(2), 
                           DRAM_ADDR_OUT(1) => DRAM_ADDR_OUT(1), 
                           DRAM_ADDR_OUT(0) => DRAM_ADDR_OUT(0), 
                           DRAM_DATA_OUT(31) => DATA_OUT(31), DRAM_DATA_OUT(30)
                           => DATA_OUT(30), DRAM_DATA_OUT(29) => DATA_OUT(29), 
                           DRAM_DATA_OUT(28) => DATA_OUT(28), DRAM_DATA_OUT(27)
                           => DATA_OUT(27), DRAM_DATA_OUT(26) => DATA_OUT(26), 
                           DRAM_DATA_OUT(25) => DATA_OUT(25), DRAM_DATA_OUT(24)
                           => DATA_OUT(24), DRAM_DATA_OUT(23) => DATA_OUT(23), 
                           DRAM_DATA_OUT(22) => DATA_OUT(22), DRAM_DATA_OUT(21)
                           => DATA_OUT(21), DRAM_DATA_OUT(20) => DATA_OUT(20), 
                           DRAM_DATA_OUT(19) => DATA_OUT(19), DRAM_DATA_OUT(18)
                           => DATA_OUT(18), DRAM_DATA_OUT(17) => DATA_OUT(17), 
                           DRAM_DATA_OUT(16) => DATA_OUT(16), DRAM_DATA_OUT(15)
                           => DATA_OUT(15), DRAM_DATA_OUT(14) => DATA_OUT(14), 
                           DRAM_DATA_OUT(13) => DATA_OUT(13), DRAM_DATA_OUT(12)
                           => DATA_OUT(12), DRAM_DATA_OUT(11) => DATA_OUT(11), 
                           DRAM_DATA_OUT(10) => DATA_OUT(10), DRAM_DATA_OUT(9) 
                           => DATA_OUT(9), DRAM_DATA_OUT(8) => DATA_OUT(8), 
                           DRAM_DATA_OUT(7) => DATA_OUT(7), DRAM_DATA_OUT(6) =>
                           DATA_OUT(6), DRAM_DATA_OUT(5) => DATA_OUT(5), 
                           DRAM_DATA_OUT(4) => DATA_OUT(4), DRAM_DATA_OUT(3) =>
                           DATA_OUT(3), DRAM_DATA_OUT(2) => DATA_OUT(2), 
                           DRAM_DATA_OUT(1) => DATA_OUT(1), DRAM_DATA_OUT(0) =>
                           DATA_OUT(0), DATA_OUT(31) => DATA_MEM_OUT_31_port, 
                           DATA_OUT(30) => DATA_MEM_OUT_30_port, DATA_OUT(29) 
                           => DATA_MEM_OUT_29_port, DATA_OUT(28) => 
                           DATA_MEM_OUT_28_port, DATA_OUT(27) => 
                           DATA_MEM_OUT_27_port, DATA_OUT(26) => 
                           DATA_MEM_OUT_26_port, DATA_OUT(25) => 
                           DATA_MEM_OUT_25_port, DATA_OUT(24) => 
                           DATA_MEM_OUT_24_port, DATA_OUT(23) => 
                           DATA_MEM_OUT_23_port, DATA_OUT(22) => 
                           DATA_MEM_OUT_22_port, DATA_OUT(21) => 
                           DATA_MEM_OUT_21_port, DATA_OUT(20) => 
                           DATA_MEM_OUT_20_port, DATA_OUT(19) => 
                           DATA_MEM_OUT_19_port, DATA_OUT(18) => 
                           DATA_MEM_OUT_18_port, DATA_OUT(17) => 
                           DATA_MEM_OUT_17_port, DATA_OUT(16) => 
                           DATA_MEM_OUT_16_port, DATA_OUT(15) => 
                           DATA_MEM_OUT_15_port, DATA_OUT(14) => 
                           DATA_MEM_OUT_14_port, DATA_OUT(13) => 
                           DATA_MEM_OUT_13_port, DATA_OUT(12) => 
                           DATA_MEM_OUT_12_port, DATA_OUT(11) => 
                           DATA_MEM_OUT_11_port, DATA_OUT(10) => 
                           DATA_MEM_OUT_10_port, DATA_OUT(9) => 
                           DATA_MEM_OUT_9_port, DATA_OUT(8) => 
                           DATA_MEM_OUT_8_port, DATA_OUT(7) => 
                           DATA_MEM_OUT_7_port, DATA_OUT(6) => 
                           DATA_MEM_OUT_6_port, DATA_OUT(5) => 
                           DATA_MEM_OUT_5_port, DATA_OUT(4) => 
                           DATA_MEM_OUT_4_port, DATA_OUT(3) => 
                           DATA_MEM_OUT_3_port, DATA_OUT(2) => 
                           DATA_MEM_OUT_2_port, DATA_OUT(1) => 
                           DATA_MEM_OUT_1_port, DATA_OUT(0) => 
                           DATA_MEM_OUT_0_port, ALU_RES_OUT(31) => 
                           ALU_RES_MEM_31_port, ALU_RES_OUT(30) => 
                           ALU_RES_MEM_30_port, ALU_RES_OUT(29) => 
                           ALU_RES_MEM_29_port, ALU_RES_OUT(28) => 
                           ALU_RES_MEM_28_port, ALU_RES_OUT(27) => 
                           ALU_RES_MEM_27_port, ALU_RES_OUT(26) => 
                           ALU_RES_MEM_26_port, ALU_RES_OUT(25) => 
                           ALU_RES_MEM_25_port, ALU_RES_OUT(24) => 
                           ALU_RES_MEM_24_port, ALU_RES_OUT(23) => 
                           ALU_RES_MEM_23_port, ALU_RES_OUT(22) => 
                           ALU_RES_MEM_22_port, ALU_RES_OUT(21) => 
                           ALU_RES_MEM_21_port, ALU_RES_OUT(20) => 
                           ALU_RES_MEM_20_port, ALU_RES_OUT(19) => 
                           ALU_RES_MEM_19_port, ALU_RES_OUT(18) => 
                           ALU_RES_MEM_18_port, ALU_RES_OUT(17) => 
                           ALU_RES_MEM_17_port, ALU_RES_OUT(16) => 
                           ALU_RES_MEM_16_port, ALU_RES_OUT(15) => 
                           ALU_RES_MEM_15_port, ALU_RES_OUT(14) => 
                           ALU_RES_MEM_14_port, ALU_RES_OUT(13) => 
                           ALU_RES_MEM_13_port, ALU_RES_OUT(12) => 
                           ALU_RES_MEM_12_port, ALU_RES_OUT(11) => 
                           ALU_RES_MEM_11_port, ALU_RES_OUT(10) => 
                           ALU_RES_MEM_10_port, ALU_RES_OUT(9) => 
                           ALU_RES_MEM_9_port, ALU_RES_OUT(8) => 
                           ALU_RES_MEM_8_port, ALU_RES_OUT(7) => 
                           ALU_RES_MEM_7_port, ALU_RES_OUT(6) => 
                           ALU_RES_MEM_6_port, ALU_RES_OUT(5) => 
                           ALU_RES_MEM_5_port, ALU_RES_OUT(4) => 
                           ALU_RES_MEM_4_port, ALU_RES_OUT(3) => 
                           ALU_RES_MEM_3_port, ALU_RES_OUT(2) => 
                           ALU_RES_MEM_2_port, ALU_RES_OUT(1) => 
                           ALU_RES_MEM_1_port, ALU_RES_OUT(0) => 
                           ALU_RES_MEM_0_port, OP_MEM(31) => OP_MEM_31_port, 
                           OP_MEM(30) => OP_MEM_30_port, OP_MEM(29) => 
                           OP_MEM_29_port, OP_MEM(28) => OP_MEM_28_port, 
                           OP_MEM(27) => OP_MEM_27_port, OP_MEM(26) => 
                           OP_MEM_26_port, OP_MEM(25) => OP_MEM_25_port, 
                           OP_MEM(24) => OP_MEM_24_port, OP_MEM(23) => 
                           OP_MEM_23_port, OP_MEM(22) => OP_MEM_22_port, 
                           OP_MEM(21) => OP_MEM_21_port, OP_MEM(20) => 
                           OP_MEM_20_port, OP_MEM(19) => OP_MEM_19_port, 
                           OP_MEM(18) => OP_MEM_18_port, OP_MEM(17) => 
                           OP_MEM_17_port, OP_MEM(16) => OP_MEM_16_port, 
                           OP_MEM(15) => OP_MEM_15_port, OP_MEM(14) => 
                           OP_MEM_14_port, OP_MEM(13) => OP_MEM_13_port, 
                           OP_MEM(12) => OP_MEM_12_port, OP_MEM(11) => 
                           OP_MEM_11_port, OP_MEM(10) => OP_MEM_10_port, 
                           OP_MEM(9) => OP_MEM_9_port, OP_MEM(8) => 
                           OP_MEM_8_port, OP_MEM(7) => OP_MEM_7_port, OP_MEM(6)
                           => OP_MEM_6_port, OP_MEM(5) => OP_MEM_5_port, 
                           OP_MEM(4) => OP_MEM_4_port, OP_MEM(3) => 
                           OP_MEM_3_port, OP_MEM(2) => OP_MEM_2_port, OP_MEM(1)
                           => OP_MEM_1_port, OP_MEM(0) => OP_MEM_0_port, 
                           ADD_WR_MEM(4) => ADD_WR_MEM_4_port, ADD_WR_MEM(3) =>
                           ADD_WR_MEM_3_port, ADD_WR_MEM(2) => 
                           ADD_WR_MEM_2_port, ADD_WR_MEM(1) => 
                           ADD_WR_MEM_1_port, ADD_WR_MEM(0) => 
                           ADD_WR_MEM_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_MEM_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_MEM_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_MEM_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_MEM_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_MEM_OUT_0_port);
   RF_WE_ff : ff_2 port map( D => RF_WE, CLK => CLK, EN => n1, RST => RST, Q =>
                           RF_WE_WB);
   WritebackStage : Writeback port map( WB_MUX_SEL => WB_MUX_SEL, DATA_IN(31) 
                           => DATA_MEM_OUT_31_port, DATA_IN(30) => 
                           DATA_MEM_OUT_30_port, DATA_IN(29) => 
                           DATA_MEM_OUT_29_port, DATA_IN(28) => 
                           DATA_MEM_OUT_28_port, DATA_IN(27) => 
                           DATA_MEM_OUT_27_port, DATA_IN(26) => 
                           DATA_MEM_OUT_26_port, DATA_IN(25) => 
                           DATA_MEM_OUT_25_port, DATA_IN(24) => 
                           DATA_MEM_OUT_24_port, DATA_IN(23) => 
                           DATA_MEM_OUT_23_port, DATA_IN(22) => 
                           DATA_MEM_OUT_22_port, DATA_IN(21) => 
                           DATA_MEM_OUT_21_port, DATA_IN(20) => 
                           DATA_MEM_OUT_20_port, DATA_IN(19) => 
                           DATA_MEM_OUT_19_port, DATA_IN(18) => 
                           DATA_MEM_OUT_18_port, DATA_IN(17) => 
                           DATA_MEM_OUT_17_port, DATA_IN(16) => 
                           DATA_MEM_OUT_16_port, DATA_IN(15) => 
                           DATA_MEM_OUT_15_port, DATA_IN(14) => 
                           DATA_MEM_OUT_14_port, DATA_IN(13) => 
                           DATA_MEM_OUT_13_port, DATA_IN(12) => 
                           DATA_MEM_OUT_12_port, DATA_IN(11) => 
                           DATA_MEM_OUT_11_port, DATA_IN(10) => 
                           DATA_MEM_OUT_10_port, DATA_IN(9) => 
                           DATA_MEM_OUT_9_port, DATA_IN(8) => 
                           DATA_MEM_OUT_8_port, DATA_IN(7) => 
                           DATA_MEM_OUT_7_port, DATA_IN(6) => 
                           DATA_MEM_OUT_6_port, DATA_IN(5) => 
                           DATA_MEM_OUT_5_port, DATA_IN(4) => 
                           DATA_MEM_OUT_4_port, DATA_IN(3) => 
                           DATA_MEM_OUT_3_port, DATA_IN(2) => 
                           DATA_MEM_OUT_2_port, DATA_IN(1) => 
                           DATA_MEM_OUT_1_port, DATA_IN(0) => 
                           DATA_MEM_OUT_0_port, ALU_RES_IN(31) => 
                           ALU_RES_MEM_31_port, ALU_RES_IN(30) => 
                           ALU_RES_MEM_30_port, ALU_RES_IN(29) => 
                           ALU_RES_MEM_29_port, ALU_RES_IN(28) => 
                           ALU_RES_MEM_28_port, ALU_RES_IN(27) => 
                           ALU_RES_MEM_27_port, ALU_RES_IN(26) => 
                           ALU_RES_MEM_26_port, ALU_RES_IN(25) => 
                           ALU_RES_MEM_25_port, ALU_RES_IN(24) => 
                           ALU_RES_MEM_24_port, ALU_RES_IN(23) => 
                           ALU_RES_MEM_23_port, ALU_RES_IN(22) => 
                           ALU_RES_MEM_22_port, ALU_RES_IN(21) => 
                           ALU_RES_MEM_21_port, ALU_RES_IN(20) => 
                           ALU_RES_MEM_20_port, ALU_RES_IN(19) => 
                           ALU_RES_MEM_19_port, ALU_RES_IN(18) => 
                           ALU_RES_MEM_18_port, ALU_RES_IN(17) => 
                           ALU_RES_MEM_17_port, ALU_RES_IN(16) => 
                           ALU_RES_MEM_16_port, ALU_RES_IN(15) => 
                           ALU_RES_MEM_15_port, ALU_RES_IN(14) => 
                           ALU_RES_MEM_14_port, ALU_RES_IN(13) => 
                           ALU_RES_MEM_13_port, ALU_RES_IN(12) => 
                           ALU_RES_MEM_12_port, ALU_RES_IN(11) => 
                           ALU_RES_MEM_11_port, ALU_RES_IN(10) => 
                           ALU_RES_MEM_10_port, ALU_RES_IN(9) => 
                           ALU_RES_MEM_9_port, ALU_RES_IN(8) => 
                           ALU_RES_MEM_8_port, ALU_RES_IN(7) => 
                           ALU_RES_MEM_7_port, ALU_RES_IN(6) => 
                           ALU_RES_MEM_6_port, ALU_RES_IN(5) => 
                           ALU_RES_MEM_5_port, ALU_RES_IN(4) => 
                           ALU_RES_MEM_4_port, ALU_RES_IN(3) => 
                           ALU_RES_MEM_3_port, ALU_RES_IN(2) => 
                           ALU_RES_MEM_2_port, ALU_RES_IN(1) => 
                           ALU_RES_MEM_1_port, ALU_RES_IN(0) => 
                           ALU_RES_MEM_0_port, ADD_WR_IN(4) => 
                           ADD_WR_MEM_OUT_4_port, ADD_WR_IN(3) => 
                           ADD_WR_MEM_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_MEM_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_MEM_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_MEM_OUT_0_port, DATA_OUT(31) => OP_WB_31_port
                           , DATA_OUT(30) => OP_WB_30_port, DATA_OUT(29) => 
                           OP_WB_29_port, DATA_OUT(28) => OP_WB_28_port, 
                           DATA_OUT(27) => OP_WB_27_port, DATA_OUT(26) => 
                           OP_WB_26_port, DATA_OUT(25) => OP_WB_25_port, 
                           DATA_OUT(24) => OP_WB_24_port, DATA_OUT(23) => 
                           OP_WB_23_port, DATA_OUT(22) => OP_WB_22_port, 
                           DATA_OUT(21) => OP_WB_21_port, DATA_OUT(20) => 
                           OP_WB_20_port, DATA_OUT(19) => OP_WB_19_port, 
                           DATA_OUT(18) => OP_WB_18_port, DATA_OUT(17) => 
                           OP_WB_17_port, DATA_OUT(16) => OP_WB_16_port, 
                           DATA_OUT(15) => OP_WB_15_port, DATA_OUT(14) => 
                           OP_WB_14_port, DATA_OUT(13) => OP_WB_13_port, 
                           DATA_OUT(12) => OP_WB_12_port, DATA_OUT(11) => 
                           OP_WB_11_port, DATA_OUT(10) => OP_WB_10_port, 
                           DATA_OUT(9) => OP_WB_9_port, DATA_OUT(8) => 
                           OP_WB_8_port, DATA_OUT(7) => OP_WB_7_port, 
                           DATA_OUT(6) => OP_WB_6_port, DATA_OUT(5) => 
                           OP_WB_5_port, DATA_OUT(4) => OP_WB_4_port, 
                           DATA_OUT(3) => OP_WB_3_port, DATA_OUT(2) => 
                           OP_WB_2_port, DATA_OUT(1) => OP_WB_1_port, 
                           DATA_OUT(0) => OP_WB_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_WB_4_port, ADD_WR_OUT(3) => ADD_WR_WB_3_port,
                           ADD_WR_OUT(2) => ADD_WR_WB_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_WB_1_port, ADD_WR_OUT(0) => ADD_WR_WB_0_port)
                           ;
   HDU : HazardDetection port map( RST => RST, ADD_RS1(4) => ADD_RS1_HDU_4_port
                           , ADD_RS1(3) => ADD_RS1_HDU_3_port, ADD_RS1(2) => 
                           ADD_RS1_HDU_2_port, ADD_RS1(1) => ADD_RS1_HDU_1_port
                           , ADD_RS1(0) => ADD_RS1_HDU_0_port, ADD_RS2(4) => 
                           ADD_RS2_HDU_4_port, ADD_RS2(3) => ADD_RS2_HDU_3_port
                           , ADD_RS2(2) => ADD_RS2_HDU_2_port, ADD_RS2(1) => 
                           ADD_RS2_HDU_1_port, ADD_RS2(0) => ADD_RS2_HDU_0_port
                           , ADD_WR(4) => ADD_WR_DECODE_OUT_4_port, ADD_WR(3) 
                           => ADD_WR_DECODE_OUT_3_port, ADD_WR(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR(0) => 
                           ADD_WR_DECODE_OUT_0_port, DRAM_R => DRAM_R_IN, 
                           INS_IN(31) => INS_OUT_31_port, INS_IN(30) => 
                           INS_OUT_30_port, INS_IN(29) => INS_OUT_29_port, 
                           INS_IN(28) => INS_OUT_28_port, INS_IN(27) => 
                           INS_OUT_27_port, INS_IN(26) => INS_OUT_26_port, 
                           INS_IN(25) => INS_OUT_25_port, INS_IN(24) => 
                           INS_OUT_24_port, INS_IN(23) => INS_OUT_23_port, 
                           INS_IN(22) => INS_OUT_22_port, INS_IN(21) => 
                           INS_OUT_21_port, INS_IN(20) => INS_OUT_20_port, 
                           INS_IN(19) => INS_OUT_19_port, INS_IN(18) => 
                           INS_OUT_18_port, INS_IN(17) => INS_OUT_17_port, 
                           INS_IN(16) => INS_OUT_16_port, INS_IN(15) => 
                           INS_OUT_15_port, INS_IN(14) => INS_OUT_14_port, 
                           INS_IN(13) => INS_OUT_13_port, INS_IN(12) => 
                           INS_OUT_12_port, INS_IN(11) => INS_OUT_11_port, 
                           INS_IN(10) => INS_OUT_10_port, INS_IN(9) => 
                           INS_OUT_9_port, INS_IN(8) => INS_OUT_8_port, 
                           INS_IN(7) => INS_OUT_7_port, INS_IN(6) => 
                           INS_OUT_6_port, INS_IN(5) => INS_OUT_5_port, 
                           INS_IN(4) => INS_OUT_4_port, INS_IN(3) => 
                           INS_OUT_3_port, INS_IN(2) => INS_OUT_2_port, 
                           INS_IN(1) => INS_OUT_1_port, INS_IN(0) => 
                           INS_OUT_0_port, PC_IN(31) => PC_FETCH_OUT_31_port, 
                           PC_IN(30) => PC_FETCH_OUT_30_port, PC_IN(29) => 
                           PC_FETCH_OUT_29_port, PC_IN(28) => 
                           PC_FETCH_OUT_28_port, PC_IN(27) => 
                           PC_FETCH_OUT_27_port, PC_IN(26) => 
                           PC_FETCH_OUT_26_port, PC_IN(25) => 
                           PC_FETCH_OUT_25_port, PC_IN(24) => 
                           PC_FETCH_OUT_24_port, PC_IN(23) => 
                           PC_FETCH_OUT_23_port, PC_IN(22) => 
                           PC_FETCH_OUT_22_port, PC_IN(21) => 
                           PC_FETCH_OUT_21_port, PC_IN(20) => 
                           PC_FETCH_OUT_20_port, PC_IN(19) => 
                           PC_FETCH_OUT_19_port, PC_IN(18) => 
                           PC_FETCH_OUT_18_port, PC_IN(17) => 
                           PC_FETCH_OUT_17_port, PC_IN(16) => 
                           PC_FETCH_OUT_16_port, PC_IN(15) => 
                           PC_FETCH_OUT_15_port, PC_IN(14) => 
                           PC_FETCH_OUT_14_port, PC_IN(13) => 
                           PC_FETCH_OUT_13_port, PC_IN(12) => 
                           PC_FETCH_OUT_12_port, PC_IN(11) => 
                           PC_FETCH_OUT_11_port, PC_IN(10) => 
                           PC_FETCH_OUT_10_port, PC_IN(9) => 
                           PC_FETCH_OUT_9_port, PC_IN(8) => PC_FETCH_OUT_8_port
                           , PC_IN(7) => PC_FETCH_OUT_7_port, PC_IN(6) => 
                           PC_FETCH_OUT_6_port, PC_IN(5) => PC_FETCH_OUT_5_port
                           , PC_IN(4) => PC_FETCH_OUT_4_port, PC_IN(3) => 
                           PC_FETCH_OUT_3_port, PC_IN(2) => PC_FETCH_OUT_2_port
                           , PC_IN(1) => PC_FETCH_OUT_1_port, PC_IN(0) => 
                           PC_FETCH_OUT_0_port, Bubble => Bubble_out_port, 
                           HDU_INS_OUT(31) => sig_HDU_INS_OUT_31_port, 
                           HDU_INS_OUT(30) => sig_HDU_INS_OUT_30_port, 
                           HDU_INS_OUT(29) => sig_HDU_INS_OUT_29_port, 
                           HDU_INS_OUT(28) => sig_HDU_INS_OUT_28_port, 
                           HDU_INS_OUT(27) => sig_HDU_INS_OUT_27_port, 
                           HDU_INS_OUT(26) => sig_HDU_INS_OUT_26_port, 
                           HDU_INS_OUT(25) => sig_HDU_INS_OUT_25_port, 
                           HDU_INS_OUT(24) => sig_HDU_INS_OUT_24_port, 
                           HDU_INS_OUT(23) => sig_HDU_INS_OUT_23_port, 
                           HDU_INS_OUT(22) => sig_HDU_INS_OUT_22_port, 
                           HDU_INS_OUT(21) => sig_HDU_INS_OUT_21_port, 
                           HDU_INS_OUT(20) => sig_HDU_INS_OUT_20_port, 
                           HDU_INS_OUT(19) => sig_HDU_INS_OUT_19_port, 
                           HDU_INS_OUT(18) => sig_HDU_INS_OUT_18_port, 
                           HDU_INS_OUT(17) => sig_HDU_INS_OUT_17_port, 
                           HDU_INS_OUT(16) => sig_HDU_INS_OUT_16_port, 
                           HDU_INS_OUT(15) => sig_HDU_INS_OUT_15_port, 
                           HDU_INS_OUT(14) => sig_HDU_INS_OUT_14_port, 
                           HDU_INS_OUT(13) => sig_HDU_INS_OUT_13_port, 
                           HDU_INS_OUT(12) => sig_HDU_INS_OUT_12_port, 
                           HDU_INS_OUT(11) => sig_HDU_INS_OUT_11_port, 
                           HDU_INS_OUT(10) => sig_HDU_INS_OUT_10_port, 
                           HDU_INS_OUT(9) => sig_HDU_INS_OUT_9_port, 
                           HDU_INS_OUT(8) => sig_HDU_INS_OUT_8_port, 
                           HDU_INS_OUT(7) => sig_HDU_INS_OUT_7_port, 
                           HDU_INS_OUT(6) => sig_HDU_INS_OUT_6_port, 
                           HDU_INS_OUT(5) => sig_HDU_INS_OUT_5_port, 
                           HDU_INS_OUT(4) => sig_HDU_INS_OUT_4_port, 
                           HDU_INS_OUT(3) => sig_HDU_INS_OUT_3_port, 
                           HDU_INS_OUT(2) => sig_HDU_INS_OUT_2_port, 
                           HDU_INS_OUT(1) => sig_HDU_INS_OUT_1_port, 
                           HDU_INS_OUT(0) => sig_HDU_INS_OUT_0_port, 
                           HDU_PC_OUT(31) => sig_HDU_PC_OUT_31_port, 
                           HDU_PC_OUT(30) => sig_HDU_PC_OUT_30_port, 
                           HDU_PC_OUT(29) => sig_HDU_PC_OUT_29_port, 
                           HDU_PC_OUT(28) => sig_HDU_PC_OUT_28_port, 
                           HDU_PC_OUT(27) => sig_HDU_PC_OUT_27_port, 
                           HDU_PC_OUT(26) => sig_HDU_PC_OUT_26_port, 
                           HDU_PC_OUT(25) => sig_HDU_PC_OUT_25_port, 
                           HDU_PC_OUT(24) => sig_HDU_PC_OUT_24_port, 
                           HDU_PC_OUT(23) => sig_HDU_PC_OUT_23_port, 
                           HDU_PC_OUT(22) => sig_HDU_PC_OUT_22_port, 
                           HDU_PC_OUT(21) => sig_HDU_PC_OUT_21_port, 
                           HDU_PC_OUT(20) => sig_HDU_PC_OUT_20_port, 
                           HDU_PC_OUT(19) => sig_HDU_PC_OUT_19_port, 
                           HDU_PC_OUT(18) => sig_HDU_PC_OUT_18_port, 
                           HDU_PC_OUT(17) => sig_HDU_PC_OUT_17_port, 
                           HDU_PC_OUT(16) => sig_HDU_PC_OUT_16_port, 
                           HDU_PC_OUT(15) => sig_HDU_PC_OUT_15_port, 
                           HDU_PC_OUT(14) => sig_HDU_PC_OUT_14_port, 
                           HDU_PC_OUT(13) => sig_HDU_PC_OUT_13_port, 
                           HDU_PC_OUT(12) => sig_HDU_PC_OUT_12_port, 
                           HDU_PC_OUT(11) => sig_HDU_PC_OUT_11_port, 
                           HDU_PC_OUT(10) => sig_HDU_PC_OUT_10_port, 
                           HDU_PC_OUT(9) => sig_HDU_PC_OUT_9_port, 
                           HDU_PC_OUT(8) => sig_HDU_PC_OUT_8_port, 
                           HDU_PC_OUT(7) => sig_HDU_PC_OUT_7_port, 
                           HDU_PC_OUT(6) => sig_HDU_PC_OUT_6_port, 
                           HDU_PC_OUT(5) => sig_HDU_PC_OUT_5_port, 
                           HDU_PC_OUT(4) => sig_HDU_PC_OUT_4_port, 
                           HDU_PC_OUT(3) => sig_HDU_PC_OUT_3_port, 
                           HDU_PC_OUT(2) => sig_HDU_PC_OUT_2_port, 
                           HDU_PC_OUT(1) => sig_HDU_PC_OUT_1_port, 
                           HDU_PC_OUT(0) => sig_HDU_PC_OUT_0_port, 
                           HDU_NPC_OUT(31) => sig_HDU_NPC_OUT_31_port, 
                           HDU_NPC_OUT(30) => sig_HDU_NPC_OUT_30_port, 
                           HDU_NPC_OUT(29) => sig_HDU_NPC_OUT_29_port, 
                           HDU_NPC_OUT(28) => sig_HDU_NPC_OUT_28_port, 
                           HDU_NPC_OUT(27) => sig_HDU_NPC_OUT_27_port, 
                           HDU_NPC_OUT(26) => sig_HDU_NPC_OUT_26_port, 
                           HDU_NPC_OUT(25) => sig_HDU_NPC_OUT_25_port, 
                           HDU_NPC_OUT(24) => sig_HDU_NPC_OUT_24_port, 
                           HDU_NPC_OUT(23) => sig_HDU_NPC_OUT_23_port, 
                           HDU_NPC_OUT(22) => sig_HDU_NPC_OUT_22_port, 
                           HDU_NPC_OUT(21) => sig_HDU_NPC_OUT_21_port, 
                           HDU_NPC_OUT(20) => sig_HDU_NPC_OUT_20_port, 
                           HDU_NPC_OUT(19) => sig_HDU_NPC_OUT_19_port, 
                           HDU_NPC_OUT(18) => sig_HDU_NPC_OUT_18_port, 
                           HDU_NPC_OUT(17) => sig_HDU_NPC_OUT_17_port, 
                           HDU_NPC_OUT(16) => sig_HDU_NPC_OUT_16_port, 
                           HDU_NPC_OUT(15) => sig_HDU_NPC_OUT_15_port, 
                           HDU_NPC_OUT(14) => sig_HDU_NPC_OUT_14_port, 
                           HDU_NPC_OUT(13) => sig_HDU_NPC_OUT_13_port, 
                           HDU_NPC_OUT(12) => sig_HDU_NPC_OUT_12_port, 
                           HDU_NPC_OUT(11) => sig_HDU_NPC_OUT_11_port, 
                           HDU_NPC_OUT(10) => sig_HDU_NPC_OUT_10_port, 
                           HDU_NPC_OUT(9) => sig_HDU_NPC_OUT_9_port, 
                           HDU_NPC_OUT(8) => sig_HDU_NPC_OUT_8_port, 
                           HDU_NPC_OUT(7) => sig_HDU_NPC_OUT_7_port, 
                           HDU_NPC_OUT(6) => sig_HDU_NPC_OUT_6_port, 
                           HDU_NPC_OUT(5) => sig_HDU_NPC_OUT_5_port, 
                           HDU_NPC_OUT(4) => sig_HDU_NPC_OUT_4_port, 
                           HDU_NPC_OUT(3) => sig_HDU_NPC_OUT_3_port, 
                           HDU_NPC_OUT(2) => sig_HDU_NPC_OUT_2_port, 
                           HDU_NPC_OUT(1) => sig_HDU_NPC_OUT_1_port, 
                           HDU_NPC_OUT(0) => sig_HDU_NPC_OUT_0_port);
   n1 <= '1';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( Clk, Rst : in std_logic);

end DLX;

architecture SYN_dlx_rtl of DLX is

   component DRAM
      port( En, Rst : in std_logic;  ADDR_IN, DATA_IN : in std_logic_vector (31
            downto 0);  DRAM_W, DRAM_R : in std_logic;  DATA_OUT : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component IRAM
      port( Rst : in std_logic;  Addr : in std_logic_vector (31 downto 0);  
            Iout : out std_logic_vector (31 downto 0));
   end component;
   
   component hardwired_cu_NBIT32
      port( REG_LATCH_EN, RD1, RD2, MUX_A_SEL : out std_logic;  MUX_B_SEL : out
            std_logic_vector (1 downto 0);  ALU_OPC : out std_logic_vector (0 
            to 3);  ALU_OUTREG_EN, DRAM_R_IN : out std_logic;  JUMP_TYPE : out 
            std_logic_vector (1 downto 0);  MEM_EN_IN, DRAM_W_IN, RF_WE, 
            DRAM_EN_IN, WB_MUX_SEL : out std_logic;  INS_IN : in 
            std_logic_vector (31 downto 0);  Bubble, Clk, Rst : in std_logic);
   end component;
   
   component Datapath
      port( CLK, RST : in std_logic;  INS_IN, DATA_IN : in std_logic_vector (31
            downto 0);  REG_LATCH_EN, RD1, RD2, MUX_A_SEL : in std_logic;  
            MUX_B_SEL : in std_logic_vector (1 downto 0);  ALU_OPC : in 
            std_logic_vector (0 to 3);  ALU_OUTREG_EN : in std_logic;  
            JUMP_TYPE : in std_logic_vector (1 downto 0);  DRAM_R_IN, MEM_EN_IN
            , DRAM_W_IN, RF_WE, DRAM_EN_IN, WB_MUX_SEL : in std_logic;  INS_OUT
            , IRAM_ADDR_OUT, DRAM_ADDR_OUT, DATA_OUT : out std_logic_vector (31
            downto 0);  DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble_out : out 
            std_logic);
   end component;
   
   signal INS_IN_31_port, INS_IN_30_port, INS_IN_29_port, INS_IN_28_port, 
      INS_IN_27_port, INS_IN_26_port, INS_IN_25_port, INS_IN_24_port, 
      INS_IN_23_port, INS_IN_22_port, INS_IN_21_port, INS_IN_20_port, 
      INS_IN_19_port, INS_IN_18_port, INS_IN_17_port, INS_IN_16_port, 
      INS_IN_15_port, INS_IN_14_port, INS_IN_13_port, INS_IN_12_port, 
      INS_IN_11_port, INS_IN_10_port, INS_IN_9_port, INS_IN_8_port, 
      INS_IN_7_port, INS_IN_6_port, INS_IN_5_port, INS_IN_4_port, INS_IN_3_port
      , INS_IN_2_port, INS_IN_1_port, INS_IN_0_port, DATA_IN_31_port, 
      DATA_IN_30_port, DATA_IN_29_port, DATA_IN_28_port, DATA_IN_27_port, 
      DATA_IN_26_port, DATA_IN_25_port, DATA_IN_24_port, DATA_IN_23_port, 
      DATA_IN_22_port, DATA_IN_21_port, DATA_IN_20_port, DATA_IN_19_port, 
      DATA_IN_18_port, DATA_IN_17_port, DATA_IN_16_port, DATA_IN_15_port, 
      DATA_IN_14_port, DATA_IN_13_port, DATA_IN_12_port, DATA_IN_11_port, 
      DATA_IN_10_port, DATA_IN_9_port, DATA_IN_8_port, DATA_IN_7_port, 
      DATA_IN_6_port, DATA_IN_5_port, DATA_IN_4_port, DATA_IN_3_port, 
      DATA_IN_2_port, DATA_IN_1_port, DATA_IN_0_port, REG_LATCH_EN, RD1, RD2, 
      MUX_A_SEL, MUX_B_SEL_1_port, MUX_B_SEL_0_port, ALU_OPC_3_port, 
      ALU_OPC_2_port, ALU_OPC_1_port, ALU_OPC_0_port, ALU_OUTREG_EN, 
      JUMP_TYPE_1_port, JUMP_TYPE_0_port, DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, 
      RF_WE, DRAM_EN_IN, WB_MUX_SEL, IRAM_ADDR_OUT_31_port, 
      IRAM_ADDR_OUT_30_port, IRAM_ADDR_OUT_29_port, IRAM_ADDR_OUT_28_port, 
      IRAM_ADDR_OUT_27_port, IRAM_ADDR_OUT_26_port, IRAM_ADDR_OUT_25_port, 
      IRAM_ADDR_OUT_24_port, IRAM_ADDR_OUT_23_port, IRAM_ADDR_OUT_22_port, 
      IRAM_ADDR_OUT_21_port, IRAM_ADDR_OUT_20_port, IRAM_ADDR_OUT_19_port, 
      IRAM_ADDR_OUT_18_port, IRAM_ADDR_OUT_17_port, IRAM_ADDR_OUT_16_port, 
      IRAM_ADDR_OUT_15_port, IRAM_ADDR_OUT_14_port, IRAM_ADDR_OUT_13_port, 
      IRAM_ADDR_OUT_12_port, IRAM_ADDR_OUT_11_port, IRAM_ADDR_OUT_10_port, 
      IRAM_ADDR_OUT_9_port, IRAM_ADDR_OUT_8_port, IRAM_ADDR_OUT_7_port, 
      IRAM_ADDR_OUT_6_port, IRAM_ADDR_OUT_5_port, IRAM_ADDR_OUT_4_port, 
      IRAM_ADDR_OUT_3_port, IRAM_ADDR_OUT_2_port, IRAM_ADDR_OUT_1_port, 
      IRAM_ADDR_OUT_0_port, DRAM_ADDR_OUT_31_port, DRAM_ADDR_OUT_30_port, 
      DRAM_ADDR_OUT_29_port, DRAM_ADDR_OUT_28_port, DRAM_ADDR_OUT_27_port, 
      DRAM_ADDR_OUT_26_port, DRAM_ADDR_OUT_25_port, DRAM_ADDR_OUT_24_port, 
      DRAM_ADDR_OUT_23_port, DRAM_ADDR_OUT_22_port, DRAM_ADDR_OUT_21_port, 
      DRAM_ADDR_OUT_20_port, DRAM_ADDR_OUT_19_port, DRAM_ADDR_OUT_18_port, 
      DRAM_ADDR_OUT_17_port, DRAM_ADDR_OUT_16_port, DRAM_ADDR_OUT_15_port, 
      DRAM_ADDR_OUT_14_port, DRAM_ADDR_OUT_13_port, DRAM_ADDR_OUT_12_port, 
      DRAM_ADDR_OUT_11_port, DRAM_ADDR_OUT_10_port, DRAM_ADDR_OUT_9_port, 
      DRAM_ADDR_OUT_8_port, DRAM_ADDR_OUT_7_port, DRAM_ADDR_OUT_6_port, 
      DRAM_ADDR_OUT_5_port, DRAM_ADDR_OUT_4_port, DRAM_ADDR_OUT_3_port, 
      DRAM_ADDR_OUT_2_port, DRAM_ADDR_OUT_1_port, DRAM_ADDR_OUT_0_port, 
      DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, DATA_OUT_28_port, 
      DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, DATA_OUT_24_port, 
      DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, DATA_OUT_20_port, 
      DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, DATA_OUT_16_port, 
      DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, DATA_OUT_12_port, 
      DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, DATA_OUT_8_port, 
      DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, DATA_OUT_4_port, 
      DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, DATA_OUT_0_port, 
      DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble, n_1182, n_1183, n_1184, 
      n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, 
      n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, 
      n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, 
      n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, 
      n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228 : 
      std_logic;

begin
   
   DP : Datapath port map( CLK => Clk, RST => Rst, INS_IN(31) => INS_IN_31_port
                           , INS_IN(30) => INS_IN_30_port, INS_IN(29) => 
                           INS_IN_29_port, INS_IN(28) => INS_IN_28_port, 
                           INS_IN(27) => INS_IN_27_port, INS_IN(26) => 
                           INS_IN_26_port, INS_IN(25) => INS_IN_25_port, 
                           INS_IN(24) => INS_IN_24_port, INS_IN(23) => 
                           INS_IN_23_port, INS_IN(22) => INS_IN_22_port, 
                           INS_IN(21) => INS_IN_21_port, INS_IN(20) => 
                           INS_IN_20_port, INS_IN(19) => INS_IN_19_port, 
                           INS_IN(18) => INS_IN_18_port, INS_IN(17) => 
                           INS_IN_17_port, INS_IN(16) => INS_IN_16_port, 
                           INS_IN(15) => INS_IN_15_port, INS_IN(14) => 
                           INS_IN_14_port, INS_IN(13) => INS_IN_13_port, 
                           INS_IN(12) => INS_IN_12_port, INS_IN(11) => 
                           INS_IN_11_port, INS_IN(10) => INS_IN_10_port, 
                           INS_IN(9) => INS_IN_9_port, INS_IN(8) => 
                           INS_IN_8_port, INS_IN(7) => INS_IN_7_port, INS_IN(6)
                           => INS_IN_6_port, INS_IN(5) => INS_IN_5_port, 
                           INS_IN(4) => INS_IN_4_port, INS_IN(3) => 
                           INS_IN_3_port, INS_IN(2) => INS_IN_2_port, INS_IN(1)
                           => INS_IN_1_port, INS_IN(0) => INS_IN_0_port, 
                           DATA_IN(31) => DATA_IN_31_port, DATA_IN(30) => 
                           DATA_IN_30_port, DATA_IN(29) => DATA_IN_29_port, 
                           DATA_IN(28) => DATA_IN_28_port, DATA_IN(27) => 
                           DATA_IN_27_port, DATA_IN(26) => DATA_IN_26_port, 
                           DATA_IN(25) => DATA_IN_25_port, DATA_IN(24) => 
                           DATA_IN_24_port, DATA_IN(23) => DATA_IN_23_port, 
                           DATA_IN(22) => DATA_IN_22_port, DATA_IN(21) => 
                           DATA_IN_21_port, DATA_IN(20) => DATA_IN_20_port, 
                           DATA_IN(19) => DATA_IN_19_port, DATA_IN(18) => 
                           DATA_IN_18_port, DATA_IN(17) => DATA_IN_17_port, 
                           DATA_IN(16) => DATA_IN_16_port, DATA_IN(15) => 
                           DATA_IN_15_port, DATA_IN(14) => DATA_IN_14_port, 
                           DATA_IN(13) => DATA_IN_13_port, DATA_IN(12) => 
                           DATA_IN_12_port, DATA_IN(11) => DATA_IN_11_port, 
                           DATA_IN(10) => DATA_IN_10_port, DATA_IN(9) => 
                           DATA_IN_9_port, DATA_IN(8) => DATA_IN_8_port, 
                           DATA_IN(7) => DATA_IN_7_port, DATA_IN(6) => 
                           DATA_IN_6_port, DATA_IN(5) => DATA_IN_5_port, 
                           DATA_IN(4) => DATA_IN_4_port, DATA_IN(3) => 
                           DATA_IN_3_port, DATA_IN(2) => DATA_IN_2_port, 
                           DATA_IN(1) => DATA_IN_1_port, DATA_IN(0) => 
                           DATA_IN_0_port, REG_LATCH_EN => REG_LATCH_EN, RD1 =>
                           RD1, RD2 => RD2, MUX_A_SEL => MUX_A_SEL, 
                           MUX_B_SEL(1) => MUX_B_SEL_1_port, MUX_B_SEL(0) => 
                           MUX_B_SEL_0_port, ALU_OPC(0) => ALU_OPC_3_port, 
                           ALU_OPC(1) => ALU_OPC_2_port, ALU_OPC(2) => 
                           ALU_OPC_1_port, ALU_OPC(3) => ALU_OPC_0_port, 
                           ALU_OUTREG_EN => ALU_OUTREG_EN, JUMP_TYPE(1) => 
                           JUMP_TYPE_1_port, JUMP_TYPE(0) => JUMP_TYPE_0_port, 
                           DRAM_R_IN => DRAM_R_IN, MEM_EN_IN => MEM_EN_IN, 
                           DRAM_W_IN => DRAM_W_IN, RF_WE => RF_WE, DRAM_EN_IN 
                           => DRAM_EN_IN, WB_MUX_SEL => WB_MUX_SEL, INS_OUT(31)
                           => n_1182, INS_OUT(30) => n_1183, INS_OUT(29) => 
                           n_1184, INS_OUT(28) => n_1185, INS_OUT(27) => n_1186
                           , INS_OUT(26) => n_1187, INS_OUT(25) => n_1188, 
                           INS_OUT(24) => n_1189, INS_OUT(23) => n_1190, 
                           INS_OUT(22) => n_1191, INS_OUT(21) => n_1192, 
                           INS_OUT(20) => n_1193, INS_OUT(19) => n_1194, 
                           INS_OUT(18) => n_1195, INS_OUT(17) => n_1196, 
                           INS_OUT(16) => n_1197, INS_OUT(15) => n_1198, 
                           INS_OUT(14) => n_1199, INS_OUT(13) => n_1200, 
                           INS_OUT(12) => n_1201, INS_OUT(11) => n_1202, 
                           INS_OUT(10) => n_1203, INS_OUT(9) => n_1204, 
                           INS_OUT(8) => n_1205, INS_OUT(7) => n_1206, 
                           INS_OUT(6) => n_1207, INS_OUT(5) => n_1208, 
                           INS_OUT(4) => n_1209, INS_OUT(3) => n_1210, 
                           INS_OUT(2) => n_1211, INS_OUT(1) => n_1212, 
                           INS_OUT(0) => n_1213, IRAM_ADDR_OUT(31) => 
                           IRAM_ADDR_OUT_31_port, IRAM_ADDR_OUT(30) => 
                           IRAM_ADDR_OUT_30_port, IRAM_ADDR_OUT(29) => 
                           IRAM_ADDR_OUT_29_port, IRAM_ADDR_OUT(28) => 
                           IRAM_ADDR_OUT_28_port, IRAM_ADDR_OUT(27) => 
                           IRAM_ADDR_OUT_27_port, IRAM_ADDR_OUT(26) => 
                           IRAM_ADDR_OUT_26_port, IRAM_ADDR_OUT(25) => 
                           IRAM_ADDR_OUT_25_port, IRAM_ADDR_OUT(24) => 
                           IRAM_ADDR_OUT_24_port, IRAM_ADDR_OUT(23) => 
                           IRAM_ADDR_OUT_23_port, IRAM_ADDR_OUT(22) => 
                           IRAM_ADDR_OUT_22_port, IRAM_ADDR_OUT(21) => 
                           IRAM_ADDR_OUT_21_port, IRAM_ADDR_OUT(20) => 
                           IRAM_ADDR_OUT_20_port, IRAM_ADDR_OUT(19) => 
                           IRAM_ADDR_OUT_19_port, IRAM_ADDR_OUT(18) => 
                           IRAM_ADDR_OUT_18_port, IRAM_ADDR_OUT(17) => 
                           IRAM_ADDR_OUT_17_port, IRAM_ADDR_OUT(16) => 
                           IRAM_ADDR_OUT_16_port, IRAM_ADDR_OUT(15) => 
                           IRAM_ADDR_OUT_15_port, IRAM_ADDR_OUT(14) => 
                           IRAM_ADDR_OUT_14_port, IRAM_ADDR_OUT(13) => 
                           IRAM_ADDR_OUT_13_port, IRAM_ADDR_OUT(12) => 
                           IRAM_ADDR_OUT_12_port, IRAM_ADDR_OUT(11) => 
                           IRAM_ADDR_OUT_11_port, IRAM_ADDR_OUT(10) => 
                           IRAM_ADDR_OUT_10_port, IRAM_ADDR_OUT(9) => 
                           IRAM_ADDR_OUT_9_port, IRAM_ADDR_OUT(8) => 
                           IRAM_ADDR_OUT_8_port, IRAM_ADDR_OUT(7) => 
                           IRAM_ADDR_OUT_7_port, IRAM_ADDR_OUT(6) => 
                           IRAM_ADDR_OUT_6_port, IRAM_ADDR_OUT(5) => 
                           IRAM_ADDR_OUT_5_port, IRAM_ADDR_OUT(4) => 
                           IRAM_ADDR_OUT_4_port, IRAM_ADDR_OUT(3) => 
                           IRAM_ADDR_OUT_3_port, IRAM_ADDR_OUT(2) => 
                           IRAM_ADDR_OUT_2_port, IRAM_ADDR_OUT(1) => 
                           IRAM_ADDR_OUT_1_port, IRAM_ADDR_OUT(0) => 
                           IRAM_ADDR_OUT_0_port, DRAM_ADDR_OUT(31) => 
                           DRAM_ADDR_OUT_31_port, DRAM_ADDR_OUT(30) => 
                           DRAM_ADDR_OUT_30_port, DRAM_ADDR_OUT(29) => 
                           DRAM_ADDR_OUT_29_port, DRAM_ADDR_OUT(28) => 
                           DRAM_ADDR_OUT_28_port, DRAM_ADDR_OUT(27) => 
                           DRAM_ADDR_OUT_27_port, DRAM_ADDR_OUT(26) => 
                           DRAM_ADDR_OUT_26_port, DRAM_ADDR_OUT(25) => 
                           DRAM_ADDR_OUT_25_port, DRAM_ADDR_OUT(24) => 
                           DRAM_ADDR_OUT_24_port, DRAM_ADDR_OUT(23) => 
                           DRAM_ADDR_OUT_23_port, DRAM_ADDR_OUT(22) => 
                           DRAM_ADDR_OUT_22_port, DRAM_ADDR_OUT(21) => 
                           DRAM_ADDR_OUT_21_port, DRAM_ADDR_OUT(20) => 
                           DRAM_ADDR_OUT_20_port, DRAM_ADDR_OUT(19) => 
                           DRAM_ADDR_OUT_19_port, DRAM_ADDR_OUT(18) => 
                           DRAM_ADDR_OUT_18_port, DRAM_ADDR_OUT(17) => 
                           DRAM_ADDR_OUT_17_port, DRAM_ADDR_OUT(16) => 
                           DRAM_ADDR_OUT_16_port, DRAM_ADDR_OUT(15) => 
                           DRAM_ADDR_OUT_15_port, DRAM_ADDR_OUT(14) => 
                           DRAM_ADDR_OUT_14_port, DRAM_ADDR_OUT(13) => 
                           DRAM_ADDR_OUT_13_port, DRAM_ADDR_OUT(12) => 
                           DRAM_ADDR_OUT_12_port, DRAM_ADDR_OUT(11) => 
                           DRAM_ADDR_OUT_11_port, DRAM_ADDR_OUT(10) => 
                           DRAM_ADDR_OUT_10_port, DRAM_ADDR_OUT(9) => 
                           DRAM_ADDR_OUT_9_port, DRAM_ADDR_OUT(8) => 
                           DRAM_ADDR_OUT_8_port, DRAM_ADDR_OUT(7) => 
                           DRAM_ADDR_OUT_7_port, DRAM_ADDR_OUT(6) => 
                           DRAM_ADDR_OUT_6_port, DRAM_ADDR_OUT(5) => 
                           DRAM_ADDR_OUT_5_port, DRAM_ADDR_OUT(4) => 
                           DRAM_ADDR_OUT_4_port, DRAM_ADDR_OUT(3) => 
                           DRAM_ADDR_OUT_3_port, DRAM_ADDR_OUT(2) => 
                           DRAM_ADDR_OUT_2_port, DRAM_ADDR_OUT(1) => 
                           DRAM_ADDR_OUT_1_port, DRAM_ADDR_OUT(0) => 
                           DRAM_ADDR_OUT_0_port, DATA_OUT(31) => 
                           DATA_OUT_31_port, DATA_OUT(30) => DATA_OUT_30_port, 
                           DATA_OUT(29) => DATA_OUT_29_port, DATA_OUT(28) => 
                           DATA_OUT_28_port, DATA_OUT(27) => DATA_OUT_27_port, 
                           DATA_OUT(26) => DATA_OUT_26_port, DATA_OUT(25) => 
                           DATA_OUT_25_port, DATA_OUT(24) => DATA_OUT_24_port, 
                           DATA_OUT(23) => DATA_OUT_23_port, DATA_OUT(22) => 
                           DATA_OUT_22_port, DATA_OUT(21) => DATA_OUT_21_port, 
                           DATA_OUT(20) => DATA_OUT_20_port, DATA_OUT(19) => 
                           DATA_OUT_19_port, DATA_OUT(18) => DATA_OUT_18_port, 
                           DATA_OUT(17) => DATA_OUT_17_port, DATA_OUT(16) => 
                           DATA_OUT_16_port, DATA_OUT(15) => DATA_OUT_15_port, 
                           DATA_OUT(14) => DATA_OUT_14_port, DATA_OUT(13) => 
                           DATA_OUT_13_port, DATA_OUT(12) => DATA_OUT_12_port, 
                           DATA_OUT(11) => DATA_OUT_11_port, DATA_OUT(10) => 
                           DATA_OUT_10_port, DATA_OUT(9) => DATA_OUT_9_port, 
                           DATA_OUT(8) => DATA_OUT_8_port, DATA_OUT(7) => 
                           DATA_OUT_7_port, DATA_OUT(6) => DATA_OUT_6_port, 
                           DATA_OUT(5) => DATA_OUT_5_port, DATA_OUT(4) => 
                           DATA_OUT_4_port, DATA_OUT(3) => DATA_OUT_3_port, 
                           DATA_OUT(2) => DATA_OUT_2_port, DATA_OUT(1) => 
                           DATA_OUT_1_port, DATA_OUT(0) => DATA_OUT_0_port, 
                           DRAM_EN_OUT => DRAM_EN_OUT, DRAM_R_OUT => DRAM_R_OUT
                           , DRAM_W_OUT => DRAM_W_OUT, Bubble_out => Bubble);
   CU : hardwired_cu_NBIT32 port map( REG_LATCH_EN => n_1214, RD1 => n_1215, 
                           RD2 => n_1216, MUX_A_SEL => n_1217, MUX_B_SEL(1) => 
                           n_1218, MUX_B_SEL(0) => n_1219, ALU_OPC(0) => 
                           ALU_OPC_3_port, ALU_OPC(1) => ALU_OPC_2_port, 
                           ALU_OPC(2) => ALU_OPC_1_port, ALU_OPC(3) => 
                           ALU_OPC_0_port, ALU_OUTREG_EN => n_1220, DRAM_R_IN 
                           => n_1221, JUMP_TYPE(1) => n_1222, JUMP_TYPE(0) => 
                           n_1223, MEM_EN_IN => n_1224, DRAM_W_IN => n_1225, 
                           RF_WE => n_1226, DRAM_EN_IN => n_1227, WB_MUX_SEL =>
                           n_1228, INS_IN(31) => INS_IN_31_port, INS_IN(30) => 
                           INS_IN_30_port, INS_IN(29) => INS_IN_29_port, 
                           INS_IN(28) => INS_IN_28_port, INS_IN(27) => 
                           INS_IN_27_port, INS_IN(26) => INS_IN_26_port, 
                           INS_IN(25) => INS_IN_25_port, INS_IN(24) => 
                           INS_IN_24_port, INS_IN(23) => INS_IN_23_port, 
                           INS_IN(22) => INS_IN_22_port, INS_IN(21) => 
                           INS_IN_21_port, INS_IN(20) => INS_IN_20_port, 
                           INS_IN(19) => INS_IN_19_port, INS_IN(18) => 
                           INS_IN_18_port, INS_IN(17) => INS_IN_17_port, 
                           INS_IN(16) => INS_IN_16_port, INS_IN(15) => 
                           INS_IN_15_port, INS_IN(14) => INS_IN_14_port, 
                           INS_IN(13) => INS_IN_13_port, INS_IN(12) => 
                           INS_IN_12_port, INS_IN(11) => INS_IN_11_port, 
                           INS_IN(10) => INS_IN_10_port, INS_IN(9) => 
                           INS_IN_9_port, INS_IN(8) => INS_IN_8_port, INS_IN(7)
                           => INS_IN_7_port, INS_IN(6) => INS_IN_6_port, 
                           INS_IN(5) => INS_IN_5_port, INS_IN(4) => 
                           INS_IN_4_port, INS_IN(3) => INS_IN_3_port, INS_IN(2)
                           => INS_IN_2_port, INS_IN(1) => INS_IN_1_port, 
                           INS_IN(0) => INS_IN_0_port, Bubble => Bubble, Clk =>
                           Clk, Rst => Rst);
   IRAM_I : IRAM port map( Rst => Rst, Addr(31) => IRAM_ADDR_OUT_31_port, 
                           Addr(30) => IRAM_ADDR_OUT_30_port, Addr(29) => 
                           IRAM_ADDR_OUT_29_port, Addr(28) => 
                           IRAM_ADDR_OUT_28_port, Addr(27) => 
                           IRAM_ADDR_OUT_27_port, Addr(26) => 
                           IRAM_ADDR_OUT_26_port, Addr(25) => 
                           IRAM_ADDR_OUT_25_port, Addr(24) => 
                           IRAM_ADDR_OUT_24_port, Addr(23) => 
                           IRAM_ADDR_OUT_23_port, Addr(22) => 
                           IRAM_ADDR_OUT_22_port, Addr(21) => 
                           IRAM_ADDR_OUT_21_port, Addr(20) => 
                           IRAM_ADDR_OUT_20_port, Addr(19) => 
                           IRAM_ADDR_OUT_19_port, Addr(18) => 
                           IRAM_ADDR_OUT_18_port, Addr(17) => 
                           IRAM_ADDR_OUT_17_port, Addr(16) => 
                           IRAM_ADDR_OUT_16_port, Addr(15) => 
                           IRAM_ADDR_OUT_15_port, Addr(14) => 
                           IRAM_ADDR_OUT_14_port, Addr(13) => 
                           IRAM_ADDR_OUT_13_port, Addr(12) => 
                           IRAM_ADDR_OUT_12_port, Addr(11) => 
                           IRAM_ADDR_OUT_11_port, Addr(10) => 
                           IRAM_ADDR_OUT_10_port, Addr(9) => 
                           IRAM_ADDR_OUT_9_port, Addr(8) => 
                           IRAM_ADDR_OUT_8_port, Addr(7) => 
                           IRAM_ADDR_OUT_7_port, Addr(6) => 
                           IRAM_ADDR_OUT_6_port, Addr(5) => 
                           IRAM_ADDR_OUT_5_port, Addr(4) => 
                           IRAM_ADDR_OUT_4_port, Addr(3) => 
                           IRAM_ADDR_OUT_3_port, Addr(2) => 
                           IRAM_ADDR_OUT_2_port, Addr(1) => 
                           IRAM_ADDR_OUT_1_port, Addr(0) => 
                           IRAM_ADDR_OUT_0_port, Iout(31) => INS_IN_31_port, 
                           Iout(30) => INS_IN_30_port, Iout(29) => 
                           INS_IN_29_port, Iout(28) => INS_IN_28_port, Iout(27)
                           => INS_IN_27_port, Iout(26) => INS_IN_26_port, 
                           Iout(25) => INS_IN_25_port, Iout(24) => 
                           INS_IN_24_port, Iout(23) => INS_IN_23_port, Iout(22)
                           => INS_IN_22_port, Iout(21) => INS_IN_21_port, 
                           Iout(20) => INS_IN_20_port, Iout(19) => 
                           INS_IN_19_port, Iout(18) => INS_IN_18_port, Iout(17)
                           => INS_IN_17_port, Iout(16) => INS_IN_16_port, 
                           Iout(15) => INS_IN_15_port, Iout(14) => 
                           INS_IN_14_port, Iout(13) => INS_IN_13_port, Iout(12)
                           => INS_IN_12_port, Iout(11) => INS_IN_11_port, 
                           Iout(10) => INS_IN_10_port, Iout(9) => INS_IN_9_port
                           , Iout(8) => INS_IN_8_port, Iout(7) => INS_IN_7_port
                           , Iout(6) => INS_IN_6_port, Iout(5) => INS_IN_5_port
                           , Iout(4) => INS_IN_4_port, Iout(3) => INS_IN_3_port
                           , Iout(2) => INS_IN_2_port, Iout(1) => INS_IN_1_port
                           , Iout(0) => INS_IN_0_port);
   DRAM_I : DRAM port map( En => DRAM_EN_OUT, Rst => Rst, ADDR_IN(31) => 
                           DRAM_ADDR_OUT_31_port, ADDR_IN(30) => 
                           DRAM_ADDR_OUT_30_port, ADDR_IN(29) => 
                           DRAM_ADDR_OUT_29_port, ADDR_IN(28) => 
                           DRAM_ADDR_OUT_28_port, ADDR_IN(27) => 
                           DRAM_ADDR_OUT_27_port, ADDR_IN(26) => 
                           DRAM_ADDR_OUT_26_port, ADDR_IN(25) => 
                           DRAM_ADDR_OUT_25_port, ADDR_IN(24) => 
                           DRAM_ADDR_OUT_24_port, ADDR_IN(23) => 
                           DRAM_ADDR_OUT_23_port, ADDR_IN(22) => 
                           DRAM_ADDR_OUT_22_port, ADDR_IN(21) => 
                           DRAM_ADDR_OUT_21_port, ADDR_IN(20) => 
                           DRAM_ADDR_OUT_20_port, ADDR_IN(19) => 
                           DRAM_ADDR_OUT_19_port, ADDR_IN(18) => 
                           DRAM_ADDR_OUT_18_port, ADDR_IN(17) => 
                           DRAM_ADDR_OUT_17_port, ADDR_IN(16) => 
                           DRAM_ADDR_OUT_16_port, ADDR_IN(15) => 
                           DRAM_ADDR_OUT_15_port, ADDR_IN(14) => 
                           DRAM_ADDR_OUT_14_port, ADDR_IN(13) => 
                           DRAM_ADDR_OUT_13_port, ADDR_IN(12) => 
                           DRAM_ADDR_OUT_12_port, ADDR_IN(11) => 
                           DRAM_ADDR_OUT_11_port, ADDR_IN(10) => 
                           DRAM_ADDR_OUT_10_port, ADDR_IN(9) => 
                           DRAM_ADDR_OUT_9_port, ADDR_IN(8) => 
                           DRAM_ADDR_OUT_8_port, ADDR_IN(7) => 
                           DRAM_ADDR_OUT_7_port, ADDR_IN(6) => 
                           DRAM_ADDR_OUT_6_port, ADDR_IN(5) => 
                           DRAM_ADDR_OUT_5_port, ADDR_IN(4) => 
                           DRAM_ADDR_OUT_4_port, ADDR_IN(3) => 
                           DRAM_ADDR_OUT_3_port, ADDR_IN(2) => 
                           DRAM_ADDR_OUT_2_port, ADDR_IN(1) => 
                           DRAM_ADDR_OUT_1_port, ADDR_IN(0) => 
                           DRAM_ADDR_OUT_0_port, DATA_IN(31) => 
                           DATA_OUT_31_port, DATA_IN(30) => DATA_OUT_30_port, 
                           DATA_IN(29) => DATA_OUT_29_port, DATA_IN(28) => 
                           DATA_OUT_28_port, DATA_IN(27) => DATA_OUT_27_port, 
                           DATA_IN(26) => DATA_OUT_26_port, DATA_IN(25) => 
                           DATA_OUT_25_port, DATA_IN(24) => DATA_OUT_24_port, 
                           DATA_IN(23) => DATA_OUT_23_port, DATA_IN(22) => 
                           DATA_OUT_22_port, DATA_IN(21) => DATA_OUT_21_port, 
                           DATA_IN(20) => DATA_OUT_20_port, DATA_IN(19) => 
                           DATA_OUT_19_port, DATA_IN(18) => DATA_OUT_18_port, 
                           DATA_IN(17) => DATA_OUT_17_port, DATA_IN(16) => 
                           DATA_OUT_16_port, DATA_IN(15) => DATA_OUT_15_port, 
                           DATA_IN(14) => DATA_OUT_14_port, DATA_IN(13) => 
                           DATA_OUT_13_port, DATA_IN(12) => DATA_OUT_12_port, 
                           DATA_IN(11) => DATA_OUT_11_port, DATA_IN(10) => 
                           DATA_OUT_10_port, DATA_IN(9) => DATA_OUT_9_port, 
                           DATA_IN(8) => DATA_OUT_8_port, DATA_IN(7) => 
                           DATA_OUT_7_port, DATA_IN(6) => DATA_OUT_6_port, 
                           DATA_IN(5) => DATA_OUT_5_port, DATA_IN(4) => 
                           DATA_OUT_4_port, DATA_IN(3) => DATA_OUT_3_port, 
                           DATA_IN(2) => DATA_OUT_2_port, DATA_IN(1) => 
                           DATA_OUT_1_port, DATA_IN(0) => DATA_OUT_0_port, 
                           DRAM_W => DRAM_W_OUT, DRAM_R => DRAM_R_OUT, 
                           DATA_OUT(31) => DATA_IN_31_port, DATA_OUT(30) => 
                           DATA_IN_30_port, DATA_OUT(29) => DATA_IN_29_port, 
                           DATA_OUT(28) => DATA_IN_28_port, DATA_OUT(27) => 
                           DATA_IN_27_port, DATA_OUT(26) => DATA_IN_26_port, 
                           DATA_OUT(25) => DATA_IN_25_port, DATA_OUT(24) => 
                           DATA_IN_24_port, DATA_OUT(23) => DATA_IN_23_port, 
                           DATA_OUT(22) => DATA_IN_22_port, DATA_OUT(21) => 
                           DATA_IN_21_port, DATA_OUT(20) => DATA_IN_20_port, 
                           DATA_OUT(19) => DATA_IN_19_port, DATA_OUT(18) => 
                           DATA_IN_18_port, DATA_OUT(17) => DATA_IN_17_port, 
                           DATA_OUT(16) => DATA_IN_16_port, DATA_OUT(15) => 
                           DATA_IN_15_port, DATA_OUT(14) => DATA_IN_14_port, 
                           DATA_OUT(13) => DATA_IN_13_port, DATA_OUT(12) => 
                           DATA_IN_12_port, DATA_OUT(11) => DATA_IN_11_port, 
                           DATA_OUT(10) => DATA_IN_10_port, DATA_OUT(9) => 
                           DATA_IN_9_port, DATA_OUT(8) => DATA_IN_8_port, 
                           DATA_OUT(7) => DATA_IN_7_port, DATA_OUT(6) => 
                           DATA_IN_6_port, DATA_OUT(5) => DATA_IN_5_port, 
                           DATA_OUT(4) => DATA_IN_4_port, DATA_OUT(3) => 
                           DATA_IN_3_port, DATA_OUT(2) => DATA_IN_2_port, 
                           DATA_OUT(1) => DATA_IN_1_port, DATA_OUT(0) => 
                           DATA_IN_0_port);
   WB_MUX_SEL <= '0';
   DRAM_EN_IN <= '0';
   RF_WE <= '0';
   DRAM_W_IN <= '0';
   MEM_EN_IN <= '0';
   JUMP_TYPE_0_port <= '0';
   JUMP_TYPE_1_port <= '0';
   DRAM_R_IN <= '0';
   ALU_OUTREG_EN <= '0';
   MUX_B_SEL_0_port <= '0';
   MUX_B_SEL_1_port <= '0';
   MUX_A_SEL <= '0';
   RD2 <= '0';
   RD1 <= '0';
   REG_LATCH_EN <= '0';

end SYN_dlx_rtl;
