
module mux21_NBIT32_0 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n36, n37, n38, n39, n40, n43, n54, n65, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19;

  NAND2_X1 U1 ( .A1(B[19]), .A2(n16), .ZN(n5) );
  NAND2_X1 U2 ( .A1(B[15]), .A2(n16), .ZN(n8) );
  INV_X1 U3 ( .A(n17), .ZN(n16) );
  INV_X1 U4 ( .A(n19), .ZN(n15) );
  NAND2_X1 U5 ( .A1(A[23]), .A2(n19), .ZN(n9) );
  NAND2_X1 U6 ( .A1(A[31]), .A2(n18), .ZN(n1) );
  NAND2_X1 U7 ( .A1(B[31]), .A2(n15), .ZN(n2) );
  NAND2_X1 U8 ( .A1(n1), .A2(n2), .ZN(Z[31]) );
  NAND2_X1 U9 ( .A1(B[23]), .A2(n16), .ZN(n10) );
  NAND2_X1 U10 ( .A1(A[19]), .A2(n3), .ZN(n4) );
  NAND2_X1 U11 ( .A1(n4), .A2(n5), .ZN(Z[19]) );
  INV_X1 U12 ( .A(n16), .ZN(n3) );
  NAND2_X1 U13 ( .A1(A[15]), .A2(n6), .ZN(n7) );
  NAND2_X1 U14 ( .A1(n7), .A2(n8), .ZN(Z[15]) );
  INV_X1 U15 ( .A(n16), .ZN(n6) );
  NAND2_X1 U16 ( .A1(n10), .A2(n9), .ZN(Z[23]) );
  AOI22_X1 U17 ( .A1(A[7]), .A2(n19), .B1(B[7]), .B2(n15), .ZN(n36) );
  INV_X1 U18 ( .A(n37), .ZN(Z[6]) );
  AOI22_X1 U19 ( .A1(A[6]), .A2(n19), .B1(B[6]), .B2(n15), .ZN(n37) );
  INV_X1 U20 ( .A(n38), .ZN(Z[5]) );
  AOI22_X1 U21 ( .A1(A[5]), .A2(n18), .B1(B[5]), .B2(n15), .ZN(n38) );
  INV_X1 U22 ( .A(n43), .ZN(Z[2]) );
  AOI22_X1 U23 ( .A1(A[2]), .A2(n17), .B1(B[2]), .B2(n15), .ZN(n43) );
  INV_X1 U24 ( .A(n54), .ZN(Z[1]) );
  AOI22_X1 U25 ( .A1(A[1]), .A2(n18), .B1(B[1]), .B2(n15), .ZN(n54) );
  INV_X1 U26 ( .A(n65), .ZN(Z[0]) );
  AOI22_X1 U27 ( .A1(A[0]), .A2(n19), .B1(B[0]), .B2(n15), .ZN(n65) );
  INV_X1 U28 ( .A(n40), .ZN(Z[3]) );
  AOI22_X1 U29 ( .A1(A[3]), .A2(n17), .B1(B[3]), .B2(n15), .ZN(n40) );
  INV_X1 U30 ( .A(n39), .ZN(Z[4]) );
  AOI22_X1 U31 ( .A1(A[4]), .A2(n18), .B1(B[4]), .B2(n15), .ZN(n39) );
  NAND2_X1 U32 ( .A1(A[27]), .A2(n18), .ZN(n11) );
  NAND2_X1 U33 ( .A1(B[27]), .A2(n15), .ZN(n12) );
  NAND2_X1 U34 ( .A1(n11), .A2(n12), .ZN(Z[27]) );
  NAND2_X1 U35 ( .A1(A[25]), .A2(n17), .ZN(n13) );
  NAND2_X1 U36 ( .A1(B[25]), .A2(n16), .ZN(n14) );
  NAND2_X1 U37 ( .A1(n13), .A2(n14), .ZN(Z[25]) );
  INV_X1 U38 ( .A(n36), .ZN(Z[7]) );
  INV_X1 U39 ( .A(S), .ZN(n17) );
  INV_X1 U40 ( .A(S), .ZN(n18) );
  INV_X1 U41 ( .A(S), .ZN(n19) );
  MUX2_X1 U42 ( .A(A[8]), .B(B[8]), .S(n16), .Z(Z[8]) );
  MUX2_X1 U43 ( .A(A[9]), .B(B[9]), .S(n16), .Z(Z[9]) );
  MUX2_X1 U44 ( .A(A[10]), .B(B[10]), .S(n16), .Z(Z[10]) );
  MUX2_X1 U45 ( .A(A[11]), .B(B[11]), .S(n16), .Z(Z[11]) );
  MUX2_X1 U46 ( .A(A[12]), .B(B[12]), .S(n16), .Z(Z[12]) );
  MUX2_X1 U47 ( .A(A[13]), .B(B[13]), .S(n16), .Z(Z[13]) );
  MUX2_X1 U48 ( .A(A[14]), .B(B[14]), .S(n16), .Z(Z[14]) );
  MUX2_X1 U49 ( .A(A[16]), .B(B[16]), .S(n16), .Z(Z[16]) );
  MUX2_X1 U50 ( .A(A[17]), .B(B[17]), .S(n16), .Z(Z[17]) );
  MUX2_X1 U51 ( .A(A[18]), .B(B[18]), .S(n16), .Z(Z[18]) );
  MUX2_X1 U52 ( .A(A[20]), .B(B[20]), .S(n16), .Z(Z[20]) );
  MUX2_X1 U53 ( .A(A[21]), .B(B[21]), .S(n16), .Z(Z[21]) );
  MUX2_X1 U54 ( .A(A[22]), .B(B[22]), .S(n16), .Z(Z[22]) );
  MUX2_X1 U55 ( .A(A[24]), .B(B[24]), .S(n16), .Z(Z[24]) );
  MUX2_X1 U56 ( .A(A[26]), .B(B[26]), .S(n15), .Z(Z[26]) );
  MUX2_X1 U57 ( .A(A[28]), .B(B[28]), .S(n15), .Z(Z[28]) );
  MUX2_X1 U58 ( .A(A[29]), .B(B[29]), .S(n15), .Z(Z[29]) );
  MUX2_X1 U59 ( .A(A[30]), .B(B[30]), .S(n15), .Z(Z[30]) );
endmodule


module mux21_NBIT32_5 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111;

  INV_X1 U1 ( .A(n15), .ZN(n5) );
  INV_X1 U2 ( .A(n15), .ZN(n4) );
  BUF_X1 U3 ( .A(n3), .Z(n15) );
  BUF_X1 U4 ( .A(n2), .Z(n11) );
  BUF_X1 U5 ( .A(n1), .Z(n8) );
  BUF_X1 U6 ( .A(n2), .Z(n10) );
  BUF_X1 U7 ( .A(n1), .Z(n9) );
  BUF_X1 U8 ( .A(n3), .Z(n14) );
  BUF_X1 U9 ( .A(n1), .Z(n7) );
  BUF_X1 U10 ( .A(n3), .Z(n13) );
  BUF_X1 U11 ( .A(n2), .Z(n12) );
  BUF_X1 U12 ( .A(S), .Z(n3) );
  BUF_X1 U13 ( .A(S), .Z(n2) );
  BUF_X1 U14 ( .A(S), .Z(n1) );
  INV_X1 U15 ( .A(n107), .ZN(Z[5]) );
  INV_X1 U16 ( .A(n99), .ZN(Z[27]) );
  INV_X1 U17 ( .A(n82), .ZN(Z[11]) );
  INV_X1 U18 ( .A(n83), .ZN(Z[12]) );
  INV_X1 U19 ( .A(n84), .ZN(Z[13]) );
  INV_X1 U20 ( .A(n87), .ZN(Z[16]) );
  INV_X1 U21 ( .A(n88), .ZN(Z[17]) );
  INV_X1 U22 ( .A(n89), .ZN(Z[18]) );
  INV_X1 U23 ( .A(n92), .ZN(Z[20]) );
  INV_X1 U24 ( .A(n96), .ZN(Z[24]) );
  INV_X1 U25 ( .A(n98), .ZN(Z[26]) );
  INV_X1 U26 ( .A(n108), .ZN(Z[6]) );
  INV_X1 U27 ( .A(n81), .ZN(Z[10]) );
  INV_X1 U28 ( .A(n102), .ZN(Z[2]) );
  AOI22_X1 U29 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n8), .ZN(n102) );
  INV_X1 U30 ( .A(n110), .ZN(Z[8]) );
  INV_X1 U31 ( .A(n91), .ZN(Z[1]) );
  AOI22_X1 U32 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(n11), .ZN(n91) );
  INV_X1 U33 ( .A(n80), .ZN(Z[0]) );
  AOI22_X1 U34 ( .A1(A[0]), .A2(n4), .B1(B[0]), .B2(n14), .ZN(n80) );
  INV_X1 U35 ( .A(n85), .ZN(Z[14]) );
  INV_X1 U36 ( .A(n90), .ZN(Z[19]) );
  INV_X1 U37 ( .A(n105), .ZN(Z[3]) );
  INV_X1 U38 ( .A(n109), .ZN(Z[7]) );
  INV_X1 U39 ( .A(n111), .ZN(Z[9]) );
  INV_X1 U40 ( .A(n86), .ZN(Z[15]) );
  INV_X1 U41 ( .A(n97), .ZN(Z[25]) );
  INV_X1 U42 ( .A(n106), .ZN(Z[4]) );
  AOI22_X1 U43 ( .A1(A[4]), .A2(n6), .B1(B[4]), .B2(n8), .ZN(n106) );
  INV_X1 U44 ( .A(n93), .ZN(Z[21]) );
  AOI22_X1 U45 ( .A1(A[21]), .A2(n5), .B1(B[21]), .B2(n11), .ZN(n93) );
  INV_X1 U46 ( .A(n94), .ZN(Z[22]) );
  AOI22_X1 U47 ( .A1(A[22]), .A2(n5), .B1(B[22]), .B2(n10), .ZN(n94) );
  INV_X1 U48 ( .A(n95), .ZN(Z[23]) );
  AOI22_X1 U49 ( .A1(A[23]), .A2(n5), .B1(B[23]), .B2(n10), .ZN(n95) );
  INV_X1 U50 ( .A(n100), .ZN(Z[28]) );
  AOI22_X1 U51 ( .A1(A[28]), .A2(n5), .B1(B[28]), .B2(n9), .ZN(n100) );
  INV_X1 U52 ( .A(n101), .ZN(Z[29]) );
  AOI22_X1 U53 ( .A1(A[29]), .A2(n5), .B1(B[29]), .B2(n9), .ZN(n101) );
  INV_X1 U54 ( .A(n103), .ZN(Z[30]) );
  AOI22_X1 U55 ( .A1(A[30]), .A2(n5), .B1(B[30]), .B2(n11), .ZN(n103) );
  INV_X1 U56 ( .A(n104), .ZN(Z[31]) );
  AOI22_X1 U57 ( .A1(A[31]), .A2(n6), .B1(B[31]), .B2(n8), .ZN(n104) );
  AOI22_X1 U58 ( .A1(A[20]), .A2(n5), .B1(B[20]), .B2(n11), .ZN(n92) );
  AOI22_X1 U59 ( .A1(A[27]), .A2(n5), .B1(B[27]), .B2(n9), .ZN(n99) );
  AOI22_X1 U60 ( .A1(A[24]), .A2(n5), .B1(B[24]), .B2(n10), .ZN(n96) );
  AOI22_X1 U61 ( .A1(A[25]), .A2(n5), .B1(B[25]), .B2(n10), .ZN(n97) );
  AOI22_X1 U62 ( .A1(A[26]), .A2(n5), .B1(B[26]), .B2(n9), .ZN(n98) );
  AOI22_X1 U63 ( .A1(A[15]), .A2(n4), .B1(B[15]), .B2(n13), .ZN(n86) );
  AOI22_X1 U64 ( .A1(A[11]), .A2(n4), .B1(B[11]), .B2(n14), .ZN(n82) );
  AOI22_X1 U65 ( .A1(A[13]), .A2(n4), .B1(B[13]), .B2(n13), .ZN(n84) );
  AOI22_X1 U66 ( .A1(A[12]), .A2(n4), .B1(B[12]), .B2(n13), .ZN(n83) );
  AOI22_X1 U67 ( .A1(A[19]), .A2(n4), .B1(B[19]), .B2(n12), .ZN(n90) );
  AOI22_X1 U68 ( .A1(A[17]), .A2(n4), .B1(B[17]), .B2(n12), .ZN(n88) );
  AOI22_X1 U69 ( .A1(A[18]), .A2(n4), .B1(B[18]), .B2(n12), .ZN(n89) );
  AOI22_X1 U70 ( .A1(A[16]), .A2(n4), .B1(B[16]), .B2(n12), .ZN(n87) );
  AOI22_X1 U71 ( .A1(A[14]), .A2(n4), .B1(B[14]), .B2(n13), .ZN(n85) );
  AOI22_X1 U72 ( .A1(A[5]), .A2(n6), .B1(B[5]), .B2(n7), .ZN(n107) );
  AOI22_X1 U73 ( .A1(A[7]), .A2(n6), .B1(B[7]), .B2(n7), .ZN(n109) );
  AOI22_X1 U74 ( .A1(A[10]), .A2(n4), .B1(B[10]), .B2(n14), .ZN(n81) );
  AOI22_X1 U75 ( .A1(A[3]), .A2(n6), .B1(B[3]), .B2(n8), .ZN(n105) );
  AOI22_X1 U76 ( .A1(A[6]), .A2(n6), .B1(B[6]), .B2(n7), .ZN(n108) );
  AOI22_X1 U77 ( .A1(A[8]), .A2(n6), .B1(B[8]), .B2(n7), .ZN(n110) );
  AOI22_X1 U78 ( .A1(A[9]), .A2(n6), .B1(n14), .B2(B[9]), .ZN(n111) );
  INV_X1 U79 ( .A(n15), .ZN(n6) );
endmodule


module mux21_NBIT32_4 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n11) );
  BUF_X1 U6 ( .A(n2), .Z(n9) );
  BUF_X1 U7 ( .A(n1), .Z(n8) );
  BUF_X1 U8 ( .A(n2), .Z(n10) );
  BUF_X1 U9 ( .A(n1), .Z(n7) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(S), .Z(n3) );
  BUF_X1 U13 ( .A(S), .Z(n2) );
  BUF_X1 U14 ( .A(S), .Z(n1) );
  INV_X1 U15 ( .A(n90), .ZN(Z[1]) );
  AOI22_X1 U16 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(n10), .ZN(n90) );
  INV_X1 U17 ( .A(n101), .ZN(Z[2]) );
  AOI22_X1 U18 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n7), .ZN(n101) );
  INV_X1 U19 ( .A(n104), .ZN(Z[3]) );
  AOI22_X1 U20 ( .A1(A[3]), .A2(n4), .B1(B[3]), .B2(n7), .ZN(n104) );
  INV_X1 U21 ( .A(n105), .ZN(Z[4]) );
  AOI22_X1 U22 ( .A1(A[4]), .A2(n5), .B1(B[4]), .B2(n7), .ZN(n105) );
  INV_X1 U23 ( .A(n106), .ZN(Z[5]) );
  AOI22_X1 U24 ( .A1(A[5]), .A2(n4), .B1(B[5]), .B2(n6), .ZN(n106) );
  INV_X1 U25 ( .A(n107), .ZN(Z[6]) );
  AOI22_X1 U26 ( .A1(A[6]), .A2(n5), .B1(B[6]), .B2(n6), .ZN(n107) );
  INV_X1 U27 ( .A(n108), .ZN(Z[7]) );
  AOI22_X1 U28 ( .A1(A[7]), .A2(n4), .B1(B[7]), .B2(n6), .ZN(n108) );
  INV_X1 U29 ( .A(n109), .ZN(Z[8]) );
  AOI22_X1 U30 ( .A1(A[8]), .A2(n5), .B1(B[8]), .B2(n6), .ZN(n109) );
  INV_X1 U31 ( .A(n80), .ZN(Z[10]) );
  AOI22_X1 U32 ( .A1(A[10]), .A2(n4), .B1(B[10]), .B2(n13), .ZN(n80) );
  INV_X1 U33 ( .A(n81), .ZN(Z[11]) );
  AOI22_X1 U34 ( .A1(A[11]), .A2(n4), .B1(B[11]), .B2(n13), .ZN(n81) );
  INV_X1 U35 ( .A(n82), .ZN(Z[12]) );
  AOI22_X1 U36 ( .A1(A[12]), .A2(n4), .B1(B[12]), .B2(n12), .ZN(n82) );
  INV_X1 U37 ( .A(n83), .ZN(Z[13]) );
  AOI22_X1 U38 ( .A1(A[13]), .A2(n4), .B1(B[13]), .B2(n12), .ZN(n83) );
  INV_X1 U39 ( .A(n84), .ZN(Z[14]) );
  AOI22_X1 U40 ( .A1(A[14]), .A2(n4), .B1(B[14]), .B2(n12), .ZN(n84) );
  INV_X1 U41 ( .A(n85), .ZN(Z[15]) );
  AOI22_X1 U42 ( .A1(A[15]), .A2(n4), .B1(B[15]), .B2(n12), .ZN(n85) );
  INV_X1 U43 ( .A(n86), .ZN(Z[16]) );
  AOI22_X1 U44 ( .A1(A[16]), .A2(n4), .B1(B[16]), .B2(n11), .ZN(n86) );
  INV_X1 U45 ( .A(n87), .ZN(Z[17]) );
  AOI22_X1 U46 ( .A1(A[17]), .A2(n4), .B1(B[17]), .B2(n11), .ZN(n87) );
  INV_X1 U47 ( .A(n88), .ZN(Z[18]) );
  AOI22_X1 U48 ( .A1(A[18]), .A2(n4), .B1(B[18]), .B2(n11), .ZN(n88) );
  INV_X1 U49 ( .A(n89), .ZN(Z[19]) );
  AOI22_X1 U50 ( .A1(A[19]), .A2(n4), .B1(B[19]), .B2(n11), .ZN(n89) );
  INV_X1 U51 ( .A(n91), .ZN(Z[20]) );
  AOI22_X1 U52 ( .A1(A[20]), .A2(n5), .B1(B[20]), .B2(n10), .ZN(n91) );
  INV_X1 U53 ( .A(n92), .ZN(Z[21]) );
  AOI22_X1 U54 ( .A1(A[21]), .A2(n5), .B1(B[21]), .B2(n10), .ZN(n92) );
  INV_X1 U55 ( .A(n93), .ZN(Z[22]) );
  AOI22_X1 U56 ( .A1(A[22]), .A2(n5), .B1(B[22]), .B2(n9), .ZN(n93) );
  INV_X1 U57 ( .A(n94), .ZN(Z[23]) );
  AOI22_X1 U58 ( .A1(A[23]), .A2(n5), .B1(B[23]), .B2(n9), .ZN(n94) );
  INV_X1 U59 ( .A(n95), .ZN(Z[24]) );
  AOI22_X1 U60 ( .A1(A[24]), .A2(n5), .B1(B[24]), .B2(n9), .ZN(n95) );
  INV_X1 U61 ( .A(n96), .ZN(Z[25]) );
  AOI22_X1 U62 ( .A1(A[25]), .A2(n5), .B1(B[25]), .B2(n9), .ZN(n96) );
  INV_X1 U63 ( .A(n97), .ZN(Z[26]) );
  AOI22_X1 U64 ( .A1(A[26]), .A2(n5), .B1(B[26]), .B2(n8), .ZN(n97) );
  INV_X1 U65 ( .A(n98), .ZN(Z[27]) );
  AOI22_X1 U66 ( .A1(A[27]), .A2(n5), .B1(B[27]), .B2(n8), .ZN(n98) );
  INV_X1 U67 ( .A(n99), .ZN(Z[28]) );
  AOI22_X1 U68 ( .A1(A[28]), .A2(n5), .B1(B[28]), .B2(n8), .ZN(n99) );
  INV_X1 U69 ( .A(n100), .ZN(Z[29]) );
  AOI22_X1 U70 ( .A1(A[29]), .A2(n5), .B1(B[29]), .B2(n8), .ZN(n100) );
  INV_X1 U71 ( .A(n102), .ZN(Z[30]) );
  AOI22_X1 U72 ( .A1(A[30]), .A2(n5), .B1(B[30]), .B2(n10), .ZN(n102) );
  INV_X1 U73 ( .A(n103), .ZN(Z[31]) );
  AOI22_X1 U74 ( .A1(A[31]), .A2(n4), .B1(B[31]), .B2(n7), .ZN(n103) );
  INV_X1 U75 ( .A(n110), .ZN(Z[9]) );
  AOI22_X1 U76 ( .A1(A[9]), .A2(n5), .B1(n13), .B2(B[9]), .ZN(n110) );
  INV_X1 U77 ( .A(n79), .ZN(Z[0]) );
  AOI22_X1 U78 ( .A1(A[0]), .A2(n4), .B1(B[0]), .B2(n13), .ZN(n79) );
endmodule


module regn_N32_0 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n51, n52, n1, n2, n3, n4, n5, n6, n7, n8, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n53, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n9, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n49;

  DFFR_X1 \DOUT_reg[31]  ( .D(n96), .CK(CLK), .RN(n32), .Q(DOUT[31]) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n95), .CK(CLK), .RN(n32), .Q(DOUT[30]) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n94), .CK(CLK), .RN(n32), .Q(DOUT[29]) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n93), .CK(CLK), .RN(n32), .Q(DOUT[28]) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n92), .CK(CLK), .RN(n32), .Q(DOUT[27]) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n91), .CK(CLK), .RN(n32), .Q(DOUT[26]) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n90), .CK(CLK), .RN(n32), .Q(DOUT[25]) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n89), .CK(CLK), .RN(n32), .Q(DOUT[24]) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n88), .CK(CLK), .RN(n31), .Q(DOUT[23]) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n87), .CK(CLK), .RN(n31), .Q(DOUT[22]) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n86), .CK(CLK), .RN(n31), .Q(DOUT[21]) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n85), .CK(CLK), .RN(n31), .Q(DOUT[20]), .QN(n53)
         );
  DFFR_X1 \DOUT_reg[18]  ( .D(n83), .CK(CLK), .RN(n31), .Q(DOUT[18]) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n82), .CK(CLK), .RN(n31), .Q(DOUT[17]) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n81), .CK(CLK), .RN(n31), .Q(DOUT[16]) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n80), .CK(CLK), .RN(n31), .Q(DOUT[15]) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n79), .CK(CLK), .RN(n31), .Q(DOUT[14]) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n78), .CK(CLK), .RN(n31), .Q(DOUT[13]) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n77), .CK(CLK), .RN(n31), .Q(DOUT[12]) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n76), .CK(CLK), .RN(n30), .Q(DOUT[11]) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n75), .CK(CLK), .RN(n30), .Q(n9), .QN(n43) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n74), .CK(CLK), .RN(n30), .Q(n51), .QN(n42) );
  DFFR_X1 \DOUT_reg[8]  ( .D(n73), .CK(CLK), .RN(n30), .Q(n52), .QN(n41) );
  DFFR_X1 \DOUT_reg[7]  ( .D(n72), .CK(CLK), .RN(n30), .Q(DOUT[7]), .QN(n40)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n71), .CK(CLK), .RN(n30), .Q(DOUT[6]), .QN(n39)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n70), .CK(CLK), .RN(n30), .Q(DOUT[5]), .QN(n38)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n69), .CK(CLK), .RN(n30), .Q(DOUT[4]), .QN(n37)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n68), .CK(CLK), .RN(n30), .Q(DOUT[3]), .QN(n36)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n67), .CK(CLK), .RN(n30), .Q(DOUT[2]), .QN(n35)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n66), .CK(CLK), .RN(n30), .Q(DOUT[1]), .QN(n34)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n65), .CK(CLK), .RN(n30), .Q(DOUT[0]), .QN(n33)
         );
  DFFR_X1 \DOUT_reg[19]  ( .D(n84), .CK(CLK), .RN(n31), .Q(DOUT[19]) );
  INV_X1 U2 ( .A(EN), .ZN(n11) );
  INV_X1 U3 ( .A(n43), .ZN(DOUT[10]) );
  MUX2_X1 U4 ( .A(DIN[28]), .B(DOUT[28]), .S(n11), .Z(n93) );
  MUX2_X1 U5 ( .A(DIN[25]), .B(DOUT[25]), .S(n11), .Z(n90) );
  NAND2_X1 U6 ( .A1(DOUT[15]), .A2(n12), .ZN(n13) );
  NAND2_X1 U7 ( .A1(DIN[15]), .A2(EN), .ZN(n14) );
  NAND2_X1 U8 ( .A1(n13), .A2(n14), .ZN(n80) );
  INV_X1 U9 ( .A(EN), .ZN(n12) );
  BUF_X1 U10 ( .A(RST), .Z(n30) );
  BUF_X1 U11 ( .A(RST), .Z(n31) );
  BUF_X1 U12 ( .A(RST), .Z(n32) );
  NAND2_X1 U13 ( .A1(DIN[7]), .A2(EN), .ZN(n8) );
  NAND2_X1 U14 ( .A1(DIN[6]), .A2(EN), .ZN(n7) );
  NAND2_X1 U15 ( .A1(DIN[5]), .A2(EN), .ZN(n6) );
  OAI21_X1 U16 ( .B1(n35), .B2(EN), .A(n3), .ZN(n67) );
  NAND2_X1 U17 ( .A1(DIN[2]), .A2(EN), .ZN(n3) );
  OAI21_X1 U18 ( .B1(n34), .B2(EN), .A(n2), .ZN(n66) );
  NAND2_X1 U19 ( .A1(DIN[1]), .A2(EN), .ZN(n2) );
  OAI21_X1 U20 ( .B1(n33), .B2(EN), .A(n1), .ZN(n65) );
  NAND2_X1 U21 ( .A1(EN), .A2(DIN[0]), .ZN(n1) );
  NAND2_X1 U22 ( .A1(DIN[3]), .A2(EN), .ZN(n4) );
  NAND2_X1 U23 ( .A1(DIN[4]), .A2(EN), .ZN(n5) );
  INV_X1 U24 ( .A(EN), .ZN(n27) );
  INV_X1 U25 ( .A(EN), .ZN(n18) );
  INV_X1 U26 ( .A(EN), .ZN(n21) );
  OAI21_X1 U27 ( .B1(n37), .B2(EN), .A(n5), .ZN(n69) );
  OAI21_X1 U28 ( .B1(n38), .B2(EN), .A(n6), .ZN(n70) );
  OAI21_X1 U29 ( .B1(n40), .B2(EN), .A(n8), .ZN(n72) );
  NAND2_X1 U30 ( .A1(DIN[29]), .A2(n15), .ZN(n16) );
  NAND2_X1 U31 ( .A1(DOUT[29]), .A2(n18), .ZN(n17) );
  NAND2_X1 U32 ( .A1(n16), .A2(n17), .ZN(n94) );
  INV_X1 U33 ( .A(n18), .ZN(n15) );
  OAI21_X1 U34 ( .B1(n39), .B2(EN), .A(n7), .ZN(n71) );
  NAND2_X1 U35 ( .A1(DIN[31]), .A2(n24), .ZN(n19) );
  NAND2_X1 U36 ( .A1(DOUT[31]), .A2(n21), .ZN(n20) );
  NAND2_X1 U37 ( .A1(n19), .A2(n20), .ZN(n96) );
  OAI21_X1 U38 ( .B1(n36), .B2(EN), .A(n4), .ZN(n68) );
  NAND2_X1 U39 ( .A1(DIN[27]), .A2(n15), .ZN(n22) );
  NAND2_X1 U40 ( .A1(DOUT[27]), .A2(n12), .ZN(n23) );
  NAND2_X1 U41 ( .A1(n22), .A2(n23), .ZN(n92) );
  NAND2_X1 U42 ( .A1(DIN[23]), .A2(n24), .ZN(n25) );
  NAND2_X1 U43 ( .A1(DOUT[23]), .A2(n27), .ZN(n26) );
  NAND2_X1 U44 ( .A1(n25), .A2(n26), .ZN(n88) );
  INV_X1 U45 ( .A(n27), .ZN(n24) );
  NAND2_X1 U46 ( .A1(DIN[19]), .A2(n24), .ZN(n28) );
  NAND2_X1 U47 ( .A1(DOUT[19]), .A2(n12), .ZN(n29) );
  NAND2_X1 U48 ( .A1(n28), .A2(n29), .ZN(n84) );
  INV_X1 U49 ( .A(n41), .ZN(DOUT[8]) );
  MUX2_X1 U50 ( .A(n52), .B(DIN[8]), .S(EN), .Z(n73) );
  INV_X1 U51 ( .A(n42), .ZN(DOUT[9]) );
  MUX2_X1 U52 ( .A(n51), .B(DIN[9]), .S(EN), .Z(n74) );
  MUX2_X1 U53 ( .A(n9), .B(DIN[10]), .S(EN), .Z(n75) );
  MUX2_X1 U54 ( .A(DOUT[11]), .B(DIN[11]), .S(EN), .Z(n76) );
  MUX2_X1 U55 ( .A(DOUT[12]), .B(DIN[12]), .S(EN), .Z(n77) );
  MUX2_X1 U56 ( .A(DOUT[13]), .B(DIN[13]), .S(EN), .Z(n78) );
  MUX2_X1 U57 ( .A(DOUT[14]), .B(DIN[14]), .S(EN), .Z(n79) );
  MUX2_X1 U58 ( .A(DOUT[16]), .B(DIN[16]), .S(EN), .Z(n81) );
  MUX2_X1 U59 ( .A(DOUT[17]), .B(DIN[17]), .S(EN), .Z(n82) );
  MUX2_X1 U60 ( .A(DOUT[18]), .B(DIN[18]), .S(EN), .Z(n83) );
  INV_X1 U61 ( .A(n53), .ZN(n49) );
  MUX2_X1 U62 ( .A(n49), .B(DIN[20]), .S(EN), .Z(n85) );
  MUX2_X1 U63 ( .A(DOUT[21]), .B(DIN[21]), .S(EN), .Z(n86) );
  MUX2_X1 U64 ( .A(DOUT[22]), .B(DIN[22]), .S(EN), .Z(n87) );
  MUX2_X1 U65 ( .A(DOUT[24]), .B(DIN[24]), .S(EN), .Z(n89) );
  MUX2_X1 U66 ( .A(DOUT[26]), .B(DIN[26]), .S(EN), .Z(n91) );
  MUX2_X1 U67 ( .A(DOUT[30]), .B(DIN[30]), .S(EN), .Z(n95) );
endmodule


module regn_N32_10 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U6 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U7 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U8 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U9 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U10 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U11 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U12 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U13 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U14 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U15 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U16 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U17 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U18 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U19 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U20 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U21 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U22 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U23 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U24 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U25 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U26 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U27 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U28 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U29 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U30 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U31 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U32 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U33 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U34 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U35 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U36 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U37 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U38 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U39 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U40 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U41 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U42 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U43 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U44 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U45 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U46 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U47 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U48 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U49 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U50 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U51 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U52 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U53 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U54 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U55 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U56 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U57 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U58 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U59 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U60 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U61 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
endmodule


module regn_N32_9 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U6 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U7 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U8 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U9 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U10 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U11 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U12 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U13 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U14 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U15 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U16 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U17 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U18 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U19 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U20 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U21 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U22 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U23 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U24 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U25 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U26 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U27 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U28 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U29 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U30 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U31 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U32 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U33 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U34 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U35 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U36 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U37 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U38 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U39 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U40 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U41 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U42 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U43 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U44 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U45 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U46 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U47 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U48 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U49 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U50 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U51 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U52 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U53 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U54 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U55 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U56 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U57 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U58 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U59 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U60 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U61 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U62 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U63 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U64 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
  OAI21_X1 U65 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U66 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U67 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U68 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
endmodule


module Fetch_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AND2_X1 U2 ( .A1(n11), .A2(n42), .ZN(n36) );
  AND2_X1 U3 ( .A1(n54), .A2(n92), .ZN(n49) );
  AND3_X1 U4 ( .A1(A[11]), .A2(A[13]), .A3(A[12]), .ZN(n1) );
  AND2_X1 U5 ( .A1(A[25]), .A2(A[24]), .ZN(n2) );
  AND3_X1 U6 ( .A1(n12), .A2(A[14]), .A3(A[15]), .ZN(n3) );
  NOR2_X1 U7 ( .A1(n27), .A2(n70), .ZN(n4) );
  AND2_X1 U8 ( .A1(n10), .A2(n42), .ZN(n5) );
  AND4_X1 U9 ( .A1(A[25]), .A2(A[24]), .A3(n10), .A4(n42), .ZN(n73) );
  AND3_X1 U10 ( .A1(n37), .A2(n14), .A3(n4), .ZN(n30) );
  NOR2_X1 U11 ( .A1(n95), .A2(n94), .ZN(n52) );
  AND4_X1 U12 ( .A1(A[26]), .A2(n22), .A3(n5), .A4(n2), .ZN(n72) );
  AND4_X1 U13 ( .A1(n83), .A2(n84), .A3(A[16]), .A4(A[17]), .ZN(n47) );
  AND4_X1 U14 ( .A1(n67), .A2(n34), .A3(n36), .A4(A[30]), .ZN(n15) );
  AND3_X1 U15 ( .A1(n54), .A2(n92), .A3(A[13]), .ZN(n90) );
  AND3_X2 U16 ( .A1(n23), .A2(n3), .A3(n1), .ZN(n22) );
  XOR2_X1 U17 ( .A(A[25]), .B(n51), .Z(SUM[25]) );
  AND3_X1 U18 ( .A1(n14), .A2(n36), .A3(n6), .ZN(n41) );
  INV_X1 U19 ( .A(n27), .ZN(n6) );
  NAND4_X1 U20 ( .A1(A[10]), .A2(A[6]), .A3(A[8]), .A4(A[9]), .ZN(n87) );
  BUF_X1 U21 ( .A(A[6]), .Z(n7) );
  AND2_X1 U22 ( .A1(A[22]), .A2(A[23]), .ZN(n8) );
  AND2_X1 U23 ( .A1(A[22]), .A2(A[23]), .ZN(n24) );
  AND2_X2 U24 ( .A1(n61), .A2(n9), .ZN(n56) );
  AND4_X1 U25 ( .A1(n32), .A2(A[5]), .A3(n7), .A4(A[4]), .ZN(n9) );
  XNOR2_X1 U26 ( .A(n44), .B(n98), .ZN(SUM[10]) );
  AND2_X1 U27 ( .A1(n8), .A2(n25), .ZN(n10) );
  AND2_X1 U28 ( .A1(n24), .A2(n25), .ZN(n11) );
  AND2_X1 U29 ( .A1(n8), .A2(n25), .ZN(n74) );
  AND2_X1 U30 ( .A1(A[3]), .A2(A[7]), .ZN(n12) );
  CLKBUF_X1 U31 ( .A(n7), .Z(n13) );
  AND2_X1 U32 ( .A1(n84), .A2(n83), .ZN(n14) );
  AND2_X1 U33 ( .A1(n83), .A2(n84), .ZN(n34) );
  XOR2_X1 U34 ( .A(A[31]), .B(n15), .Z(SUM[31]) );
  XOR2_X1 U35 ( .A(n16), .B(A[21]), .Z(SUM[21]) );
  AND2_X1 U36 ( .A1(n78), .A2(n22), .ZN(n16) );
  CLKBUF_X1 U37 ( .A(n22), .Z(n17) );
  AND3_X1 U38 ( .A1(n34), .A2(n67), .A3(n36), .ZN(n48) );
  XNOR2_X1 U39 ( .A(A[23]), .B(n18), .ZN(SUM[23]) );
  NAND2_X1 U40 ( .A1(n22), .A2(n31), .ZN(n18) );
  AND3_X1 U41 ( .A1(A[5]), .A2(A[6]), .A3(A[4]), .ZN(n19) );
  AND2_X1 U42 ( .A1(n32), .A2(n19), .ZN(n28) );
  CLKBUF_X1 U43 ( .A(A[7]), .Z(n32) );
  AND2_X1 U44 ( .A1(A[22]), .A2(n20), .ZN(n21) );
  INV_X1 U45 ( .A(n76), .ZN(n20) );
  NOR2_X1 U46 ( .A1(n87), .A2(n88), .ZN(n23) );
  AND2_X1 U47 ( .A1(A[20]), .A2(A[21]), .ZN(n25) );
  OR2_X1 U48 ( .A1(n69), .A2(n70), .ZN(n26) );
  NAND4_X1 U49 ( .A1(A[24]), .A2(A[25]), .A3(A[26]), .A4(A[27]), .ZN(n27) );
  AND2_X1 U50 ( .A1(n37), .A2(A[24]), .ZN(n29) );
  XOR2_X1 U51 ( .A(A[29]), .B(n30), .Z(SUM[29]) );
  AND2_X1 U52 ( .A1(n42), .A2(n21), .ZN(n31) );
  AND2_X1 U53 ( .A1(n22), .A2(n75), .ZN(n33) );
  AND2_X1 U54 ( .A1(n56), .A2(n35), .ZN(n99) );
  NOR2_X1 U55 ( .A1(n96), .A2(n97), .ZN(n35) );
  AND2_X1 U56 ( .A1(n74), .A2(n42), .ZN(n37) );
  NOR2_X1 U57 ( .A1(n66), .A2(SUM[2]), .ZN(n38) );
  NOR2_X1 U58 ( .A1(n66), .A2(SUM[2]), .ZN(n61) );
  AND2_X1 U59 ( .A1(n37), .A2(n22), .ZN(n39) );
  AND2_X1 U60 ( .A1(A[3]), .A2(A[7]), .ZN(n40) );
  AND4_X2 U61 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(A[19]), .ZN(n42) );
  NOR2_X1 U62 ( .A1(n26), .A2(n27), .ZN(n67) );
  NAND3_X1 U63 ( .A1(n40), .A2(A[14]), .A3(A[15]), .ZN(n85) );
  AND2_X1 U64 ( .A1(n47), .A2(A[18]), .ZN(n81) );
  XOR2_X1 U65 ( .A(A[19]), .B(n81), .Z(SUM[19]) );
  XNOR2_X1 U66 ( .A(n41), .B(n70), .ZN(SUM[28]) );
  XOR2_X1 U67 ( .A(n43), .B(A[11]), .Z(SUM[11]) );
  AND2_X1 U68 ( .A1(A[10]), .A2(n99), .ZN(n43) );
  NOR2_X1 U69 ( .A1(n55), .A2(n97), .ZN(n44) );
  AND2_X1 U70 ( .A1(n45), .A2(A[5]), .ZN(n59) );
  NAND4_X1 U71 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(A[19]), .ZN(n77) );
  AND2_X1 U72 ( .A1(n61), .A2(n62), .ZN(n45) );
  AND2_X1 U73 ( .A1(n73), .A2(n22), .ZN(n46) );
  INV_X1 U74 ( .A(n66), .ZN(n65) );
  AND2_X1 U75 ( .A1(n28), .A2(n38), .ZN(n54) );
  INV_X1 U76 ( .A(n64), .ZN(n62) );
  INV_X1 U77 ( .A(n96), .ZN(n57) );
  NAND2_X1 U78 ( .A1(A[21]), .A2(A[20]), .ZN(n76) );
  AND2_X1 U79 ( .A1(n13), .A2(n59), .ZN(n50) );
  AND2_X1 U80 ( .A1(n22), .A2(n29), .ZN(n51) );
  INV_X1 U81 ( .A(A[27]), .ZN(n71) );
  INV_X1 U82 ( .A(A[2]), .ZN(SUM[2]) );
  INV_X1 U83 ( .A(A[14]), .ZN(n91) );
  XOR2_X1 U84 ( .A(A[22]), .B(n33), .Z(SUM[22]) );
  XNOR2_X1 U85 ( .A(n52), .B(n93), .ZN(SUM[12]) );
  XOR2_X1 U86 ( .A(n55), .B(n97), .Z(SUM[9]) );
  XOR2_X1 U87 ( .A(A[13]), .B(n49), .Z(SUM[13]) );
  XOR2_X1 U88 ( .A(n46), .B(A[26]), .Z(SUM[26]) );
  XOR2_X1 U89 ( .A(n48), .B(A[30]), .Z(SUM[30]) );
  XOR2_X1 U90 ( .A(n47), .B(A[18]), .Z(SUM[18]) );
  XNOR2_X1 U91 ( .A(n53), .B(n89), .ZN(SUM[15]) );
  AND2_X1 U92 ( .A1(A[14]), .A2(n90), .ZN(n53) );
  XOR2_X1 U93 ( .A(n39), .B(A[24]), .Z(SUM[24]) );
  XOR2_X1 U94 ( .A(n17), .B(A[16]), .Z(SUM[16]) );
  XOR2_X1 U95 ( .A(n56), .B(n57), .Z(SUM[8]) );
  XNOR2_X1 U96 ( .A(n80), .B(A[20]), .ZN(SUM[20]) );
  XNOR2_X1 U97 ( .A(n82), .B(A[17]), .ZN(SUM[17]) );
  INV_X1 U98 ( .A(A[28]), .ZN(n70) );
  XNOR2_X1 U99 ( .A(n63), .B(n45), .ZN(SUM[5]) );
  XNOR2_X1 U100 ( .A(SUM[2]), .B(n65), .ZN(SUM[3]) );
  INV_X1 U101 ( .A(A[29]), .ZN(n69) );
  INV_X1 U102 ( .A(n32), .ZN(n58) );
  NOR2_X1 U103 ( .A1(n93), .A2(n94), .ZN(n92) );
  INV_X1 U104 ( .A(n54), .ZN(n95) );
  INV_X1 U105 ( .A(A[4]), .ZN(n64) );
  NOR2_X1 U106 ( .A1(n87), .A2(n88), .ZN(n83) );
  XNOR2_X1 U107 ( .A(n58), .B(n50), .ZN(SUM[7]) );
  NOR2_X1 U108 ( .A1(n77), .A2(n76), .ZN(n75) );
  NOR2_X1 U109 ( .A1(n79), .A2(n77), .ZN(n78) );
  NOR2_X1 U110 ( .A1(n85), .A2(n86), .ZN(n84) );
  NAND4_X1 U111 ( .A1(A[10]), .A2(A[9]), .A3(A[8]), .A4(A[11]), .ZN(n94) );
  INV_X1 U112 ( .A(A[5]), .ZN(n63) );
  INV_X1 U113 ( .A(A[10]), .ZN(n98) );
  NAND2_X1 U114 ( .A1(n56), .A2(n57), .ZN(n55) );
  INV_X1 U115 ( .A(n13), .ZN(n60) );
  XNOR2_X1 U116 ( .A(n60), .B(n59), .ZN(SUM[6]) );
  XNOR2_X1 U117 ( .A(n64), .B(n38), .ZN(SUM[4]) );
  INV_X1 U118 ( .A(A[8]), .ZN(n96) );
  NAND2_X1 U119 ( .A1(n22), .A2(n42), .ZN(n80) );
  NAND2_X1 U120 ( .A1(n22), .A2(A[16]), .ZN(n82) );
  INV_X1 U121 ( .A(A[9]), .ZN(n97) );
  XNOR2_X1 U122 ( .A(n72), .B(n71), .ZN(SUM[27]) );
  INV_X1 U123 ( .A(A[20]), .ZN(n79) );
  NAND3_X1 U124 ( .A1(A[11]), .A2(A[13]), .A3(A[12]), .ZN(n86) );
  NAND3_X1 U125 ( .A1(A[5]), .A2(A[2]), .A3(A[4]), .ZN(n88) );
  INV_X1 U126 ( .A(A[15]), .ZN(n89) );
  XNOR2_X1 U127 ( .A(n91), .B(n90), .ZN(SUM[14]) );
  INV_X1 U128 ( .A(A[12]), .ZN(n93) );
  INV_X1 U129 ( .A(A[3]), .ZN(n66) );
endmodule


module Fetch ( CLK, RST, ZERO_FLAG, PC_EXT, INS_IN, Bubble_in, HDU_INS_IN, 
        HDU_PC_IN, HDU_NPC_IN, PC_OUT, ADDR_OUT, NPC_OUT, INS_OUT );
  input [31:0] PC_EXT;
  input [31:0] INS_IN;
  input [31:0] HDU_INS_IN;
  input [31:0] HDU_PC_IN;
  input [31:0] HDU_NPC_IN;
  output [31:0] PC_OUT;
  output [31:0] ADDR_OUT;
  output [31:0] NPC_OUT;
  output [31:0] INS_OUT;
  input CLK, RST, ZERO_FLAG, Bubble_in;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         sig_RST, n18;
  wire   [31:0] sig_NPC;
  wire   [31:0] PC_MUX_OUT;
  wire   [31:0] sig_INS;

  mux21_NBIT32_0 NPC_or_NPC_HDU ( .A(PC_EXT), .B(HDU_NPC_IN), .S(Bubble_in), 
        .Z(sig_NPC) );
  mux21_NBIT32_5 PC_or_PC_HDU ( .A(ADDR_OUT), .B(HDU_PC_IN), .S(Bubble_in), 
        .Z(PC_MUX_OUT) );
  mux21_NBIT32_4 INS_or_HDU_INS ( .A(INS_IN), .B(HDU_INS_IN), .S(Bubble_in), 
        .Z(sig_INS) );
  regn_N32_0 PC ( .DIN(sig_NPC), .CLK(CLK), .EN(1'b1), .RST(RST), .DOUT({
        ADDR_OUT[31:30], n19, ADDR_OUT[28:24], n20, ADDR_OUT[22:18], n21, n22, 
        ADDR_OUT[15], n23, ADDR_OUT[13], n24, ADDR_OUT[11:10], n25, n26, n27, 
        n28, n29, n30, n31, n32, ADDR_OUT[1:0]}) );
  regn_N32_10 PC_reg ( .DIN(PC_MUX_OUT), .CLK(CLK), .EN(1'b1), .RST(sig_RST), 
        .DOUT(PC_OUT) );
  regn_N32_9 IR ( .DIN(sig_INS), .CLK(CLK), .EN(1'b1), .RST(sig_RST), .DOUT(
        INS_OUT) );
  Fetch_DW01_add_1 add_54 ( .A({ADDR_OUT[31:30], n19, ADDR_OUT[28:24], n20, 
        ADDR_OUT[22:18], n21, n22, ADDR_OUT[15], n23, ADDR_OUT[13], n24, 
        ADDR_OUT[11:10], n25, n26, n27, n28, n29, n30, n31, n32, ADDR_OUT[1:0]}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(
        NPC_OUT) );
  CLKBUF_X1 U6 ( .A(n26), .Z(ADDR_OUT[8]) );
  CLKBUF_X1 U7 ( .A(n19), .Z(ADDR_OUT[29]) );
  CLKBUF_X1 U8 ( .A(n27), .Z(ADDR_OUT[7]) );
  CLKBUF_X1 U9 ( .A(n32), .Z(ADDR_OUT[2]) );
  CLKBUF_X1 U10 ( .A(n20), .Z(ADDR_OUT[23]) );
  CLKBUF_X1 U11 ( .A(n24), .Z(ADDR_OUT[12]) );
  CLKBUF_X1 U12 ( .A(n28), .Z(ADDR_OUT[6]) );
  CLKBUF_X1 U13 ( .A(n31), .Z(ADDR_OUT[3]) );
  CLKBUF_X1 U14 ( .A(n21), .Z(ADDR_OUT[17]) );
  CLKBUF_X1 U15 ( .A(n22), .Z(ADDR_OUT[16]) );
  NOR2_X1 U16 ( .A1(ZERO_FLAG), .A2(n18), .ZN(sig_RST) );
  CLKBUF_X1 U17 ( .A(n29), .Z(ADDR_OUT[5]) );
  CLKBUF_X1 U18 ( .A(n23), .Z(ADDR_OUT[14]) );
  CLKBUF_X1 U19 ( .A(n30), .Z(ADDR_OUT[4]) );
  CLKBUF_X1 U20 ( .A(n25), .Z(ADDR_OUT[9]) );
  INV_X1 U21 ( .A(RST), .ZN(n18) );
endmodule


module instruction_type ( INST_IN, Rtype, Itype, Jtype );
  input [31:0] INST_IN;
  output Rtype, Itype, Jtype;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n1, n2, n3, n4, n5,
         n6, n7, n8;

  OAI33_X1 U21 ( .A1(n5), .A2(INST_IN[29]), .A3(n2), .B1(n4), .B2(INST_IN[30]), 
        .B3(INST_IN[26]), .ZN(n17) );
  NOR2_X1 U1 ( .A1(n9), .A2(n10), .ZN(Rtype) );
  OAI22_X1 U2 ( .A1(n10), .A2(n5), .B1(n7), .B2(n4), .ZN(n16) );
  NOR2_X1 U3 ( .A1(n9), .A2(n6), .ZN(Jtype) );
  NAND4_X1 U4 ( .A1(n5), .A2(n4), .A3(n3), .A4(n1), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n6), .A2(n8), .ZN(n10) );
  INV_X1 U6 ( .A(n14), .ZN(n7) );
  INV_X1 U7 ( .A(n18), .ZN(n2) );
  OAI221_X1 U8 ( .B1(n7), .B2(INST_IN[30]), .C1(n3), .C2(INST_IN[26]), .A(n10), 
        .ZN(n18) );
  OAI211_X1 U9 ( .C1(INST_IN[31]), .C2(n11), .A(n12), .B(n13), .ZN(Itype) );
  NAND4_X1 U10 ( .A1(INST_IN[29]), .A2(INST_IN[28]), .A3(n14), .A4(n1), .ZN(
        n13) );
  NAND4_X1 U11 ( .A1(INST_IN[31]), .A2(INST_IN[27]), .A3(n15), .A4(INST_IN[26]), .ZN(n12) );
  AOI21_X1 U12 ( .B1(INST_IN[30]), .B2(n16), .A(n17), .ZN(n11) );
  NOR2_X1 U13 ( .A1(n8), .A2(INST_IN[27]), .ZN(n14) );
  NOR2_X1 U14 ( .A1(INST_IN[30]), .A2(INST_IN[28]), .ZN(n15) );
  INV_X1 U15 ( .A(INST_IN[30]), .ZN(n3) );
  INV_X1 U16 ( .A(INST_IN[28]), .ZN(n5) );
  INV_X1 U17 ( .A(INST_IN[29]), .ZN(n4) );
  INV_X1 U18 ( .A(INST_IN[26]), .ZN(n8) );
  INV_X1 U19 ( .A(INST_IN[31]), .ZN(n1) );
  INV_X1 U20 ( .A(INST_IN[27]), .ZN(n6) );
endmodule


module instruction_decomposition ( INST_IN, Rtype, Itype, Jtype, ADD_RS1, 
        ADD_RS2, ADD_WR, IMM );
  input [31:0] INST_IN;
  output [4:0] ADD_RS1;
  output [4:0] ADD_RS2;
  output [4:0] ADD_WR;
  output [31:0] IMM;
  input Rtype, Itype, Jtype;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n1, n2,
         \IMM[31] , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20;
  assign IMM[25] = \IMM[31] ;
  assign IMM[26] = \IMM[31] ;
  assign IMM[27] = \IMM[31] ;
  assign IMM[28] = \IMM[31] ;
  assign IMM[29] = \IMM[31] ;
  assign IMM[30] = \IMM[31] ;
  assign IMM[31] = \IMM[31] ;

  NAND3_X1 U72 ( .A1(INST_IN[29]), .A2(INST_IN[27]), .A3(INST_IN[31]), .ZN(n31) );
  NAND3_X1 U73 ( .A1(INST_IN[26]), .A2(Itype), .A3(n32), .ZN(n30) );
  INV_X1 U2 ( .A(Rtype), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n28), .A2(Jtype), .ZN(n24) );
  INV_X1 U4 ( .A(n27), .ZN(n2) );
  OAI21_X1 U5 ( .B1(Itype), .B2(Jtype), .A(n4), .ZN(n27) );
  NOR2_X1 U6 ( .A1(Rtype), .A2(Itype), .ZN(n28) );
  NOR2_X1 U7 ( .A1(n28), .A2(n10), .ZN(ADD_RS1[0]) );
  NOR2_X1 U8 ( .A1(n1), .A2(n15), .ZN(ADD_RS2[0]) );
  NOR2_X1 U9 ( .A1(n28), .A2(n7), .ZN(ADD_RS1[3]) );
  NOR2_X1 U10 ( .A1(n1), .A2(n12), .ZN(ADD_RS2[3]) );
  NOR2_X1 U11 ( .A1(n1), .A2(n11), .ZN(ADD_RS2[4]) );
  NOR2_X1 U12 ( .A1(n28), .A2(n8), .ZN(ADD_RS1[2]) );
  NOR2_X1 U13 ( .A1(n1), .A2(n13), .ZN(ADD_RS2[2]) );
  OR2_X1 U14 ( .A1(n26), .A2(n16), .ZN(n25) );
  NOR2_X1 U15 ( .A1(n28), .A2(n9), .ZN(ADD_RS1[1]) );
  NOR2_X1 U16 ( .A1(n1), .A2(n14), .ZN(ADD_RS2[1]) );
  NAND2_X1 U17 ( .A1(Itype), .A2(n4), .ZN(n26) );
  INV_X1 U18 ( .A(Itype), .ZN(n5) );
  AND2_X1 U19 ( .A1(INST_IN[0]), .A2(n2), .ZN(IMM[0]) );
  AND2_X1 U20 ( .A1(INST_IN[1]), .A2(n2), .ZN(IMM[1]) );
  AND2_X1 U21 ( .A1(INST_IN[2]), .A2(n2), .ZN(IMM[2]) );
  AND2_X1 U22 ( .A1(INST_IN[3]), .A2(n2), .ZN(IMM[3]) );
  AND2_X1 U23 ( .A1(INST_IN[4]), .A2(n2), .ZN(IMM[4]) );
  AND2_X1 U24 ( .A1(INST_IN[5]), .A2(n2), .ZN(IMM[5]) );
  AND2_X1 U25 ( .A1(INST_IN[6]), .A2(n2), .ZN(IMM[6]) );
  AND2_X1 U26 ( .A1(INST_IN[7]), .A2(n2), .ZN(IMM[7]) );
  AND2_X1 U27 ( .A1(INST_IN[8]), .A2(n2), .ZN(IMM[8]) );
  AND2_X1 U28 ( .A1(INST_IN[9]), .A2(n2), .ZN(IMM[9]) );
  AND2_X1 U29 ( .A1(INST_IN[10]), .A2(n2), .ZN(IMM[10]) );
  NOR2_X1 U30 ( .A1(n27), .A2(n20), .ZN(IMM[11]) );
  NOR2_X1 U31 ( .A1(n27), .A2(n19), .ZN(IMM[12]) );
  NOR2_X1 U32 ( .A1(n27), .A2(n18), .ZN(IMM[13]) );
  NOR2_X1 U33 ( .A1(n27), .A2(n17), .ZN(IMM[14]) );
  NOR2_X1 U34 ( .A1(n27), .A2(n16), .ZN(IMM[15]) );
  OAI21_X1 U35 ( .B1(n24), .B2(n15), .A(n25), .ZN(IMM[16]) );
  OAI21_X1 U36 ( .B1(n24), .B2(n14), .A(n25), .ZN(IMM[17]) );
  OAI21_X1 U37 ( .B1(n24), .B2(n13), .A(n25), .ZN(IMM[18]) );
  OAI21_X1 U38 ( .B1(n24), .B2(n12), .A(n25), .ZN(IMM[19]) );
  OAI21_X1 U39 ( .B1(n24), .B2(n11), .A(n25), .ZN(IMM[20]) );
  OAI21_X1 U40 ( .B1(n24), .B2(n10), .A(n25), .ZN(IMM[21]) );
  OAI21_X1 U41 ( .B1(n24), .B2(n9), .A(n25), .ZN(IMM[22]) );
  OAI21_X1 U42 ( .B1(n24), .B2(n8), .A(n25), .ZN(IMM[23]) );
  OAI21_X1 U43 ( .B1(n24), .B2(n7), .A(n25), .ZN(IMM[24]) );
  OAI221_X1 U44 ( .B1(n26), .B2(n15), .C1(n20), .C2(n4), .A(n24), .ZN(
        ADD_WR[0]) );
  OAI221_X1 U45 ( .B1(n26), .B2(n14), .C1(n19), .C2(n4), .A(n24), .ZN(
        ADD_WR[1]) );
  OAI221_X1 U46 ( .B1(n26), .B2(n13), .C1(n18), .C2(n4), .A(n24), .ZN(
        ADD_WR[2]) );
  OAI221_X1 U47 ( .B1(n26), .B2(n12), .C1(n17), .C2(n4), .A(n24), .ZN(
        ADD_WR[3]) );
  OAI221_X1 U48 ( .B1(n26), .B2(n11), .C1(n16), .C2(n4), .A(n24), .ZN(
        ADD_WR[4]) );
  NOR2_X1 U49 ( .A1(n28), .A2(n6), .ZN(ADD_RS1[4]) );
  INV_X1 U50 ( .A(INST_IN[25]), .ZN(n6) );
  INV_X1 U51 ( .A(n21), .ZN(\IMM[31] ) );
  OAI21_X1 U52 ( .B1(n22), .B2(n23), .A(n4), .ZN(n21) );
  AND3_X1 U53 ( .A1(Jtype), .A2(n5), .A3(INST_IN[25]), .ZN(n22) );
  NOR2_X1 U54 ( .A1(n16), .A2(n5), .ZN(n23) );
  INV_X1 U55 ( .A(n29), .ZN(n1) );
  OAI21_X1 U56 ( .B1(n30), .B2(n31), .A(n4), .ZN(n29) );
  INV_X1 U57 ( .A(INST_IN[15]), .ZN(n16) );
  INV_X1 U58 ( .A(INST_IN[16]), .ZN(n15) );
  INV_X1 U59 ( .A(INST_IN[17]), .ZN(n14) );
  INV_X1 U60 ( .A(INST_IN[19]), .ZN(n12) );
  INV_X1 U61 ( .A(INST_IN[18]), .ZN(n13) );
  INV_X1 U62 ( .A(INST_IN[20]), .ZN(n11) );
  NOR2_X1 U63 ( .A1(INST_IN[30]), .A2(INST_IN[28]), .ZN(n32) );
  INV_X1 U64 ( .A(INST_IN[21]), .ZN(n10) );
  INV_X1 U65 ( .A(INST_IN[22]), .ZN(n9) );
  INV_X1 U66 ( .A(INST_IN[24]), .ZN(n7) );
  INV_X1 U67 ( .A(INST_IN[23]), .ZN(n8) );
  INV_X1 U68 ( .A(INST_IN[11]), .ZN(n20) );
  INV_X1 U69 ( .A(INST_IN[12]), .ZN(n19) );
  INV_X1 U70 ( .A(INST_IN[13]), .ZN(n18) );
  INV_X1 U71 ( .A(INST_IN[14]), .ZN(n17) );
endmodule


module regn_N32_8 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U6 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U7 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U8 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U9 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U10 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U11 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U12 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U13 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U14 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U15 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U16 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U17 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U18 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U19 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U20 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U21 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U22 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U23 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U24 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U25 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U26 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U27 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U28 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U29 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U30 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U31 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U32 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U33 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U34 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U35 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U36 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U37 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U38 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U39 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U40 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U41 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U42 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U43 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U44 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U45 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U46 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U47 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U48 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U49 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U50 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U51 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U52 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U53 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U54 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U55 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U56 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U57 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U58 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U59 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U60 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U61 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U62 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U63 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U64 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
  OAI21_X1 U65 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U66 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U67 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U68 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
endmodule


module regn_N32_7 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
endmodule


module regn_N5_0 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  DFFR_X1 \DOUT_reg[4]  ( .D(n15), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n10)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n14), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n9) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n13), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n8) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n12), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n7) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n11), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n6) );
  OAI21_X1 U2 ( .B1(n6), .B2(EN), .A(n1), .ZN(n11) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n1) );
  OAI21_X1 U4 ( .B1(n7), .B2(EN), .A(n2), .ZN(n12) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n2) );
  OAI21_X1 U6 ( .B1(n8), .B2(EN), .A(n3), .ZN(n13) );
  NAND2_X1 U7 ( .A1(DIN[2]), .A2(EN), .ZN(n3) );
  OAI21_X1 U8 ( .B1(n9), .B2(EN), .A(n4), .ZN(n14) );
  NAND2_X1 U9 ( .A1(DIN[3]), .A2(EN), .ZN(n4) );
  OAI21_X1 U10 ( .B1(n10), .B2(EN), .A(n5), .ZN(n15) );
  NAND2_X1 U11 ( .A1(DIN[4]), .A2(EN), .ZN(n5) );
endmodule


module regn_N5_4 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 \DOUT_reg[4]  ( .D(n16), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n21)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n17), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n22)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n18), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n23)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n19), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n24)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n20), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n25)
         );
  OAI21_X1 U2 ( .B1(n25), .B2(EN), .A(n30), .ZN(n20) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n30) );
  OAI21_X1 U4 ( .B1(n24), .B2(EN), .A(n29), .ZN(n19) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n29) );
  OAI21_X1 U6 ( .B1(n23), .B2(EN), .A(n28), .ZN(n18) );
  NAND2_X1 U7 ( .A1(DIN[2]), .A2(EN), .ZN(n28) );
  OAI21_X1 U8 ( .B1(n22), .B2(EN), .A(n27), .ZN(n17) );
  NAND2_X1 U9 ( .A1(DIN[3]), .A2(EN), .ZN(n27) );
  OAI21_X1 U10 ( .B1(n21), .B2(EN), .A(n26), .ZN(n16) );
  NAND2_X1 U11 ( .A1(DIN[4]), .A2(EN), .ZN(n26) );
endmodule


module regn_N5_3 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 \DOUT_reg[4]  ( .D(n16), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n21)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n17), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n22)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n18), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n23)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n19), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n24)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n20), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n25)
         );
  OAI21_X1 U2 ( .B1(n25), .B2(EN), .A(n30), .ZN(n20) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n30) );
  OAI21_X1 U4 ( .B1(n24), .B2(EN), .A(n29), .ZN(n19) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n29) );
  OAI21_X1 U6 ( .B1(n23), .B2(EN), .A(n28), .ZN(n18) );
  NAND2_X1 U7 ( .A1(DIN[2]), .A2(EN), .ZN(n28) );
  OAI21_X1 U8 ( .B1(n22), .B2(EN), .A(n27), .ZN(n17) );
  NAND2_X1 U9 ( .A1(DIN[3]), .A2(EN), .ZN(n27) );
  OAI21_X1 U10 ( .B1(n21), .B2(EN), .A(n26), .ZN(n16) );
  NAND2_X1 U11 ( .A1(DIN[4]), .A2(EN), .ZN(n26) );
endmodule


module register_file_NBIT_ADD5_NBIT_DATA32 ( CLK, RST, ENABLE, RD1, RD2, WR, 
        ADD_WR, ADD_RS1, ADD_RS2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RST, ENABLE, RD1, RD2, WR;
  wire   n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344;

  DFFR_X1 \REGISTERS_reg[1][31]  ( .D(n4024), .CK(CLK), .RN(n378), .Q(n603) );
  DFFR_X1 \REGISTERS_reg[1][30]  ( .D(n4023), .CK(CLK), .RN(n337), .Q(n602) );
  DFFR_X1 \REGISTERS_reg[1][29]  ( .D(n4022), .CK(CLK), .RN(n368), .Q(n601) );
  DFFR_X1 \REGISTERS_reg[1][28]  ( .D(n4021), .CK(CLK), .RN(n367), .Q(n600) );
  DFFR_X1 \REGISTERS_reg[1][27]  ( .D(n4020), .CK(CLK), .RN(n367), .Q(n599) );
  DFFR_X1 \REGISTERS_reg[1][26]  ( .D(n4019), .CK(CLK), .RN(n367), .Q(n598) );
  DFFR_X1 \REGISTERS_reg[1][25]  ( .D(n4018), .CK(CLK), .RN(n367), .Q(n597) );
  DFFR_X1 \REGISTERS_reg[1][24]  ( .D(n4017), .CK(CLK), .RN(n367), .Q(n596) );
  DFFR_X1 \REGISTERS_reg[1][23]  ( .D(n4016), .CK(CLK), .RN(n367), .Q(n595) );
  DFFR_X1 \REGISTERS_reg[1][22]  ( .D(n4015), .CK(CLK), .RN(n367), .Q(n594) );
  DFFR_X1 \REGISTERS_reg[1][21]  ( .D(n4014), .CK(CLK), .RN(n367), .Q(n593) );
  DFFR_X1 \REGISTERS_reg[1][20]  ( .D(n4013), .CK(CLK), .RN(n367), .Q(n592) );
  DFFR_X1 \REGISTERS_reg[1][19]  ( .D(n4012), .CK(CLK), .RN(n367), .Q(n591) );
  DFFR_X1 \REGISTERS_reg[1][18]  ( .D(n4011), .CK(CLK), .RN(n367), .Q(n590) );
  DFFR_X1 \REGISTERS_reg[1][17]  ( .D(n4010), .CK(CLK), .RN(n367), .Q(n589) );
  DFFR_X1 \REGISTERS_reg[1][16]  ( .D(n4009), .CK(CLK), .RN(n366), .Q(n588) );
  DFFR_X1 \REGISTERS_reg[1][15]  ( .D(n4008), .CK(CLK), .RN(n366), .Q(n587) );
  DFFR_X1 \REGISTERS_reg[1][14]  ( .D(n4007), .CK(CLK), .RN(n366), .Q(n586) );
  DFFR_X1 \REGISTERS_reg[1][13]  ( .D(n4006), .CK(CLK), .RN(n366), .Q(n585) );
  DFFR_X1 \REGISTERS_reg[1][12]  ( .D(n4005), .CK(CLK), .RN(n366), .Q(n584) );
  DFFR_X1 \REGISTERS_reg[1][11]  ( .D(n4004), .CK(CLK), .RN(n366), .Q(n583) );
  DFFR_X1 \REGISTERS_reg[1][10]  ( .D(n4003), .CK(CLK), .RN(n366), .Q(n582) );
  DFFR_X1 \REGISTERS_reg[1][9]  ( .D(n4002), .CK(CLK), .RN(n366), .Q(n581) );
  DFFR_X1 \REGISTERS_reg[1][8]  ( .D(n4001), .CK(CLK), .RN(n366), .Q(n580) );
  DFFR_X1 \REGISTERS_reg[1][7]  ( .D(n4000), .CK(CLK), .RN(n366), .Q(n579) );
  DFFR_X1 \REGISTERS_reg[1][6]  ( .D(n3999), .CK(CLK), .RN(n366), .Q(n578) );
  DFFR_X1 \REGISTERS_reg[1][5]  ( .D(n3998), .CK(CLK), .RN(n366), .Q(n577) );
  DFFR_X1 \REGISTERS_reg[1][4]  ( .D(n3997), .CK(CLK), .RN(n365), .Q(n576) );
  DFFR_X1 \REGISTERS_reg[1][3]  ( .D(n3996), .CK(CLK), .RN(n365), .Q(n575) );
  DFFR_X1 \REGISTERS_reg[1][2]  ( .D(n3995), .CK(CLK), .RN(n365), .Q(n574) );
  DFFR_X1 \REGISTERS_reg[1][1]  ( .D(n3994), .CK(CLK), .RN(n365), .Q(n573) );
  DFFR_X1 \REGISTERS_reg[1][0]  ( .D(n3993), .CK(CLK), .RN(n365), .Q(n571) );
  DFFR_X1 \REGISTERS_reg[4][31]  ( .D(n4056), .CK(CLK), .RN(n360), .Q(n637) );
  DFFR_X1 \REGISTERS_reg[4][30]  ( .D(n4055), .CK(CLK), .RN(n360), .Q(n636) );
  DFFR_X1 \REGISTERS_reg[4][29]  ( .D(n4054), .CK(CLK), .RN(n359), .Q(n635) );
  DFFR_X1 \REGISTERS_reg[4][28]  ( .D(n4053), .CK(CLK), .RN(n359), .Q(n634) );
  DFFR_X1 \REGISTERS_reg[4][27]  ( .D(n4052), .CK(CLK), .RN(n359), .Q(n633) );
  DFFR_X1 \REGISTERS_reg[4][26]  ( .D(n4051), .CK(CLK), .RN(n359), .Q(n632) );
  DFFR_X1 \REGISTERS_reg[4][25]  ( .D(n4050), .CK(CLK), .RN(n359), .Q(n631) );
  DFFR_X1 \REGISTERS_reg[4][24]  ( .D(n4049), .CK(CLK), .RN(n359), .Q(n630) );
  DFFR_X1 \REGISTERS_reg[4][23]  ( .D(n4048), .CK(CLK), .RN(n359), .Q(n629) );
  DFFR_X1 \REGISTERS_reg[4][22]  ( .D(n4047), .CK(CLK), .RN(n359), .Q(n628) );
  DFFR_X1 \REGISTERS_reg[4][21]  ( .D(n4046), .CK(CLK), .RN(n359), .Q(n627) );
  DFFR_X1 \REGISTERS_reg[4][20]  ( .D(n4045), .CK(CLK), .RN(n359), .Q(n626) );
  DFFR_X1 \REGISTERS_reg[4][19]  ( .D(n4044), .CK(CLK), .RN(n359), .Q(n625) );
  DFFR_X1 \REGISTERS_reg[4][18]  ( .D(n4043), .CK(CLK), .RN(n359), .Q(n624) );
  DFFR_X1 \REGISTERS_reg[4][17]  ( .D(n4042), .CK(CLK), .RN(n358), .Q(n623) );
  DFFR_X1 \REGISTERS_reg[4][16]  ( .D(n4041), .CK(CLK), .RN(n358), .Q(n622) );
  DFFR_X1 \REGISTERS_reg[4][15]  ( .D(n4040), .CK(CLK), .RN(n358), .Q(n621) );
  DFFR_X1 \REGISTERS_reg[4][14]  ( .D(n4039), .CK(CLK), .RN(n358), .Q(n620) );
  DFFR_X1 \REGISTERS_reg[4][13]  ( .D(n4038), .CK(CLK), .RN(n358), .Q(n619) );
  DFFR_X1 \REGISTERS_reg[4][12]  ( .D(n4037), .CK(CLK), .RN(n358), .Q(n618) );
  DFFR_X1 \REGISTERS_reg[4][11]  ( .D(n4036), .CK(CLK), .RN(n358), .Q(n617) );
  DFFR_X1 \REGISTERS_reg[4][10]  ( .D(n4035), .CK(CLK), .RN(n358), .Q(n616) );
  DFFR_X1 \REGISTERS_reg[4][9]  ( .D(n4034), .CK(CLK), .RN(n358), .Q(n615) );
  DFFR_X1 \REGISTERS_reg[4][8]  ( .D(n4033), .CK(CLK), .RN(n358), .Q(n614) );
  DFFR_X1 \REGISTERS_reg[4][7]  ( .D(n4032), .CK(CLK), .RN(n358), .Q(n613) );
  DFFR_X1 \REGISTERS_reg[4][6]  ( .D(n4031), .CK(CLK), .RN(n358), .Q(n612) );
  DFFR_X1 \REGISTERS_reg[4][5]  ( .D(n4030), .CK(CLK), .RN(n357), .Q(n611) );
  DFFR_X1 \REGISTERS_reg[4][4]  ( .D(n4029), .CK(CLK), .RN(n357), .Q(n610) );
  DFFR_X1 \REGISTERS_reg[4][3]  ( .D(n4028), .CK(CLK), .RN(n357), .Q(n609) );
  DFFR_X1 \REGISTERS_reg[4][2]  ( .D(n4027), .CK(CLK), .RN(n362), .Q(n608) );
  DFFR_X1 \REGISTERS_reg[4][1]  ( .D(n4026), .CK(CLK), .RN(n378), .Q(n607) );
  DFFR_X1 \REGISTERS_reg[4][0]  ( .D(n4025), .CK(CLK), .RN(n378), .Q(n605) );
  DFFR_X1 \REGISTERS_reg[5][31]  ( .D(n4088), .CK(CLK), .RN(n378), .Q(n670) );
  DFFR_X1 \REGISTERS_reg[5][30]  ( .D(n4087), .CK(CLK), .RN(n378), .Q(n669) );
  DFFR_X1 \REGISTERS_reg[5][29]  ( .D(n4086), .CK(CLK), .RN(n377), .Q(n668) );
  DFFR_X1 \REGISTERS_reg[5][28]  ( .D(n4085), .CK(CLK), .RN(n377), .Q(n667) );
  DFFR_X1 \REGISTERS_reg[5][27]  ( .D(n4084), .CK(CLK), .RN(n377), .Q(n666) );
  DFFR_X1 \REGISTERS_reg[5][26]  ( .D(n4083), .CK(CLK), .RN(n377), .Q(n665) );
  DFFR_X1 \REGISTERS_reg[5][25]  ( .D(n4082), .CK(CLK), .RN(n377), .Q(n664) );
  DFFR_X1 \REGISTERS_reg[5][24]  ( .D(n4081), .CK(CLK), .RN(n377), .Q(n663) );
  DFFR_X1 \REGISTERS_reg[5][23]  ( .D(n4080), .CK(CLK), .RN(n377), .Q(n662) );
  DFFR_X1 \REGISTERS_reg[5][22]  ( .D(n4079), .CK(CLK), .RN(n377), .Q(n661) );
  DFFR_X1 \REGISTERS_reg[5][21]  ( .D(n4078), .CK(CLK), .RN(n377), .Q(n660) );
  DFFR_X1 \REGISTERS_reg[5][20]  ( .D(n4077), .CK(CLK), .RN(n377), .Q(n659) );
  DFFR_X1 \REGISTERS_reg[5][19]  ( .D(n4076), .CK(CLK), .RN(n377), .Q(n658) );
  DFFR_X1 \REGISTERS_reg[5][18]  ( .D(n4075), .CK(CLK), .RN(n377), .Q(n657) );
  DFFR_X1 \REGISTERS_reg[5][17]  ( .D(n4074), .CK(CLK), .RN(n376), .Q(n656) );
  DFFR_X1 \REGISTERS_reg[5][16]  ( .D(n4073), .CK(CLK), .RN(n376), .Q(n655) );
  DFFR_X1 \REGISTERS_reg[5][15]  ( .D(n4072), .CK(CLK), .RN(n376), .Q(n654) );
  DFFR_X1 \REGISTERS_reg[5][14]  ( .D(n4071), .CK(CLK), .RN(n376), .Q(n653) );
  DFFR_X1 \REGISTERS_reg[5][13]  ( .D(n4070), .CK(CLK), .RN(n376), .Q(n652) );
  DFFR_X1 \REGISTERS_reg[5][12]  ( .D(n4069), .CK(CLK), .RN(n376), .Q(n651) );
  DFFR_X1 \REGISTERS_reg[5][11]  ( .D(n4068), .CK(CLK), .RN(n376), .Q(n650) );
  DFFR_X1 \REGISTERS_reg[5][10]  ( .D(n4067), .CK(CLK), .RN(n376), .Q(n649) );
  DFFR_X1 \REGISTERS_reg[5][9]  ( .D(n4066), .CK(CLK), .RN(n376), .Q(n648) );
  DFFR_X1 \REGISTERS_reg[5][8]  ( .D(n4065), .CK(CLK), .RN(n376), .Q(n647) );
  DFFR_X1 \REGISTERS_reg[5][7]  ( .D(n4064), .CK(CLK), .RN(n376), .Q(n646) );
  DFFR_X1 \REGISTERS_reg[5][6]  ( .D(n4063), .CK(CLK), .RN(n376), .Q(n645) );
  DFFR_X1 \REGISTERS_reg[5][5]  ( .D(n4062), .CK(CLK), .RN(n375), .Q(n644) );
  DFFR_X1 \REGISTERS_reg[5][4]  ( .D(n4061), .CK(CLK), .RN(n375), .Q(n643) );
  DFFR_X1 \REGISTERS_reg[5][3]  ( .D(n4060), .CK(CLK), .RN(n375), .Q(n642) );
  DFFR_X1 \REGISTERS_reg[5][2]  ( .D(n4059), .CK(CLK), .RN(n375), .Q(n641) );
  DFFR_X1 \REGISTERS_reg[5][1]  ( .D(n4058), .CK(CLK), .RN(n375), .Q(n640) );
  DFFR_X1 \REGISTERS_reg[5][0]  ( .D(n4057), .CK(CLK), .RN(n375), .Q(n638) );
  DFFR_X1 \REGISTERS_reg[8][31]  ( .D(n3896), .CK(CLK), .RN(n370), .QN(n2494)
         );
  DFFR_X1 \REGISTERS_reg[8][30]  ( .D(n3895), .CK(CLK), .RN(n369), .QN(n2515)
         );
  DFFR_X1 \REGISTERS_reg[8][29]  ( .D(n3894), .CK(CLK), .RN(n369), .QN(n2536)
         );
  DFFR_X1 \REGISTERS_reg[8][28]  ( .D(n3893), .CK(CLK), .RN(n369), .QN(n2557)
         );
  DFFR_X1 \REGISTERS_reg[8][27]  ( .D(n3892), .CK(CLK), .RN(n369), .QN(n2578)
         );
  DFFR_X1 \REGISTERS_reg[8][26]  ( .D(n3891), .CK(CLK), .RN(n369), .QN(n2599)
         );
  DFFR_X1 \REGISTERS_reg[8][25]  ( .D(n3890), .CK(CLK), .RN(n369), .QN(n2620)
         );
  DFFR_X1 \REGISTERS_reg[8][24]  ( .D(n3889), .CK(CLK), .RN(n369), .QN(n2641)
         );
  DFFR_X1 \REGISTERS_reg[8][23]  ( .D(n3888), .CK(CLK), .RN(n369), .QN(n2662)
         );
  DFFR_X1 \REGISTERS_reg[8][22]  ( .D(n3887), .CK(CLK), .RN(n369), .QN(n2683)
         );
  DFFR_X1 \REGISTERS_reg[8][21]  ( .D(n3886), .CK(CLK), .RN(n369), .QN(n2704)
         );
  DFFR_X1 \REGISTERS_reg[8][20]  ( .D(n3885), .CK(CLK), .RN(n369), .QN(n2725)
         );
  DFFR_X1 \REGISTERS_reg[8][19]  ( .D(n3884), .CK(CLK), .RN(n369), .QN(n2746)
         );
  DFFR_X1 \REGISTERS_reg[8][18]  ( .D(n3883), .CK(CLK), .RN(n368), .QN(n2767)
         );
  DFFR_X1 \REGISTERS_reg[8][17]  ( .D(n3882), .CK(CLK), .RN(n368), .QN(n2788)
         );
  DFFR_X1 \REGISTERS_reg[8][16]  ( .D(n3881), .CK(CLK), .RN(n368), .QN(n2809)
         );
  DFFR_X1 \REGISTERS_reg[8][15]  ( .D(n3880), .CK(CLK), .RN(n368), .QN(n2830)
         );
  DFFR_X1 \REGISTERS_reg[8][14]  ( .D(n3879), .CK(CLK), .RN(n368), .QN(n2851)
         );
  DFFR_X1 \REGISTERS_reg[8][13]  ( .D(n3878), .CK(CLK), .RN(n368), .QN(n2872)
         );
  DFFR_X1 \REGISTERS_reg[8][12]  ( .D(n3877), .CK(CLK), .RN(n368), .QN(n2893)
         );
  DFFR_X1 \REGISTERS_reg[8][11]  ( .D(n3876), .CK(CLK), .RN(n368), .QN(n2914)
         );
  DFFR_X1 \REGISTERS_reg[8][10]  ( .D(n3875), .CK(CLK), .RN(n368), .QN(n2935)
         );
  DFFR_X1 \REGISTERS_reg[8][9]  ( .D(n3874), .CK(CLK), .RN(n368), .QN(n2956)
         );
  DFFR_X1 \REGISTERS_reg[8][8]  ( .D(n3873), .CK(CLK), .RN(n368), .QN(n2977)
         );
  DFFR_X1 \REGISTERS_reg[8][7]  ( .D(n3872), .CK(CLK), .RN(n373), .QN(n3574)
         );
  DFFR_X1 \REGISTERS_reg[8][6]  ( .D(n3871), .CK(CLK), .RN(n347), .QN(n3595)
         );
  DFFR_X1 \REGISTERS_reg[8][5]  ( .D(n3870), .CK(CLK), .RN(n347), .QN(n3616)
         );
  DFFR_X1 \REGISTERS_reg[8][4]  ( .D(n3869), .CK(CLK), .RN(n347), .QN(n3637)
         );
  DFFR_X1 \REGISTERS_reg[8][3]  ( .D(n3868), .CK(CLK), .RN(n347), .QN(n3658)
         );
  DFFR_X1 \REGISTERS_reg[8][2]  ( .D(n3867), .CK(CLK), .RN(n347), .QN(n3679)
         );
  DFFR_X1 \REGISTERS_reg[8][1]  ( .D(n3866), .CK(CLK), .RN(n346), .QN(n3700)
         );
  DFFR_X1 \REGISTERS_reg[8][0]  ( .D(n3865), .CK(CLK), .RN(n346), .QN(n3721)
         );
  DFFR_X1 \REGISTERS_reg[9][31]  ( .D(n3928), .CK(CLK), .RN(n346), .QN(n2495)
         );
  DFFR_X1 \REGISTERS_reg[9][30]  ( .D(n3927), .CK(CLK), .RN(n346), .QN(n2516)
         );
  DFFR_X1 \REGISTERS_reg[9][29]  ( .D(n3926), .CK(CLK), .RN(n346), .QN(n2537)
         );
  DFFR_X1 \REGISTERS_reg[9][28]  ( .D(n3925), .CK(CLK), .RN(n346), .QN(n2558)
         );
  DFFR_X1 \REGISTERS_reg[9][27]  ( .D(n3924), .CK(CLK), .RN(n346), .QN(n2579)
         );
  DFFR_X1 \REGISTERS_reg[9][26]  ( .D(n3923), .CK(CLK), .RN(n346), .QN(n2600)
         );
  DFFR_X1 \REGISTERS_reg[9][25]  ( .D(n3922), .CK(CLK), .RN(n346), .QN(n2621)
         );
  DFFR_X1 \REGISTERS_reg[9][24]  ( .D(n3921), .CK(CLK), .RN(n346), .QN(n2642)
         );
  DFFR_X1 \REGISTERS_reg[9][23]  ( .D(n3920), .CK(CLK), .RN(n346), .QN(n2663)
         );
  DFFR_X1 \REGISTERS_reg[9][22]  ( .D(n3919), .CK(CLK), .RN(n346), .QN(n2684)
         );
  DFFR_X1 \REGISTERS_reg[9][21]  ( .D(n3918), .CK(CLK), .RN(n345), .QN(n2705)
         );
  DFFR_X1 \REGISTERS_reg[9][20]  ( .D(n3917), .CK(CLK), .RN(n345), .QN(n2726)
         );
  DFFR_X1 \REGISTERS_reg[9][19]  ( .D(n3916), .CK(CLK), .RN(n345), .QN(n2747)
         );
  DFFR_X1 \REGISTERS_reg[9][18]  ( .D(n3915), .CK(CLK), .RN(n345), .QN(n2768)
         );
  DFFR_X1 \REGISTERS_reg[9][17]  ( .D(n3914), .CK(CLK), .RN(n345), .QN(n2789)
         );
  DFFR_X1 \REGISTERS_reg[9][16]  ( .D(n3913), .CK(CLK), .RN(n345), .QN(n2810)
         );
  DFFR_X1 \REGISTERS_reg[9][15]  ( .D(n3912), .CK(CLK), .RN(n345), .QN(n2831)
         );
  DFFR_X1 \REGISTERS_reg[9][14]  ( .D(n3911), .CK(CLK), .RN(n345), .QN(n2852)
         );
  DFFR_X1 \REGISTERS_reg[9][13]  ( .D(n3910), .CK(CLK), .RN(n345), .QN(n2873)
         );
  DFFR_X1 \REGISTERS_reg[9][12]  ( .D(n3909), .CK(CLK), .RN(n345), .QN(n2894)
         );
  DFFR_X1 \REGISTERS_reg[9][11]  ( .D(n3908), .CK(CLK), .RN(n345), .QN(n2915)
         );
  DFFR_X1 \REGISTERS_reg[9][10]  ( .D(n3907), .CK(CLK), .RN(n345), .QN(n2936)
         );
  DFFR_X1 \REGISTERS_reg[9][9]  ( .D(n3906), .CK(CLK), .RN(n344), .QN(n2957)
         );
  DFFR_X1 \REGISTERS_reg[9][8]  ( .D(n3905), .CK(CLK), .RN(n344), .QN(n2978)
         );
  DFFR_X1 \REGISTERS_reg[9][7]  ( .D(n3904), .CK(CLK), .RN(n344), .QN(n3575)
         );
  DFFR_X1 \REGISTERS_reg[9][6]  ( .D(n3903), .CK(CLK), .RN(n344), .QN(n3596)
         );
  DFFR_X1 \REGISTERS_reg[9][5]  ( .D(n3902), .CK(CLK), .RN(n344), .QN(n3617)
         );
  DFFR_X1 \REGISTERS_reg[9][4]  ( .D(n3901), .CK(CLK), .RN(n344), .QN(n3638)
         );
  DFFR_X1 \REGISTERS_reg[9][3]  ( .D(n3900), .CK(CLK), .RN(n344), .QN(n3659)
         );
  DFFR_X1 \REGISTERS_reg[9][2]  ( .D(n3899), .CK(CLK), .RN(n344), .QN(n3680)
         );
  DFFR_X1 \REGISTERS_reg[9][1]  ( .D(n3898), .CK(CLK), .RN(n344), .QN(n3701)
         );
  DFFR_X1 \REGISTERS_reg[9][0]  ( .D(n3897), .CK(CLK), .RN(n344), .QN(n3722)
         );
  DFFR_X1 \REGISTERS_reg[10][31]  ( .D(n3430), .CK(CLK), .RN(n344), .Q(n2497)
         );
  DFFR_X1 \REGISTERS_reg[10][30]  ( .D(n3429), .CK(CLK), .RN(n344), .Q(n2518)
         );
  DFFR_X1 \REGISTERS_reg[10][29]  ( .D(n3428), .CK(CLK), .RN(n343), .Q(n2539)
         );
  DFFR_X1 \REGISTERS_reg[10][28]  ( .D(n3427), .CK(CLK), .RN(n343), .Q(n2560)
         );
  DFFR_X1 \REGISTERS_reg[10][27]  ( .D(n3426), .CK(CLK), .RN(n343), .Q(n2581)
         );
  DFFR_X1 \REGISTERS_reg[10][26]  ( .D(n3425), .CK(CLK), .RN(n343), .Q(n2602)
         );
  DFFR_X1 \REGISTERS_reg[10][25]  ( .D(n3424), .CK(CLK), .RN(n343), .Q(n2623)
         );
  DFFR_X1 \REGISTERS_reg[10][24]  ( .D(n3423), .CK(CLK), .RN(n343), .Q(n2644)
         );
  DFFR_X1 \REGISTERS_reg[10][23]  ( .D(n3422), .CK(CLK), .RN(n343), .Q(n2665)
         );
  DFFR_X1 \REGISTERS_reg[10][22]  ( .D(n3421), .CK(CLK), .RN(n343), .Q(n2686)
         );
  DFFR_X1 \REGISTERS_reg[10][21]  ( .D(n3420), .CK(CLK), .RN(n343), .Q(n2707)
         );
  DFFR_X1 \REGISTERS_reg[10][20]  ( .D(n3419), .CK(CLK), .RN(n343), .Q(n2728)
         );
  DFFR_X1 \REGISTERS_reg[10][19]  ( .D(n3418), .CK(CLK), .RN(n343), .Q(n2749)
         );
  DFFR_X1 \REGISTERS_reg[10][18]  ( .D(n3417), .CK(CLK), .RN(n343), .Q(n2770)
         );
  DFFR_X1 \REGISTERS_reg[10][17]  ( .D(n3416), .CK(CLK), .RN(n342), .Q(n2791)
         );
  DFFR_X1 \REGISTERS_reg[10][16]  ( .D(n3415), .CK(CLK), .RN(n342), .Q(n2812)
         );
  DFFR_X1 \REGISTERS_reg[10][15]  ( .D(n3414), .CK(CLK), .RN(n342), .Q(n2833)
         );
  DFFR_X1 \REGISTERS_reg[10][14]  ( .D(n3413), .CK(CLK), .RN(n342), .Q(n2854)
         );
  DFFR_X1 \REGISTERS_reg[10][13]  ( .D(n3412), .CK(CLK), .RN(n342), .Q(n2875)
         );
  DFFR_X1 \REGISTERS_reg[10][12]  ( .D(n3411), .CK(CLK), .RN(n342), .Q(n2896)
         );
  DFFR_X1 \REGISTERS_reg[10][11]  ( .D(n3410), .CK(CLK), .RN(n342), .Q(n2917)
         );
  DFFR_X1 \REGISTERS_reg[10][10]  ( .D(n3409), .CK(CLK), .RN(n342), .Q(n2938)
         );
  DFFR_X1 \REGISTERS_reg[10][9]  ( .D(n3408), .CK(CLK), .RN(n342), .Q(n2959)
         );
  DFFR_X1 \REGISTERS_reg[10][8]  ( .D(n3407), .CK(CLK), .RN(n342), .Q(n2980)
         );
  DFFR_X1 \REGISTERS_reg[10][7]  ( .D(n3406), .CK(CLK), .RN(n342), .Q(n3577)
         );
  DFFR_X1 \REGISTERS_reg[10][6]  ( .D(n3405), .CK(CLK), .RN(n341), .Q(n3598)
         );
  DFFR_X1 \REGISTERS_reg[10][5]  ( .D(n3404), .CK(CLK), .RN(n341), .Q(n3619)
         );
  DFFR_X1 \REGISTERS_reg[10][4]  ( .D(n3403), .CK(CLK), .RN(n341), .Q(n3640)
         );
  DFFR_X1 \REGISTERS_reg[10][3]  ( .D(n3402), .CK(CLK), .RN(n341), .Q(n3661)
         );
  DFFR_X1 \REGISTERS_reg[10][2]  ( .D(n3401), .CK(CLK), .RN(n341), .Q(n3682)
         );
  DFFR_X1 \REGISTERS_reg[10][1]  ( .D(n3400), .CK(CLK), .RN(n341), .Q(n3703)
         );
  DFFR_X1 \REGISTERS_reg[10][0]  ( .D(n3399), .CK(CLK), .RN(n341), .Q(n3724)
         );
  DFFR_X1 \REGISTERS_reg[11][31]  ( .D(n3398), .CK(CLK), .RN(n341), .Q(n2496)
         );
  DFFR_X1 \REGISTERS_reg[11][30]  ( .D(n3397), .CK(CLK), .RN(n341), .Q(n2517)
         );
  DFFR_X1 \REGISTERS_reg[11][29]  ( .D(n3396), .CK(CLK), .RN(n341), .Q(n2538)
         );
  DFFR_X1 \REGISTERS_reg[11][28]  ( .D(n3395), .CK(CLK), .RN(n341), .Q(n2559)
         );
  DFFR_X1 \REGISTERS_reg[11][27]  ( .D(n3394), .CK(CLK), .RN(n341), .Q(n2580)
         );
  DFFR_X1 \REGISTERS_reg[11][26]  ( .D(n3393), .CK(CLK), .RN(n340), .Q(n2601)
         );
  DFFR_X1 \REGISTERS_reg[11][25]  ( .D(n3392), .CK(CLK), .RN(n340), .Q(n2622)
         );
  DFFR_X1 \REGISTERS_reg[11][24]  ( .D(n3391), .CK(CLK), .RN(n340), .Q(n2643)
         );
  DFFR_X1 \REGISTERS_reg[11][23]  ( .D(n3390), .CK(CLK), .RN(n340), .Q(n2664)
         );
  DFFR_X1 \REGISTERS_reg[11][22]  ( .D(n3389), .CK(CLK), .RN(n340), .Q(n2685)
         );
  DFFR_X1 \REGISTERS_reg[11][21]  ( .D(n3388), .CK(CLK), .RN(n340), .Q(n2706)
         );
  DFFR_X1 \REGISTERS_reg[11][20]  ( .D(n3387), .CK(CLK), .RN(n340), .Q(n2727)
         );
  DFFR_X1 \REGISTERS_reg[11][19]  ( .D(n3386), .CK(CLK), .RN(n340), .Q(n2748)
         );
  DFFR_X1 \REGISTERS_reg[11][18]  ( .D(n3385), .CK(CLK), .RN(n340), .Q(n2769)
         );
  DFFR_X1 \REGISTERS_reg[11][17]  ( .D(n3384), .CK(CLK), .RN(n340), .Q(n2790)
         );
  DFFR_X1 \REGISTERS_reg[11][16]  ( .D(n3383), .CK(CLK), .RN(n340), .Q(n2811)
         );
  DFFR_X1 \REGISTERS_reg[11][15]  ( .D(n3382), .CK(CLK), .RN(n340), .Q(n2832)
         );
  DFFR_X1 \REGISTERS_reg[11][14]  ( .D(n3381), .CK(CLK), .RN(n339), .Q(n2853)
         );
  DFFR_X1 \REGISTERS_reg[11][13]  ( .D(n3380), .CK(CLK), .RN(n339), .Q(n2874)
         );
  DFFR_X1 \REGISTERS_reg[11][12]  ( .D(n3379), .CK(CLK), .RN(n339), .Q(n2895)
         );
  DFFR_X1 \REGISTERS_reg[11][11]  ( .D(n3378), .CK(CLK), .RN(n339), .Q(n2916)
         );
  DFFR_X1 \REGISTERS_reg[11][10]  ( .D(n3377), .CK(CLK), .RN(n339), .Q(n2937)
         );
  DFFR_X1 \REGISTERS_reg[11][9]  ( .D(n3376), .CK(CLK), .RN(n339), .Q(n2958)
         );
  DFFR_X1 \REGISTERS_reg[11][8]  ( .D(n3375), .CK(CLK), .RN(n339), .Q(n2979)
         );
  DFFR_X1 \REGISTERS_reg[11][7]  ( .D(n3374), .CK(CLK), .RN(n339), .Q(n3576)
         );
  DFFR_X1 \REGISTERS_reg[11][6]  ( .D(n3373), .CK(CLK), .RN(n339), .Q(n3597)
         );
  DFFR_X1 \REGISTERS_reg[11][5]  ( .D(n3372), .CK(CLK), .RN(n339), .Q(n3618)
         );
  DFFR_X1 \REGISTERS_reg[11][4]  ( .D(n3371), .CK(CLK), .RN(n339), .Q(n3639)
         );
  DFFR_X1 \REGISTERS_reg[11][3]  ( .D(n3370), .CK(CLK), .RN(n339), .Q(n3660)
         );
  DFFR_X1 \REGISTERS_reg[11][2]  ( .D(n3369), .CK(CLK), .RN(n338), .Q(n3681)
         );
  DFFR_X1 \REGISTERS_reg[11][1]  ( .D(n3368), .CK(CLK), .RN(n338), .Q(n3702)
         );
  DFFR_X1 \REGISTERS_reg[11][0]  ( .D(n3367), .CK(CLK), .RN(n338), .Q(n3723)
         );
  DFFR_X1 \REGISTERS_reg[12][31]  ( .D(n3960), .CK(CLK), .RN(n338), .QN(n2490)
         );
  DFFR_X1 \REGISTERS_reg[12][30]  ( .D(n3959), .CK(CLK), .RN(n338), .QN(n2511)
         );
  DFFR_X1 \REGISTERS_reg[12][29]  ( .D(n3958), .CK(CLK), .RN(n338), .QN(n2532)
         );
  DFFR_X1 \REGISTERS_reg[12][28]  ( .D(n3957), .CK(CLK), .RN(n338), .QN(n2553)
         );
  DFFR_X1 \REGISTERS_reg[12][27]  ( .D(n3956), .CK(CLK), .RN(n338), .QN(n2574)
         );
  DFFR_X1 \REGISTERS_reg[12][26]  ( .D(n3955), .CK(CLK), .RN(n338), .QN(n2595)
         );
  DFFR_X1 \REGISTERS_reg[12][25]  ( .D(n3954), .CK(CLK), .RN(n338), .QN(n2616)
         );
  DFFR_X1 \REGISTERS_reg[12][24]  ( .D(n3953), .CK(CLK), .RN(n338), .QN(n2637)
         );
  DFFR_X1 \REGISTERS_reg[12][23]  ( .D(n3952), .CK(CLK), .RN(n338), .QN(n2658)
         );
  DFFR_X1 \REGISTERS_reg[12][22]  ( .D(n3951), .CK(CLK), .RN(n337), .QN(n2679)
         );
  DFFR_X1 \REGISTERS_reg[12][21]  ( .D(n3950), .CK(CLK), .RN(n337), .QN(n2700)
         );
  DFFR_X1 \REGISTERS_reg[12][20]  ( .D(n3949), .CK(CLK), .RN(n337), .QN(n2721)
         );
  DFFR_X1 \REGISTERS_reg[12][19]  ( .D(n3948), .CK(CLK), .RN(n337), .QN(n2742)
         );
  DFFR_X1 \REGISTERS_reg[12][18]  ( .D(n3947), .CK(CLK), .RN(n337), .QN(n2763)
         );
  DFFR_X1 \REGISTERS_reg[12][17]  ( .D(n3946), .CK(CLK), .RN(n337), .QN(n2784)
         );
  DFFR_X1 \REGISTERS_reg[12][16]  ( .D(n3945), .CK(CLK), .RN(n337), .QN(n2805)
         );
  DFFR_X1 \REGISTERS_reg[12][15]  ( .D(n3944), .CK(CLK), .RN(n337), .QN(n2826)
         );
  DFFR_X1 \REGISTERS_reg[12][14]  ( .D(n3943), .CK(CLK), .RN(n337), .QN(n2847)
         );
  DFFR_X1 \REGISTERS_reg[12][13]  ( .D(n3942), .CK(CLK), .RN(n337), .QN(n2868)
         );
  DFFR_X1 \REGISTERS_reg[12][12]  ( .D(n3941), .CK(CLK), .RN(n337), .QN(n2889)
         );
  DFFR_X1 \REGISTERS_reg[12][11]  ( .D(n3940), .CK(CLK), .RN(n342), .QN(n2910)
         );
  DFFR_X1 \REGISTERS_reg[12][10]  ( .D(n3939), .CK(CLK), .RN(n357), .QN(n2931)
         );
  DFFR_X1 \REGISTERS_reg[12][9]  ( .D(n3938), .CK(CLK), .RN(n357), .QN(n2952)
         );
  DFFR_X1 \REGISTERS_reg[12][8]  ( .D(n3937), .CK(CLK), .RN(n357), .QN(n2973)
         );
  DFFR_X1 \REGISTERS_reg[12][7]  ( .D(n3936), .CK(CLK), .RN(n357), .QN(n3570)
         );
  DFFR_X1 \REGISTERS_reg[12][6]  ( .D(n3935), .CK(CLK), .RN(n357), .QN(n3591)
         );
  DFFR_X1 \REGISTERS_reg[12][5]  ( .D(n3934), .CK(CLK), .RN(n357), .QN(n3612)
         );
  DFFR_X1 \REGISTERS_reg[12][4]  ( .D(n3933), .CK(CLK), .RN(n357), .QN(n3633)
         );
  DFFR_X1 \REGISTERS_reg[12][3]  ( .D(n3932), .CK(CLK), .RN(n357), .QN(n3654)
         );
  DFFR_X1 \REGISTERS_reg[12][2]  ( .D(n3931), .CK(CLK), .RN(n356), .QN(n3675)
         );
  DFFR_X1 \REGISTERS_reg[12][1]  ( .D(n3930), .CK(CLK), .RN(n356), .QN(n3696)
         );
  DFFR_X1 \REGISTERS_reg[12][0]  ( .D(n3929), .CK(CLK), .RN(n356), .QN(n3717)
         );
  DFFR_X1 \REGISTERS_reg[13][31]  ( .D(n3992), .CK(CLK), .RN(n356), .QN(n2491)
         );
  DFFR_X1 \REGISTERS_reg[13][30]  ( .D(n3991), .CK(CLK), .RN(n356), .QN(n2512)
         );
  DFFR_X1 \REGISTERS_reg[13][29]  ( .D(n3990), .CK(CLK), .RN(n356), .QN(n2533)
         );
  DFFR_X1 \REGISTERS_reg[13][28]  ( .D(n3989), .CK(CLK), .RN(n356), .QN(n2554)
         );
  DFFR_X1 \REGISTERS_reg[13][27]  ( .D(n3988), .CK(CLK), .RN(n356), .QN(n2575)
         );
  DFFR_X1 \REGISTERS_reg[13][26]  ( .D(n3987), .CK(CLK), .RN(n356), .QN(n2596)
         );
  DFFR_X1 \REGISTERS_reg[13][25]  ( .D(n3986), .CK(CLK), .RN(n356), .QN(n2617)
         );
  DFFR_X1 \REGISTERS_reg[13][24]  ( .D(n3985), .CK(CLK), .RN(n356), .QN(n2638)
         );
  DFFR_X1 \REGISTERS_reg[13][23]  ( .D(n3984), .CK(CLK), .RN(n356), .QN(n2659)
         );
  DFFR_X1 \REGISTERS_reg[13][22]  ( .D(n3983), .CK(CLK), .RN(n355), .QN(n2680)
         );
  DFFR_X1 \REGISTERS_reg[13][21]  ( .D(n3982), .CK(CLK), .RN(n355), .QN(n2701)
         );
  DFFR_X1 \REGISTERS_reg[13][20]  ( .D(n3981), .CK(CLK), .RN(n355), .QN(n2722)
         );
  DFFR_X1 \REGISTERS_reg[13][19]  ( .D(n3980), .CK(CLK), .RN(n355), .QN(n2743)
         );
  DFFR_X1 \REGISTERS_reg[13][18]  ( .D(n3979), .CK(CLK), .RN(n355), .QN(n2764)
         );
  DFFR_X1 \REGISTERS_reg[13][17]  ( .D(n3978), .CK(CLK), .RN(n355), .QN(n2785)
         );
  DFFR_X1 \REGISTERS_reg[13][16]  ( .D(n3977), .CK(CLK), .RN(n355), .QN(n2806)
         );
  DFFR_X1 \REGISTERS_reg[13][15]  ( .D(n3976), .CK(CLK), .RN(n355), .QN(n2827)
         );
  DFFR_X1 \REGISTERS_reg[13][14]  ( .D(n3975), .CK(CLK), .RN(n355), .QN(n2848)
         );
  DFFR_X1 \REGISTERS_reg[13][13]  ( .D(n3974), .CK(CLK), .RN(n355), .QN(n2869)
         );
  DFFR_X1 \REGISTERS_reg[13][12]  ( .D(n3973), .CK(CLK), .RN(n355), .QN(n2890)
         );
  DFFR_X1 \REGISTERS_reg[13][11]  ( .D(n3972), .CK(CLK), .RN(n355), .QN(n2911)
         );
  DFFR_X1 \REGISTERS_reg[13][10]  ( .D(n3971), .CK(CLK), .RN(n354), .QN(n2932)
         );
  DFFR_X1 \REGISTERS_reg[13][9]  ( .D(n3970), .CK(CLK), .RN(n354), .QN(n2953)
         );
  DFFR_X1 \REGISTERS_reg[13][8]  ( .D(n3969), .CK(CLK), .RN(n354), .QN(n2974)
         );
  DFFR_X1 \REGISTERS_reg[13][7]  ( .D(n3968), .CK(CLK), .RN(n354), .QN(n3571)
         );
  DFFR_X1 \REGISTERS_reg[13][6]  ( .D(n3967), .CK(CLK), .RN(n354), .QN(n3592)
         );
  DFFR_X1 \REGISTERS_reg[13][5]  ( .D(n3966), .CK(CLK), .RN(n354), .QN(n3613)
         );
  DFFR_X1 \REGISTERS_reg[13][4]  ( .D(n3965), .CK(CLK), .RN(n354), .QN(n3634)
         );
  DFFR_X1 \REGISTERS_reg[13][3]  ( .D(n3964), .CK(CLK), .RN(n354), .QN(n3655)
         );
  DFFR_X1 \REGISTERS_reg[13][2]  ( .D(n3963), .CK(CLK), .RN(n354), .QN(n3676)
         );
  DFFR_X1 \REGISTERS_reg[13][1]  ( .D(n3962), .CK(CLK), .RN(n354), .QN(n3697)
         );
  DFFR_X1 \REGISTERS_reg[13][0]  ( .D(n3961), .CK(CLK), .RN(n354), .QN(n3718)
         );
  DFFR_X1 \REGISTERS_reg[14][31]  ( .D(n3366), .CK(CLK), .RN(n354), .Q(n2493)
         );
  DFFR_X1 \REGISTERS_reg[14][30]  ( .D(n3365), .CK(CLK), .RN(n353), .Q(n2514)
         );
  DFFR_X1 \REGISTERS_reg[14][29]  ( .D(n3364), .CK(CLK), .RN(n353), .Q(n2535)
         );
  DFFR_X1 \REGISTERS_reg[14][28]  ( .D(n3363), .CK(CLK), .RN(n353), .Q(n2556)
         );
  DFFR_X1 \REGISTERS_reg[14][27]  ( .D(n3362), .CK(CLK), .RN(n353), .Q(n2577)
         );
  DFFR_X1 \REGISTERS_reg[14][26]  ( .D(n3361), .CK(CLK), .RN(n353), .Q(n2598)
         );
  DFFR_X1 \REGISTERS_reg[14][25]  ( .D(n3360), .CK(CLK), .RN(n353), .Q(n2619)
         );
  DFFR_X1 \REGISTERS_reg[14][24]  ( .D(n3359), .CK(CLK), .RN(n353), .Q(n2640)
         );
  DFFR_X1 \REGISTERS_reg[14][23]  ( .D(n3358), .CK(CLK), .RN(n353), .Q(n2661)
         );
  DFFR_X1 \REGISTERS_reg[14][22]  ( .D(n3357), .CK(CLK), .RN(n353), .Q(n2682)
         );
  DFFR_X1 \REGISTERS_reg[14][21]  ( .D(n3356), .CK(CLK), .RN(n353), .Q(n2703)
         );
  DFFR_X1 \REGISTERS_reg[14][20]  ( .D(n3355), .CK(CLK), .RN(n353), .Q(n2724)
         );
  DFFR_X1 \REGISTERS_reg[14][19]  ( .D(n3354), .CK(CLK), .RN(n353), .Q(n2745)
         );
  DFFR_X1 \REGISTERS_reg[14][18]  ( .D(n3353), .CK(CLK), .RN(n352), .Q(n2766)
         );
  DFFR_X1 \REGISTERS_reg[14][17]  ( .D(n3352), .CK(CLK), .RN(n352), .Q(n2787)
         );
  DFFR_X1 \REGISTERS_reg[14][16]  ( .D(n3351), .CK(CLK), .RN(n352), .Q(n2808)
         );
  DFFR_X1 \REGISTERS_reg[14][15]  ( .D(n3350), .CK(CLK), .RN(n352), .Q(n2829)
         );
  DFFR_X1 \REGISTERS_reg[14][14]  ( .D(n3349), .CK(CLK), .RN(n352), .Q(n2850)
         );
  DFFR_X1 \REGISTERS_reg[14][13]  ( .D(n3348), .CK(CLK), .RN(n352), .Q(n2871)
         );
  DFFR_X1 \REGISTERS_reg[14][12]  ( .D(n3347), .CK(CLK), .RN(n352), .Q(n2892)
         );
  DFFR_X1 \REGISTERS_reg[14][11]  ( .D(n3346), .CK(CLK), .RN(n352), .Q(n2913)
         );
  DFFR_X1 \REGISTERS_reg[14][10]  ( .D(n3345), .CK(CLK), .RN(n352), .Q(n2934)
         );
  DFFR_X1 \REGISTERS_reg[14][9]  ( .D(n3344), .CK(CLK), .RN(n352), .Q(n2955)
         );
  DFFR_X1 \REGISTERS_reg[14][8]  ( .D(n3343), .CK(CLK), .RN(n352), .Q(n2976)
         );
  DFFR_X1 \REGISTERS_reg[14][7]  ( .D(n3342), .CK(CLK), .RN(n351), .Q(n3573)
         );
  DFFR_X1 \REGISTERS_reg[14][6]  ( .D(n3341), .CK(CLK), .RN(n351), .Q(n3594)
         );
  DFFR_X1 \REGISTERS_reg[14][5]  ( .D(n3340), .CK(CLK), .RN(n351), .Q(n3615)
         );
  DFFR_X1 \REGISTERS_reg[14][4]  ( .D(n3339), .CK(CLK), .RN(n351), .Q(n3636)
         );
  DFFR_X1 \REGISTERS_reg[14][3]  ( .D(n3338), .CK(CLK), .RN(n351), .Q(n3657)
         );
  DFFR_X1 \REGISTERS_reg[14][2]  ( .D(n3337), .CK(CLK), .RN(n351), .Q(n3678)
         );
  DFFR_X1 \REGISTERS_reg[14][1]  ( .D(n3336), .CK(CLK), .RN(n351), .Q(n3699)
         );
  DFFR_X1 \REGISTERS_reg[14][0]  ( .D(n3335), .CK(CLK), .RN(n351), .Q(n3720)
         );
  DFFR_X1 \REGISTERS_reg[15][31]  ( .D(n3334), .CK(CLK), .RN(n351), .Q(n2492)
         );
  DFFR_X1 \REGISTERS_reg[15][30]  ( .D(n3333), .CK(CLK), .RN(n351), .Q(n2513)
         );
  DFFR_X1 \REGISTERS_reg[15][29]  ( .D(n3332), .CK(CLK), .RN(n351), .Q(n2534)
         );
  DFFR_X1 \REGISTERS_reg[15][28]  ( .D(n3331), .CK(CLK), .RN(n351), .Q(n2555)
         );
  DFFR_X1 \REGISTERS_reg[15][27]  ( .D(n3330), .CK(CLK), .RN(n350), .Q(n2576)
         );
  DFFR_X1 \REGISTERS_reg[15][26]  ( .D(n3329), .CK(CLK), .RN(n350), .Q(n2597)
         );
  DFFR_X1 \REGISTERS_reg[15][25]  ( .D(n3328), .CK(CLK), .RN(n350), .Q(n2618)
         );
  DFFR_X1 \REGISTERS_reg[15][24]  ( .D(n3327), .CK(CLK), .RN(n350), .Q(n2639)
         );
  DFFR_X1 \REGISTERS_reg[15][23]  ( .D(n3326), .CK(CLK), .RN(n350), .Q(n2660)
         );
  DFFR_X1 \REGISTERS_reg[15][22]  ( .D(n3325), .CK(CLK), .RN(n350), .Q(n2681)
         );
  DFFR_X1 \REGISTERS_reg[15][21]  ( .D(n3324), .CK(CLK), .RN(n350), .Q(n2702)
         );
  DFFR_X1 \REGISTERS_reg[15][20]  ( .D(n3323), .CK(CLK), .RN(n350), .Q(n2723)
         );
  DFFR_X1 \REGISTERS_reg[15][19]  ( .D(n3322), .CK(CLK), .RN(n350), .Q(n2744)
         );
  DFFR_X1 \REGISTERS_reg[15][18]  ( .D(n3321), .CK(CLK), .RN(n350), .Q(n2765)
         );
  DFFR_X1 \REGISTERS_reg[15][17]  ( .D(n3320), .CK(CLK), .RN(n350), .Q(n2786)
         );
  DFFR_X1 \REGISTERS_reg[15][16]  ( .D(n3319), .CK(CLK), .RN(n350), .Q(n2807)
         );
  DFFR_X1 \REGISTERS_reg[15][15]  ( .D(n3318), .CK(CLK), .RN(n349), .Q(n2828)
         );
  DFFR_X1 \REGISTERS_reg[15][14]  ( .D(n3317), .CK(CLK), .RN(n349), .Q(n2849)
         );
  DFFR_X1 \REGISTERS_reg[15][13]  ( .D(n3316), .CK(CLK), .RN(n349), .Q(n2870)
         );
  DFFR_X1 \REGISTERS_reg[15][12]  ( .D(n3315), .CK(CLK), .RN(n349), .Q(n2891)
         );
  DFFR_X1 \REGISTERS_reg[15][11]  ( .D(n3314), .CK(CLK), .RN(n349), .Q(n2912)
         );
  DFFR_X1 \REGISTERS_reg[15][10]  ( .D(n3313), .CK(CLK), .RN(n349), .Q(n2933)
         );
  DFFR_X1 \REGISTERS_reg[15][9]  ( .D(n3312), .CK(CLK), .RN(n349), .Q(n2954)
         );
  DFFR_X1 \REGISTERS_reg[15][8]  ( .D(n3311), .CK(CLK), .RN(n349), .Q(n2975)
         );
  DFFR_X1 \REGISTERS_reg[15][7]  ( .D(n3310), .CK(CLK), .RN(n349), .Q(n3572)
         );
  DFFR_X1 \REGISTERS_reg[15][6]  ( .D(n3309), .CK(CLK), .RN(n349), .Q(n3593)
         );
  DFFR_X1 \REGISTERS_reg[15][5]  ( .D(n3308), .CK(CLK), .RN(n349), .Q(n3614)
         );
  DFFR_X1 \REGISTERS_reg[15][4]  ( .D(n3307), .CK(CLK), .RN(n349), .Q(n3635)
         );
  DFFR_X1 \REGISTERS_reg[15][3]  ( .D(n3306), .CK(CLK), .RN(n348), .Q(n3656)
         );
  DFFR_X1 \REGISTERS_reg[15][2]  ( .D(n3305), .CK(CLK), .RN(n348), .Q(n3677)
         );
  DFFR_X1 \REGISTERS_reg[15][1]  ( .D(n3304), .CK(CLK), .RN(n348), .Q(n3698)
         );
  DFFR_X1 \REGISTERS_reg[15][0]  ( .D(n3303), .CK(CLK), .RN(n348), .Q(n3719)
         );
  DFFR_X1 \REGISTERS_reg[16][31]  ( .D(n4248), .CK(CLK), .RN(n348), .Q(n840)
         );
  DFFR_X1 \REGISTERS_reg[16][30]  ( .D(n4247), .CK(CLK), .RN(n348), .Q(n839)
         );
  DFFR_X1 \REGISTERS_reg[16][29]  ( .D(n4246), .CK(CLK), .RN(n348), .Q(n838)
         );
  DFFR_X1 \REGISTERS_reg[16][28]  ( .D(n4245), .CK(CLK), .RN(n348), .Q(n837)
         );
  DFFR_X1 \REGISTERS_reg[16][27]  ( .D(n4244), .CK(CLK), .RN(n348), .Q(n836)
         );
  DFFR_X1 \REGISTERS_reg[16][26]  ( .D(n4243), .CK(CLK), .RN(n348), .Q(n835)
         );
  DFFR_X1 \REGISTERS_reg[16][25]  ( .D(n4242), .CK(CLK), .RN(n348), .Q(n834)
         );
  DFFR_X1 \REGISTERS_reg[16][24]  ( .D(n4241), .CK(CLK), .RN(n348), .Q(n833)
         );
  DFFR_X1 \REGISTERS_reg[16][23]  ( .D(n4240), .CK(CLK), .RN(n347), .Q(n832)
         );
  DFFR_X1 \REGISTERS_reg[16][22]  ( .D(n4239), .CK(CLK), .RN(n347), .Q(n831)
         );
  DFFR_X1 \REGISTERS_reg[16][21]  ( .D(n4238), .CK(CLK), .RN(n347), .Q(n830)
         );
  DFFR_X1 \REGISTERS_reg[16][20]  ( .D(n4237), .CK(CLK), .RN(n347), .Q(n829)
         );
  DFFR_X1 \REGISTERS_reg[16][19]  ( .D(n4236), .CK(CLK), .RN(n347), .Q(n828)
         );
  DFFR_X1 \REGISTERS_reg[16][18]  ( .D(n4235), .CK(CLK), .RN(n347), .Q(n827)
         );
  DFFR_X1 \REGISTERS_reg[16][17]  ( .D(n4234), .CK(CLK), .RN(n347), .Q(n826)
         );
  DFFR_X1 \REGISTERS_reg[16][16]  ( .D(n4233), .CK(CLK), .RN(n352), .Q(n825)
         );
  DFFR_X1 \REGISTERS_reg[16][15]  ( .D(n4232), .CK(CLK), .RN(n357), .Q(n824)
         );
  DFFR_X1 \REGISTERS_reg[16][14]  ( .D(n4231), .CK(CLK), .RN(n409), .Q(n823)
         );
  DFFR_X1 \REGISTERS_reg[16][13]  ( .D(n4230), .CK(CLK), .RN(n409), .Q(n822)
         );
  DFFR_X1 \REGISTERS_reg[16][12]  ( .D(n4229), .CK(CLK), .RN(n409), .Q(n821)
         );
  DFFR_X1 \REGISTERS_reg[16][11]  ( .D(n4228), .CK(CLK), .RN(n409), .Q(n820)
         );
  DFFR_X1 \REGISTERS_reg[16][10]  ( .D(n4227), .CK(CLK), .RN(n409), .Q(n819)
         );
  DFFR_X1 \REGISTERS_reg[16][9]  ( .D(n4226), .CK(CLK), .RN(n408), .Q(n818) );
  DFFR_X1 \REGISTERS_reg[16][8]  ( .D(n4225), .CK(CLK), .RN(n408), .Q(n817) );
  DFFR_X1 \REGISTERS_reg[16][7]  ( .D(n4224), .CK(CLK), .RN(n408), .Q(n816) );
  DFFR_X1 \REGISTERS_reg[16][6]  ( .D(n4223), .CK(CLK), .RN(n408), .Q(n815) );
  DFFR_X1 \REGISTERS_reg[16][5]  ( .D(n4222), .CK(CLK), .RN(n408), .Q(n814) );
  DFFR_X1 \REGISTERS_reg[16][4]  ( .D(n4221), .CK(CLK), .RN(n408), .Q(n813) );
  DFFR_X1 \REGISTERS_reg[16][3]  ( .D(n4220), .CK(CLK), .RN(n408), .Q(n812) );
  DFFR_X1 \REGISTERS_reg[16][2]  ( .D(n4219), .CK(CLK), .RN(n408), .Q(n811) );
  DFFR_X1 \REGISTERS_reg[16][1]  ( .D(n4218), .CK(CLK), .RN(n408), .Q(n810) );
  DFFR_X1 \REGISTERS_reg[16][0]  ( .D(n4217), .CK(CLK), .RN(n408), .Q(n808) );
  DFFR_X1 \REGISTERS_reg[17][31]  ( .D(n4280), .CK(CLK), .RN(n408), .QN(n2507)
         );
  DFFR_X1 \REGISTERS_reg[17][30]  ( .D(n4279), .CK(CLK), .RN(n408), .QN(n2528)
         );
  DFFR_X1 \REGISTERS_reg[17][29]  ( .D(n4278), .CK(CLK), .RN(n407), .QN(n2549)
         );
  DFFR_X1 \REGISTERS_reg[17][28]  ( .D(n4277), .CK(CLK), .RN(n407), .QN(n2570)
         );
  DFFR_X1 \REGISTERS_reg[17][27]  ( .D(n4276), .CK(CLK), .RN(n407), .QN(n2591)
         );
  DFFR_X1 \REGISTERS_reg[17][26]  ( .D(n4275), .CK(CLK), .RN(n407), .QN(n2612)
         );
  DFFR_X1 \REGISTERS_reg[17][25]  ( .D(n4274), .CK(CLK), .RN(n407), .QN(n2633)
         );
  DFFR_X1 \REGISTERS_reg[17][24]  ( .D(n4273), .CK(CLK), .RN(n407), .QN(n2654)
         );
  DFFR_X1 \REGISTERS_reg[17][23]  ( .D(n4272), .CK(CLK), .RN(n407), .QN(n2675)
         );
  DFFR_X1 \REGISTERS_reg[17][22]  ( .D(n4271), .CK(CLK), .RN(n407), .QN(n2696)
         );
  DFFR_X1 \REGISTERS_reg[17][21]  ( .D(n4270), .CK(CLK), .RN(n407), .QN(n2717)
         );
  DFFR_X1 \REGISTERS_reg[17][20]  ( .D(n4269), .CK(CLK), .RN(n407), .QN(n2738)
         );
  DFFR_X1 \REGISTERS_reg[17][19]  ( .D(n4268), .CK(CLK), .RN(n407), .QN(n2759)
         );
  DFFR_X1 \REGISTERS_reg[17][18]  ( .D(n4267), .CK(CLK), .RN(n407), .QN(n2780)
         );
  DFFR_X1 \REGISTERS_reg[17][17]  ( .D(n4266), .CK(CLK), .RN(n406), .QN(n2801)
         );
  DFFR_X1 \REGISTERS_reg[17][16]  ( .D(n4265), .CK(CLK), .RN(n406), .QN(n2822)
         );
  DFFR_X1 \REGISTERS_reg[17][15]  ( .D(n4264), .CK(CLK), .RN(n406), .QN(n2843)
         );
  DFFR_X1 \REGISTERS_reg[17][14]  ( .D(n4263), .CK(CLK), .RN(n406), .QN(n2864)
         );
  DFFR_X1 \REGISTERS_reg[17][13]  ( .D(n4262), .CK(CLK), .RN(n406), .QN(n2885)
         );
  DFFR_X1 \REGISTERS_reg[17][12]  ( .D(n4261), .CK(CLK), .RN(n406), .QN(n2906)
         );
  DFFR_X1 \REGISTERS_reg[17][11]  ( .D(n4260), .CK(CLK), .RN(n406), .QN(n2927)
         );
  DFFR_X1 \REGISTERS_reg[17][10]  ( .D(n4259), .CK(CLK), .RN(n406), .QN(n2948)
         );
  DFFR_X1 \REGISTERS_reg[17][9]  ( .D(n4258), .CK(CLK), .RN(n406), .QN(n2969)
         );
  DFFR_X1 \REGISTERS_reg[17][8]  ( .D(n4257), .CK(CLK), .RN(n406), .QN(n3566)
         );
  DFFR_X1 \REGISTERS_reg[17][7]  ( .D(n4256), .CK(CLK), .RN(n406), .QN(n3587)
         );
  DFFR_X1 \REGISTERS_reg[17][6]  ( .D(n4255), .CK(CLK), .RN(n406), .QN(n3608)
         );
  DFFR_X1 \REGISTERS_reg[17][5]  ( .D(n4254), .CK(CLK), .RN(n405), .QN(n3629)
         );
  DFFR_X1 \REGISTERS_reg[17][4]  ( .D(n4253), .CK(CLK), .RN(n405), .QN(n3650)
         );
  DFFR_X1 \REGISTERS_reg[17][3]  ( .D(n4252), .CK(CLK), .RN(n405), .QN(n3671)
         );
  DFFR_X1 \REGISTERS_reg[17][2]  ( .D(n4251), .CK(CLK), .RN(n405), .QN(n3692)
         );
  DFFR_X1 \REGISTERS_reg[17][1]  ( .D(n4250), .CK(CLK), .RN(n405), .QN(n3713)
         );
  DFFR_X1 \REGISTERS_reg[17][0]  ( .D(n4249), .CK(CLK), .RN(n405), .QN(n3734)
         );
  DFFR_X1 \REGISTERS_reg[18][31]  ( .D(n3302), .CK(CLK), .RN(n405), .Q(n2509)
         );
  DFFR_X1 \REGISTERS_reg[18][30]  ( .D(n3301), .CK(CLK), .RN(n405), .Q(n2530)
         );
  DFFR_X1 \REGISTERS_reg[18][29]  ( .D(n3300), .CK(CLK), .RN(n405), .Q(n2551)
         );
  DFFR_X1 \REGISTERS_reg[18][28]  ( .D(n3299), .CK(CLK), .RN(n405), .Q(n2572)
         );
  DFFR_X1 \REGISTERS_reg[18][27]  ( .D(n3298), .CK(CLK), .RN(n405), .Q(n2593)
         );
  DFFR_X1 \REGISTERS_reg[18][26]  ( .D(n3297), .CK(CLK), .RN(n405), .Q(n2614)
         );
  DFFR_X1 \REGISTERS_reg[18][25]  ( .D(n3296), .CK(CLK), .RN(n404), .Q(n2635)
         );
  DFFR_X1 \REGISTERS_reg[18][24]  ( .D(n3295), .CK(CLK), .RN(n404), .Q(n2656)
         );
  DFFR_X1 \REGISTERS_reg[18][23]  ( .D(n3294), .CK(CLK), .RN(n404), .Q(n2677)
         );
  DFFR_X1 \REGISTERS_reg[18][22]  ( .D(n3293), .CK(CLK), .RN(n404), .Q(n2698)
         );
  DFFR_X1 \REGISTERS_reg[18][21]  ( .D(n3292), .CK(CLK), .RN(n404), .Q(n2719)
         );
  DFFR_X1 \REGISTERS_reg[18][20]  ( .D(n3291), .CK(CLK), .RN(n404), .Q(n2740)
         );
  DFFR_X1 \REGISTERS_reg[18][19]  ( .D(n3290), .CK(CLK), .RN(n404), .Q(n2761)
         );
  DFFR_X1 \REGISTERS_reg[18][18]  ( .D(n3289), .CK(CLK), .RN(n404), .Q(n2782)
         );
  DFFR_X1 \REGISTERS_reg[18][17]  ( .D(n3288), .CK(CLK), .RN(n404), .Q(n2803)
         );
  DFFR_X1 \REGISTERS_reg[18][16]  ( .D(n3287), .CK(CLK), .RN(n404), .Q(n2824)
         );
  DFFR_X1 \REGISTERS_reg[18][15]  ( .D(n3286), .CK(CLK), .RN(n404), .Q(n2845)
         );
  DFFR_X1 \REGISTERS_reg[18][14]  ( .D(n3285), .CK(CLK), .RN(n403), .Q(n2866)
         );
  DFFR_X1 \REGISTERS_reg[18][13]  ( .D(n3284), .CK(CLK), .RN(n403), .Q(n2887)
         );
  DFFR_X1 \REGISTERS_reg[18][12]  ( .D(n3283), .CK(CLK), .RN(n403), .Q(n2908)
         );
  DFFR_X1 \REGISTERS_reg[18][11]  ( .D(n3282), .CK(CLK), .RN(n403), .Q(n2929)
         );
  DFFR_X1 \REGISTERS_reg[18][10]  ( .D(n3281), .CK(CLK), .RN(n403), .Q(n2950)
         );
  DFFR_X1 \REGISTERS_reg[18][9]  ( .D(n3280), .CK(CLK), .RN(n403), .Q(n2971)
         );
  DFFR_X1 \REGISTERS_reg[18][8]  ( .D(n3279), .CK(CLK), .RN(n403), .Q(n3568)
         );
  DFFR_X1 \REGISTERS_reg[18][7]  ( .D(n3278), .CK(CLK), .RN(n403), .Q(n3589)
         );
  DFFR_X1 \REGISTERS_reg[18][6]  ( .D(n3277), .CK(CLK), .RN(n403), .Q(n3610)
         );
  DFFR_X1 \REGISTERS_reg[18][5]  ( .D(n3276), .CK(CLK), .RN(n403), .Q(n3631)
         );
  DFFR_X1 \REGISTERS_reg[18][4]  ( .D(n3275), .CK(CLK), .RN(n403), .Q(n3652)
         );
  DFFR_X1 \REGISTERS_reg[18][3]  ( .D(n3274), .CK(CLK), .RN(n403), .Q(n3673)
         );
  DFFR_X1 \REGISTERS_reg[18][2]  ( .D(n3273), .CK(CLK), .RN(n402), .Q(n3694)
         );
  DFFR_X1 \REGISTERS_reg[18][1]  ( .D(n3272), .CK(CLK), .RN(n402), .Q(n3715)
         );
  DFFR_X1 \REGISTERS_reg[18][0]  ( .D(n3271), .CK(CLK), .RN(n402), .Q(n3736)
         );
  DFFR_X1 \REGISTERS_reg[19][31]  ( .D(n3270), .CK(CLK), .RN(n402), .Q(n2508)
         );
  DFFR_X1 \REGISTERS_reg[19][30]  ( .D(n3269), .CK(CLK), .RN(n402), .Q(n2529)
         );
  DFFR_X1 \REGISTERS_reg[19][29]  ( .D(n3268), .CK(CLK), .RN(n402), .Q(n2550)
         );
  DFFR_X1 \REGISTERS_reg[19][28]  ( .D(n3267), .CK(CLK), .RN(n402), .Q(n2571)
         );
  DFFR_X1 \REGISTERS_reg[19][27]  ( .D(n3266), .CK(CLK), .RN(n402), .Q(n2592)
         );
  DFFR_X1 \REGISTERS_reg[19][26]  ( .D(n3265), .CK(CLK), .RN(n402), .Q(n2613)
         );
  DFFR_X1 \REGISTERS_reg[19][25]  ( .D(n3264), .CK(CLK), .RN(n402), .Q(n2634)
         );
  DFFR_X1 \REGISTERS_reg[19][24]  ( .D(n3263), .CK(CLK), .RN(n402), .Q(n2655)
         );
  DFFR_X1 \REGISTERS_reg[19][23]  ( .D(n3262), .CK(CLK), .RN(n402), .Q(n2676)
         );
  DFFR_X1 \REGISTERS_reg[19][22]  ( .D(n3261), .CK(CLK), .RN(n401), .Q(n2697)
         );
  DFFR_X1 \REGISTERS_reg[19][21]  ( .D(n3260), .CK(CLK), .RN(n401), .Q(n2718)
         );
  DFFR_X1 \REGISTERS_reg[19][20]  ( .D(n3259), .CK(CLK), .RN(n401), .Q(n2739)
         );
  DFFR_X1 \REGISTERS_reg[19][19]  ( .D(n3258), .CK(CLK), .RN(n401), .Q(n2760)
         );
  DFFR_X1 \REGISTERS_reg[19][18]  ( .D(n3257), .CK(CLK), .RN(n401), .Q(n2781)
         );
  DFFR_X1 \REGISTERS_reg[19][17]  ( .D(n3256), .CK(CLK), .RN(n401), .Q(n2802)
         );
  DFFR_X1 \REGISTERS_reg[19][16]  ( .D(n3255), .CK(CLK), .RN(n401), .Q(n2823)
         );
  DFFR_X1 \REGISTERS_reg[19][15]  ( .D(n3254), .CK(CLK), .RN(n401), .Q(n2844)
         );
  DFFR_X1 \REGISTERS_reg[19][14]  ( .D(n3253), .CK(CLK), .RN(n401), .Q(n2865)
         );
  DFFR_X1 \REGISTERS_reg[19][13]  ( .D(n3252), .CK(CLK), .RN(n401), .Q(n2886)
         );
  DFFR_X1 \REGISTERS_reg[19][12]  ( .D(n3251), .CK(CLK), .RN(n401), .Q(n2907)
         );
  DFFR_X1 \REGISTERS_reg[19][11]  ( .D(n3250), .CK(CLK), .RN(n401), .Q(n2928)
         );
  DFFR_X1 \REGISTERS_reg[19][10]  ( .D(n3249), .CK(CLK), .RN(n400), .Q(n2949)
         );
  DFFR_X1 \REGISTERS_reg[19][9]  ( .D(n3248), .CK(CLK), .RN(n400), .Q(n2970)
         );
  DFFR_X1 \REGISTERS_reg[19][8]  ( .D(n3247), .CK(CLK), .RN(n400), .Q(n3567)
         );
  DFFR_X1 \REGISTERS_reg[19][7]  ( .D(n3246), .CK(CLK), .RN(n400), .Q(n3588)
         );
  DFFR_X1 \REGISTERS_reg[19][6]  ( .D(n3245), .CK(CLK), .RN(n400), .Q(n3609)
         );
  DFFR_X1 \REGISTERS_reg[19][5]  ( .D(n3244), .CK(CLK), .RN(n400), .Q(n3630)
         );
  DFFR_X1 \REGISTERS_reg[19][4]  ( .D(n3243), .CK(CLK), .RN(n400), .Q(n3651)
         );
  DFFR_X1 \REGISTERS_reg[19][3]  ( .D(n3242), .CK(CLK), .RN(n400), .Q(n3672)
         );
  DFFR_X1 \REGISTERS_reg[19][2]  ( .D(n3241), .CK(CLK), .RN(n400), .Q(n3693)
         );
  DFFR_X1 \REGISTERS_reg[19][1]  ( .D(n3240), .CK(CLK), .RN(n400), .Q(n3714)
         );
  DFFR_X1 \REGISTERS_reg[19][0]  ( .D(n3239), .CK(CLK), .RN(n400), .Q(n3735)
         );
  DFFR_X1 \REGISTERS_reg[20][31]  ( .D(n4312), .CK(CLK), .RN(n400), .QN(n2504)
         );
  DFFR_X1 \REGISTERS_reg[20][30]  ( .D(n4311), .CK(CLK), .RN(n399), .QN(n2525)
         );
  DFFR_X1 \REGISTERS_reg[20][29]  ( .D(n4310), .CK(CLK), .RN(n399), .QN(n2546)
         );
  DFFR_X1 \REGISTERS_reg[20][28]  ( .D(n4309), .CK(CLK), .RN(n399), .QN(n2567)
         );
  DFFR_X1 \REGISTERS_reg[20][27]  ( .D(n4308), .CK(CLK), .RN(n399), .QN(n2588)
         );
  DFFR_X1 \REGISTERS_reg[20][26]  ( .D(n4307), .CK(CLK), .RN(n399), .QN(n2609)
         );
  DFFR_X1 \REGISTERS_reg[20][25]  ( .D(n4306), .CK(CLK), .RN(n399), .QN(n2630)
         );
  DFFR_X1 \REGISTERS_reg[20][24]  ( .D(n4305), .CK(CLK), .RN(n399), .QN(n2651)
         );
  DFFR_X1 \REGISTERS_reg[20][23]  ( .D(n4304), .CK(CLK), .RN(n399), .QN(n2672)
         );
  DFFR_X1 \REGISTERS_reg[20][22]  ( .D(n4303), .CK(CLK), .RN(n399), .QN(n2693)
         );
  DFFR_X1 \REGISTERS_reg[20][21]  ( .D(n4302), .CK(CLK), .RN(n399), .QN(n2714)
         );
  DFFR_X1 \REGISTERS_reg[20][20]  ( .D(n4301), .CK(CLK), .RN(n399), .QN(n2735)
         );
  DFFR_X1 \REGISTERS_reg[20][19]  ( .D(n4300), .CK(CLK), .RN(n404), .QN(n2756)
         );
  DFFR_X1 \REGISTERS_reg[20][18]  ( .D(n4299), .CK(CLK), .RN(n419), .QN(n2777)
         );
  DFFR_X1 \REGISTERS_reg[20][17]  ( .D(n4298), .CK(CLK), .RN(n419), .QN(n2798)
         );
  DFFR_X1 \REGISTERS_reg[20][16]  ( .D(n4297), .CK(CLK), .RN(n419), .QN(n2819)
         );
  DFFR_X1 \REGISTERS_reg[20][15]  ( .D(n4296), .CK(CLK), .RN(n419), .QN(n2840)
         );
  DFFR_X1 \REGISTERS_reg[20][14]  ( .D(n4295), .CK(CLK), .RN(n419), .QN(n2861)
         );
  DFFR_X1 \REGISTERS_reg[20][13]  ( .D(n4294), .CK(CLK), .RN(n419), .QN(n2882)
         );
  DFFR_X1 \REGISTERS_reg[20][12]  ( .D(n4293), .CK(CLK), .RN(n419), .QN(n2903)
         );
  DFFR_X1 \REGISTERS_reg[20][11]  ( .D(n4292), .CK(CLK), .RN(n419), .QN(n2924)
         );
  DFFR_X1 \REGISTERS_reg[20][10]  ( .D(n4291), .CK(CLK), .RN(n418), .QN(n2945)
         );
  DFFR_X1 \REGISTERS_reg[20][9]  ( .D(n4290), .CK(CLK), .RN(n418), .QN(n2966)
         );
  DFFR_X1 \REGISTERS_reg[20][8]  ( .D(n4289), .CK(CLK), .RN(n418), .QN(n3563)
         );
  DFFR_X1 \REGISTERS_reg[20][7]  ( .D(n4288), .CK(CLK), .RN(n418), .QN(n3584)
         );
  DFFR_X1 \REGISTERS_reg[20][6]  ( .D(n4287), .CK(CLK), .RN(n418), .QN(n3605)
         );
  DFFR_X1 \REGISTERS_reg[20][5]  ( .D(n4286), .CK(CLK), .RN(n418), .QN(n3626)
         );
  DFFR_X1 \REGISTERS_reg[20][4]  ( .D(n4285), .CK(CLK), .RN(n418), .QN(n3647)
         );
  DFFR_X1 \REGISTERS_reg[20][3]  ( .D(n4284), .CK(CLK), .RN(n418), .QN(n3668)
         );
  DFFR_X1 \REGISTERS_reg[20][2]  ( .D(n4283), .CK(CLK), .RN(n418), .QN(n3689)
         );
  DFFR_X1 \REGISTERS_reg[20][1]  ( .D(n4282), .CK(CLK), .RN(n418), .QN(n3710)
         );
  DFFR_X1 \REGISTERS_reg[20][0]  ( .D(n4281), .CK(CLK), .RN(n418), .QN(n3731)
         );
  DFFR_X1 \REGISTERS_reg[21][31]  ( .D(n4344), .CK(CLK), .RN(n418), .Q(n940)
         );
  DFFR_X1 \REGISTERS_reg[21][30]  ( .D(n4343), .CK(CLK), .RN(n417), .Q(n939)
         );
  DFFR_X1 \REGISTERS_reg[21][29]  ( .D(n4342), .CK(CLK), .RN(n417), .Q(n938)
         );
  DFFR_X1 \REGISTERS_reg[21][28]  ( .D(n4341), .CK(CLK), .RN(n417), .Q(n937)
         );
  DFFR_X1 \REGISTERS_reg[21][27]  ( .D(n4340), .CK(CLK), .RN(n417), .Q(n936)
         );
  DFFR_X1 \REGISTERS_reg[21][26]  ( .D(n4339), .CK(CLK), .RN(n417), .Q(n935)
         );
  DFFR_X1 \REGISTERS_reg[21][25]  ( .D(n4338), .CK(CLK), .RN(n417), .Q(n934)
         );
  DFFR_X1 \REGISTERS_reg[21][24]  ( .D(n4337), .CK(CLK), .RN(n417), .Q(n933)
         );
  DFFR_X1 \REGISTERS_reg[21][23]  ( .D(n4336), .CK(CLK), .RN(n417), .Q(n932)
         );
  DFFR_X1 \REGISTERS_reg[21][22]  ( .D(n4335), .CK(CLK), .RN(n417), .Q(n931)
         );
  DFFR_X1 \REGISTERS_reg[21][21]  ( .D(n4334), .CK(CLK), .RN(n417), .Q(n930)
         );
  DFFR_X1 \REGISTERS_reg[21][20]  ( .D(n4333), .CK(CLK), .RN(n417), .Q(n929)
         );
  DFFR_X1 \REGISTERS_reg[21][19]  ( .D(n4332), .CK(CLK), .RN(n417), .Q(n928)
         );
  DFFR_X1 \REGISTERS_reg[21][18]  ( .D(n4331), .CK(CLK), .RN(n416), .Q(n927)
         );
  DFFR_X1 \REGISTERS_reg[21][17]  ( .D(n4330), .CK(CLK), .RN(n416), .Q(n926)
         );
  DFFR_X1 \REGISTERS_reg[21][16]  ( .D(n4329), .CK(CLK), .RN(n416), .Q(n925)
         );
  DFFR_X1 \REGISTERS_reg[21][15]  ( .D(n4328), .CK(CLK), .RN(n416), .Q(n924)
         );
  DFFR_X1 \REGISTERS_reg[21][14]  ( .D(n4327), .CK(CLK), .RN(n416), .Q(n923)
         );
  DFFR_X1 \REGISTERS_reg[21][13]  ( .D(n4326), .CK(CLK), .RN(n416), .Q(n922)
         );
  DFFR_X1 \REGISTERS_reg[21][12]  ( .D(n4325), .CK(CLK), .RN(n416), .Q(n921)
         );
  DFFR_X1 \REGISTERS_reg[21][11]  ( .D(n4324), .CK(CLK), .RN(n416), .Q(n920)
         );
  DFFR_X1 \REGISTERS_reg[21][10]  ( .D(n4323), .CK(CLK), .RN(n416), .Q(n919)
         );
  DFFR_X1 \REGISTERS_reg[21][9]  ( .D(n4322), .CK(CLK), .RN(n416), .Q(n918) );
  DFFR_X1 \REGISTERS_reg[21][8]  ( .D(n4321), .CK(CLK), .RN(n416), .Q(n917) );
  DFFR_X1 \REGISTERS_reg[21][7]  ( .D(n4320), .CK(CLK), .RN(n416), .Q(n916) );
  DFFR_X1 \REGISTERS_reg[21][6]  ( .D(n4319), .CK(CLK), .RN(n415), .Q(n915) );
  DFFR_X1 \REGISTERS_reg[21][5]  ( .D(n4318), .CK(CLK), .RN(n415), .Q(n914) );
  DFFR_X1 \REGISTERS_reg[21][4]  ( .D(n4317), .CK(CLK), .RN(n415), .Q(n913) );
  DFFR_X1 \REGISTERS_reg[21][3]  ( .D(n4316), .CK(CLK), .RN(n415), .Q(n912) );
  DFFR_X1 \REGISTERS_reg[21][2]  ( .D(n4315), .CK(CLK), .RN(n415), .Q(n911) );
  DFFR_X1 \REGISTERS_reg[21][1]  ( .D(n4314), .CK(CLK), .RN(n415), .Q(n910) );
  DFFR_X1 \REGISTERS_reg[21][0]  ( .D(n4313), .CK(CLK), .RN(n415), .Q(n908) );
  DFFR_X1 \REGISTERS_reg[24][31]  ( .D(n3174), .CK(CLK), .RN(n409), .Q(n2503)
         );
  DFFR_X1 \REGISTERS_reg[24][30]  ( .D(n3173), .CK(CLK), .RN(n409), .Q(n2524)
         );
  DFFR_X1 \REGISTERS_reg[24][29]  ( .D(n3172), .CK(CLK), .RN(n409), .Q(n2545)
         );
  DFFR_X1 \REGISTERS_reg[24][28]  ( .D(n3171), .CK(CLK), .RN(n409), .Q(n2566)
         );
  DFFR_X1 \REGISTERS_reg[24][27]  ( .D(n3170), .CK(CLK), .RN(n409), .Q(n2587)
         );
  DFFR_X1 \REGISTERS_reg[24][26]  ( .D(n3169), .CK(CLK), .RN(n409), .Q(n2608)
         );
  DFFR_X1 \REGISTERS_reg[24][25]  ( .D(n3168), .CK(CLK), .RN(n409), .Q(n2629)
         );
  DFFR_X1 \REGISTERS_reg[24][24]  ( .D(n3167), .CK(CLK), .RN(n414), .Q(n2650)
         );
  DFFR_X1 \REGISTERS_reg[24][23]  ( .D(n3166), .CK(CLK), .RN(n388), .Q(n2671)
         );
  DFFR_X1 \REGISTERS_reg[24][22]  ( .D(n3165), .CK(CLK), .RN(n388), .Q(n2692)
         );
  DFFR_X1 \REGISTERS_reg[24][21]  ( .D(n3164), .CK(CLK), .RN(n388), .Q(n2713)
         );
  DFFR_X1 \REGISTERS_reg[24][20]  ( .D(n3163), .CK(CLK), .RN(n388), .Q(n2734)
         );
  DFFR_X1 \REGISTERS_reg[24][19]  ( .D(n3162), .CK(CLK), .RN(n388), .Q(n2755)
         );
  DFFR_X1 \REGISTERS_reg[24][18]  ( .D(n3161), .CK(CLK), .RN(n388), .Q(n2776)
         );
  DFFR_X1 \REGISTERS_reg[24][17]  ( .D(n3160), .CK(CLK), .RN(n388), .Q(n2797)
         );
  DFFR_X1 \REGISTERS_reg[24][16]  ( .D(n3159), .CK(CLK), .RN(n388), .Q(n2818)
         );
  DFFR_X1 \REGISTERS_reg[24][15]  ( .D(n3158), .CK(CLK), .RN(n388), .Q(n2839)
         );
  DFFR_X1 \REGISTERS_reg[24][14]  ( .D(n3157), .CK(CLK), .RN(n387), .Q(n2860)
         );
  DFFR_X1 \REGISTERS_reg[24][13]  ( .D(n3156), .CK(CLK), .RN(n387), .Q(n2881)
         );
  DFFR_X1 \REGISTERS_reg[24][12]  ( .D(n3155), .CK(CLK), .RN(n387), .Q(n2902)
         );
  DFFR_X1 \REGISTERS_reg[24][11]  ( .D(n3154), .CK(CLK), .RN(n387), .Q(n2923)
         );
  DFFR_X1 \REGISTERS_reg[24][10]  ( .D(n3153), .CK(CLK), .RN(n387), .Q(n2944)
         );
  DFFR_X1 \REGISTERS_reg[24][9]  ( .D(n3152), .CK(CLK), .RN(n387), .Q(n2965)
         );
  DFFR_X1 \REGISTERS_reg[24][8]  ( .D(n3151), .CK(CLK), .RN(n387), .Q(n3562)
         );
  DFFR_X1 \REGISTERS_reg[24][7]  ( .D(n3150), .CK(CLK), .RN(n387), .Q(n3583)
         );
  DFFR_X1 \REGISTERS_reg[24][6]  ( .D(n3149), .CK(CLK), .RN(n387), .Q(n3604)
         );
  DFFR_X1 \REGISTERS_reg[24][5]  ( .D(n3148), .CK(CLK), .RN(n387), .Q(n3625)
         );
  DFFR_X1 \REGISTERS_reg[24][4]  ( .D(n3147), .CK(CLK), .RN(n387), .Q(n3646)
         );
  DFFR_X1 \REGISTERS_reg[24][3]  ( .D(n3146), .CK(CLK), .RN(n387), .Q(n3667)
         );
  DFFR_X1 \REGISTERS_reg[24][2]  ( .D(n3145), .CK(CLK), .RN(n386), .Q(n3688)
         );
  DFFR_X1 \REGISTERS_reg[24][1]  ( .D(n3144), .CK(CLK), .RN(n386), .Q(n3709)
         );
  DFFR_X1 \REGISTERS_reg[24][0]  ( .D(n3143), .CK(CLK), .RN(n386), .Q(n3730)
         );
  DFFR_X1 \REGISTERS_reg[25][3]  ( .D(n3114), .CK(CLK), .RN(n384), .Q(n3666)
         );
  DFFR_X1 \REGISTERS_reg[25][2]  ( .D(n3113), .CK(CLK), .RN(n384), .Q(n3687)
         );
  DFFR_X1 \REGISTERS_reg[25][1]  ( .D(n3112), .CK(CLK), .RN(n384), .Q(n3708)
         );
  DFFR_X1 \REGISTERS_reg[25][0]  ( .D(n3111), .CK(CLK), .RN(n384), .Q(n3729)
         );
  DFFR_X1 \REGISTERS_reg[26][31]  ( .D(n4089), .CK(CLK), .RN(n384), .Q(n671)
         );
  DFFR_X1 \REGISTERS_reg[26][30]  ( .D(n4120), .CK(CLK), .RN(n383), .Q(n703)
         );
  DFFR_X1 \REGISTERS_reg[26][29]  ( .D(n4119), .CK(CLK), .RN(n383), .Q(n702)
         );
  DFFR_X1 \REGISTERS_reg[26][28]  ( .D(n4118), .CK(CLK), .RN(n383), .Q(n701)
         );
  DFFR_X1 \REGISTERS_reg[26][27]  ( .D(n4117), .CK(CLK), .RN(n383), .Q(n700)
         );
  DFFR_X1 \REGISTERS_reg[26][26]  ( .D(n4116), .CK(CLK), .RN(n383), .Q(n699)
         );
  DFFR_X1 \REGISTERS_reg[26][25]  ( .D(n4115), .CK(CLK), .RN(n383), .Q(n698)
         );
  DFFR_X1 \REGISTERS_reg[26][24]  ( .D(n4114), .CK(CLK), .RN(n383), .Q(n697)
         );
  DFFR_X1 \REGISTERS_reg[26][23]  ( .D(n4113), .CK(CLK), .RN(n383), .Q(n696)
         );
  DFFR_X1 \REGISTERS_reg[26][22]  ( .D(n4112), .CK(CLK), .RN(n383), .Q(n695)
         );
  DFFR_X1 \REGISTERS_reg[26][21]  ( .D(n4111), .CK(CLK), .RN(n383), .Q(n694)
         );
  DFFR_X1 \REGISTERS_reg[26][20]  ( .D(n4110), .CK(CLK), .RN(n383), .Q(n693)
         );
  DFFR_X1 \REGISTERS_reg[26][19]  ( .D(n4109), .CK(CLK), .RN(n382), .Q(n692)
         );
  DFFR_X1 \REGISTERS_reg[26][18]  ( .D(n4108), .CK(CLK), .RN(n382), .Q(n691)
         );
  DFFR_X1 \REGISTERS_reg[26][17]  ( .D(n4107), .CK(CLK), .RN(n382), .Q(n690)
         );
  DFFR_X1 \REGISTERS_reg[26][16]  ( .D(n4106), .CK(CLK), .RN(n382), .Q(n689)
         );
  DFFR_X1 \REGISTERS_reg[26][15]  ( .D(n4105), .CK(CLK), .RN(n382), .Q(n688)
         );
  DFFR_X1 \REGISTERS_reg[26][14]  ( .D(n4104), .CK(CLK), .RN(n382), .Q(n687)
         );
  DFFR_X1 \REGISTERS_reg[26][13]  ( .D(n4103), .CK(CLK), .RN(n382), .Q(n686)
         );
  DFFR_X1 \REGISTERS_reg[26][12]  ( .D(n4102), .CK(CLK), .RN(n382), .Q(n685)
         );
  DFFR_X1 \REGISTERS_reg[26][11]  ( .D(n4101), .CK(CLK), .RN(n382), .Q(n684)
         );
  DFFR_X1 \REGISTERS_reg[26][10]  ( .D(n4100), .CK(CLK), .RN(n382), .Q(n683)
         );
  DFFR_X1 \REGISTERS_reg[26][9]  ( .D(n4099), .CK(CLK), .RN(n382), .Q(n682) );
  DFFR_X1 \REGISTERS_reg[26][8]  ( .D(n4098), .CK(CLK), .RN(n382), .Q(n681) );
  DFFR_X1 \REGISTERS_reg[26][7]  ( .D(n4097), .CK(CLK), .RN(n381), .Q(n680) );
  DFFR_X1 \REGISTERS_reg[26][6]  ( .D(n4096), .CK(CLK), .RN(n381), .Q(n679) );
  DFFR_X1 \REGISTERS_reg[26][5]  ( .D(n4095), .CK(CLK), .RN(n381), .Q(n678) );
  DFFR_X1 \REGISTERS_reg[26][4]  ( .D(n4094), .CK(CLK), .RN(n381), .Q(n677) );
  DFFR_X1 \REGISTERS_reg[26][3]  ( .D(n4093), .CK(CLK), .RN(n381), .Q(n676) );
  DFFR_X1 \REGISTERS_reg[26][2]  ( .D(n4092), .CK(CLK), .RN(n381), .Q(n675) );
  DFFR_X1 \REGISTERS_reg[26][1]  ( .D(n4091), .CK(CLK), .RN(n381), .Q(n674) );
  DFFR_X1 \REGISTERS_reg[26][0]  ( .D(n4090), .CK(CLK), .RN(n381), .Q(n673) );
  DFFR_X1 \REGISTERS_reg[27][31]  ( .D(n4152), .CK(CLK), .RN(n381), .QN(n3864)
         );
  DFFR_X1 \REGISTERS_reg[27][30]  ( .D(n4151), .CK(CLK), .RN(n381), .QN(n3863)
         );
  DFFR_X1 \REGISTERS_reg[27][29]  ( .D(n4150), .CK(CLK), .RN(n381), .QN(n3862)
         );
  DFFR_X1 \REGISTERS_reg[27][28]  ( .D(n4149), .CK(CLK), .RN(n381), .QN(n3861)
         );
  DFFR_X1 \REGISTERS_reg[27][27]  ( .D(n4148), .CK(CLK), .RN(n380), .QN(n3860)
         );
  DFFR_X1 \REGISTERS_reg[27][26]  ( .D(n4147), .CK(CLK), .RN(n380), .QN(n3859)
         );
  DFFR_X1 \REGISTERS_reg[27][25]  ( .D(n4146), .CK(CLK), .RN(n380), .QN(n3858)
         );
  DFFR_X1 \REGISTERS_reg[27][24]  ( .D(n4145), .CK(CLK), .RN(n380), .QN(n3857)
         );
  DFFR_X1 \REGISTERS_reg[27][23]  ( .D(n4144), .CK(CLK), .RN(n380), .QN(n3856)
         );
  DFFR_X1 \REGISTERS_reg[27][22]  ( .D(n4143), .CK(CLK), .RN(n380), .QN(n3855)
         );
  DFFR_X1 \REGISTERS_reg[27][21]  ( .D(n4142), .CK(CLK), .RN(n380), .QN(n3854)
         );
  DFFR_X1 \REGISTERS_reg[27][20]  ( .D(n4141), .CK(CLK), .RN(n380), .QN(n3853)
         );
  DFFR_X1 \REGISTERS_reg[27][19]  ( .D(n4140), .CK(CLK), .RN(n380), .QN(n3852)
         );
  DFFR_X1 \REGISTERS_reg[27][18]  ( .D(n4139), .CK(CLK), .RN(n380), .QN(n3851)
         );
  DFFR_X1 \REGISTERS_reg[27][17]  ( .D(n4138), .CK(CLK), .RN(n380), .QN(n3850)
         );
  DFFR_X1 \REGISTERS_reg[27][16]  ( .D(n4137), .CK(CLK), .RN(n380), .QN(n3849)
         );
  DFFR_X1 \REGISTERS_reg[27][15]  ( .D(n4136), .CK(CLK), .RN(n379), .QN(n3848)
         );
  DFFR_X1 \REGISTERS_reg[27][14]  ( .D(n4135), .CK(CLK), .RN(n379), .QN(n3847)
         );
  DFFR_X1 \REGISTERS_reg[27][13]  ( .D(n4134), .CK(CLK), .RN(n379), .QN(n3846)
         );
  DFFR_X1 \REGISTERS_reg[27][12]  ( .D(n4133), .CK(CLK), .RN(n379), .QN(n3845)
         );
  DFFR_X1 \REGISTERS_reg[27][11]  ( .D(n4132), .CK(CLK), .RN(n379), .QN(n3844)
         );
  DFFR_X1 \REGISTERS_reg[27][10]  ( .D(n4131), .CK(CLK), .RN(n379), .QN(n3843)
         );
  DFFR_X1 \REGISTERS_reg[27][9]  ( .D(n4130), .CK(CLK), .RN(n379), .QN(n3842)
         );
  DFFR_X1 \REGISTERS_reg[27][8]  ( .D(n4129), .CK(CLK), .RN(n379), .QN(n3841)
         );
  DFFR_X1 \REGISTERS_reg[27][7]  ( .D(n4128), .CK(CLK), .RN(n379), .QN(n3840)
         );
  DFFR_X1 \REGISTERS_reg[27][6]  ( .D(n4127), .CK(CLK), .RN(n379), .QN(n3839)
         );
  DFFR_X1 \REGISTERS_reg[27][5]  ( .D(n4126), .CK(CLK), .RN(n379), .QN(n3838)
         );
  DFFR_X1 \REGISTERS_reg[27][4]  ( .D(n4125), .CK(CLK), .RN(n379), .QN(n3837)
         );
  DFFR_X1 \REGISTERS_reg[27][3]  ( .D(n4124), .CK(CLK), .RN(n378), .QN(n3836)
         );
  DFFR_X1 \REGISTERS_reg[27][2]  ( .D(n4123), .CK(CLK), .RN(n378), .QN(n3835)
         );
  DFFR_X1 \REGISTERS_reg[27][1]  ( .D(n4122), .CK(CLK), .RN(n378), .QN(n3834)
         );
  DFFR_X1 \REGISTERS_reg[27][0]  ( .D(n4121), .CK(CLK), .RN(n378), .QN(n3833)
         );
  DFFR_X1 \REGISTERS_reg[29][31]  ( .D(n3078), .CK(CLK), .RN(n396), .Q(n3800)
         );
  DFFR_X1 \REGISTERS_reg[29][30]  ( .D(n3077), .CK(CLK), .RN(n396), .Q(n3799)
         );
  DFFR_X1 \REGISTERS_reg[29][29]  ( .D(n3076), .CK(CLK), .RN(n396), .Q(n3798)
         );
  DFFR_X1 \REGISTERS_reg[29][28]  ( .D(n3075), .CK(CLK), .RN(n396), .Q(n3797)
         );
  DFFR_X1 \REGISTERS_reg[29][27]  ( .D(n3074), .CK(CLK), .RN(n396), .Q(n3796)
         );
  DFFR_X1 \REGISTERS_reg[29][26]  ( .D(n3073), .CK(CLK), .RN(n396), .Q(n3795)
         );
  DFFR_X1 \REGISTERS_reg[29][25]  ( .D(n3072), .CK(CLK), .RN(n396), .Q(n3794)
         );
  DFFR_X1 \REGISTERS_reg[29][24]  ( .D(n3071), .CK(CLK), .RN(n396), .Q(n3793)
         );
  DFFR_X1 \REGISTERS_reg[29][23]  ( .D(n3070), .CK(CLK), .RN(n396), .Q(n3792)
         );
  DFFR_X1 \REGISTERS_reg[29][22]  ( .D(n3069), .CK(CLK), .RN(n395), .Q(n3791)
         );
  DFFR_X1 \REGISTERS_reg[29][21]  ( .D(n3068), .CK(CLK), .RN(n395), .Q(n3790)
         );
  DFFR_X1 \REGISTERS_reg[29][20]  ( .D(n3067), .CK(CLK), .RN(n395), .Q(n3789)
         );
  DFFR_X1 \REGISTERS_reg[29][19]  ( .D(n3066), .CK(CLK), .RN(n395), .Q(n3788)
         );
  DFFR_X1 \REGISTERS_reg[29][18]  ( .D(n3065), .CK(CLK), .RN(n395), .Q(n3787)
         );
  DFFR_X1 \REGISTERS_reg[29][17]  ( .D(n3064), .CK(CLK), .RN(n395), .Q(n3786)
         );
  DFFR_X1 \REGISTERS_reg[29][16]  ( .D(n3063), .CK(CLK), .RN(n395), .Q(n3785)
         );
  DFFR_X1 \REGISTERS_reg[29][15]  ( .D(n3062), .CK(CLK), .RN(n395), .Q(n3784)
         );
  DFFR_X1 \REGISTERS_reg[29][14]  ( .D(n3061), .CK(CLK), .RN(n395), .Q(n3783)
         );
  DFFR_X1 \REGISTERS_reg[29][13]  ( .D(n3060), .CK(CLK), .RN(n395), .Q(n3782)
         );
  DFFR_X1 \REGISTERS_reg[29][12]  ( .D(n3059), .CK(CLK), .RN(n395), .Q(n3781)
         );
  DFFR_X1 \REGISTERS_reg[29][11]  ( .D(n3058), .CK(CLK), .RN(n395), .Q(n3780)
         );
  DFFR_X1 \REGISTERS_reg[29][10]  ( .D(n3057), .CK(CLK), .RN(n394), .Q(n3779)
         );
  DFFR_X1 \REGISTERS_reg[29][9]  ( .D(n3056), .CK(CLK), .RN(n394), .Q(n3778)
         );
  DFFR_X1 \REGISTERS_reg[29][8]  ( .D(n3055), .CK(CLK), .RN(n394), .Q(n3777)
         );
  DFFR_X1 \REGISTERS_reg[29][7]  ( .D(n3054), .CK(CLK), .RN(n394), .Q(n3776)
         );
  DFFR_X1 \REGISTERS_reg[29][6]  ( .D(n3053), .CK(CLK), .RN(n394), .Q(n3775)
         );
  DFFR_X1 \REGISTERS_reg[29][5]  ( .D(n3052), .CK(CLK), .RN(n394), .Q(n3774)
         );
  DFFR_X1 \REGISTERS_reg[29][4]  ( .D(n3051), .CK(CLK), .RN(n394), .Q(n3773)
         );
  DFFR_X1 \REGISTERS_reg[29][3]  ( .D(n3050), .CK(CLK), .RN(n394), .Q(n3772)
         );
  DFFR_X1 \REGISTERS_reg[29][2]  ( .D(n3049), .CK(CLK), .RN(n394), .Q(n3771)
         );
  DFFR_X1 \REGISTERS_reg[29][1]  ( .D(n3048), .CK(CLK), .RN(n394), .Q(n3770)
         );
  DFFR_X1 \REGISTERS_reg[29][0]  ( .D(n3047), .CK(CLK), .RN(n394), .Q(n3769)
         );
  DFFR_X1 \REGISTERS_reg[30][31]  ( .D(n4184), .CK(CLK), .RN(n394), .QN(n3768)
         );
  DFFR_X1 \REGISTERS_reg[30][30]  ( .D(n4183), .CK(CLK), .RN(n393), .QN(n3767)
         );
  DFFR_X1 \REGISTERS_reg[30][29]  ( .D(n4182), .CK(CLK), .RN(n393), .QN(n3766)
         );
  DFFR_X1 \REGISTERS_reg[30][28]  ( .D(n4181), .CK(CLK), .RN(n393), .QN(n3765)
         );
  DFFR_X1 \REGISTERS_reg[30][27]  ( .D(n4180), .CK(CLK), .RN(n393), .QN(n3764)
         );
  DFFR_X1 \REGISTERS_reg[30][26]  ( .D(n4179), .CK(CLK), .RN(n393), .QN(n3763)
         );
  DFFR_X1 \REGISTERS_reg[30][25]  ( .D(n4178), .CK(CLK), .RN(n393), .QN(n3762)
         );
  DFFR_X1 \REGISTERS_reg[30][24]  ( .D(n4177), .CK(CLK), .RN(n393), .QN(n3761)
         );
  DFFR_X1 \REGISTERS_reg[30][23]  ( .D(n4176), .CK(CLK), .RN(n393), .QN(n3760)
         );
  DFFR_X1 \REGISTERS_reg[30][22]  ( .D(n4175), .CK(CLK), .RN(n393), .QN(n3759)
         );
  DFFR_X1 \REGISTERS_reg[30][21]  ( .D(n4174), .CK(CLK), .RN(n393), .QN(n3758)
         );
  DFFR_X1 \REGISTERS_reg[30][20]  ( .D(n4173), .CK(CLK), .RN(n393), .QN(n3757)
         );
  DFFR_X1 \REGISTERS_reg[30][19]  ( .D(n4172), .CK(CLK), .RN(n392), .QN(n3756)
         );
  DFFR_X1 \REGISTERS_reg[30][18]  ( .D(n4171), .CK(CLK), .RN(n392), .QN(n3755)
         );
  DFFR_X1 \REGISTERS_reg[30][17]  ( .D(n4170), .CK(CLK), .RN(n392), .QN(n3754)
         );
  DFFR_X1 \REGISTERS_reg[30][16]  ( .D(n4169), .CK(CLK), .RN(n392), .QN(n3753)
         );
  DFFR_X1 \REGISTERS_reg[30][15]  ( .D(n4168), .CK(CLK), .RN(n392), .QN(n3752)
         );
  DFFR_X1 \REGISTERS_reg[30][14]  ( .D(n4167), .CK(CLK), .RN(n392), .QN(n3751)
         );
  DFFR_X1 \REGISTERS_reg[30][13]  ( .D(n4166), .CK(CLK), .RN(n392), .QN(n3750)
         );
  DFFR_X1 \REGISTERS_reg[30][12]  ( .D(n4165), .CK(CLK), .RN(n392), .QN(n3749)
         );
  DFFR_X1 \REGISTERS_reg[30][11]  ( .D(n4164), .CK(CLK), .RN(n392), .QN(n3748)
         );
  DFFR_X1 \REGISTERS_reg[30][10]  ( .D(n4163), .CK(CLK), .RN(n392), .QN(n3747)
         );
  DFFR_X1 \REGISTERS_reg[30][9]  ( .D(n4162), .CK(CLK), .RN(n392), .QN(n3746)
         );
  DFFR_X1 \REGISTERS_reg[30][8]  ( .D(n4161), .CK(CLK), .RN(n392), .QN(n3745)
         );
  DFFR_X1 \REGISTERS_reg[30][7]  ( .D(n4160), .CK(CLK), .RN(n391), .QN(n3744)
         );
  DFFR_X1 \REGISTERS_reg[30][6]  ( .D(n4159), .CK(CLK), .RN(n391), .QN(n3743)
         );
  DFFR_X1 \REGISTERS_reg[30][5]  ( .D(n4158), .CK(CLK), .RN(n391), .QN(n3742)
         );
  DFFR_X1 \REGISTERS_reg[30][4]  ( .D(n4157), .CK(CLK), .RN(n391), .QN(n3741)
         );
  DFFR_X1 \REGISTERS_reg[30][3]  ( .D(n4156), .CK(CLK), .RN(n391), .QN(n3740)
         );
  DFFR_X1 \REGISTERS_reg[30][2]  ( .D(n4155), .CK(CLK), .RN(n391), .QN(n3739)
         );
  DFFR_X1 \REGISTERS_reg[30][1]  ( .D(n4154), .CK(CLK), .RN(n391), .QN(n3738)
         );
  DFFR_X1 \REGISTERS_reg[30][0]  ( .D(n4153), .CK(CLK), .RN(n391), .QN(n3737)
         );
  DFFR_X1 \REGISTERS_reg[31][31]  ( .D(n4216), .CK(CLK), .RN(n391), .Q(n806)
         );
  DFF_X1 \OUT2_reg[31]  ( .D(n3015), .CK(CLK), .Q(OUT2[31]), .QN(n2489) );
  DFFR_X1 \REGISTERS_reg[31][30]  ( .D(n4215), .CK(CLK), .RN(n391), .Q(n805)
         );
  DFF_X1 \OUT2_reg[30]  ( .D(n3016), .CK(CLK), .Q(OUT2[30]), .QN(n2510) );
  DFFR_X1 \REGISTERS_reg[31][29]  ( .D(n4214), .CK(CLK), .RN(n391), .Q(n804)
         );
  DFF_X1 \OUT2_reg[29]  ( .D(n3017), .CK(CLK), .Q(OUT2[29]), .QN(n2531) );
  DFFR_X1 \REGISTERS_reg[31][28]  ( .D(n4213), .CK(CLK), .RN(n391), .Q(n803)
         );
  DFF_X1 \OUT2_reg[28]  ( .D(n3018), .CK(CLK), .Q(OUT2[28]), .QN(n2552) );
  DFFR_X1 \REGISTERS_reg[31][27]  ( .D(n4212), .CK(CLK), .RN(n390), .Q(n802)
         );
  DFF_X1 \OUT2_reg[27]  ( .D(n3019), .CK(CLK), .Q(OUT2[27]), .QN(n2573) );
  DFFR_X1 \REGISTERS_reg[31][26]  ( .D(n4211), .CK(CLK), .RN(n390), .Q(n801)
         );
  DFF_X1 \OUT2_reg[26]  ( .D(n3020), .CK(CLK), .Q(OUT2[26]), .QN(n2594) );
  DFFR_X1 \REGISTERS_reg[31][25]  ( .D(n4210), .CK(CLK), .RN(n390), .Q(n800)
         );
  DFF_X1 \OUT2_reg[25]  ( .D(n3021), .CK(CLK), .Q(OUT2[25]), .QN(n2615) );
  DFFR_X1 \REGISTERS_reg[31][24]  ( .D(n4209), .CK(CLK), .RN(n390), .Q(n799)
         );
  DFF_X1 \OUT2_reg[24]  ( .D(n3022), .CK(CLK), .Q(OUT2[24]), .QN(n2636) );
  DFFR_X1 \REGISTERS_reg[31][23]  ( .D(n4208), .CK(CLK), .RN(n390), .Q(n798)
         );
  DFF_X1 \OUT2_reg[23]  ( .D(n3023), .CK(CLK), .Q(OUT2[23]), .QN(n2657) );
  DFFR_X1 \REGISTERS_reg[31][22]  ( .D(n4207), .CK(CLK), .RN(n390), .Q(n797)
         );
  DFF_X1 \OUT2_reg[22]  ( .D(n3024), .CK(CLK), .Q(OUT2[22]), .QN(n2678) );
  DFFR_X1 \REGISTERS_reg[31][21]  ( .D(n4206), .CK(CLK), .RN(n390), .Q(n796)
         );
  DFF_X1 \OUT2_reg[21]  ( .D(n3025), .CK(CLK), .Q(OUT2[21]), .QN(n2699) );
  DFFR_X1 \REGISTERS_reg[31][20]  ( .D(n4205), .CK(CLK), .RN(n390), .Q(n795)
         );
  DFF_X1 \OUT2_reg[20]  ( .D(n3026), .CK(CLK), .Q(OUT2[20]), .QN(n2720) );
  DFFR_X1 \REGISTERS_reg[31][19]  ( .D(n4204), .CK(CLK), .RN(n390), .Q(n794)
         );
  DFF_X1 \OUT2_reg[19]  ( .D(n3027), .CK(CLK), .Q(OUT2[19]), .QN(n2741) );
  DFFR_X1 \REGISTERS_reg[31][18]  ( .D(n4203), .CK(CLK), .RN(n390), .Q(n793)
         );
  DFF_X1 \OUT2_reg[18]  ( .D(n3028), .CK(CLK), .Q(OUT2[18]), .QN(n2762) );
  DFFR_X1 \REGISTERS_reg[31][17]  ( .D(n4202), .CK(CLK), .RN(n390), .Q(n792)
         );
  DFF_X1 \OUT2_reg[17]  ( .D(n3029), .CK(CLK), .Q(OUT2[17]), .QN(n2783) );
  DFFR_X1 \REGISTERS_reg[31][16]  ( .D(n4201), .CK(CLK), .RN(n390), .Q(n791)
         );
  DFF_X1 \OUT2_reg[16]  ( .D(n3030), .CK(CLK), .Q(OUT2[16]), .QN(n2804) );
  DFFR_X1 \REGISTERS_reg[31][15]  ( .D(n4200), .CK(CLK), .RN(n389), .Q(n790)
         );
  DFF_X1 \OUT2_reg[15]  ( .D(n3031), .CK(CLK), .Q(OUT2[15]), .QN(n2825) );
  DFFR_X1 \REGISTERS_reg[31][14]  ( .D(n4199), .CK(CLK), .RN(n389), .Q(n789)
         );
  DFF_X1 \OUT2_reg[14]  ( .D(n3032), .CK(CLK), .Q(OUT2[14]), .QN(n2846) );
  DFFR_X1 \REGISTERS_reg[31][13]  ( .D(n4198), .CK(CLK), .RN(n389), .Q(n788)
         );
  DFF_X1 \OUT2_reg[13]  ( .D(n3033), .CK(CLK), .Q(OUT2[13]), .QN(n2867) );
  DFFR_X1 \REGISTERS_reg[31][12]  ( .D(n4197), .CK(CLK), .RN(n389), .Q(n787)
         );
  DFF_X1 \OUT2_reg[12]  ( .D(n3034), .CK(CLK), .Q(OUT2[12]), .QN(n2888) );
  DFFR_X1 \REGISTERS_reg[31][11]  ( .D(n4196), .CK(CLK), .RN(n389), .Q(n786)
         );
  DFF_X1 \OUT2_reg[11]  ( .D(n3035), .CK(CLK), .Q(OUT2[11]), .QN(n2909) );
  DFFR_X1 \REGISTERS_reg[31][10]  ( .D(n4195), .CK(CLK), .RN(n389), .Q(n785)
         );
  DFF_X1 \OUT2_reg[10]  ( .D(n3036), .CK(CLK), .Q(OUT2[10]), .QN(n2930) );
  DFFR_X1 \REGISTERS_reg[31][9]  ( .D(n4194), .CK(CLK), .RN(n389), .Q(n784) );
  DFF_X1 \OUT2_reg[9]  ( .D(n3037), .CK(CLK), .Q(OUT2[9]), .QN(n2951) );
  DFFR_X1 \REGISTERS_reg[31][8]  ( .D(n4193), .CK(CLK), .RN(n389), .Q(n783) );
  DFF_X1 \OUT2_reg[8]  ( .D(n3038), .CK(CLK), .Q(OUT2[8]), .QN(n2972) );
  DFFR_X1 \REGISTERS_reg[31][7]  ( .D(n4192), .CK(CLK), .RN(n389), .Q(n782) );
  DFF_X1 \OUT2_reg[7]  ( .D(n3039), .CK(CLK), .Q(OUT2[7]), .QN(n3569) );
  DFFR_X1 \REGISTERS_reg[31][6]  ( .D(n4191), .CK(CLK), .RN(n389), .Q(n781) );
  DFF_X1 \OUT2_reg[6]  ( .D(n3040), .CK(CLK), .Q(OUT2[6]), .QN(n3590) );
  DFFR_X1 \REGISTERS_reg[31][5]  ( .D(n4190), .CK(CLK), .RN(n389), .Q(n780) );
  DFF_X1 \OUT2_reg[5]  ( .D(n3041), .CK(CLK), .Q(OUT2[5]), .QN(n3611) );
  DFFR_X1 \REGISTERS_reg[31][4]  ( .D(n4189), .CK(CLK), .RN(n389), .Q(n779) );
  DFF_X1 \OUT2_reg[4]  ( .D(n3042), .CK(CLK), .Q(OUT2[4]), .QN(n3632) );
  DFFR_X1 \REGISTERS_reg[31][3]  ( .D(n4188), .CK(CLK), .RN(n388), .Q(n778) );
  DFF_X1 \OUT2_reg[3]  ( .D(n3043), .CK(CLK), .Q(OUT2[3]), .QN(n3653) );
  DFFR_X1 \REGISTERS_reg[31][2]  ( .D(n4187), .CK(CLK), .RN(n388), .Q(n777) );
  DFF_X1 \OUT2_reg[2]  ( .D(n3044), .CK(CLK), .Q(OUT2[2]), .QN(n3674) );
  DFFR_X1 \REGISTERS_reg[31][1]  ( .D(n4186), .CK(CLK), .RN(n388), .Q(n776) );
  DFF_X1 \OUT2_reg[1]  ( .D(n3045), .CK(CLK), .Q(OUT2[1]), .QN(n3695) );
  DFFR_X1 \REGISTERS_reg[31][0]  ( .D(n4185), .CK(CLK), .RN(n393), .Q(n774) );
  DFF_X1 \OUT2_reg[0]  ( .D(n3046), .CK(CLK), .Q(OUT2[0]), .QN(n3716) );
  DFF_X1 \OUT1_reg[31]  ( .D(n3014), .CK(CLK), .Q(OUT1[31]), .QN(n2488) );
  DFF_X1 \OUT1_reg[30]  ( .D(n3013), .CK(CLK), .Q(OUT1[30]), .QN(n2487) );
  DFF_X1 \OUT1_reg[29]  ( .D(n3012), .CK(CLK), .Q(OUT1[29]), .QN(n2486) );
  DFF_X1 \OUT1_reg[28]  ( .D(n3011), .CK(CLK), .Q(OUT1[28]), .QN(n2485) );
  DFF_X1 \OUT1_reg[27]  ( .D(n3010), .CK(CLK), .Q(OUT1[27]), .QN(n2484) );
  DFF_X1 \OUT1_reg[26]  ( .D(n3009), .CK(CLK), .Q(OUT1[26]), .QN(n2483) );
  DFF_X1 \OUT1_reg[25]  ( .D(n3008), .CK(CLK), .Q(OUT1[25]), .QN(n2482) );
  DFF_X1 \OUT1_reg[24]  ( .D(n3007), .CK(CLK), .Q(OUT1[24]), .QN(n2481) );
  DFF_X1 \OUT1_reg[23]  ( .D(n3006), .CK(CLK), .Q(OUT1[23]), .QN(n2480) );
  DFF_X1 \OUT1_reg[22]  ( .D(n3005), .CK(CLK), .Q(OUT1[22]), .QN(n2479) );
  DFF_X1 \OUT1_reg[21]  ( .D(n3004), .CK(CLK), .Q(OUT1[21]), .QN(n2478) );
  DFF_X1 \OUT1_reg[20]  ( .D(n3003), .CK(CLK), .Q(OUT1[20]), .QN(n2477) );
  DFF_X1 \OUT1_reg[19]  ( .D(n3002), .CK(CLK), .Q(OUT1[19]), .QN(n2476) );
  DFF_X1 \OUT1_reg[18]  ( .D(n3001), .CK(CLK), .Q(OUT1[18]), .QN(n2475) );
  DFF_X1 \OUT1_reg[17]  ( .D(n3000), .CK(CLK), .Q(OUT1[17]), .QN(n2474) );
  DFF_X1 \OUT1_reg[16]  ( .D(n2999), .CK(CLK), .Q(OUT1[16]), .QN(n2473) );
  DFF_X1 \OUT1_reg[15]  ( .D(n2998), .CK(CLK), .Q(OUT1[15]), .QN(n2472) );
  DFF_X1 \OUT1_reg[14]  ( .D(n2997), .CK(CLK), .Q(OUT1[14]), .QN(n2471) );
  DFF_X1 \OUT1_reg[13]  ( .D(n2996), .CK(CLK), .Q(OUT1[13]), .QN(n2470) );
  DFF_X1 \OUT1_reg[12]  ( .D(n2995), .CK(CLK), .Q(OUT1[12]), .QN(n2469) );
  DFF_X1 \OUT1_reg[11]  ( .D(n2994), .CK(CLK), .Q(OUT1[11]), .QN(n2468) );
  DFF_X1 \OUT1_reg[10]  ( .D(n2993), .CK(CLK), .Q(OUT1[10]), .QN(n2467) );
  DFF_X1 \OUT1_reg[9]  ( .D(n2992), .CK(CLK), .Q(OUT1[9]), .QN(n2466) );
  DFF_X1 \OUT1_reg[8]  ( .D(n2991), .CK(CLK), .Q(OUT1[8]), .QN(n2465) );
  DFF_X1 \OUT1_reg[7]  ( .D(n2990), .CK(CLK), .Q(OUT1[7]), .QN(n2464) );
  DFF_X1 \OUT1_reg[6]  ( .D(n2989), .CK(CLK), .Q(OUT1[6]), .QN(n2463) );
  DFF_X1 \OUT1_reg[5]  ( .D(n2988), .CK(CLK), .Q(OUT1[5]), .QN(n2462) );
  DFF_X1 \OUT1_reg[4]  ( .D(n2987), .CK(CLK), .Q(OUT1[4]), .QN(n2461) );
  DFF_X1 \OUT1_reg[3]  ( .D(n2986), .CK(CLK), .Q(OUT1[3]), .QN(n2460) );
  DFF_X1 \OUT1_reg[2]  ( .D(n2985), .CK(CLK), .Q(OUT1[2]), .QN(n2459) );
  DFF_X1 \OUT1_reg[1]  ( .D(n2984), .CK(CLK), .Q(OUT1[1]), .QN(n2458) );
  DFF_X1 \OUT1_reg[0]  ( .D(n2983), .CK(CLK), .Q(OUT1[0]), .QN(n2457) );
  DFFR_X1 \REGISTERS_reg[28][31]  ( .D(n3110), .CK(CLK), .RN(n378), .Q(n3832), 
        .QN(n1785) );
  DFFR_X1 \REGISTERS_reg[28][30]  ( .D(n3109), .CK(CLK), .RN(n378), .Q(n3831), 
        .QN(n1753) );
  DFFR_X1 \REGISTERS_reg[28][29]  ( .D(n3108), .CK(CLK), .RN(n378), .Q(n3830), 
        .QN(n1728) );
  DFFR_X1 \REGISTERS_reg[28][28]  ( .D(n3107), .CK(CLK), .RN(n383), .Q(n3829), 
        .QN(n1703) );
  DFFR_X1 \REGISTERS_reg[28][27]  ( .D(n3106), .CK(CLK), .RN(n398), .Q(n3828), 
        .QN(n1678) );
  DFFR_X1 \REGISTERS_reg[28][26]  ( .D(n3105), .CK(CLK), .RN(n399), .Q(n3827), 
        .QN(n1653) );
  DFFR_X1 \REGISTERS_reg[28][25]  ( .D(n3104), .CK(CLK), .RN(n398), .Q(n3826), 
        .QN(n1628) );
  DFFR_X1 \REGISTERS_reg[28][24]  ( .D(n3103), .CK(CLK), .RN(n398), .Q(n3825), 
        .QN(n1603) );
  DFFR_X1 \REGISTERS_reg[28][23]  ( .D(n3102), .CK(CLK), .RN(n398), .Q(n3824), 
        .QN(n1578) );
  DFFR_X1 \REGISTERS_reg[28][22]  ( .D(n3101), .CK(CLK), .RN(n398), .Q(n3823), 
        .QN(n1553) );
  DFFR_X1 \REGISTERS_reg[28][21]  ( .D(n3100), .CK(CLK), .RN(n398), .Q(n3822), 
        .QN(n1528) );
  DFFR_X1 \REGISTERS_reg[28][20]  ( .D(n3099), .CK(CLK), .RN(n398), .Q(n3821), 
        .QN(n1503) );
  DFFR_X1 \REGISTERS_reg[28][19]  ( .D(n3098), .CK(CLK), .RN(n398), .Q(n3820), 
        .QN(n1478) );
  DFFR_X1 \REGISTERS_reg[28][18]  ( .D(n3097), .CK(CLK), .RN(n398), .Q(n3819), 
        .QN(n1453) );
  DFFR_X1 \REGISTERS_reg[28][17]  ( .D(n3096), .CK(CLK), .RN(n398), .Q(n3818), 
        .QN(n1428) );
  DFFR_X1 \REGISTERS_reg[28][16]  ( .D(n3095), .CK(CLK), .RN(n398), .Q(n3817), 
        .QN(n1403) );
  DFFR_X1 \REGISTERS_reg[28][15]  ( .D(n3094), .CK(CLK), .RN(n398), .Q(n3816), 
        .QN(n1378) );
  DFFR_X1 \REGISTERS_reg[28][14]  ( .D(n3093), .CK(CLK), .RN(n397), .Q(n3815), 
        .QN(n1353) );
  DFFR_X1 \REGISTERS_reg[28][13]  ( .D(n3092), .CK(CLK), .RN(n397), .Q(n3814), 
        .QN(n1328) );
  DFFR_X1 \REGISTERS_reg[28][12]  ( .D(n3091), .CK(CLK), .RN(n397), .Q(n3813), 
        .QN(n1303) );
  DFFR_X1 \REGISTERS_reg[28][11]  ( .D(n3090), .CK(CLK), .RN(n397), .Q(n3812), 
        .QN(n1278) );
  DFFR_X1 \REGISTERS_reg[28][10]  ( .D(n3089), .CK(CLK), .RN(n397), .Q(n3811), 
        .QN(n1253) );
  DFFR_X1 \REGISTERS_reg[28][9]  ( .D(n3088), .CK(CLK), .RN(n397), .Q(n3810), 
        .QN(n1228) );
  DFFR_X1 \REGISTERS_reg[28][8]  ( .D(n3087), .CK(CLK), .RN(n397), .Q(n3809), 
        .QN(n1203) );
  DFFR_X1 \REGISTERS_reg[28][7]  ( .D(n3086), .CK(CLK), .RN(n397), .Q(n3808), 
        .QN(n1178) );
  DFFR_X1 \REGISTERS_reg[28][6]  ( .D(n3085), .CK(CLK), .RN(n397), .Q(n3807), 
        .QN(n1153) );
  DFFR_X1 \REGISTERS_reg[28][5]  ( .D(n3084), .CK(CLK), .RN(n397), .Q(n3806), 
        .QN(n1128) );
  DFFR_X1 \REGISTERS_reg[28][4]  ( .D(n3083), .CK(CLK), .RN(n397), .Q(n3805), 
        .QN(n1103) );
  DFFR_X1 \REGISTERS_reg[28][3]  ( .D(n3082), .CK(CLK), .RN(n397), .Q(n3804), 
        .QN(n1078) );
  DFFR_X1 \REGISTERS_reg[28][2]  ( .D(n3081), .CK(CLK), .RN(n396), .Q(n3803), 
        .QN(n1053) );
  DFFR_X1 \REGISTERS_reg[28][1]  ( .D(n3080), .CK(CLK), .RN(n396), .Q(n3802), 
        .QN(n1028) );
  DFFR_X1 \REGISTERS_reg[28][0]  ( .D(n3079), .CK(CLK), .RN(n396), .Q(n3801), 
        .QN(n976) );
  DFFR_X1 \REGISTERS_reg[23][31]  ( .D(n3206), .CK(CLK), .RN(n412), .Q(n2505), 
        .QN(n1777) );
  DFFR_X1 \REGISTERS_reg[23][30]  ( .D(n3205), .CK(CLK), .RN(n412), .Q(n2526), 
        .QN(n1751) );
  DFFR_X1 \REGISTERS_reg[23][29]  ( .D(n3204), .CK(CLK), .RN(n412), .Q(n2547), 
        .QN(n1726) );
  DFFR_X1 \REGISTERS_reg[23][28]  ( .D(n3203), .CK(CLK), .RN(n412), .Q(n2568), 
        .QN(n1701) );
  DFFR_X1 \REGISTERS_reg[23][27]  ( .D(n3202), .CK(CLK), .RN(n412), .Q(n2589), 
        .QN(n1676) );
  DFFR_X1 \REGISTERS_reg[23][26]  ( .D(n3201), .CK(CLK), .RN(n412), .Q(n2610), 
        .QN(n1651) );
  DFFR_X1 \REGISTERS_reg[23][25]  ( .D(n3200), .CK(CLK), .RN(n412), .Q(n2631), 
        .QN(n1626) );
  DFFR_X1 \REGISTERS_reg[23][24]  ( .D(n3199), .CK(CLK), .RN(n412), .Q(n2652), 
        .QN(n1601) );
  DFFR_X1 \REGISTERS_reg[23][23]  ( .D(n3198), .CK(CLK), .RN(n411), .Q(n2673), 
        .QN(n1576) );
  DFFR_X1 \REGISTERS_reg[23][22]  ( .D(n3197), .CK(CLK), .RN(n411), .Q(n2694), 
        .QN(n1551) );
  DFFR_X1 \REGISTERS_reg[23][21]  ( .D(n3196), .CK(CLK), .RN(n411), .Q(n2715), 
        .QN(n1526) );
  DFFR_X1 \REGISTERS_reg[23][20]  ( .D(n3195), .CK(CLK), .RN(n411), .Q(n2736), 
        .QN(n1501) );
  DFFR_X1 \REGISTERS_reg[23][19]  ( .D(n3194), .CK(CLK), .RN(n411), .Q(n2757), 
        .QN(n1476) );
  DFFR_X1 \REGISTERS_reg[23][18]  ( .D(n3193), .CK(CLK), .RN(n411), .Q(n2778), 
        .QN(n1451) );
  DFFR_X1 \REGISTERS_reg[23][17]  ( .D(n3192), .CK(CLK), .RN(n411), .Q(n2799), 
        .QN(n1426) );
  DFFR_X1 \REGISTERS_reg[23][16]  ( .D(n3191), .CK(CLK), .RN(n411), .Q(n2820), 
        .QN(n1401) );
  DFFR_X1 \REGISTERS_reg[23][15]  ( .D(n3190), .CK(CLK), .RN(n411), .Q(n2841), 
        .QN(n1376) );
  DFFR_X1 \REGISTERS_reg[23][14]  ( .D(n3189), .CK(CLK), .RN(n411), .Q(n2862), 
        .QN(n1351) );
  DFFR_X1 \REGISTERS_reg[23][13]  ( .D(n3188), .CK(CLK), .RN(n411), .Q(n2883), 
        .QN(n1326) );
  DFFR_X1 \REGISTERS_reg[23][12]  ( .D(n3187), .CK(CLK), .RN(n411), .Q(n2904), 
        .QN(n1301) );
  DFFR_X1 \REGISTERS_reg[23][11]  ( .D(n3186), .CK(CLK), .RN(n410), .Q(n2925), 
        .QN(n1276) );
  DFFR_X1 \REGISTERS_reg[23][10]  ( .D(n3185), .CK(CLK), .RN(n410), .Q(n2946), 
        .QN(n1251) );
  DFFR_X1 \REGISTERS_reg[23][9]  ( .D(n3184), .CK(CLK), .RN(n410), .Q(n2967), 
        .QN(n1226) );
  DFFR_X1 \REGISTERS_reg[23][8]  ( .D(n3183), .CK(CLK), .RN(n410), .Q(n3564), 
        .QN(n1201) );
  DFFR_X1 \REGISTERS_reg[23][7]  ( .D(n3182), .CK(CLK), .RN(n410), .Q(n3585), 
        .QN(n1176) );
  DFFR_X1 \REGISTERS_reg[23][6]  ( .D(n3181), .CK(CLK), .RN(n410), .Q(n3606), 
        .QN(n1151) );
  DFFR_X1 \REGISTERS_reg[23][5]  ( .D(n3180), .CK(CLK), .RN(n410), .Q(n3627), 
        .QN(n1126) );
  DFFR_X1 \REGISTERS_reg[23][4]  ( .D(n3179), .CK(CLK), .RN(n410), .Q(n3648), 
        .QN(n1101) );
  DFFR_X1 \REGISTERS_reg[23][3]  ( .D(n3178), .CK(CLK), .RN(n410), .Q(n3669), 
        .QN(n1076) );
  DFFR_X1 \REGISTERS_reg[23][2]  ( .D(n3177), .CK(CLK), .RN(n410), .Q(n3690), 
        .QN(n1051) );
  DFFR_X1 \REGISTERS_reg[23][1]  ( .D(n3176), .CK(CLK), .RN(n410), .Q(n3711), 
        .QN(n1026) );
  DFFR_X1 \REGISTERS_reg[23][0]  ( .D(n3175), .CK(CLK), .RN(n410), .Q(n3732), 
        .QN(n971) );
  DFFR_X1 \REGISTERS_reg[22][31]  ( .D(n3238), .CK(CLK), .RN(n415), .Q(n2506), 
        .QN(n1793) );
  DFFR_X1 \REGISTERS_reg[22][30]  ( .D(n3237), .CK(CLK), .RN(n415), .Q(n2527), 
        .QN(n1758) );
  DFFR_X1 \REGISTERS_reg[22][29]  ( .D(n3236), .CK(CLK), .RN(n415), .Q(n2548), 
        .QN(n1733) );
  DFFR_X1 \REGISTERS_reg[22][28]  ( .D(n3235), .CK(CLK), .RN(n415), .Q(n2569), 
        .QN(n1708) );
  DFFR_X1 \REGISTERS_reg[22][27]  ( .D(n3234), .CK(CLK), .RN(n415), .Q(n2590), 
        .QN(n1683) );
  DFFR_X1 \REGISTERS_reg[22][26]  ( .D(n3233), .CK(CLK), .RN(n414), .Q(n2611), 
        .QN(n1658) );
  DFFR_X1 \REGISTERS_reg[22][25]  ( .D(n3232), .CK(CLK), .RN(n414), .Q(n2632), 
        .QN(n1633) );
  DFFR_X1 \REGISTERS_reg[22][24]  ( .D(n3231), .CK(CLK), .RN(n414), .Q(n2653), 
        .QN(n1608) );
  DFFR_X1 \REGISTERS_reg[22][23]  ( .D(n3230), .CK(CLK), .RN(n414), .Q(n2674), 
        .QN(n1583) );
  DFFR_X1 \REGISTERS_reg[22][22]  ( .D(n3229), .CK(CLK), .RN(n414), .Q(n2695), 
        .QN(n1558) );
  DFFR_X1 \REGISTERS_reg[22][21]  ( .D(n3228), .CK(CLK), .RN(n414), .Q(n2716), 
        .QN(n1533) );
  DFFR_X1 \REGISTERS_reg[22][20]  ( .D(n3227), .CK(CLK), .RN(n414), .Q(n2737), 
        .QN(n1508) );
  DFFR_X1 \REGISTERS_reg[22][19]  ( .D(n3226), .CK(CLK), .RN(n414), .Q(n2758), 
        .QN(n1483) );
  DFFR_X1 \REGISTERS_reg[22][18]  ( .D(n3225), .CK(CLK), .RN(n414), .Q(n2779), 
        .QN(n1458) );
  DFFR_X1 \REGISTERS_reg[22][17]  ( .D(n3224), .CK(CLK), .RN(n414), .Q(n2800), 
        .QN(n1433) );
  DFFR_X1 \REGISTERS_reg[22][16]  ( .D(n3223), .CK(CLK), .RN(n414), .Q(n2821), 
        .QN(n1408) );
  DFFR_X1 \REGISTERS_reg[22][15]  ( .D(n3222), .CK(CLK), .RN(n413), .Q(n2842), 
        .QN(n1383) );
  DFFR_X1 \REGISTERS_reg[22][14]  ( .D(n3221), .CK(CLK), .RN(n413), .Q(n2863), 
        .QN(n1358) );
  DFFR_X1 \REGISTERS_reg[22][13]  ( .D(n3220), .CK(CLK), .RN(n413), .Q(n2884), 
        .QN(n1333) );
  DFFR_X1 \REGISTERS_reg[22][12]  ( .D(n3219), .CK(CLK), .RN(n413), .Q(n2905), 
        .QN(n1308) );
  DFFR_X1 \REGISTERS_reg[22][11]  ( .D(n3218), .CK(CLK), .RN(n413), .Q(n2926), 
        .QN(n1283) );
  DFFR_X1 \REGISTERS_reg[22][10]  ( .D(n3217), .CK(CLK), .RN(n413), .Q(n2947), 
        .QN(n1258) );
  DFFR_X1 \REGISTERS_reg[22][9]  ( .D(n3216), .CK(CLK), .RN(n413), .Q(n2968), 
        .QN(n1233) );
  DFFR_X1 \REGISTERS_reg[22][8]  ( .D(n3215), .CK(CLK), .RN(n413), .Q(n3565), 
        .QN(n1208) );
  DFFR_X1 \REGISTERS_reg[22][7]  ( .D(n3214), .CK(CLK), .RN(n413), .Q(n3586), 
        .QN(n1183) );
  DFFR_X1 \REGISTERS_reg[22][6]  ( .D(n3213), .CK(CLK), .RN(n413), .Q(n3607), 
        .QN(n1158) );
  DFFR_X1 \REGISTERS_reg[22][5]  ( .D(n3212), .CK(CLK), .RN(n413), .Q(n3628), 
        .QN(n1133) );
  DFFR_X1 \REGISTERS_reg[22][4]  ( .D(n3211), .CK(CLK), .RN(n413), .Q(n3649), 
        .QN(n1108) );
  DFFR_X1 \REGISTERS_reg[22][3]  ( .D(n3210), .CK(CLK), .RN(n412), .Q(n3670), 
        .QN(n1083) );
  DFFR_X1 \REGISTERS_reg[22][2]  ( .D(n3209), .CK(CLK), .RN(n412), .Q(n3691), 
        .QN(n1058) );
  DFFR_X1 \REGISTERS_reg[22][1]  ( .D(n3208), .CK(CLK), .RN(n412), .Q(n3712), 
        .QN(n1033) );
  DFFR_X1 \REGISTERS_reg[22][0]  ( .D(n3207), .CK(CLK), .RN(n412), .Q(n3733), 
        .QN(n989) );
  DFFR_X1 \REGISTERS_reg[7][31]  ( .D(n3462), .CK(CLK), .RN(n372), .Q(n2498), 
        .QN(n1806) );
  DFFR_X1 \REGISTERS_reg[7][30]  ( .D(n3461), .CK(CLK), .RN(n372), .Q(n2519), 
        .QN(n1767) );
  DFFR_X1 \REGISTERS_reg[7][29]  ( .D(n3460), .CK(CLK), .RN(n372), .Q(n2540), 
        .QN(n1742) );
  DFFR_X1 \REGISTERS_reg[7][28]  ( .D(n3459), .CK(CLK), .RN(n372), .Q(n2561), 
        .QN(n1717) );
  DFFR_X1 \REGISTERS_reg[7][27]  ( .D(n3458), .CK(CLK), .RN(n372), .Q(n2582), 
        .QN(n1692) );
  DFFR_X1 \REGISTERS_reg[7][26]  ( .D(n3457), .CK(CLK), .RN(n372), .Q(n2603), 
        .QN(n1667) );
  DFFR_X1 \REGISTERS_reg[7][25]  ( .D(n3456), .CK(CLK), .RN(n372), .Q(n2624), 
        .QN(n1642) );
  DFFR_X1 \REGISTERS_reg[7][24]  ( .D(n3455), .CK(CLK), .RN(n372), .Q(n2645), 
        .QN(n1617) );
  DFFR_X1 \REGISTERS_reg[7][23]  ( .D(n3454), .CK(CLK), .RN(n372), .Q(n2666), 
        .QN(n1592) );
  DFFR_X1 \REGISTERS_reg[7][22]  ( .D(n3453), .CK(CLK), .RN(n371), .Q(n2687), 
        .QN(n1567) );
  DFFR_X1 \REGISTERS_reg[7][21]  ( .D(n3452), .CK(CLK), .RN(n371), .Q(n2708), 
        .QN(n1542) );
  DFFR_X1 \REGISTERS_reg[7][20]  ( .D(n3451), .CK(CLK), .RN(n371), .Q(n2729), 
        .QN(n1517) );
  DFFR_X1 \REGISTERS_reg[7][19]  ( .D(n3450), .CK(CLK), .RN(n371), .Q(n2750), 
        .QN(n1492) );
  DFFR_X1 \REGISTERS_reg[7][18]  ( .D(n3449), .CK(CLK), .RN(n371), .Q(n2771), 
        .QN(n1467) );
  DFFR_X1 \REGISTERS_reg[7][17]  ( .D(n3448), .CK(CLK), .RN(n371), .Q(n2792), 
        .QN(n1442) );
  DFFR_X1 \REGISTERS_reg[7][16]  ( .D(n3447), .CK(CLK), .RN(n371), .Q(n2813), 
        .QN(n1417) );
  DFFR_X1 \REGISTERS_reg[7][15]  ( .D(n3446), .CK(CLK), .RN(n371), .Q(n2834), 
        .QN(n1392) );
  DFFR_X1 \REGISTERS_reg[7][14]  ( .D(n3445), .CK(CLK), .RN(n371), .Q(n2855), 
        .QN(n1367) );
  DFFR_X1 \REGISTERS_reg[7][13]  ( .D(n3444), .CK(CLK), .RN(n371), .Q(n2876), 
        .QN(n1342) );
  DFFR_X1 \REGISTERS_reg[7][12]  ( .D(n3443), .CK(CLK), .RN(n371), .Q(n2897), 
        .QN(n1317) );
  DFFR_X1 \REGISTERS_reg[7][11]  ( .D(n3442), .CK(CLK), .RN(n371), .Q(n2918), 
        .QN(n1292) );
  DFFR_X1 \REGISTERS_reg[7][10]  ( .D(n3441), .CK(CLK), .RN(n370), .Q(n2939), 
        .QN(n1267) );
  DFFR_X1 \REGISTERS_reg[7][9]  ( .D(n3440), .CK(CLK), .RN(n370), .Q(n2960), 
        .QN(n1242) );
  DFFR_X1 \REGISTERS_reg[7][8]  ( .D(n3439), .CK(CLK), .RN(n370), .Q(n2981), 
        .QN(n1217) );
  DFFR_X1 \REGISTERS_reg[7][7]  ( .D(n3438), .CK(CLK), .RN(n370), .Q(n3578), 
        .QN(n1192) );
  DFFR_X1 \REGISTERS_reg[7][6]  ( .D(n3437), .CK(CLK), .RN(n370), .Q(n3599), 
        .QN(n1167) );
  DFFR_X1 \REGISTERS_reg[7][5]  ( .D(n3436), .CK(CLK), .RN(n370), .Q(n3620), 
        .QN(n1142) );
  DFFR_X1 \REGISTERS_reg[7][4]  ( .D(n3435), .CK(CLK), .RN(n370), .Q(n3641), 
        .QN(n1117) );
  DFFR_X1 \REGISTERS_reg[7][3]  ( .D(n3434), .CK(CLK), .RN(n370), .Q(n3662), 
        .QN(n1092) );
  DFFR_X1 \REGISTERS_reg[7][2]  ( .D(n3433), .CK(CLK), .RN(n370), .Q(n3683), 
        .QN(n1067) );
  DFFR_X1 \REGISTERS_reg[7][1]  ( .D(n3432), .CK(CLK), .RN(n370), .Q(n3704), 
        .QN(n1042) );
  DFFR_X1 \REGISTERS_reg[7][0]  ( .D(n3431), .CK(CLK), .RN(n370), .Q(n3725), 
        .QN(n1012) );
  DFFR_X1 \REGISTERS_reg[6][31]  ( .D(n3494), .CK(CLK), .RN(n375), .Q(n2499), 
        .QN(n1805) );
  DFFR_X1 \REGISTERS_reg[6][30]  ( .D(n3493), .CK(CLK), .RN(n375), .Q(n2520), 
        .QN(n1766) );
  DFFR_X1 \REGISTERS_reg[6][29]  ( .D(n3492), .CK(CLK), .RN(n375), .Q(n2541), 
        .QN(n1741) );
  DFFR_X1 \REGISTERS_reg[6][28]  ( .D(n3491), .CK(CLK), .RN(n375), .Q(n2562), 
        .QN(n1716) );
  DFFR_X1 \REGISTERS_reg[6][27]  ( .D(n3490), .CK(CLK), .RN(n375), .Q(n2583), 
        .QN(n1691) );
  DFFR_X1 \REGISTERS_reg[6][26]  ( .D(n3489), .CK(CLK), .RN(n375), .Q(n2604), 
        .QN(n1666) );
  DFFR_X1 \REGISTERS_reg[6][25]  ( .D(n3488), .CK(CLK), .RN(n374), .Q(n2625), 
        .QN(n1641) );
  DFFR_X1 \REGISTERS_reg[6][24]  ( .D(n3487), .CK(CLK), .RN(n374), .Q(n2646), 
        .QN(n1616) );
  DFFR_X1 \REGISTERS_reg[6][23]  ( .D(n3486), .CK(CLK), .RN(n374), .Q(n2667), 
        .QN(n1591) );
  DFFR_X1 \REGISTERS_reg[6][22]  ( .D(n3485), .CK(CLK), .RN(n374), .Q(n2688), 
        .QN(n1566) );
  DFFR_X1 \REGISTERS_reg[6][21]  ( .D(n3484), .CK(CLK), .RN(n374), .Q(n2709), 
        .QN(n1541) );
  DFFR_X1 \REGISTERS_reg[6][20]  ( .D(n3483), .CK(CLK), .RN(n374), .Q(n2730), 
        .QN(n1516) );
  DFFR_X1 \REGISTERS_reg[6][19]  ( .D(n3482), .CK(CLK), .RN(n374), .Q(n2751), 
        .QN(n1491) );
  DFFR_X1 \REGISTERS_reg[6][18]  ( .D(n3481), .CK(CLK), .RN(n374), .Q(n2772), 
        .QN(n1466) );
  DFFR_X1 \REGISTERS_reg[6][17]  ( .D(n3480), .CK(CLK), .RN(n374), .Q(n2793), 
        .QN(n1441) );
  DFFR_X1 \REGISTERS_reg[6][16]  ( .D(n3479), .CK(CLK), .RN(n374), .Q(n2814), 
        .QN(n1416) );
  DFFR_X1 \REGISTERS_reg[6][15]  ( .D(n3478), .CK(CLK), .RN(n374), .Q(n2835), 
        .QN(n1391) );
  DFFR_X1 \REGISTERS_reg[6][14]  ( .D(n3477), .CK(CLK), .RN(n374), .Q(n2856), 
        .QN(n1366) );
  DFFR_X1 \REGISTERS_reg[6][13]  ( .D(n3476), .CK(CLK), .RN(n373), .Q(n2877), 
        .QN(n1341) );
  DFFR_X1 \REGISTERS_reg[6][12]  ( .D(n3475), .CK(CLK), .RN(n373), .Q(n2898), 
        .QN(n1316) );
  DFFR_X1 \REGISTERS_reg[6][11]  ( .D(n3474), .CK(CLK), .RN(n373), .Q(n2919), 
        .QN(n1291) );
  DFFR_X1 \REGISTERS_reg[6][10]  ( .D(n3473), .CK(CLK), .RN(n373), .Q(n2940), 
        .QN(n1266) );
  DFFR_X1 \REGISTERS_reg[6][9]  ( .D(n3472), .CK(CLK), .RN(n373), .Q(n2961), 
        .QN(n1241) );
  DFFR_X1 \REGISTERS_reg[6][8]  ( .D(n3471), .CK(CLK), .RN(n373), .Q(n2982), 
        .QN(n1216) );
  DFFR_X1 \REGISTERS_reg[6][7]  ( .D(n3470), .CK(CLK), .RN(n373), .Q(n3579), 
        .QN(n1191) );
  DFFR_X1 \REGISTERS_reg[6][6]  ( .D(n3469), .CK(CLK), .RN(n373), .Q(n3600), 
        .QN(n1166) );
  DFFR_X1 \REGISTERS_reg[6][5]  ( .D(n3468), .CK(CLK), .RN(n373), .Q(n3621), 
        .QN(n1141) );
  DFFR_X1 \REGISTERS_reg[6][4]  ( .D(n3467), .CK(CLK), .RN(n373), .Q(n3642), 
        .QN(n1116) );
  DFFR_X1 \REGISTERS_reg[6][3]  ( .D(n3466), .CK(CLK), .RN(n373), .Q(n3663), 
        .QN(n1091) );
  DFFR_X1 \REGISTERS_reg[6][2]  ( .D(n3465), .CK(CLK), .RN(n372), .Q(n3684), 
        .QN(n1066) );
  DFFR_X1 \REGISTERS_reg[6][1]  ( .D(n3464), .CK(CLK), .RN(n372), .Q(n3705), 
        .QN(n1041) );
  DFFR_X1 \REGISTERS_reg[6][0]  ( .D(n3463), .CK(CLK), .RN(n372), .Q(n3726), 
        .QN(n1010) );
  DFFR_X1 \REGISTERS_reg[3][31]  ( .D(n3526), .CK(CLK), .RN(n362), .Q(n2500), 
        .QN(n1813) );
  DFFR_X1 \REGISTERS_reg[3][30]  ( .D(n3525), .CK(CLK), .RN(n362), .Q(n2521), 
        .QN(n1770) );
  DFFR_X1 \REGISTERS_reg[3][29]  ( .D(n3524), .CK(CLK), .RN(n362), .Q(n2542), 
        .QN(n1745) );
  DFFR_X1 \REGISTERS_reg[3][28]  ( .D(n3523), .CK(CLK), .RN(n362), .Q(n2563), 
        .QN(n1720) );
  DFFR_X1 \REGISTERS_reg[3][27]  ( .D(n3522), .CK(CLK), .RN(n362), .Q(n2584), 
        .QN(n1695) );
  DFFR_X1 \REGISTERS_reg[3][26]  ( .D(n3521), .CK(CLK), .RN(n362), .Q(n2605), 
        .QN(n1670) );
  DFFR_X1 \REGISTERS_reg[3][25]  ( .D(n3520), .CK(CLK), .RN(n362), .Q(n2626), 
        .QN(n1645) );
  DFFR_X1 \REGISTERS_reg[3][24]  ( .D(n3519), .CK(CLK), .RN(n362), .Q(n2647), 
        .QN(n1620) );
  DFFR_X1 \REGISTERS_reg[3][23]  ( .D(n3518), .CK(CLK), .RN(n362), .Q(n2668), 
        .QN(n1595) );
  DFFR_X1 \REGISTERS_reg[3][22]  ( .D(n3517), .CK(CLK), .RN(n362), .Q(n2689), 
        .QN(n1570) );
  DFFR_X1 \REGISTERS_reg[3][21]  ( .D(n3516), .CK(CLK), .RN(n361), .Q(n2710), 
        .QN(n1545) );
  DFFR_X1 \REGISTERS_reg[3][20]  ( .D(n3515), .CK(CLK), .RN(n361), .Q(n2731), 
        .QN(n1520) );
  DFFR_X1 \REGISTERS_reg[3][19]  ( .D(n3514), .CK(CLK), .RN(n361), .Q(n2752), 
        .QN(n1495) );
  DFFR_X1 \REGISTERS_reg[3][18]  ( .D(n3513), .CK(CLK), .RN(n361), .Q(n2773), 
        .QN(n1470) );
  DFFR_X1 \REGISTERS_reg[3][17]  ( .D(n3512), .CK(CLK), .RN(n361), .Q(n2794), 
        .QN(n1445) );
  DFFR_X1 \REGISTERS_reg[3][16]  ( .D(n3511), .CK(CLK), .RN(n361), .Q(n2815), 
        .QN(n1420) );
  DFFR_X1 \REGISTERS_reg[3][15]  ( .D(n3510), .CK(CLK), .RN(n361), .Q(n2836), 
        .QN(n1395) );
  DFFR_X1 \REGISTERS_reg[3][14]  ( .D(n3509), .CK(CLK), .RN(n361), .Q(n2857), 
        .QN(n1370) );
  DFFR_X1 \REGISTERS_reg[3][13]  ( .D(n3508), .CK(CLK), .RN(n361), .Q(n2878), 
        .QN(n1345) );
  DFFR_X1 \REGISTERS_reg[3][12]  ( .D(n3507), .CK(CLK), .RN(n361), .Q(n2899), 
        .QN(n1320) );
  DFFR_X1 \REGISTERS_reg[3][11]  ( .D(n3506), .CK(CLK), .RN(n361), .Q(n2920), 
        .QN(n1295) );
  DFFR_X1 \REGISTERS_reg[3][10]  ( .D(n3505), .CK(CLK), .RN(n361), .Q(n2941), 
        .QN(n1270) );
  DFFR_X1 \REGISTERS_reg[3][9]  ( .D(n3504), .CK(CLK), .RN(n360), .Q(n2962), 
        .QN(n1245) );
  DFFR_X1 \REGISTERS_reg[3][8]  ( .D(n3503), .CK(CLK), .RN(n360), .Q(n3559), 
        .QN(n1220) );
  DFFR_X1 \REGISTERS_reg[3][7]  ( .D(n3502), .CK(CLK), .RN(n360), .Q(n3580), 
        .QN(n1195) );
  DFFR_X1 \REGISTERS_reg[3][6]  ( .D(n3501), .CK(CLK), .RN(n360), .Q(n3601), 
        .QN(n1170) );
  DFFR_X1 \REGISTERS_reg[3][5]  ( .D(n3500), .CK(CLK), .RN(n360), .Q(n3622), 
        .QN(n1145) );
  DFFR_X1 \REGISTERS_reg[3][4]  ( .D(n3499), .CK(CLK), .RN(n360), .Q(n3643), 
        .QN(n1120) );
  DFFR_X1 \REGISTERS_reg[3][3]  ( .D(n3498), .CK(CLK), .RN(n360), .Q(n3664), 
        .QN(n1095) );
  DFFR_X1 \REGISTERS_reg[3][2]  ( .D(n3497), .CK(CLK), .RN(n360), .Q(n3685), 
        .QN(n1070) );
  DFFR_X1 \REGISTERS_reg[3][1]  ( .D(n3496), .CK(CLK), .RN(n360), .Q(n3706), 
        .QN(n1045) );
  DFFR_X1 \REGISTERS_reg[3][0]  ( .D(n3495), .CK(CLK), .RN(n360), .Q(n3727), 
        .QN(n1019) );
  DFFR_X1 \REGISTERS_reg[2][31]  ( .D(n3558), .CK(CLK), .RN(n365), .Q(n2501), 
        .QN(n1812) );
  DFFR_X1 \REGISTERS_reg[2][30]  ( .D(n3557), .CK(CLK), .RN(n365), .Q(n2522), 
        .QN(n1769) );
  DFFR_X1 \REGISTERS_reg[2][29]  ( .D(n3556), .CK(CLK), .RN(n365), .Q(n2543), 
        .QN(n1744) );
  DFFR_X1 \REGISTERS_reg[2][28]  ( .D(n3555), .CK(CLK), .RN(n365), .Q(n2564), 
        .QN(n1719) );
  DFFR_X1 \REGISTERS_reg[2][27]  ( .D(n3554), .CK(CLK), .RN(n365), .Q(n2585), 
        .QN(n1694) );
  DFFR_X1 \REGISTERS_reg[2][26]  ( .D(n3553), .CK(CLK), .RN(n365), .Q(n2606), 
        .QN(n1669) );
  DFFR_X1 \REGISTERS_reg[2][25]  ( .D(n3552), .CK(CLK), .RN(n365), .Q(n2627), 
        .QN(n1644) );
  DFFR_X1 \REGISTERS_reg[2][24]  ( .D(n3551), .CK(CLK), .RN(n364), .Q(n2648), 
        .QN(n1619) );
  DFFR_X1 \REGISTERS_reg[2][23]  ( .D(n3550), .CK(CLK), .RN(n364), .Q(n2669), 
        .QN(n1594) );
  DFFR_X1 \REGISTERS_reg[2][22]  ( .D(n3549), .CK(CLK), .RN(n364), .Q(n2690), 
        .QN(n1569) );
  DFFR_X1 \REGISTERS_reg[2][21]  ( .D(n3548), .CK(CLK), .RN(n364), .Q(n2711), 
        .QN(n1544) );
  DFFR_X1 \REGISTERS_reg[2][20]  ( .D(n3547), .CK(CLK), .RN(n364), .Q(n2732), 
        .QN(n1519) );
  DFFR_X1 \REGISTERS_reg[2][19]  ( .D(n3546), .CK(CLK), .RN(n364), .Q(n2753), 
        .QN(n1494) );
  DFFR_X1 \REGISTERS_reg[2][18]  ( .D(n3545), .CK(CLK), .RN(n364), .Q(n2774), 
        .QN(n1469) );
  DFFR_X1 \REGISTERS_reg[2][17]  ( .D(n3544), .CK(CLK), .RN(n364), .Q(n2795), 
        .QN(n1444) );
  DFFR_X1 \REGISTERS_reg[2][16]  ( .D(n3543), .CK(CLK), .RN(n364), .Q(n2816), 
        .QN(n1419) );
  DFFR_X1 \REGISTERS_reg[2][15]  ( .D(n3542), .CK(CLK), .RN(n364), .Q(n2837), 
        .QN(n1394) );
  DFFR_X1 \REGISTERS_reg[2][14]  ( .D(n3541), .CK(CLK), .RN(n364), .Q(n2858), 
        .QN(n1369) );
  DFFR_X1 \REGISTERS_reg[2][13]  ( .D(n3540), .CK(CLK), .RN(n364), .Q(n2879), 
        .QN(n1344) );
  DFFR_X1 \REGISTERS_reg[2][12]  ( .D(n3539), .CK(CLK), .RN(n363), .Q(n2900), 
        .QN(n1319) );
  DFFR_X1 \REGISTERS_reg[2][11]  ( .D(n3538), .CK(CLK), .RN(n363), .Q(n2921), 
        .QN(n1294) );
  DFFR_X1 \REGISTERS_reg[2][10]  ( .D(n3537), .CK(CLK), .RN(n363), .Q(n2942), 
        .QN(n1269) );
  DFFR_X1 \REGISTERS_reg[2][9]  ( .D(n3536), .CK(CLK), .RN(n363), .Q(n2963), 
        .QN(n1244) );
  DFFR_X1 \REGISTERS_reg[2][8]  ( .D(n3535), .CK(CLK), .RN(n363), .Q(n3560), 
        .QN(n1219) );
  DFFR_X1 \REGISTERS_reg[2][7]  ( .D(n3534), .CK(CLK), .RN(n363), .Q(n3581), 
        .QN(n1194) );
  DFFR_X1 \REGISTERS_reg[2][6]  ( .D(n3533), .CK(CLK), .RN(n363), .Q(n3602), 
        .QN(n1169) );
  DFFR_X1 \REGISTERS_reg[2][5]  ( .D(n3532), .CK(CLK), .RN(n363), .Q(n3623), 
        .QN(n1144) );
  DFFR_X1 \REGISTERS_reg[2][4]  ( .D(n3531), .CK(CLK), .RN(n363), .Q(n3644), 
        .QN(n1119) );
  DFFR_X1 \REGISTERS_reg[2][3]  ( .D(n3530), .CK(CLK), .RN(n363), .Q(n3665), 
        .QN(n1094) );
  DFFR_X1 \REGISTERS_reg[2][2]  ( .D(n3529), .CK(CLK), .RN(n363), .Q(n3686), 
        .QN(n1069) );
  DFFR_X1 \REGISTERS_reg[2][1]  ( .D(n3528), .CK(CLK), .RN(n363), .Q(n3707), 
        .QN(n1044) );
  DFFR_X1 \REGISTERS_reg[2][0]  ( .D(n3527), .CK(CLK), .RN(n362), .Q(n3728), 
        .QN(n1017) );
  DFFR_X1 \REGISTERS_reg[25][31]  ( .D(n3142), .CK(CLK), .RN(n386), .Q(n2502)
         );
  DFFR_X1 \REGISTERS_reg[25][30]  ( .D(n3141), .CK(CLK), .RN(n386), .Q(n2523)
         );
  DFFR_X1 \REGISTERS_reg[25][29]  ( .D(n3140), .CK(CLK), .RN(n386), .Q(n2544)
         );
  DFFR_X1 \REGISTERS_reg[25][28]  ( .D(n3139), .CK(CLK), .RN(n386), .Q(n2565)
         );
  DFFR_X1 \REGISTERS_reg[25][27]  ( .D(n3138), .CK(CLK), .RN(n386), .Q(n2586)
         );
  DFFR_X1 \REGISTERS_reg[25][26]  ( .D(n3137), .CK(CLK), .RN(n386), .Q(n2607)
         );
  DFFR_X1 \REGISTERS_reg[25][25]  ( .D(n3136), .CK(CLK), .RN(n386), .Q(n2628)
         );
  DFFR_X1 \REGISTERS_reg[25][24]  ( .D(n3135), .CK(CLK), .RN(n386), .Q(n2649)
         );
  DFFR_X1 \REGISTERS_reg[25][23]  ( .D(n3134), .CK(CLK), .RN(n386), .Q(n2670)
         );
  DFFR_X1 \REGISTERS_reg[25][22]  ( .D(n3133), .CK(CLK), .RN(n385), .Q(n2691)
         );
  DFFR_X1 \REGISTERS_reg[25][21]  ( .D(n3132), .CK(CLK), .RN(n385), .Q(n2712)
         );
  DFFR_X1 \REGISTERS_reg[25][20]  ( .D(n3131), .CK(CLK), .RN(n385), .Q(n2733)
         );
  DFFR_X1 \REGISTERS_reg[25][19]  ( .D(n3130), .CK(CLK), .RN(n385), .Q(n2754)
         );
  DFFR_X1 \REGISTERS_reg[25][18]  ( .D(n3129), .CK(CLK), .RN(n385), .Q(n2775)
         );
  DFFR_X1 \REGISTERS_reg[25][17]  ( .D(n3128), .CK(CLK), .RN(n385), .Q(n2796)
         );
  DFFR_X1 \REGISTERS_reg[25][16]  ( .D(n3127), .CK(CLK), .RN(n385), .Q(n2817)
         );
  DFFR_X1 \REGISTERS_reg[25][15]  ( .D(n3126), .CK(CLK), .RN(n385), .Q(n2838)
         );
  DFFR_X1 \REGISTERS_reg[25][14]  ( .D(n3125), .CK(CLK), .RN(n385), .Q(n2859)
         );
  DFFR_X1 \REGISTERS_reg[25][13]  ( .D(n3124), .CK(CLK), .RN(n385), .Q(n2880)
         );
  DFFR_X1 \REGISTERS_reg[25][12]  ( .D(n3123), .CK(CLK), .RN(n385), .Q(n2901)
         );
  DFFR_X1 \REGISTERS_reg[25][11]  ( .D(n3122), .CK(CLK), .RN(n385), .Q(n2922)
         );
  DFFR_X1 \REGISTERS_reg[25][10]  ( .D(n3121), .CK(CLK), .RN(n384), .Q(n2943)
         );
  DFFR_X1 \REGISTERS_reg[25][9]  ( .D(n3120), .CK(CLK), .RN(n384), .Q(n2964)
         );
  DFFR_X1 \REGISTERS_reg[25][8]  ( .D(n3119), .CK(CLK), .RN(n384), .Q(n3561)
         );
  DFFR_X1 \REGISTERS_reg[25][7]  ( .D(n3118), .CK(CLK), .RN(n384), .Q(n3582)
         );
  DFFR_X1 \REGISTERS_reg[25][6]  ( .D(n3117), .CK(CLK), .RN(n384), .Q(n3603)
         );
  DFFR_X1 \REGISTERS_reg[25][5]  ( .D(n3116), .CK(CLK), .RN(n384), .Q(n3624)
         );
  DFFR_X1 \REGISTERS_reg[25][4]  ( .D(n3115), .CK(CLK), .RN(n384), .Q(n3645)
         );
  BUF_X1 U2 ( .A(n420), .Z(n419) );
  BUF_X1 U3 ( .A(n980), .Z(n122) );
  BUF_X1 U4 ( .A(n980), .Z(n121) );
  BUF_X1 U5 ( .A(n980), .Z(n123) );
  BUF_X1 U6 ( .A(n1838), .Z(n223) );
  BUF_X1 U7 ( .A(n1833), .Z(n211) );
  BUF_X1 U8 ( .A(n1848), .Z(n244) );
  BUF_X1 U9 ( .A(n1838), .Z(n224) );
  BUF_X1 U10 ( .A(n1833), .Z(n212) );
  BUF_X1 U11 ( .A(n1848), .Z(n245) );
  BUF_X1 U12 ( .A(n974), .Z(n110) );
  BUF_X1 U13 ( .A(n991), .Z(n143) );
  BUF_X1 U14 ( .A(n974), .Z(n109) );
  BUF_X1 U15 ( .A(n991), .Z(n142) );
  BUF_X1 U16 ( .A(n1003), .Z(n164) );
  BUF_X1 U17 ( .A(n1003), .Z(n163) );
  BUF_X1 U18 ( .A(n1844), .Z(n235) );
  BUF_X1 U19 ( .A(n1870), .Z(n289) );
  BUF_X1 U20 ( .A(n1844), .Z(n236) );
  BUF_X1 U21 ( .A(n1870), .Z(n290) );
  BUF_X1 U22 ( .A(n986), .Z(n134) );
  BUF_X1 U23 ( .A(n998), .Z(n152) );
  BUF_X1 U24 ( .A(n1008), .Z(n176) );
  BUF_X1 U25 ( .A(n1015), .Z(n188) );
  BUF_X1 U26 ( .A(n986), .Z(n133) );
  BUF_X1 U27 ( .A(n998), .Z(n151) );
  BUF_X1 U28 ( .A(n1008), .Z(n175) );
  BUF_X1 U29 ( .A(n1015), .Z(n187) );
  BUF_X1 U30 ( .A(n1020), .Z(n194) );
  BUF_X1 U31 ( .A(n1020), .Z(n193) );
  BUF_X1 U32 ( .A(n1001), .Z(n158) );
  BUF_X1 U33 ( .A(n1006), .Z(n170) );
  BUF_X1 U34 ( .A(n1001), .Z(n157) );
  BUF_X1 U35 ( .A(n1006), .Z(n169) );
  BUF_X1 U36 ( .A(n1847), .Z(n241) );
  BUF_X1 U37 ( .A(n1847), .Z(n242) );
  BUF_X1 U38 ( .A(n990), .Z(n140) );
  BUF_X1 U39 ( .A(n1013), .Z(n182) );
  BUF_X1 U40 ( .A(n990), .Z(n139) );
  BUF_X1 U41 ( .A(n1013), .Z(n181) );
  BUF_X1 U42 ( .A(n1830), .Z(n205) );
  BUF_X1 U43 ( .A(n1830), .Z(n206) );
  BUF_X1 U44 ( .A(n970), .Z(n104) );
  BUF_X1 U45 ( .A(n970), .Z(n103) );
  BUF_X1 U46 ( .A(n1835), .Z(n217) );
  BUF_X1 U47 ( .A(n1835), .Z(n218) );
  BUF_X1 U48 ( .A(n977), .Z(n116) );
  BUF_X1 U49 ( .A(n977), .Z(n115) );
  BUF_X1 U50 ( .A(n1018), .Z(n191) );
  BUF_X1 U51 ( .A(n1018), .Z(n190) );
  BUF_X1 U52 ( .A(n1846), .Z(n238) );
  BUF_X1 U53 ( .A(n1846), .Z(n239) );
  BUF_X1 U54 ( .A(n988), .Z(n137) );
  BUF_X1 U55 ( .A(n988), .Z(n136) );
  BUF_X1 U56 ( .A(n1000), .Z(n155) );
  BUF_X1 U57 ( .A(n1005), .Z(n167) );
  BUF_X1 U58 ( .A(n1000), .Z(n154) );
  BUF_X1 U59 ( .A(n1005), .Z(n166) );
  BUF_X1 U60 ( .A(n1011), .Z(n179) );
  BUF_X1 U61 ( .A(n1011), .Z(n178) );
  BUF_X1 U62 ( .A(n1836), .Z(n220) );
  BUF_X1 U63 ( .A(n1831), .Z(n208) );
  BUF_X1 U64 ( .A(n1836), .Z(n221) );
  BUF_X1 U65 ( .A(n1831), .Z(n209) );
  BUF_X1 U66 ( .A(n978), .Z(n119) );
  BUF_X1 U67 ( .A(n972), .Z(n107) );
  BUF_X1 U68 ( .A(n978), .Z(n118) );
  BUF_X1 U69 ( .A(n972), .Z(n106) );
  BUF_X1 U70 ( .A(n1839), .Z(n226) );
  BUF_X1 U71 ( .A(n1834), .Z(n214) );
  BUF_X1 U72 ( .A(n1849), .Z(n247) );
  BUF_X1 U73 ( .A(n1839), .Z(n227) );
  BUF_X1 U74 ( .A(n1834), .Z(n215) );
  BUF_X1 U75 ( .A(n1849), .Z(n248) );
  BUF_X1 U76 ( .A(n981), .Z(n125) );
  BUF_X1 U77 ( .A(n975), .Z(n113) );
  BUF_X1 U78 ( .A(n992), .Z(n146) );
  BUF_X1 U79 ( .A(n981), .Z(n124) );
  BUF_X1 U80 ( .A(n975), .Z(n112) );
  BUF_X1 U81 ( .A(n992), .Z(n145) );
  BUF_X1 U82 ( .A(n997), .Z(n149) );
  BUF_X1 U83 ( .A(n997), .Z(n148) );
  BUF_X1 U84 ( .A(n1002), .Z(n161) );
  BUF_X1 U85 ( .A(n1002), .Z(n160) );
  BUF_X1 U86 ( .A(n1843), .Z(n232) );
  BUF_X1 U87 ( .A(n1843), .Z(n233) );
  BUF_X1 U88 ( .A(n985), .Z(n131) );
  BUF_X1 U89 ( .A(n1007), .Z(n173) );
  BUF_X1 U90 ( .A(n1014), .Z(n185) );
  BUF_X1 U91 ( .A(n985), .Z(n130) );
  BUF_X1 U92 ( .A(n1007), .Z(n172) );
  BUF_X1 U93 ( .A(n1014), .Z(n184) );
  BUF_X1 U94 ( .A(n1840), .Z(n229) );
  BUF_X1 U95 ( .A(n1840), .Z(n230) );
  BUF_X1 U96 ( .A(n982), .Z(n128) );
  BUF_X1 U97 ( .A(n982), .Z(n127) );
  BUF_X1 U98 ( .A(n1838), .Z(n225) );
  BUF_X1 U99 ( .A(n1833), .Z(n213) );
  BUF_X1 U100 ( .A(n1848), .Z(n246) );
  BUF_X1 U101 ( .A(n974), .Z(n111) );
  BUF_X1 U102 ( .A(n991), .Z(n144) );
  BUF_X1 U103 ( .A(n1003), .Z(n165) );
  BUF_X1 U104 ( .A(n998), .Z(n153) );
  BUF_X1 U105 ( .A(n1844), .Z(n237) );
  BUF_X1 U106 ( .A(n1870), .Z(n291) );
  BUF_X1 U107 ( .A(n986), .Z(n135) );
  BUF_X1 U108 ( .A(n1008), .Z(n177) );
  BUF_X1 U109 ( .A(n1015), .Z(n189) );
  BUF_X1 U110 ( .A(n1020), .Z(n195) );
  BUF_X1 U111 ( .A(n1001), .Z(n159) );
  BUF_X1 U112 ( .A(n1006), .Z(n171) );
  BUF_X1 U113 ( .A(n1847), .Z(n243) );
  BUF_X1 U114 ( .A(n990), .Z(n141) );
  BUF_X1 U115 ( .A(n1013), .Z(n183) );
  BUF_X1 U116 ( .A(n1830), .Z(n207) );
  BUF_X1 U117 ( .A(n970), .Z(n105) );
  BUF_X1 U118 ( .A(n1835), .Z(n219) );
  BUF_X1 U119 ( .A(n977), .Z(n117) );
  BUF_X1 U120 ( .A(n1018), .Z(n192) );
  BUF_X1 U121 ( .A(n1846), .Z(n240) );
  BUF_X1 U122 ( .A(n988), .Z(n138) );
  BUF_X1 U123 ( .A(n1000), .Z(n156) );
  BUF_X1 U124 ( .A(n1005), .Z(n168) );
  BUF_X1 U125 ( .A(n1011), .Z(n180) );
  BUF_X1 U126 ( .A(n1836), .Z(n222) );
  BUF_X1 U127 ( .A(n1831), .Z(n210) );
  BUF_X1 U128 ( .A(n978), .Z(n120) );
  BUF_X1 U129 ( .A(n972), .Z(n108) );
  BUF_X1 U130 ( .A(n1839), .Z(n228) );
  BUF_X1 U131 ( .A(n1834), .Z(n216) );
  BUF_X1 U132 ( .A(n1849), .Z(n249) );
  BUF_X1 U133 ( .A(n981), .Z(n126) );
  BUF_X1 U134 ( .A(n975), .Z(n114) );
  BUF_X1 U135 ( .A(n992), .Z(n147) );
  BUF_X1 U136 ( .A(n997), .Z(n150) );
  BUF_X1 U137 ( .A(n1002), .Z(n162) );
  BUF_X1 U138 ( .A(n1843), .Z(n234) );
  BUF_X1 U139 ( .A(n985), .Z(n132) );
  BUF_X1 U140 ( .A(n1007), .Z(n174) );
  BUF_X1 U141 ( .A(n1014), .Z(n186) );
  BUF_X1 U142 ( .A(n1840), .Z(n231) );
  BUF_X1 U143 ( .A(n982), .Z(n129) );
  BUF_X1 U144 ( .A(n330), .Z(n420) );
  BUF_X1 U145 ( .A(n331), .Z(n424) );
  BUF_X1 U146 ( .A(n331), .Z(n425) );
  BUF_X1 U147 ( .A(n331), .Z(n423) );
  BUF_X1 U148 ( .A(n330), .Z(n422) );
  BUF_X1 U149 ( .A(n330), .Z(n421) );
  BUF_X1 U150 ( .A(n333), .Z(n431) );
  BUF_X1 U151 ( .A(n332), .Z(n427) );
  BUF_X1 U152 ( .A(n333), .Z(n430) );
  BUF_X1 U153 ( .A(n333), .Z(n429) );
  BUF_X1 U154 ( .A(n332), .Z(n428) );
  BUF_X1 U155 ( .A(n332), .Z(n426) );
  BUF_X1 U156 ( .A(n334), .Z(n432) );
  BUF_X1 U157 ( .A(n334), .Z(n433) );
  BUF_X1 U158 ( .A(n1860), .Z(n265) );
  BUF_X1 U159 ( .A(n1860), .Z(n266) );
  BUF_X1 U160 ( .A(n1855), .Z(n253) );
  BUF_X1 U161 ( .A(n1865), .Z(n277) );
  BUF_X1 U162 ( .A(n1855), .Z(n254) );
  BUF_X1 U163 ( .A(n1865), .Z(n278) );
  BUF_X1 U164 ( .A(n1873), .Z(n295) );
  BUF_X1 U165 ( .A(n1873), .Z(n296) );
  BUF_X1 U166 ( .A(n1858), .Z(n259) );
  BUF_X1 U167 ( .A(n1863), .Z(n271) );
  BUF_X1 U168 ( .A(n1858), .Z(n260) );
  BUF_X1 U169 ( .A(n1863), .Z(n272) );
  BUF_X1 U170 ( .A(n1868), .Z(n283) );
  BUF_X1 U171 ( .A(n1868), .Z(n284) );
  BUF_X1 U172 ( .A(n1872), .Z(n292) );
  BUF_X1 U173 ( .A(n1872), .Z(n293) );
  BUF_X1 U174 ( .A(n1857), .Z(n256) );
  BUF_X1 U175 ( .A(n1862), .Z(n268) );
  BUF_X1 U176 ( .A(n1857), .Z(n257) );
  BUF_X1 U177 ( .A(n1862), .Z(n269) );
  BUF_X1 U178 ( .A(n1867), .Z(n280) );
  BUF_X1 U179 ( .A(n1867), .Z(n281) );
  BUF_X1 U180 ( .A(n1854), .Z(n250) );
  BUF_X1 U181 ( .A(n1854), .Z(n251) );
  BUF_X1 U182 ( .A(n1859), .Z(n262) );
  BUF_X1 U183 ( .A(n1859), .Z(n263) );
  BUF_X1 U184 ( .A(n1864), .Z(n274) );
  BUF_X1 U185 ( .A(n1869), .Z(n286) );
  BUF_X1 U186 ( .A(n1864), .Z(n275) );
  BUF_X1 U187 ( .A(n1869), .Z(n287) );
  BUF_X1 U188 ( .A(n1860), .Z(n267) );
  BUF_X1 U189 ( .A(n1855), .Z(n255) );
  BUF_X1 U190 ( .A(n1865), .Z(n279) );
  BUF_X1 U191 ( .A(n1873), .Z(n297) );
  BUF_X1 U192 ( .A(n1858), .Z(n261) );
  BUF_X1 U193 ( .A(n1863), .Z(n273) );
  BUF_X1 U194 ( .A(n1868), .Z(n285) );
  BUF_X1 U195 ( .A(n1872), .Z(n294) );
  BUF_X1 U196 ( .A(n1857), .Z(n258) );
  BUF_X1 U197 ( .A(n1862), .Z(n270) );
  BUF_X1 U198 ( .A(n1867), .Z(n282) );
  BUF_X1 U199 ( .A(n1854), .Z(n252) );
  BUF_X1 U200 ( .A(n1859), .Z(n264) );
  BUF_X1 U201 ( .A(n1864), .Z(n276) );
  BUF_X1 U202 ( .A(n1869), .Z(n288) );
  BUF_X1 U203 ( .A(n335), .Z(n333) );
  BUF_X1 U204 ( .A(n335), .Z(n332) );
  BUF_X1 U205 ( .A(n336), .Z(n331) );
  BUF_X1 U206 ( .A(n336), .Z(n330) );
  BUF_X1 U207 ( .A(n335), .Z(n334) );
  BUF_X1 U208 ( .A(n741), .Z(n29) );
  BUF_X1 U209 ( .A(n741), .Z(n28) );
  BUF_X1 U210 ( .A(n707), .Z(n26) );
  BUF_X1 U211 ( .A(n707), .Z(n25) );
  BUF_X1 U212 ( .A(n876), .Z(n41) );
  BUF_X1 U213 ( .A(n876), .Z(n40) );
  BUF_X1 U214 ( .A(n843), .Z(n38) );
  BUF_X1 U215 ( .A(n843), .Z(n37) );
  BUF_X1 U216 ( .A(n538), .Z(n11) );
  BUF_X1 U217 ( .A(n538), .Z(n10) );
  BUF_X1 U218 ( .A(n504), .Z(n8) );
  BUF_X1 U219 ( .A(n504), .Z(n7) );
  BUF_X1 U220 ( .A(n470), .Z(n5) );
  BUF_X1 U221 ( .A(n470), .Z(n4) );
  BUF_X1 U222 ( .A(n435), .Z(n2) );
  BUF_X1 U223 ( .A(n435), .Z(n1) );
  BUF_X1 U224 ( .A(n775), .Z(n32) );
  BUF_X1 U225 ( .A(n775), .Z(n31) );
  BUF_X1 U226 ( .A(n961), .Z(n91) );
  BUF_X1 U227 ( .A(n961), .Z(n92) );
  BUF_X1 U228 ( .A(n960), .Z(n88) );
  BUF_X1 U229 ( .A(n960), .Z(n89) );
  BUF_X1 U230 ( .A(n672), .Z(n23) );
  BUF_X1 U231 ( .A(n672), .Z(n22) );
  BUF_X1 U232 ( .A(n959), .Z(n85) );
  BUF_X1 U233 ( .A(n959), .Z(n86) );
  BUF_X1 U234 ( .A(n958), .Z(n82) );
  BUF_X1 U235 ( .A(n958), .Z(n83) );
  BUF_X1 U236 ( .A(n957), .Z(n79) );
  BUF_X1 U237 ( .A(n957), .Z(n80) );
  BUF_X1 U238 ( .A(n956), .Z(n76) );
  BUF_X1 U239 ( .A(n956), .Z(n77) );
  BUF_X1 U240 ( .A(n909), .Z(n44) );
  BUF_X1 U241 ( .A(n909), .Z(n43) );
  BUF_X1 U242 ( .A(n955), .Z(n73) );
  BUF_X1 U243 ( .A(n955), .Z(n74) );
  BUF_X1 U244 ( .A(n952), .Z(n70) );
  BUF_X1 U245 ( .A(n952), .Z(n71) );
  BUF_X1 U246 ( .A(n809), .Z(n35) );
  BUF_X1 U247 ( .A(n809), .Z(n34) );
  BUF_X1 U248 ( .A(n951), .Z(n67) );
  BUF_X1 U249 ( .A(n951), .Z(n68) );
  BUF_X1 U250 ( .A(n950), .Z(n64) );
  BUF_X1 U251 ( .A(n950), .Z(n65) );
  BUF_X1 U252 ( .A(n949), .Z(n61) );
  BUF_X1 U253 ( .A(n949), .Z(n62) );
  BUF_X1 U254 ( .A(n948), .Z(n58) );
  BUF_X1 U255 ( .A(n948), .Z(n59) );
  BUF_X1 U256 ( .A(n944), .Z(n55) );
  BUF_X1 U257 ( .A(n944), .Z(n56) );
  BUF_X1 U258 ( .A(n943), .Z(n52) );
  BUF_X1 U259 ( .A(n943), .Z(n53) );
  BUF_X1 U260 ( .A(n639), .Z(n20) );
  BUF_X1 U261 ( .A(n639), .Z(n19) );
  BUF_X1 U262 ( .A(n606), .Z(n17) );
  BUF_X1 U263 ( .A(n606), .Z(n16) );
  BUF_X1 U264 ( .A(n942), .Z(n49) );
  BUF_X1 U265 ( .A(n942), .Z(n50) );
  BUF_X1 U266 ( .A(n941), .Z(n46) );
  BUF_X1 U267 ( .A(n941), .Z(n47) );
  BUF_X1 U268 ( .A(n572), .Z(n14) );
  BUF_X1 U269 ( .A(n572), .Z(n13) );
  BUF_X1 U270 ( .A(n1824), .Z(n199) );
  BUF_X1 U271 ( .A(n1824), .Z(n200) );
  BUF_X1 U272 ( .A(n964), .Z(n98) );
  BUF_X1 U273 ( .A(n964), .Z(n97) );
  BUF_X1 U274 ( .A(n1822), .Z(n196) );
  BUF_X1 U275 ( .A(n1822), .Z(n197) );
  BUF_X1 U276 ( .A(n962), .Z(n95) );
  BUF_X1 U277 ( .A(n962), .Z(n94) );
  BUF_X1 U278 ( .A(n876), .Z(n42) );
  BUF_X1 U279 ( .A(n843), .Z(n39) );
  BUF_X1 U280 ( .A(n538), .Z(n12) );
  BUF_X1 U281 ( .A(n504), .Z(n9) );
  BUF_X1 U282 ( .A(n470), .Z(n6) );
  BUF_X1 U283 ( .A(n435), .Z(n3) );
  BUF_X1 U284 ( .A(n961), .Z(n93) );
  BUF_X1 U285 ( .A(n960), .Z(n90) );
  BUF_X1 U286 ( .A(n959), .Z(n87) );
  BUF_X1 U287 ( .A(n707), .Z(n27) );
  BUF_X1 U288 ( .A(n775), .Z(n33) );
  BUF_X1 U289 ( .A(n672), .Z(n24) );
  BUF_X1 U290 ( .A(n958), .Z(n84) );
  BUF_X1 U291 ( .A(n957), .Z(n81) );
  BUF_X1 U292 ( .A(n956), .Z(n78) );
  BUF_X1 U293 ( .A(n909), .Z(n45) );
  BUF_X1 U294 ( .A(n955), .Z(n75) );
  BUF_X1 U295 ( .A(n952), .Z(n72) );
  BUF_X1 U296 ( .A(n809), .Z(n36) );
  BUF_X1 U297 ( .A(n639), .Z(n21) );
  BUF_X1 U298 ( .A(n606), .Z(n18) );
  BUF_X1 U299 ( .A(n572), .Z(n15) );
  BUF_X1 U300 ( .A(n741), .Z(n30) );
  BUF_X1 U301 ( .A(n951), .Z(n69) );
  BUF_X1 U302 ( .A(n950), .Z(n66) );
  BUF_X1 U303 ( .A(n949), .Z(n63) );
  BUF_X1 U304 ( .A(n948), .Z(n60) );
  BUF_X1 U305 ( .A(n944), .Z(n57) );
  BUF_X1 U306 ( .A(n943), .Z(n54) );
  BUF_X1 U307 ( .A(n942), .Z(n51) );
  BUF_X1 U308 ( .A(n941), .Z(n48) );
  BUF_X1 U309 ( .A(n1824), .Z(n201) );
  BUF_X1 U310 ( .A(n964), .Z(n99) );
  BUF_X1 U311 ( .A(n1822), .Z(n198) );
  BUF_X1 U312 ( .A(n962), .Z(n96) );
  BUF_X1 U313 ( .A(RST), .Z(n335) );
  BUF_X1 U314 ( .A(RST), .Z(n336) );
  BUF_X1 U315 ( .A(n1825), .Z(n202) );
  BUF_X1 U316 ( .A(n965), .Z(n100) );
  BUF_X1 U317 ( .A(n1825), .Z(n203) );
  BUF_X1 U318 ( .A(n965), .Z(n101) );
  BUF_X1 U319 ( .A(n1825), .Z(n204) );
  BUF_X1 U320 ( .A(n965), .Z(n102) );
  INV_X1 U321 ( .A(DATAIN[0]), .ZN(n298) );
  INV_X1 U322 ( .A(DATAIN[1]), .ZN(n299) );
  INV_X1 U323 ( .A(DATAIN[2]), .ZN(n300) );
  INV_X1 U324 ( .A(DATAIN[3]), .ZN(n301) );
  INV_X1 U325 ( .A(DATAIN[4]), .ZN(n302) );
  INV_X1 U326 ( .A(DATAIN[5]), .ZN(n303) );
  INV_X1 U327 ( .A(DATAIN[6]), .ZN(n304) );
  INV_X1 U328 ( .A(DATAIN[7]), .ZN(n305) );
  INV_X1 U329 ( .A(DATAIN[8]), .ZN(n306) );
  INV_X1 U330 ( .A(DATAIN[10]), .ZN(n308) );
  INV_X1 U331 ( .A(DATAIN[11]), .ZN(n309) );
  INV_X1 U332 ( .A(DATAIN[12]), .ZN(n310) );
  INV_X1 U333 ( .A(DATAIN[13]), .ZN(n311) );
  INV_X1 U334 ( .A(DATAIN[14]), .ZN(n312) );
  INV_X1 U335 ( .A(DATAIN[15]), .ZN(n313) );
  INV_X1 U336 ( .A(DATAIN[16]), .ZN(n314) );
  INV_X1 U337 ( .A(DATAIN[17]), .ZN(n315) );
  INV_X1 U338 ( .A(DATAIN[18]), .ZN(n316) );
  INV_X1 U339 ( .A(DATAIN[19]), .ZN(n317) );
  INV_X1 U340 ( .A(DATAIN[20]), .ZN(n318) );
  INV_X1 U341 ( .A(DATAIN[21]), .ZN(n319) );
  INV_X1 U342 ( .A(DATAIN[22]), .ZN(n320) );
  INV_X1 U343 ( .A(DATAIN[23]), .ZN(n321) );
  INV_X1 U344 ( .A(DATAIN[24]), .ZN(n322) );
  INV_X1 U345 ( .A(DATAIN[25]), .ZN(n323) );
  INV_X1 U346 ( .A(DATAIN[26]), .ZN(n324) );
  INV_X1 U347 ( .A(DATAIN[27]), .ZN(n325) );
  INV_X1 U348 ( .A(DATAIN[28]), .ZN(n326) );
  INV_X1 U349 ( .A(DATAIN[29]), .ZN(n327) );
  INV_X1 U350 ( .A(DATAIN[30]), .ZN(n328) );
  INV_X1 U351 ( .A(DATAIN[31]), .ZN(n329) );
  INV_X1 U352 ( .A(DATAIN[9]), .ZN(n307) );
  CLKBUF_X1 U353 ( .A(n433), .Z(n337) );
  CLKBUF_X1 U354 ( .A(n433), .Z(n338) );
  CLKBUF_X1 U355 ( .A(n433), .Z(n339) );
  CLKBUF_X1 U356 ( .A(n433), .Z(n340) );
  CLKBUF_X1 U357 ( .A(n433), .Z(n341) );
  CLKBUF_X1 U358 ( .A(n432), .Z(n342) );
  CLKBUF_X1 U359 ( .A(n432), .Z(n343) );
  CLKBUF_X1 U360 ( .A(n432), .Z(n344) );
  CLKBUF_X1 U361 ( .A(n432), .Z(n345) );
  CLKBUF_X1 U362 ( .A(n432), .Z(n346) );
  CLKBUF_X1 U363 ( .A(n432), .Z(n347) );
  CLKBUF_X1 U364 ( .A(n431), .Z(n348) );
  CLKBUF_X1 U365 ( .A(n431), .Z(n349) );
  CLKBUF_X1 U366 ( .A(n431), .Z(n350) );
  CLKBUF_X1 U367 ( .A(n431), .Z(n351) );
  CLKBUF_X1 U368 ( .A(n431), .Z(n352) );
  CLKBUF_X1 U369 ( .A(n431), .Z(n353) );
  CLKBUF_X1 U370 ( .A(n430), .Z(n354) );
  CLKBUF_X1 U371 ( .A(n430), .Z(n355) );
  CLKBUF_X1 U372 ( .A(n430), .Z(n356) );
  CLKBUF_X1 U373 ( .A(n430), .Z(n357) );
  CLKBUF_X1 U374 ( .A(n430), .Z(n358) );
  CLKBUF_X1 U375 ( .A(n430), .Z(n359) );
  CLKBUF_X1 U376 ( .A(n429), .Z(n360) );
  CLKBUF_X1 U377 ( .A(n429), .Z(n361) );
  CLKBUF_X1 U378 ( .A(n429), .Z(n362) );
  CLKBUF_X1 U379 ( .A(n429), .Z(n363) );
  CLKBUF_X1 U380 ( .A(n429), .Z(n364) );
  CLKBUF_X1 U381 ( .A(n429), .Z(n365) );
  CLKBUF_X1 U382 ( .A(n428), .Z(n366) );
  CLKBUF_X1 U383 ( .A(n428), .Z(n367) );
  CLKBUF_X1 U384 ( .A(n428), .Z(n368) );
  CLKBUF_X1 U385 ( .A(n428), .Z(n369) );
  CLKBUF_X1 U386 ( .A(n428), .Z(n370) );
  CLKBUF_X1 U387 ( .A(n428), .Z(n371) );
  CLKBUF_X1 U388 ( .A(n427), .Z(n372) );
  CLKBUF_X1 U389 ( .A(n427), .Z(n373) );
  CLKBUF_X1 U390 ( .A(n427), .Z(n374) );
  CLKBUF_X1 U391 ( .A(n427), .Z(n375) );
  CLKBUF_X1 U392 ( .A(n427), .Z(n376) );
  CLKBUF_X1 U393 ( .A(n427), .Z(n377) );
  CLKBUF_X1 U394 ( .A(n426), .Z(n378) );
  CLKBUF_X1 U395 ( .A(n426), .Z(n379) );
  CLKBUF_X1 U396 ( .A(n426), .Z(n380) );
  CLKBUF_X1 U397 ( .A(n426), .Z(n381) );
  CLKBUF_X1 U398 ( .A(n426), .Z(n382) );
  CLKBUF_X1 U399 ( .A(n426), .Z(n383) );
  CLKBUF_X1 U400 ( .A(n425), .Z(n384) );
  CLKBUF_X1 U401 ( .A(n425), .Z(n385) );
  CLKBUF_X1 U402 ( .A(n425), .Z(n386) );
  CLKBUF_X1 U403 ( .A(n425), .Z(n387) );
  CLKBUF_X1 U404 ( .A(n425), .Z(n388) );
  CLKBUF_X1 U405 ( .A(n425), .Z(n389) );
  CLKBUF_X1 U406 ( .A(n424), .Z(n390) );
  CLKBUF_X1 U407 ( .A(n424), .Z(n391) );
  CLKBUF_X1 U408 ( .A(n424), .Z(n392) );
  CLKBUF_X1 U409 ( .A(n424), .Z(n393) );
  CLKBUF_X1 U410 ( .A(n424), .Z(n394) );
  CLKBUF_X1 U411 ( .A(n424), .Z(n395) );
  CLKBUF_X1 U412 ( .A(n423), .Z(n396) );
  CLKBUF_X1 U413 ( .A(n423), .Z(n397) );
  CLKBUF_X1 U414 ( .A(n423), .Z(n398) );
  CLKBUF_X1 U415 ( .A(n423), .Z(n399) );
  CLKBUF_X1 U416 ( .A(n423), .Z(n400) );
  CLKBUF_X1 U417 ( .A(n423), .Z(n401) );
  CLKBUF_X1 U418 ( .A(n422), .Z(n402) );
  CLKBUF_X1 U419 ( .A(n422), .Z(n403) );
  CLKBUF_X1 U420 ( .A(n422), .Z(n404) );
  CLKBUF_X1 U421 ( .A(n422), .Z(n405) );
  CLKBUF_X1 U422 ( .A(n422), .Z(n406) );
  CLKBUF_X1 U423 ( .A(n422), .Z(n407) );
  CLKBUF_X1 U424 ( .A(n421), .Z(n408) );
  CLKBUF_X1 U425 ( .A(n421), .Z(n409) );
  CLKBUF_X1 U426 ( .A(n421), .Z(n410) );
  CLKBUF_X1 U427 ( .A(n421), .Z(n411) );
  CLKBUF_X1 U428 ( .A(n421), .Z(n412) );
  CLKBUF_X1 U429 ( .A(n421), .Z(n413) );
  CLKBUF_X1 U430 ( .A(n420), .Z(n414) );
  CLKBUF_X1 U431 ( .A(n420), .Z(n415) );
  CLKBUF_X1 U432 ( .A(n420), .Z(n416) );
  CLKBUF_X1 U433 ( .A(n420), .Z(n417) );
  CLKBUF_X1 U434 ( .A(n420), .Z(n418) );
  INV_X1 U435 ( .A(n434), .ZN(n3865) );
  MUX2_X1 U436 ( .A(n3721), .B(n298), .S(n3), .Z(n434) );
  INV_X1 U437 ( .A(n436), .ZN(n3866) );
  MUX2_X1 U438 ( .A(n3700), .B(n299), .S(n3), .Z(n436) );
  INV_X1 U439 ( .A(n437), .ZN(n3867) );
  MUX2_X1 U440 ( .A(n3679), .B(n300), .S(n3), .Z(n437) );
  INV_X1 U441 ( .A(n438), .ZN(n3868) );
  MUX2_X1 U442 ( .A(n3658), .B(n301), .S(n3), .Z(n438) );
  INV_X1 U443 ( .A(n439), .ZN(n3869) );
  MUX2_X1 U444 ( .A(n3637), .B(n302), .S(n3), .Z(n439) );
  INV_X1 U445 ( .A(n440), .ZN(n3870) );
  MUX2_X1 U446 ( .A(n3616), .B(n303), .S(n3), .Z(n440) );
  INV_X1 U447 ( .A(n441), .ZN(n3871) );
  MUX2_X1 U448 ( .A(n3595), .B(n304), .S(n3), .Z(n441) );
  INV_X1 U449 ( .A(n442), .ZN(n3872) );
  MUX2_X1 U450 ( .A(n3574), .B(n305), .S(n3), .Z(n442) );
  INV_X1 U451 ( .A(n443), .ZN(n3873) );
  MUX2_X1 U452 ( .A(n2977), .B(n306), .S(n2), .Z(n443) );
  INV_X1 U453 ( .A(n444), .ZN(n3874) );
  MUX2_X1 U454 ( .A(n2956), .B(n307), .S(n2), .Z(n444) );
  INV_X1 U455 ( .A(n445), .ZN(n3875) );
  MUX2_X1 U456 ( .A(n2935), .B(n308), .S(n2), .Z(n445) );
  INV_X1 U457 ( .A(n446), .ZN(n3876) );
  MUX2_X1 U458 ( .A(n2914), .B(n309), .S(n2), .Z(n446) );
  INV_X1 U459 ( .A(n447), .ZN(n3877) );
  MUX2_X1 U460 ( .A(n2893), .B(n310), .S(n2), .Z(n447) );
  INV_X1 U461 ( .A(n448), .ZN(n3878) );
  MUX2_X1 U462 ( .A(n2872), .B(n311), .S(n2), .Z(n448) );
  INV_X1 U463 ( .A(n449), .ZN(n3879) );
  MUX2_X1 U464 ( .A(n2851), .B(n312), .S(n2), .Z(n449) );
  INV_X1 U465 ( .A(n450), .ZN(n3880) );
  MUX2_X1 U466 ( .A(n2830), .B(n313), .S(n2), .Z(n450) );
  INV_X1 U467 ( .A(n451), .ZN(n3881) );
  MUX2_X1 U468 ( .A(n2809), .B(n314), .S(n2), .Z(n451) );
  INV_X1 U469 ( .A(n452), .ZN(n3882) );
  MUX2_X1 U470 ( .A(n2788), .B(n315), .S(n2), .Z(n452) );
  INV_X1 U471 ( .A(n453), .ZN(n3883) );
  MUX2_X1 U472 ( .A(n2767), .B(n316), .S(n2), .Z(n453) );
  INV_X1 U473 ( .A(n454), .ZN(n3884) );
  MUX2_X1 U474 ( .A(n2746), .B(n317), .S(n2), .Z(n454) );
  INV_X1 U475 ( .A(n455), .ZN(n3885) );
  MUX2_X1 U476 ( .A(n2725), .B(n318), .S(n1), .Z(n455) );
  INV_X1 U477 ( .A(n456), .ZN(n3886) );
  MUX2_X1 U478 ( .A(n2704), .B(n319), .S(n1), .Z(n456) );
  INV_X1 U479 ( .A(n457), .ZN(n3887) );
  MUX2_X1 U480 ( .A(n2683), .B(n320), .S(n1), .Z(n457) );
  INV_X1 U481 ( .A(n458), .ZN(n3888) );
  MUX2_X1 U482 ( .A(n2662), .B(n321), .S(n1), .Z(n458) );
  INV_X1 U483 ( .A(n459), .ZN(n3889) );
  MUX2_X1 U484 ( .A(n2641), .B(n322), .S(n1), .Z(n459) );
  INV_X1 U485 ( .A(n460), .ZN(n3890) );
  MUX2_X1 U486 ( .A(n2620), .B(n323), .S(n1), .Z(n460) );
  INV_X1 U487 ( .A(n461), .ZN(n3891) );
  MUX2_X1 U488 ( .A(n2599), .B(n324), .S(n1), .Z(n461) );
  INV_X1 U489 ( .A(n462), .ZN(n3892) );
  MUX2_X1 U490 ( .A(n2578), .B(n325), .S(n1), .Z(n462) );
  INV_X1 U491 ( .A(n463), .ZN(n3893) );
  MUX2_X1 U492 ( .A(n2557), .B(n326), .S(n1), .Z(n463) );
  INV_X1 U493 ( .A(n464), .ZN(n3894) );
  MUX2_X1 U494 ( .A(n2536), .B(n327), .S(n1), .Z(n464) );
  INV_X1 U495 ( .A(n465), .ZN(n3895) );
  MUX2_X1 U496 ( .A(n2515), .B(n328), .S(n1), .Z(n465) );
  INV_X1 U497 ( .A(n466), .ZN(n3896) );
  MUX2_X1 U498 ( .A(n2494), .B(n329), .S(n1), .Z(n466) );
  AND2_X1 U499 ( .A1(n467), .A2(n468), .ZN(n435) );
  INV_X1 U500 ( .A(n469), .ZN(n3897) );
  MUX2_X1 U501 ( .A(n3722), .B(n298), .S(n6), .Z(n469) );
  INV_X1 U502 ( .A(n471), .ZN(n3898) );
  MUX2_X1 U503 ( .A(n3701), .B(n299), .S(n6), .Z(n471) );
  INV_X1 U504 ( .A(n472), .ZN(n3899) );
  MUX2_X1 U505 ( .A(n3680), .B(n300), .S(n6), .Z(n472) );
  INV_X1 U506 ( .A(n473), .ZN(n3900) );
  MUX2_X1 U507 ( .A(n3659), .B(n301), .S(n6), .Z(n473) );
  INV_X1 U508 ( .A(n474), .ZN(n3901) );
  MUX2_X1 U509 ( .A(n3638), .B(n302), .S(n6), .Z(n474) );
  INV_X1 U510 ( .A(n475), .ZN(n3902) );
  MUX2_X1 U511 ( .A(n3617), .B(n303), .S(n6), .Z(n475) );
  INV_X1 U512 ( .A(n476), .ZN(n3903) );
  MUX2_X1 U513 ( .A(n3596), .B(n304), .S(n6), .Z(n476) );
  INV_X1 U514 ( .A(n477), .ZN(n3904) );
  MUX2_X1 U515 ( .A(n3575), .B(n305), .S(n6), .Z(n477) );
  INV_X1 U516 ( .A(n478), .ZN(n3905) );
  MUX2_X1 U517 ( .A(n2978), .B(n306), .S(n5), .Z(n478) );
  INV_X1 U518 ( .A(n479), .ZN(n3906) );
  MUX2_X1 U519 ( .A(n2957), .B(n307), .S(n5), .Z(n479) );
  INV_X1 U520 ( .A(n480), .ZN(n3907) );
  MUX2_X1 U521 ( .A(n2936), .B(n308), .S(n5), .Z(n480) );
  INV_X1 U522 ( .A(n481), .ZN(n3908) );
  MUX2_X1 U523 ( .A(n2915), .B(n309), .S(n5), .Z(n481) );
  INV_X1 U524 ( .A(n482), .ZN(n3909) );
  MUX2_X1 U525 ( .A(n2894), .B(n310), .S(n5), .Z(n482) );
  INV_X1 U526 ( .A(n483), .ZN(n3910) );
  MUX2_X1 U527 ( .A(n2873), .B(n311), .S(n5), .Z(n483) );
  INV_X1 U528 ( .A(n484), .ZN(n3911) );
  MUX2_X1 U529 ( .A(n2852), .B(n312), .S(n5), .Z(n484) );
  INV_X1 U530 ( .A(n485), .ZN(n3912) );
  MUX2_X1 U531 ( .A(n2831), .B(n313), .S(n5), .Z(n485) );
  INV_X1 U532 ( .A(n486), .ZN(n3913) );
  MUX2_X1 U533 ( .A(n2810), .B(n314), .S(n5), .Z(n486) );
  INV_X1 U534 ( .A(n487), .ZN(n3914) );
  MUX2_X1 U535 ( .A(n2789), .B(n315), .S(n5), .Z(n487) );
  INV_X1 U536 ( .A(n488), .ZN(n3915) );
  MUX2_X1 U537 ( .A(n2768), .B(n316), .S(n5), .Z(n488) );
  INV_X1 U538 ( .A(n489), .ZN(n3916) );
  MUX2_X1 U539 ( .A(n2747), .B(n317), .S(n5), .Z(n489) );
  INV_X1 U540 ( .A(n490), .ZN(n3917) );
  MUX2_X1 U541 ( .A(n2726), .B(n318), .S(n4), .Z(n490) );
  INV_X1 U542 ( .A(n491), .ZN(n3918) );
  MUX2_X1 U543 ( .A(n2705), .B(n319), .S(n4), .Z(n491) );
  INV_X1 U544 ( .A(n492), .ZN(n3919) );
  MUX2_X1 U545 ( .A(n2684), .B(n320), .S(n4), .Z(n492) );
  INV_X1 U546 ( .A(n493), .ZN(n3920) );
  MUX2_X1 U547 ( .A(n2663), .B(n321), .S(n4), .Z(n493) );
  INV_X1 U548 ( .A(n494), .ZN(n3921) );
  MUX2_X1 U549 ( .A(n2642), .B(n322), .S(n4), .Z(n494) );
  INV_X1 U550 ( .A(n495), .ZN(n3922) );
  MUX2_X1 U551 ( .A(n2621), .B(n323), .S(n4), .Z(n495) );
  INV_X1 U552 ( .A(n496), .ZN(n3923) );
  MUX2_X1 U553 ( .A(n2600), .B(n324), .S(n4), .Z(n496) );
  INV_X1 U554 ( .A(n497), .ZN(n3924) );
  MUX2_X1 U555 ( .A(n2579), .B(n325), .S(n4), .Z(n497) );
  INV_X1 U556 ( .A(n498), .ZN(n3925) );
  MUX2_X1 U557 ( .A(n2558), .B(n326), .S(n4), .Z(n498) );
  INV_X1 U558 ( .A(n499), .ZN(n3926) );
  MUX2_X1 U559 ( .A(n2537), .B(n327), .S(n4), .Z(n499) );
  INV_X1 U560 ( .A(n500), .ZN(n3927) );
  MUX2_X1 U561 ( .A(n2516), .B(n328), .S(n4), .Z(n500) );
  INV_X1 U562 ( .A(n501), .ZN(n3928) );
  MUX2_X1 U563 ( .A(n2495), .B(n329), .S(n4), .Z(n501) );
  AND2_X1 U564 ( .A1(n502), .A2(n467), .ZN(n470) );
  INV_X1 U565 ( .A(n503), .ZN(n3929) );
  MUX2_X1 U566 ( .A(n3717), .B(n298), .S(n9), .Z(n503) );
  INV_X1 U567 ( .A(n505), .ZN(n3930) );
  MUX2_X1 U568 ( .A(n3696), .B(n299), .S(n9), .Z(n505) );
  INV_X1 U569 ( .A(n506), .ZN(n3931) );
  MUX2_X1 U570 ( .A(n3675), .B(n300), .S(n9), .Z(n506) );
  INV_X1 U571 ( .A(n507), .ZN(n3932) );
  MUX2_X1 U572 ( .A(n3654), .B(n301), .S(n9), .Z(n507) );
  INV_X1 U573 ( .A(n508), .ZN(n3933) );
  MUX2_X1 U574 ( .A(n3633), .B(n302), .S(n9), .Z(n508) );
  INV_X1 U575 ( .A(n509), .ZN(n3934) );
  MUX2_X1 U576 ( .A(n3612), .B(n303), .S(n9), .Z(n509) );
  INV_X1 U577 ( .A(n510), .ZN(n3935) );
  MUX2_X1 U578 ( .A(n3591), .B(n304), .S(n9), .Z(n510) );
  INV_X1 U579 ( .A(n511), .ZN(n3936) );
  MUX2_X1 U580 ( .A(n3570), .B(n305), .S(n9), .Z(n511) );
  INV_X1 U581 ( .A(n512), .ZN(n3937) );
  MUX2_X1 U582 ( .A(n2973), .B(n306), .S(n8), .Z(n512) );
  INV_X1 U583 ( .A(n513), .ZN(n3938) );
  MUX2_X1 U584 ( .A(n2952), .B(n307), .S(n8), .Z(n513) );
  INV_X1 U585 ( .A(n514), .ZN(n3939) );
  MUX2_X1 U586 ( .A(n2931), .B(n308), .S(n8), .Z(n514) );
  INV_X1 U587 ( .A(n515), .ZN(n3940) );
  MUX2_X1 U588 ( .A(n2910), .B(n309), .S(n8), .Z(n515) );
  INV_X1 U589 ( .A(n516), .ZN(n3941) );
  MUX2_X1 U590 ( .A(n2889), .B(n310), .S(n8), .Z(n516) );
  INV_X1 U591 ( .A(n517), .ZN(n3942) );
  MUX2_X1 U592 ( .A(n2868), .B(n311), .S(n8), .Z(n517) );
  INV_X1 U593 ( .A(n518), .ZN(n3943) );
  MUX2_X1 U594 ( .A(n2847), .B(n312), .S(n8), .Z(n518) );
  INV_X1 U595 ( .A(n519), .ZN(n3944) );
  MUX2_X1 U596 ( .A(n2826), .B(n313), .S(n8), .Z(n519) );
  INV_X1 U597 ( .A(n520), .ZN(n3945) );
  MUX2_X1 U598 ( .A(n2805), .B(n314), .S(n8), .Z(n520) );
  INV_X1 U599 ( .A(n521), .ZN(n3946) );
  MUX2_X1 U600 ( .A(n2784), .B(n315), .S(n8), .Z(n521) );
  INV_X1 U601 ( .A(n522), .ZN(n3947) );
  MUX2_X1 U602 ( .A(n2763), .B(n316), .S(n8), .Z(n522) );
  INV_X1 U603 ( .A(n523), .ZN(n3948) );
  MUX2_X1 U604 ( .A(n2742), .B(n317), .S(n8), .Z(n523) );
  INV_X1 U605 ( .A(n524), .ZN(n3949) );
  MUX2_X1 U606 ( .A(n2721), .B(n318), .S(n7), .Z(n524) );
  INV_X1 U607 ( .A(n525), .ZN(n3950) );
  MUX2_X1 U608 ( .A(n2700), .B(n319), .S(n7), .Z(n525) );
  INV_X1 U609 ( .A(n526), .ZN(n3951) );
  MUX2_X1 U610 ( .A(n2679), .B(n320), .S(n7), .Z(n526) );
  INV_X1 U611 ( .A(n527), .ZN(n3952) );
  MUX2_X1 U612 ( .A(n2658), .B(n321), .S(n7), .Z(n527) );
  INV_X1 U613 ( .A(n528), .ZN(n3953) );
  MUX2_X1 U614 ( .A(n2637), .B(n322), .S(n7), .Z(n528) );
  INV_X1 U615 ( .A(n529), .ZN(n3954) );
  MUX2_X1 U616 ( .A(n2616), .B(n323), .S(n7), .Z(n529) );
  INV_X1 U617 ( .A(n530), .ZN(n3955) );
  MUX2_X1 U618 ( .A(n2595), .B(n324), .S(n7), .Z(n530) );
  INV_X1 U619 ( .A(n531), .ZN(n3956) );
  MUX2_X1 U620 ( .A(n2574), .B(n325), .S(n7), .Z(n531) );
  INV_X1 U621 ( .A(n532), .ZN(n3957) );
  MUX2_X1 U622 ( .A(n2553), .B(n326), .S(n7), .Z(n532) );
  INV_X1 U623 ( .A(n533), .ZN(n3958) );
  MUX2_X1 U624 ( .A(n2532), .B(n327), .S(n7), .Z(n533) );
  INV_X1 U625 ( .A(n534), .ZN(n3959) );
  MUX2_X1 U626 ( .A(n2511), .B(n328), .S(n7), .Z(n534) );
  INV_X1 U627 ( .A(n535), .ZN(n3960) );
  MUX2_X1 U628 ( .A(n2490), .B(n329), .S(n7), .Z(n535) );
  AND2_X1 U629 ( .A1(n536), .A2(n467), .ZN(n504) );
  INV_X1 U630 ( .A(n537), .ZN(n3961) );
  MUX2_X1 U631 ( .A(n3718), .B(n298), .S(n12), .Z(n537) );
  INV_X1 U632 ( .A(n539), .ZN(n3962) );
  MUX2_X1 U633 ( .A(n3697), .B(n299), .S(n12), .Z(n539) );
  INV_X1 U634 ( .A(n540), .ZN(n3963) );
  MUX2_X1 U635 ( .A(n3676), .B(n300), .S(n12), .Z(n540) );
  INV_X1 U636 ( .A(n541), .ZN(n3964) );
  MUX2_X1 U637 ( .A(n3655), .B(n301), .S(n12), .Z(n541) );
  INV_X1 U638 ( .A(n542), .ZN(n3965) );
  MUX2_X1 U639 ( .A(n3634), .B(n302), .S(n12), .Z(n542) );
  INV_X1 U640 ( .A(n543), .ZN(n3966) );
  MUX2_X1 U641 ( .A(n3613), .B(n303), .S(n12), .Z(n543) );
  INV_X1 U642 ( .A(n544), .ZN(n3967) );
  MUX2_X1 U643 ( .A(n3592), .B(n304), .S(n12), .Z(n544) );
  INV_X1 U644 ( .A(n545), .ZN(n3968) );
  MUX2_X1 U645 ( .A(n3571), .B(n305), .S(n12), .Z(n545) );
  INV_X1 U646 ( .A(n546), .ZN(n3969) );
  MUX2_X1 U647 ( .A(n2974), .B(n306), .S(n11), .Z(n546) );
  INV_X1 U648 ( .A(n547), .ZN(n3970) );
  MUX2_X1 U649 ( .A(n2953), .B(n307), .S(n11), .Z(n547) );
  INV_X1 U650 ( .A(n548), .ZN(n3971) );
  MUX2_X1 U651 ( .A(n2932), .B(n308), .S(n11), .Z(n548) );
  INV_X1 U652 ( .A(n549), .ZN(n3972) );
  MUX2_X1 U653 ( .A(n2911), .B(n309), .S(n11), .Z(n549) );
  INV_X1 U654 ( .A(n550), .ZN(n3973) );
  MUX2_X1 U655 ( .A(n2890), .B(n310), .S(n11), .Z(n550) );
  INV_X1 U656 ( .A(n551), .ZN(n3974) );
  MUX2_X1 U657 ( .A(n2869), .B(n311), .S(n11), .Z(n551) );
  INV_X1 U658 ( .A(n552), .ZN(n3975) );
  MUX2_X1 U659 ( .A(n2848), .B(n312), .S(n11), .Z(n552) );
  INV_X1 U660 ( .A(n553), .ZN(n3976) );
  MUX2_X1 U661 ( .A(n2827), .B(n313), .S(n11), .Z(n553) );
  INV_X1 U662 ( .A(n554), .ZN(n3977) );
  MUX2_X1 U663 ( .A(n2806), .B(n314), .S(n11), .Z(n554) );
  INV_X1 U664 ( .A(n555), .ZN(n3978) );
  MUX2_X1 U665 ( .A(n2785), .B(n315), .S(n11), .Z(n555) );
  INV_X1 U666 ( .A(n556), .ZN(n3979) );
  MUX2_X1 U667 ( .A(n2764), .B(n316), .S(n11), .Z(n556) );
  INV_X1 U668 ( .A(n557), .ZN(n3980) );
  MUX2_X1 U669 ( .A(n2743), .B(n317), .S(n11), .Z(n557) );
  INV_X1 U670 ( .A(n558), .ZN(n3981) );
  MUX2_X1 U671 ( .A(n2722), .B(n318), .S(n10), .Z(n558) );
  INV_X1 U672 ( .A(n559), .ZN(n3982) );
  MUX2_X1 U673 ( .A(n2701), .B(n319), .S(n10), .Z(n559) );
  INV_X1 U674 ( .A(n560), .ZN(n3983) );
  MUX2_X1 U675 ( .A(n2680), .B(n320), .S(n10), .Z(n560) );
  INV_X1 U676 ( .A(n561), .ZN(n3984) );
  MUX2_X1 U677 ( .A(n2659), .B(n321), .S(n10), .Z(n561) );
  INV_X1 U678 ( .A(n562), .ZN(n3985) );
  MUX2_X1 U679 ( .A(n2638), .B(n322), .S(n10), .Z(n562) );
  INV_X1 U680 ( .A(n563), .ZN(n3986) );
  MUX2_X1 U681 ( .A(n2617), .B(n323), .S(n10), .Z(n563) );
  INV_X1 U682 ( .A(n564), .ZN(n3987) );
  MUX2_X1 U683 ( .A(n2596), .B(n324), .S(n10), .Z(n564) );
  INV_X1 U684 ( .A(n565), .ZN(n3988) );
  MUX2_X1 U685 ( .A(n2575), .B(n325), .S(n10), .Z(n565) );
  INV_X1 U686 ( .A(n566), .ZN(n3989) );
  MUX2_X1 U687 ( .A(n2554), .B(n326), .S(n10), .Z(n566) );
  INV_X1 U688 ( .A(n567), .ZN(n3990) );
  MUX2_X1 U689 ( .A(n2533), .B(n327), .S(n10), .Z(n567) );
  INV_X1 U690 ( .A(n568), .ZN(n3991) );
  MUX2_X1 U691 ( .A(n2512), .B(n328), .S(n10), .Z(n568) );
  INV_X1 U692 ( .A(n569), .ZN(n3992) );
  MUX2_X1 U693 ( .A(n2491), .B(n329), .S(n10), .Z(n569) );
  AND2_X1 U694 ( .A1(n570), .A2(n467), .ZN(n538) );
  MUX2_X1 U695 ( .A(n571), .B(DATAIN[0]), .S(n15), .Z(n3993) );
  MUX2_X1 U696 ( .A(n573), .B(DATAIN[1]), .S(n15), .Z(n3994) );
  MUX2_X1 U697 ( .A(n574), .B(DATAIN[2]), .S(n15), .Z(n3995) );
  MUX2_X1 U698 ( .A(n575), .B(DATAIN[3]), .S(n15), .Z(n3996) );
  MUX2_X1 U699 ( .A(n576), .B(DATAIN[4]), .S(n15), .Z(n3997) );
  MUX2_X1 U700 ( .A(n577), .B(DATAIN[5]), .S(n15), .Z(n3998) );
  MUX2_X1 U701 ( .A(n578), .B(DATAIN[6]), .S(n15), .Z(n3999) );
  MUX2_X1 U702 ( .A(n579), .B(DATAIN[7]), .S(n15), .Z(n4000) );
  MUX2_X1 U703 ( .A(n580), .B(DATAIN[8]), .S(n14), .Z(n4001) );
  MUX2_X1 U704 ( .A(n581), .B(DATAIN[9]), .S(n14), .Z(n4002) );
  MUX2_X1 U705 ( .A(n582), .B(DATAIN[10]), .S(n14), .Z(n4003) );
  MUX2_X1 U706 ( .A(n583), .B(DATAIN[11]), .S(n14), .Z(n4004) );
  MUX2_X1 U707 ( .A(n584), .B(DATAIN[12]), .S(n14), .Z(n4005) );
  MUX2_X1 U708 ( .A(n585), .B(DATAIN[13]), .S(n14), .Z(n4006) );
  MUX2_X1 U709 ( .A(n586), .B(DATAIN[14]), .S(n14), .Z(n4007) );
  MUX2_X1 U710 ( .A(n587), .B(DATAIN[15]), .S(n14), .Z(n4008) );
  MUX2_X1 U711 ( .A(n588), .B(DATAIN[16]), .S(n14), .Z(n4009) );
  MUX2_X1 U712 ( .A(n589), .B(DATAIN[17]), .S(n14), .Z(n4010) );
  MUX2_X1 U713 ( .A(n590), .B(DATAIN[18]), .S(n14), .Z(n4011) );
  MUX2_X1 U714 ( .A(n591), .B(DATAIN[19]), .S(n14), .Z(n4012) );
  MUX2_X1 U715 ( .A(n592), .B(DATAIN[20]), .S(n13), .Z(n4013) );
  MUX2_X1 U716 ( .A(n593), .B(DATAIN[21]), .S(n13), .Z(n4014) );
  MUX2_X1 U717 ( .A(n594), .B(DATAIN[22]), .S(n13), .Z(n4015) );
  MUX2_X1 U718 ( .A(n595), .B(DATAIN[23]), .S(n13), .Z(n4016) );
  MUX2_X1 U719 ( .A(n596), .B(DATAIN[24]), .S(n13), .Z(n4017) );
  MUX2_X1 U720 ( .A(n597), .B(DATAIN[25]), .S(n13), .Z(n4018) );
  MUX2_X1 U721 ( .A(n598), .B(DATAIN[26]), .S(n13), .Z(n4019) );
  MUX2_X1 U722 ( .A(n599), .B(DATAIN[27]), .S(n13), .Z(n4020) );
  MUX2_X1 U723 ( .A(n600), .B(DATAIN[28]), .S(n13), .Z(n4021) );
  MUX2_X1 U724 ( .A(n601), .B(DATAIN[29]), .S(n13), .Z(n4022) );
  MUX2_X1 U725 ( .A(n602), .B(DATAIN[30]), .S(n13), .Z(n4023) );
  MUX2_X1 U726 ( .A(n603), .B(DATAIN[31]), .S(n13), .Z(n4024) );
  AND2_X1 U727 ( .A1(n604), .A2(n502), .ZN(n572) );
  MUX2_X1 U728 ( .A(n605), .B(DATAIN[0]), .S(n18), .Z(n4025) );
  MUX2_X1 U729 ( .A(n607), .B(DATAIN[1]), .S(n18), .Z(n4026) );
  MUX2_X1 U730 ( .A(n608), .B(DATAIN[2]), .S(n18), .Z(n4027) );
  MUX2_X1 U731 ( .A(n609), .B(DATAIN[3]), .S(n18), .Z(n4028) );
  MUX2_X1 U732 ( .A(n610), .B(DATAIN[4]), .S(n18), .Z(n4029) );
  MUX2_X1 U733 ( .A(n611), .B(DATAIN[5]), .S(n18), .Z(n4030) );
  MUX2_X1 U734 ( .A(n612), .B(DATAIN[6]), .S(n18), .Z(n4031) );
  MUX2_X1 U735 ( .A(n613), .B(DATAIN[7]), .S(n18), .Z(n4032) );
  MUX2_X1 U736 ( .A(n614), .B(DATAIN[8]), .S(n17), .Z(n4033) );
  MUX2_X1 U737 ( .A(n615), .B(DATAIN[9]), .S(n17), .Z(n4034) );
  MUX2_X1 U738 ( .A(n616), .B(DATAIN[10]), .S(n17), .Z(n4035) );
  MUX2_X1 U739 ( .A(n617), .B(DATAIN[11]), .S(n17), .Z(n4036) );
  MUX2_X1 U740 ( .A(n618), .B(DATAIN[12]), .S(n17), .Z(n4037) );
  MUX2_X1 U741 ( .A(n619), .B(DATAIN[13]), .S(n17), .Z(n4038) );
  MUX2_X1 U742 ( .A(n620), .B(DATAIN[14]), .S(n17), .Z(n4039) );
  MUX2_X1 U743 ( .A(n621), .B(DATAIN[15]), .S(n17), .Z(n4040) );
  MUX2_X1 U744 ( .A(n622), .B(DATAIN[16]), .S(n17), .Z(n4041) );
  MUX2_X1 U745 ( .A(n623), .B(DATAIN[17]), .S(n17), .Z(n4042) );
  MUX2_X1 U746 ( .A(n624), .B(DATAIN[18]), .S(n17), .Z(n4043) );
  MUX2_X1 U747 ( .A(n625), .B(DATAIN[19]), .S(n17), .Z(n4044) );
  MUX2_X1 U748 ( .A(n626), .B(DATAIN[20]), .S(n16), .Z(n4045) );
  MUX2_X1 U749 ( .A(n627), .B(DATAIN[21]), .S(n16), .Z(n4046) );
  MUX2_X1 U750 ( .A(n628), .B(DATAIN[22]), .S(n16), .Z(n4047) );
  MUX2_X1 U751 ( .A(n629), .B(DATAIN[23]), .S(n16), .Z(n4048) );
  MUX2_X1 U752 ( .A(n630), .B(DATAIN[24]), .S(n16), .Z(n4049) );
  MUX2_X1 U753 ( .A(n631), .B(DATAIN[25]), .S(n16), .Z(n4050) );
  MUX2_X1 U754 ( .A(n632), .B(DATAIN[26]), .S(n16), .Z(n4051) );
  MUX2_X1 U755 ( .A(n633), .B(DATAIN[27]), .S(n16), .Z(n4052) );
  MUX2_X1 U756 ( .A(n634), .B(DATAIN[28]), .S(n16), .Z(n4053) );
  MUX2_X1 U757 ( .A(n635), .B(DATAIN[29]), .S(n16), .Z(n4054) );
  MUX2_X1 U758 ( .A(n636), .B(DATAIN[30]), .S(n16), .Z(n4055) );
  MUX2_X1 U759 ( .A(n637), .B(DATAIN[31]), .S(n16), .Z(n4056) );
  AND2_X1 U760 ( .A1(n604), .A2(n536), .ZN(n606) );
  MUX2_X1 U761 ( .A(n638), .B(DATAIN[0]), .S(n21), .Z(n4057) );
  MUX2_X1 U762 ( .A(n640), .B(DATAIN[1]), .S(n21), .Z(n4058) );
  MUX2_X1 U763 ( .A(n641), .B(DATAIN[2]), .S(n21), .Z(n4059) );
  MUX2_X1 U764 ( .A(n642), .B(DATAIN[3]), .S(n21), .Z(n4060) );
  MUX2_X1 U765 ( .A(n643), .B(DATAIN[4]), .S(n21), .Z(n4061) );
  MUX2_X1 U766 ( .A(n644), .B(DATAIN[5]), .S(n21), .Z(n4062) );
  MUX2_X1 U767 ( .A(n645), .B(DATAIN[6]), .S(n21), .Z(n4063) );
  MUX2_X1 U768 ( .A(n646), .B(DATAIN[7]), .S(n21), .Z(n4064) );
  MUX2_X1 U769 ( .A(n647), .B(DATAIN[8]), .S(n20), .Z(n4065) );
  MUX2_X1 U770 ( .A(n648), .B(DATAIN[9]), .S(n20), .Z(n4066) );
  MUX2_X1 U771 ( .A(n649), .B(DATAIN[10]), .S(n20), .Z(n4067) );
  MUX2_X1 U772 ( .A(n650), .B(DATAIN[11]), .S(n20), .Z(n4068) );
  MUX2_X1 U773 ( .A(n651), .B(DATAIN[12]), .S(n20), .Z(n4069) );
  MUX2_X1 U774 ( .A(n652), .B(DATAIN[13]), .S(n20), .Z(n4070) );
  MUX2_X1 U775 ( .A(n653), .B(DATAIN[14]), .S(n20), .Z(n4071) );
  MUX2_X1 U776 ( .A(n654), .B(DATAIN[15]), .S(n20), .Z(n4072) );
  MUX2_X1 U777 ( .A(n655), .B(DATAIN[16]), .S(n20), .Z(n4073) );
  MUX2_X1 U778 ( .A(n656), .B(DATAIN[17]), .S(n20), .Z(n4074) );
  MUX2_X1 U779 ( .A(n657), .B(DATAIN[18]), .S(n20), .Z(n4075) );
  MUX2_X1 U780 ( .A(n658), .B(DATAIN[19]), .S(n20), .Z(n4076) );
  MUX2_X1 U781 ( .A(n659), .B(DATAIN[20]), .S(n19), .Z(n4077) );
  MUX2_X1 U782 ( .A(n660), .B(DATAIN[21]), .S(n19), .Z(n4078) );
  MUX2_X1 U783 ( .A(n661), .B(DATAIN[22]), .S(n19), .Z(n4079) );
  MUX2_X1 U784 ( .A(n662), .B(DATAIN[23]), .S(n19), .Z(n4080) );
  MUX2_X1 U785 ( .A(n663), .B(DATAIN[24]), .S(n19), .Z(n4081) );
  MUX2_X1 U786 ( .A(n664), .B(DATAIN[25]), .S(n19), .Z(n4082) );
  MUX2_X1 U787 ( .A(n665), .B(DATAIN[26]), .S(n19), .Z(n4083) );
  MUX2_X1 U788 ( .A(n666), .B(DATAIN[27]), .S(n19), .Z(n4084) );
  MUX2_X1 U789 ( .A(n667), .B(DATAIN[28]), .S(n19), .Z(n4085) );
  MUX2_X1 U790 ( .A(n668), .B(DATAIN[29]), .S(n19), .Z(n4086) );
  MUX2_X1 U791 ( .A(n669), .B(DATAIN[30]), .S(n19), .Z(n4087) );
  MUX2_X1 U792 ( .A(n670), .B(DATAIN[31]), .S(n19), .Z(n4088) );
  AND2_X1 U793 ( .A1(n604), .A2(n570), .ZN(n639) );
  MUX2_X1 U794 ( .A(n671), .B(DATAIN[31]), .S(n24), .Z(n4089) );
  MUX2_X1 U795 ( .A(n673), .B(DATAIN[0]), .S(n24), .Z(n4090) );
  MUX2_X1 U796 ( .A(n674), .B(DATAIN[1]), .S(n24), .Z(n4091) );
  MUX2_X1 U797 ( .A(n675), .B(DATAIN[2]), .S(n24), .Z(n4092) );
  MUX2_X1 U798 ( .A(n676), .B(DATAIN[3]), .S(n24), .Z(n4093) );
  MUX2_X1 U799 ( .A(n677), .B(DATAIN[4]), .S(n24), .Z(n4094) );
  MUX2_X1 U800 ( .A(n678), .B(DATAIN[5]), .S(n24), .Z(n4095) );
  MUX2_X1 U801 ( .A(n679), .B(DATAIN[6]), .S(n24), .Z(n4096) );
  MUX2_X1 U802 ( .A(n680), .B(DATAIN[7]), .S(n23), .Z(n4097) );
  MUX2_X1 U803 ( .A(n681), .B(DATAIN[8]), .S(n23), .Z(n4098) );
  MUX2_X1 U804 ( .A(n682), .B(DATAIN[9]), .S(n23), .Z(n4099) );
  MUX2_X1 U805 ( .A(n683), .B(DATAIN[10]), .S(n23), .Z(n4100) );
  MUX2_X1 U806 ( .A(n684), .B(DATAIN[11]), .S(n23), .Z(n4101) );
  MUX2_X1 U807 ( .A(n685), .B(DATAIN[12]), .S(n23), .Z(n4102) );
  MUX2_X1 U808 ( .A(n686), .B(DATAIN[13]), .S(n23), .Z(n4103) );
  MUX2_X1 U809 ( .A(n687), .B(DATAIN[14]), .S(n23), .Z(n4104) );
  MUX2_X1 U810 ( .A(n688), .B(DATAIN[15]), .S(n23), .Z(n4105) );
  MUX2_X1 U811 ( .A(n689), .B(DATAIN[16]), .S(n23), .Z(n4106) );
  MUX2_X1 U812 ( .A(n690), .B(DATAIN[17]), .S(n23), .Z(n4107) );
  MUX2_X1 U813 ( .A(n691), .B(DATAIN[18]), .S(n23), .Z(n4108) );
  MUX2_X1 U814 ( .A(n692), .B(DATAIN[19]), .S(n22), .Z(n4109) );
  MUX2_X1 U815 ( .A(n693), .B(DATAIN[20]), .S(n22), .Z(n4110) );
  MUX2_X1 U816 ( .A(n694), .B(DATAIN[21]), .S(n22), .Z(n4111) );
  MUX2_X1 U817 ( .A(n695), .B(DATAIN[22]), .S(n22), .Z(n4112) );
  MUX2_X1 U818 ( .A(n696), .B(DATAIN[23]), .S(n22), .Z(n4113) );
  MUX2_X1 U819 ( .A(n697), .B(DATAIN[24]), .S(n22), .Z(n4114) );
  MUX2_X1 U820 ( .A(n698), .B(DATAIN[25]), .S(n22), .Z(n4115) );
  MUX2_X1 U821 ( .A(n699), .B(DATAIN[26]), .S(n22), .Z(n4116) );
  MUX2_X1 U822 ( .A(n700), .B(DATAIN[27]), .S(n22), .Z(n4117) );
  MUX2_X1 U823 ( .A(n701), .B(DATAIN[28]), .S(n22), .Z(n4118) );
  MUX2_X1 U824 ( .A(n702), .B(DATAIN[29]), .S(n22), .Z(n4119) );
  MUX2_X1 U825 ( .A(n703), .B(DATAIN[30]), .S(n22), .Z(n4120) );
  AND2_X1 U826 ( .A1(n704), .A2(n705), .ZN(n672) );
  INV_X1 U827 ( .A(n706), .ZN(n4121) );
  MUX2_X1 U828 ( .A(n3833), .B(n298), .S(n27), .Z(n706) );
  INV_X1 U829 ( .A(n708), .ZN(n4122) );
  MUX2_X1 U830 ( .A(n3834), .B(n299), .S(n27), .Z(n708) );
  INV_X1 U831 ( .A(n709), .ZN(n4123) );
  MUX2_X1 U832 ( .A(n3835), .B(n300), .S(n27), .Z(n709) );
  INV_X1 U833 ( .A(n710), .ZN(n4124) );
  MUX2_X1 U834 ( .A(n3836), .B(n301), .S(n27), .Z(n710) );
  INV_X1 U835 ( .A(n711), .ZN(n4125) );
  MUX2_X1 U836 ( .A(n3837), .B(n302), .S(n27), .Z(n711) );
  INV_X1 U837 ( .A(n712), .ZN(n4126) );
  MUX2_X1 U838 ( .A(n3838), .B(n303), .S(n27), .Z(n712) );
  INV_X1 U839 ( .A(n713), .ZN(n4127) );
  MUX2_X1 U840 ( .A(n3839), .B(n304), .S(n27), .Z(n713) );
  INV_X1 U841 ( .A(n714), .ZN(n4128) );
  MUX2_X1 U842 ( .A(n3840), .B(n305), .S(n27), .Z(n714) );
  INV_X1 U843 ( .A(n715), .ZN(n4129) );
  MUX2_X1 U844 ( .A(n3841), .B(n306), .S(n26), .Z(n715) );
  INV_X1 U845 ( .A(n716), .ZN(n4130) );
  MUX2_X1 U846 ( .A(n3842), .B(n307), .S(n26), .Z(n716) );
  INV_X1 U847 ( .A(n717), .ZN(n4131) );
  MUX2_X1 U848 ( .A(n3843), .B(n308), .S(n26), .Z(n717) );
  INV_X1 U849 ( .A(n718), .ZN(n4132) );
  MUX2_X1 U850 ( .A(n3844), .B(n309), .S(n26), .Z(n718) );
  INV_X1 U851 ( .A(n719), .ZN(n4133) );
  MUX2_X1 U852 ( .A(n3845), .B(n310), .S(n26), .Z(n719) );
  INV_X1 U853 ( .A(n720), .ZN(n4134) );
  MUX2_X1 U854 ( .A(n3846), .B(n311), .S(n26), .Z(n720) );
  INV_X1 U855 ( .A(n721), .ZN(n4135) );
  MUX2_X1 U856 ( .A(n3847), .B(n312), .S(n26), .Z(n721) );
  INV_X1 U857 ( .A(n722), .ZN(n4136) );
  MUX2_X1 U858 ( .A(n3848), .B(n313), .S(n26), .Z(n722) );
  INV_X1 U859 ( .A(n723), .ZN(n4137) );
  MUX2_X1 U860 ( .A(n3849), .B(n314), .S(n26), .Z(n723) );
  INV_X1 U861 ( .A(n724), .ZN(n4138) );
  MUX2_X1 U862 ( .A(n3850), .B(n315), .S(n26), .Z(n724) );
  INV_X1 U863 ( .A(n725), .ZN(n4139) );
  MUX2_X1 U864 ( .A(n3851), .B(n316), .S(n26), .Z(n725) );
  INV_X1 U865 ( .A(n726), .ZN(n4140) );
  MUX2_X1 U866 ( .A(n3852), .B(n317), .S(n26), .Z(n726) );
  INV_X1 U867 ( .A(n727), .ZN(n4141) );
  MUX2_X1 U868 ( .A(n3853), .B(n318), .S(n25), .Z(n727) );
  INV_X1 U869 ( .A(n728), .ZN(n4142) );
  MUX2_X1 U870 ( .A(n3854), .B(n319), .S(n25), .Z(n728) );
  INV_X1 U871 ( .A(n729), .ZN(n4143) );
  MUX2_X1 U872 ( .A(n3855), .B(n320), .S(n25), .Z(n729) );
  INV_X1 U873 ( .A(n730), .ZN(n4144) );
  MUX2_X1 U874 ( .A(n3856), .B(n321), .S(n25), .Z(n730) );
  INV_X1 U875 ( .A(n731), .ZN(n4145) );
  MUX2_X1 U876 ( .A(n3857), .B(n322), .S(n25), .Z(n731) );
  INV_X1 U877 ( .A(n732), .ZN(n4146) );
  MUX2_X1 U878 ( .A(n3858), .B(n323), .S(n25), .Z(n732) );
  INV_X1 U879 ( .A(n733), .ZN(n4147) );
  MUX2_X1 U880 ( .A(n3859), .B(n324), .S(n25), .Z(n733) );
  INV_X1 U881 ( .A(n734), .ZN(n4148) );
  MUX2_X1 U882 ( .A(n3860), .B(n325), .S(n25), .Z(n734) );
  INV_X1 U883 ( .A(n735), .ZN(n4149) );
  MUX2_X1 U884 ( .A(n3861), .B(n326), .S(n25), .Z(n735) );
  INV_X1 U885 ( .A(n736), .ZN(n4150) );
  MUX2_X1 U886 ( .A(n3862), .B(n327), .S(n25), .Z(n736) );
  INV_X1 U887 ( .A(n737), .ZN(n4151) );
  MUX2_X1 U888 ( .A(n3863), .B(n328), .S(n25), .Z(n737) );
  INV_X1 U889 ( .A(n738), .ZN(n4152) );
  MUX2_X1 U890 ( .A(n3864), .B(n329), .S(n25), .Z(n738) );
  AND2_X1 U891 ( .A1(n739), .A2(n704), .ZN(n707) );
  INV_X1 U892 ( .A(n740), .ZN(n4153) );
  MUX2_X1 U893 ( .A(n3737), .B(n298), .S(n30), .Z(n740) );
  INV_X1 U894 ( .A(n742), .ZN(n4154) );
  MUX2_X1 U895 ( .A(n3738), .B(n299), .S(n30), .Z(n742) );
  INV_X1 U896 ( .A(n743), .ZN(n4155) );
  MUX2_X1 U897 ( .A(n3739), .B(n300), .S(n30), .Z(n743) );
  INV_X1 U898 ( .A(n744), .ZN(n4156) );
  MUX2_X1 U899 ( .A(n3740), .B(n301), .S(n30), .Z(n744) );
  INV_X1 U900 ( .A(n745), .ZN(n4157) );
  MUX2_X1 U901 ( .A(n3741), .B(n302), .S(n30), .Z(n745) );
  INV_X1 U902 ( .A(n746), .ZN(n4158) );
  MUX2_X1 U903 ( .A(n3742), .B(n303), .S(n30), .Z(n746) );
  INV_X1 U904 ( .A(n747), .ZN(n4159) );
  MUX2_X1 U905 ( .A(n3743), .B(n304), .S(n30), .Z(n747) );
  INV_X1 U906 ( .A(n748), .ZN(n4160) );
  MUX2_X1 U907 ( .A(n3744), .B(n305), .S(n30), .Z(n748) );
  INV_X1 U908 ( .A(n749), .ZN(n4161) );
  MUX2_X1 U909 ( .A(n3745), .B(n306), .S(n29), .Z(n749) );
  INV_X1 U910 ( .A(n750), .ZN(n4162) );
  MUX2_X1 U911 ( .A(n3746), .B(n307), .S(n29), .Z(n750) );
  INV_X1 U912 ( .A(n751), .ZN(n4163) );
  MUX2_X1 U913 ( .A(n3747), .B(n308), .S(n29), .Z(n751) );
  INV_X1 U914 ( .A(n752), .ZN(n4164) );
  MUX2_X1 U915 ( .A(n3748), .B(n309), .S(n29), .Z(n752) );
  INV_X1 U916 ( .A(n753), .ZN(n4165) );
  MUX2_X1 U917 ( .A(n3749), .B(n310), .S(n29), .Z(n753) );
  INV_X1 U918 ( .A(n754), .ZN(n4166) );
  MUX2_X1 U919 ( .A(n3750), .B(n311), .S(n29), .Z(n754) );
  INV_X1 U920 ( .A(n755), .ZN(n4167) );
  MUX2_X1 U921 ( .A(n3751), .B(n312), .S(n29), .Z(n755) );
  INV_X1 U922 ( .A(n756), .ZN(n4168) );
  MUX2_X1 U923 ( .A(n3752), .B(n313), .S(n29), .Z(n756) );
  INV_X1 U924 ( .A(n757), .ZN(n4169) );
  MUX2_X1 U925 ( .A(n3753), .B(n314), .S(n29), .Z(n757) );
  INV_X1 U926 ( .A(n758), .ZN(n4170) );
  MUX2_X1 U927 ( .A(n3754), .B(n315), .S(n29), .Z(n758) );
  INV_X1 U928 ( .A(n759), .ZN(n4171) );
  MUX2_X1 U929 ( .A(n3755), .B(n316), .S(n29), .Z(n759) );
  INV_X1 U930 ( .A(n760), .ZN(n4172) );
  MUX2_X1 U931 ( .A(n3756), .B(n317), .S(n29), .Z(n760) );
  INV_X1 U932 ( .A(n761), .ZN(n4173) );
  MUX2_X1 U933 ( .A(n3757), .B(n318), .S(n28), .Z(n761) );
  INV_X1 U934 ( .A(n762), .ZN(n4174) );
  MUX2_X1 U935 ( .A(n3758), .B(n319), .S(n28), .Z(n762) );
  INV_X1 U936 ( .A(n763), .ZN(n4175) );
  MUX2_X1 U937 ( .A(n3759), .B(n320), .S(n28), .Z(n763) );
  INV_X1 U938 ( .A(n764), .ZN(n4176) );
  MUX2_X1 U939 ( .A(n3760), .B(n321), .S(n28), .Z(n764) );
  INV_X1 U940 ( .A(n765), .ZN(n4177) );
  MUX2_X1 U941 ( .A(n3761), .B(n322), .S(n28), .Z(n765) );
  INV_X1 U942 ( .A(n766), .ZN(n4178) );
  MUX2_X1 U943 ( .A(n3762), .B(n323), .S(n28), .Z(n766) );
  INV_X1 U944 ( .A(n767), .ZN(n4179) );
  MUX2_X1 U945 ( .A(n3763), .B(n324), .S(n28), .Z(n767) );
  INV_X1 U946 ( .A(n768), .ZN(n4180) );
  MUX2_X1 U947 ( .A(n3764), .B(n325), .S(n28), .Z(n768) );
  INV_X1 U948 ( .A(n769), .ZN(n4181) );
  MUX2_X1 U949 ( .A(n3765), .B(n326), .S(n28), .Z(n769) );
  INV_X1 U950 ( .A(n770), .ZN(n4182) );
  MUX2_X1 U951 ( .A(n3766), .B(n327), .S(n28), .Z(n770) );
  INV_X1 U952 ( .A(n771), .ZN(n4183) );
  MUX2_X1 U953 ( .A(n3767), .B(n328), .S(n28), .Z(n771) );
  INV_X1 U954 ( .A(n772), .ZN(n4184) );
  MUX2_X1 U955 ( .A(n3768), .B(n329), .S(n28), .Z(n772) );
  AND2_X1 U956 ( .A1(n773), .A2(n704), .ZN(n741) );
  MUX2_X1 U957 ( .A(n774), .B(DATAIN[0]), .S(n33), .Z(n4185) );
  MUX2_X1 U958 ( .A(n776), .B(DATAIN[1]), .S(n33), .Z(n4186) );
  MUX2_X1 U959 ( .A(n777), .B(DATAIN[2]), .S(n33), .Z(n4187) );
  MUX2_X1 U960 ( .A(n778), .B(DATAIN[3]), .S(n33), .Z(n4188) );
  MUX2_X1 U961 ( .A(n779), .B(DATAIN[4]), .S(n33), .Z(n4189) );
  MUX2_X1 U962 ( .A(n780), .B(DATAIN[5]), .S(n33), .Z(n4190) );
  MUX2_X1 U963 ( .A(n781), .B(DATAIN[6]), .S(n33), .Z(n4191) );
  MUX2_X1 U964 ( .A(n782), .B(DATAIN[7]), .S(n33), .Z(n4192) );
  MUX2_X1 U965 ( .A(n783), .B(DATAIN[8]), .S(n32), .Z(n4193) );
  MUX2_X1 U966 ( .A(n784), .B(DATAIN[9]), .S(n32), .Z(n4194) );
  MUX2_X1 U967 ( .A(n785), .B(DATAIN[10]), .S(n32), .Z(n4195) );
  MUX2_X1 U968 ( .A(n786), .B(DATAIN[11]), .S(n32), .Z(n4196) );
  MUX2_X1 U969 ( .A(n787), .B(DATAIN[12]), .S(n32), .Z(n4197) );
  MUX2_X1 U970 ( .A(n788), .B(DATAIN[13]), .S(n32), .Z(n4198) );
  MUX2_X1 U971 ( .A(n789), .B(DATAIN[14]), .S(n32), .Z(n4199) );
  MUX2_X1 U972 ( .A(n790), .B(DATAIN[15]), .S(n32), .Z(n4200) );
  MUX2_X1 U973 ( .A(n791), .B(DATAIN[16]), .S(n32), .Z(n4201) );
  MUX2_X1 U974 ( .A(n792), .B(DATAIN[17]), .S(n32), .Z(n4202) );
  MUX2_X1 U975 ( .A(n793), .B(DATAIN[18]), .S(n32), .Z(n4203) );
  MUX2_X1 U976 ( .A(n794), .B(DATAIN[19]), .S(n32), .Z(n4204) );
  MUX2_X1 U977 ( .A(n795), .B(DATAIN[20]), .S(n31), .Z(n4205) );
  MUX2_X1 U978 ( .A(n796), .B(DATAIN[21]), .S(n31), .Z(n4206) );
  MUX2_X1 U979 ( .A(n797), .B(DATAIN[22]), .S(n31), .Z(n4207) );
  MUX2_X1 U980 ( .A(n798), .B(DATAIN[23]), .S(n31), .Z(n4208) );
  MUX2_X1 U981 ( .A(n799), .B(DATAIN[24]), .S(n31), .Z(n4209) );
  MUX2_X1 U982 ( .A(n800), .B(DATAIN[25]), .S(n31), .Z(n4210) );
  MUX2_X1 U983 ( .A(n801), .B(DATAIN[26]), .S(n31), .Z(n4211) );
  MUX2_X1 U984 ( .A(n802), .B(DATAIN[27]), .S(n31), .Z(n4212) );
  MUX2_X1 U985 ( .A(n803), .B(DATAIN[28]), .S(n31), .Z(n4213) );
  MUX2_X1 U986 ( .A(n804), .B(DATAIN[29]), .S(n31), .Z(n4214) );
  MUX2_X1 U987 ( .A(n805), .B(DATAIN[30]), .S(n31), .Z(n4215) );
  MUX2_X1 U988 ( .A(n806), .B(DATAIN[31]), .S(n31), .Z(n4216) );
  AND2_X1 U989 ( .A1(n807), .A2(n704), .ZN(n775) );
  MUX2_X1 U990 ( .A(n808), .B(DATAIN[0]), .S(n36), .Z(n4217) );
  MUX2_X1 U991 ( .A(n810), .B(DATAIN[1]), .S(n36), .Z(n4218) );
  MUX2_X1 U992 ( .A(n811), .B(DATAIN[2]), .S(n36), .Z(n4219) );
  MUX2_X1 U993 ( .A(n812), .B(DATAIN[3]), .S(n36), .Z(n4220) );
  MUX2_X1 U994 ( .A(n813), .B(DATAIN[4]), .S(n36), .Z(n4221) );
  MUX2_X1 U995 ( .A(n814), .B(DATAIN[5]), .S(n36), .Z(n4222) );
  MUX2_X1 U996 ( .A(n815), .B(DATAIN[6]), .S(n36), .Z(n4223) );
  MUX2_X1 U997 ( .A(n816), .B(DATAIN[7]), .S(n36), .Z(n4224) );
  MUX2_X1 U998 ( .A(n817), .B(DATAIN[8]), .S(n35), .Z(n4225) );
  MUX2_X1 U999 ( .A(n818), .B(DATAIN[9]), .S(n35), .Z(n4226) );
  MUX2_X1 U1000 ( .A(n819), .B(DATAIN[10]), .S(n35), .Z(n4227) );
  MUX2_X1 U1001 ( .A(n820), .B(DATAIN[11]), .S(n35), .Z(n4228) );
  MUX2_X1 U1002 ( .A(n821), .B(DATAIN[12]), .S(n35), .Z(n4229) );
  MUX2_X1 U1003 ( .A(n822), .B(DATAIN[13]), .S(n35), .Z(n4230) );
  MUX2_X1 U1004 ( .A(n823), .B(DATAIN[14]), .S(n35), .Z(n4231) );
  MUX2_X1 U1005 ( .A(n824), .B(DATAIN[15]), .S(n35), .Z(n4232) );
  MUX2_X1 U1006 ( .A(n825), .B(DATAIN[16]), .S(n35), .Z(n4233) );
  MUX2_X1 U1007 ( .A(n826), .B(DATAIN[17]), .S(n35), .Z(n4234) );
  MUX2_X1 U1008 ( .A(n827), .B(DATAIN[18]), .S(n35), .Z(n4235) );
  MUX2_X1 U1009 ( .A(n828), .B(DATAIN[19]), .S(n35), .Z(n4236) );
  MUX2_X1 U1010 ( .A(n829), .B(DATAIN[20]), .S(n34), .Z(n4237) );
  MUX2_X1 U1011 ( .A(n830), .B(DATAIN[21]), .S(n34), .Z(n4238) );
  MUX2_X1 U1012 ( .A(n831), .B(DATAIN[22]), .S(n34), .Z(n4239) );
  MUX2_X1 U1013 ( .A(n832), .B(DATAIN[23]), .S(n34), .Z(n4240) );
  MUX2_X1 U1014 ( .A(n833), .B(DATAIN[24]), .S(n34), .Z(n4241) );
  MUX2_X1 U1015 ( .A(n834), .B(DATAIN[25]), .S(n34), .Z(n4242) );
  MUX2_X1 U1016 ( .A(n835), .B(DATAIN[26]), .S(n34), .Z(n4243) );
  MUX2_X1 U1017 ( .A(n836), .B(DATAIN[27]), .S(n34), .Z(n4244) );
  MUX2_X1 U1018 ( .A(n837), .B(DATAIN[28]), .S(n34), .Z(n4245) );
  MUX2_X1 U1019 ( .A(n838), .B(DATAIN[29]), .S(n34), .Z(n4246) );
  MUX2_X1 U1020 ( .A(n839), .B(DATAIN[30]), .S(n34), .Z(n4247) );
  MUX2_X1 U1021 ( .A(n840), .B(DATAIN[31]), .S(n34), .Z(n4248) );
  AND2_X1 U1022 ( .A1(n841), .A2(n468), .ZN(n809) );
  INV_X1 U1023 ( .A(n842), .ZN(n4249) );
  MUX2_X1 U1024 ( .A(n3734), .B(n298), .S(n39), .Z(n842) );
  INV_X1 U1025 ( .A(n844), .ZN(n4250) );
  MUX2_X1 U1026 ( .A(n3713), .B(n299), .S(n39), .Z(n844) );
  INV_X1 U1027 ( .A(n845), .ZN(n4251) );
  MUX2_X1 U1028 ( .A(n3692), .B(n300), .S(n39), .Z(n845) );
  INV_X1 U1029 ( .A(n846), .ZN(n4252) );
  MUX2_X1 U1030 ( .A(n3671), .B(n301), .S(n39), .Z(n846) );
  INV_X1 U1031 ( .A(n847), .ZN(n4253) );
  MUX2_X1 U1032 ( .A(n3650), .B(n302), .S(n39), .Z(n847) );
  INV_X1 U1033 ( .A(n848), .ZN(n4254) );
  MUX2_X1 U1034 ( .A(n3629), .B(n303), .S(n39), .Z(n848) );
  INV_X1 U1035 ( .A(n849), .ZN(n4255) );
  MUX2_X1 U1036 ( .A(n3608), .B(n304), .S(n39), .Z(n849) );
  INV_X1 U1037 ( .A(n850), .ZN(n4256) );
  MUX2_X1 U1038 ( .A(n3587), .B(n305), .S(n39), .Z(n850) );
  INV_X1 U1039 ( .A(n851), .ZN(n4257) );
  MUX2_X1 U1040 ( .A(n3566), .B(n306), .S(n38), .Z(n851) );
  INV_X1 U1041 ( .A(n852), .ZN(n4258) );
  MUX2_X1 U1042 ( .A(n2969), .B(n307), .S(n38), .Z(n852) );
  INV_X1 U1043 ( .A(n853), .ZN(n4259) );
  MUX2_X1 U1044 ( .A(n2948), .B(n308), .S(n38), .Z(n853) );
  INV_X1 U1045 ( .A(n854), .ZN(n4260) );
  MUX2_X1 U1046 ( .A(n2927), .B(n309), .S(n38), .Z(n854) );
  INV_X1 U1047 ( .A(n855), .ZN(n4261) );
  MUX2_X1 U1048 ( .A(n2906), .B(n310), .S(n38), .Z(n855) );
  INV_X1 U1049 ( .A(n856), .ZN(n4262) );
  MUX2_X1 U1050 ( .A(n2885), .B(n311), .S(n38), .Z(n856) );
  INV_X1 U1051 ( .A(n857), .ZN(n4263) );
  MUX2_X1 U1052 ( .A(n2864), .B(n312), .S(n38), .Z(n857) );
  INV_X1 U1053 ( .A(n858), .ZN(n4264) );
  MUX2_X1 U1054 ( .A(n2843), .B(n313), .S(n38), .Z(n858) );
  INV_X1 U1055 ( .A(n859), .ZN(n4265) );
  MUX2_X1 U1056 ( .A(n2822), .B(n314), .S(n38), .Z(n859) );
  INV_X1 U1057 ( .A(n860), .ZN(n4266) );
  MUX2_X1 U1058 ( .A(n2801), .B(n315), .S(n38), .Z(n860) );
  INV_X1 U1059 ( .A(n861), .ZN(n4267) );
  MUX2_X1 U1060 ( .A(n2780), .B(n316), .S(n38), .Z(n861) );
  INV_X1 U1061 ( .A(n862), .ZN(n4268) );
  MUX2_X1 U1062 ( .A(n2759), .B(n317), .S(n38), .Z(n862) );
  INV_X1 U1063 ( .A(n863), .ZN(n4269) );
  MUX2_X1 U1064 ( .A(n2738), .B(n318), .S(n37), .Z(n863) );
  INV_X1 U1065 ( .A(n864), .ZN(n4270) );
  MUX2_X1 U1066 ( .A(n2717), .B(n319), .S(n37), .Z(n864) );
  INV_X1 U1067 ( .A(n865), .ZN(n4271) );
  MUX2_X1 U1068 ( .A(n2696), .B(n320), .S(n37), .Z(n865) );
  INV_X1 U1069 ( .A(n866), .ZN(n4272) );
  MUX2_X1 U1070 ( .A(n2675), .B(n321), .S(n37), .Z(n866) );
  INV_X1 U1071 ( .A(n867), .ZN(n4273) );
  MUX2_X1 U1072 ( .A(n2654), .B(n322), .S(n37), .Z(n867) );
  INV_X1 U1073 ( .A(n868), .ZN(n4274) );
  MUX2_X1 U1074 ( .A(n2633), .B(n323), .S(n37), .Z(n868) );
  INV_X1 U1075 ( .A(n869), .ZN(n4275) );
  MUX2_X1 U1076 ( .A(n2612), .B(n324), .S(n37), .Z(n869) );
  INV_X1 U1077 ( .A(n870), .ZN(n4276) );
  MUX2_X1 U1078 ( .A(n2591), .B(n325), .S(n37), .Z(n870) );
  INV_X1 U1079 ( .A(n871), .ZN(n4277) );
  MUX2_X1 U1080 ( .A(n2570), .B(n326), .S(n37), .Z(n871) );
  INV_X1 U1081 ( .A(n872), .ZN(n4278) );
  MUX2_X1 U1082 ( .A(n2549), .B(n327), .S(n37), .Z(n872) );
  INV_X1 U1083 ( .A(n873), .ZN(n4279) );
  MUX2_X1 U1084 ( .A(n2528), .B(n328), .S(n37), .Z(n873) );
  INV_X1 U1085 ( .A(n874), .ZN(n4280) );
  MUX2_X1 U1086 ( .A(n2507), .B(n329), .S(n37), .Z(n874) );
  AND2_X1 U1087 ( .A1(n841), .A2(n502), .ZN(n843) );
  INV_X1 U1088 ( .A(n875), .ZN(n4281) );
  MUX2_X1 U1089 ( .A(n3731), .B(n298), .S(n42), .Z(n875) );
  INV_X1 U1090 ( .A(n877), .ZN(n4282) );
  MUX2_X1 U1091 ( .A(n3710), .B(n299), .S(n42), .Z(n877) );
  INV_X1 U1092 ( .A(n878), .ZN(n4283) );
  MUX2_X1 U1093 ( .A(n3689), .B(n300), .S(n42), .Z(n878) );
  INV_X1 U1094 ( .A(n879), .ZN(n4284) );
  MUX2_X1 U1095 ( .A(n3668), .B(n301), .S(n42), .Z(n879) );
  INV_X1 U1096 ( .A(n880), .ZN(n4285) );
  MUX2_X1 U1097 ( .A(n3647), .B(n302), .S(n42), .Z(n880) );
  INV_X1 U1098 ( .A(n881), .ZN(n4286) );
  MUX2_X1 U1099 ( .A(n3626), .B(n303), .S(n42), .Z(n881) );
  INV_X1 U1100 ( .A(n882), .ZN(n4287) );
  MUX2_X1 U1101 ( .A(n3605), .B(n304), .S(n42), .Z(n882) );
  INV_X1 U1102 ( .A(n883), .ZN(n4288) );
  MUX2_X1 U1103 ( .A(n3584), .B(n305), .S(n42), .Z(n883) );
  INV_X1 U1104 ( .A(n884), .ZN(n4289) );
  MUX2_X1 U1105 ( .A(n3563), .B(n306), .S(n41), .Z(n884) );
  INV_X1 U1106 ( .A(n885), .ZN(n4290) );
  MUX2_X1 U1107 ( .A(n2966), .B(n307), .S(n41), .Z(n885) );
  INV_X1 U1108 ( .A(n886), .ZN(n4291) );
  MUX2_X1 U1109 ( .A(n2945), .B(n308), .S(n41), .Z(n886) );
  INV_X1 U1110 ( .A(n887), .ZN(n4292) );
  MUX2_X1 U1111 ( .A(n2924), .B(n309), .S(n41), .Z(n887) );
  INV_X1 U1112 ( .A(n888), .ZN(n4293) );
  MUX2_X1 U1113 ( .A(n2903), .B(n310), .S(n41), .Z(n888) );
  INV_X1 U1114 ( .A(n889), .ZN(n4294) );
  MUX2_X1 U1115 ( .A(n2882), .B(n311), .S(n41), .Z(n889) );
  INV_X1 U1116 ( .A(n890), .ZN(n4295) );
  MUX2_X1 U1117 ( .A(n2861), .B(n312), .S(n41), .Z(n890) );
  INV_X1 U1118 ( .A(n891), .ZN(n4296) );
  MUX2_X1 U1119 ( .A(n2840), .B(n313), .S(n41), .Z(n891) );
  INV_X1 U1120 ( .A(n892), .ZN(n4297) );
  MUX2_X1 U1121 ( .A(n2819), .B(n314), .S(n41), .Z(n892) );
  INV_X1 U1122 ( .A(n893), .ZN(n4298) );
  MUX2_X1 U1123 ( .A(n2798), .B(n315), .S(n41), .Z(n893) );
  INV_X1 U1124 ( .A(n894), .ZN(n4299) );
  MUX2_X1 U1125 ( .A(n2777), .B(n316), .S(n41), .Z(n894) );
  INV_X1 U1126 ( .A(n895), .ZN(n4300) );
  MUX2_X1 U1127 ( .A(n2756), .B(n317), .S(n41), .Z(n895) );
  INV_X1 U1128 ( .A(n896), .ZN(n4301) );
  MUX2_X1 U1129 ( .A(n2735), .B(n318), .S(n40), .Z(n896) );
  INV_X1 U1130 ( .A(n897), .ZN(n4302) );
  MUX2_X1 U1131 ( .A(n2714), .B(n319), .S(n40), .Z(n897) );
  INV_X1 U1132 ( .A(n898), .ZN(n4303) );
  MUX2_X1 U1133 ( .A(n2693), .B(n320), .S(n40), .Z(n898) );
  INV_X1 U1134 ( .A(n899), .ZN(n4304) );
  MUX2_X1 U1135 ( .A(n2672), .B(n321), .S(n40), .Z(n899) );
  INV_X1 U1136 ( .A(n900), .ZN(n4305) );
  MUX2_X1 U1137 ( .A(n2651), .B(n322), .S(n40), .Z(n900) );
  INV_X1 U1138 ( .A(n901), .ZN(n4306) );
  MUX2_X1 U1139 ( .A(n2630), .B(n323), .S(n40), .Z(n901) );
  INV_X1 U1140 ( .A(n902), .ZN(n4307) );
  MUX2_X1 U1141 ( .A(n2609), .B(n324), .S(n40), .Z(n902) );
  INV_X1 U1142 ( .A(n903), .ZN(n4308) );
  MUX2_X1 U1143 ( .A(n2588), .B(n325), .S(n40), .Z(n903) );
  INV_X1 U1144 ( .A(n904), .ZN(n4309) );
  MUX2_X1 U1145 ( .A(n2567), .B(n326), .S(n40), .Z(n904) );
  INV_X1 U1146 ( .A(n905), .ZN(n4310) );
  MUX2_X1 U1147 ( .A(n2546), .B(n327), .S(n40), .Z(n905) );
  INV_X1 U1148 ( .A(n906), .ZN(n4311) );
  MUX2_X1 U1149 ( .A(n2525), .B(n328), .S(n40), .Z(n906) );
  INV_X1 U1150 ( .A(n907), .ZN(n4312) );
  MUX2_X1 U1151 ( .A(n2504), .B(n329), .S(n40), .Z(n907) );
  AND2_X1 U1152 ( .A1(n841), .A2(n536), .ZN(n876) );
  MUX2_X1 U1153 ( .A(n908), .B(DATAIN[0]), .S(n45), .Z(n4313) );
  MUX2_X1 U1154 ( .A(n910), .B(DATAIN[1]), .S(n45), .Z(n4314) );
  MUX2_X1 U1155 ( .A(n911), .B(DATAIN[2]), .S(n45), .Z(n4315) );
  MUX2_X1 U1156 ( .A(n912), .B(DATAIN[3]), .S(n45), .Z(n4316) );
  MUX2_X1 U1157 ( .A(n913), .B(DATAIN[4]), .S(n45), .Z(n4317) );
  MUX2_X1 U1158 ( .A(n914), .B(DATAIN[5]), .S(n45), .Z(n4318) );
  MUX2_X1 U1159 ( .A(n915), .B(DATAIN[6]), .S(n45), .Z(n4319) );
  MUX2_X1 U1160 ( .A(n916), .B(DATAIN[7]), .S(n45), .Z(n4320) );
  MUX2_X1 U1161 ( .A(n917), .B(DATAIN[8]), .S(n44), .Z(n4321) );
  MUX2_X1 U1162 ( .A(n918), .B(DATAIN[9]), .S(n44), .Z(n4322) );
  MUX2_X1 U1163 ( .A(n919), .B(DATAIN[10]), .S(n44), .Z(n4323) );
  MUX2_X1 U1164 ( .A(n920), .B(DATAIN[11]), .S(n44), .Z(n4324) );
  MUX2_X1 U1165 ( .A(n921), .B(DATAIN[12]), .S(n44), .Z(n4325) );
  MUX2_X1 U1166 ( .A(n922), .B(DATAIN[13]), .S(n44), .Z(n4326) );
  MUX2_X1 U1167 ( .A(n923), .B(DATAIN[14]), .S(n44), .Z(n4327) );
  MUX2_X1 U1168 ( .A(n924), .B(DATAIN[15]), .S(n44), .Z(n4328) );
  MUX2_X1 U1169 ( .A(n925), .B(DATAIN[16]), .S(n44), .Z(n4329) );
  MUX2_X1 U1170 ( .A(n926), .B(DATAIN[17]), .S(n44), .Z(n4330) );
  MUX2_X1 U1171 ( .A(n927), .B(DATAIN[18]), .S(n44), .Z(n4331) );
  MUX2_X1 U1172 ( .A(n928), .B(DATAIN[19]), .S(n44), .Z(n4332) );
  MUX2_X1 U1173 ( .A(n929), .B(DATAIN[20]), .S(n43), .Z(n4333) );
  MUX2_X1 U1174 ( .A(n930), .B(DATAIN[21]), .S(n43), .Z(n4334) );
  MUX2_X1 U1175 ( .A(n931), .B(DATAIN[22]), .S(n43), .Z(n4335) );
  MUX2_X1 U1176 ( .A(n932), .B(DATAIN[23]), .S(n43), .Z(n4336) );
  MUX2_X1 U1177 ( .A(n933), .B(DATAIN[24]), .S(n43), .Z(n4337) );
  MUX2_X1 U1178 ( .A(n934), .B(DATAIN[25]), .S(n43), .Z(n4338) );
  MUX2_X1 U1179 ( .A(n935), .B(DATAIN[26]), .S(n43), .Z(n4339) );
  MUX2_X1 U1180 ( .A(n936), .B(DATAIN[27]), .S(n43), .Z(n4340) );
  MUX2_X1 U1181 ( .A(n937), .B(DATAIN[28]), .S(n43), .Z(n4341) );
  MUX2_X1 U1182 ( .A(n938), .B(DATAIN[29]), .S(n43), .Z(n4342) );
  MUX2_X1 U1183 ( .A(n939), .B(DATAIN[30]), .S(n43), .Z(n4343) );
  MUX2_X1 U1184 ( .A(n940), .B(DATAIN[31]), .S(n43), .Z(n4344) );
  AND2_X1 U1185 ( .A1(n841), .A2(n570), .ZN(n909) );
  MUX2_X1 U1186 ( .A(n2501), .B(DATAIN[31]), .S(n48), .Z(n3558) );
  MUX2_X1 U1187 ( .A(n2522), .B(DATAIN[30]), .S(n48), .Z(n3557) );
  MUX2_X1 U1188 ( .A(n2543), .B(DATAIN[29]), .S(n48), .Z(n3556) );
  MUX2_X1 U1189 ( .A(n2564), .B(DATAIN[28]), .S(n48), .Z(n3555) );
  MUX2_X1 U1190 ( .A(n2585), .B(DATAIN[27]), .S(n48), .Z(n3554) );
  MUX2_X1 U1191 ( .A(n2606), .B(DATAIN[26]), .S(n48), .Z(n3553) );
  MUX2_X1 U1192 ( .A(n2627), .B(DATAIN[25]), .S(n48), .Z(n3552) );
  MUX2_X1 U1193 ( .A(n2648), .B(DATAIN[24]), .S(n48), .Z(n3551) );
  MUX2_X1 U1194 ( .A(n2669), .B(DATAIN[23]), .S(n47), .Z(n3550) );
  MUX2_X1 U1195 ( .A(n2690), .B(DATAIN[22]), .S(n47), .Z(n3549) );
  MUX2_X1 U1196 ( .A(n2711), .B(DATAIN[21]), .S(n47), .Z(n3548) );
  MUX2_X1 U1197 ( .A(n2732), .B(DATAIN[20]), .S(n47), .Z(n3547) );
  MUX2_X1 U1198 ( .A(n2753), .B(DATAIN[19]), .S(n47), .Z(n3546) );
  MUX2_X1 U1199 ( .A(n2774), .B(DATAIN[18]), .S(n47), .Z(n3545) );
  MUX2_X1 U1200 ( .A(n2795), .B(DATAIN[17]), .S(n47), .Z(n3544) );
  MUX2_X1 U1201 ( .A(n2816), .B(DATAIN[16]), .S(n47), .Z(n3543) );
  MUX2_X1 U1202 ( .A(n2837), .B(DATAIN[15]), .S(n47), .Z(n3542) );
  MUX2_X1 U1203 ( .A(n2858), .B(DATAIN[14]), .S(n47), .Z(n3541) );
  MUX2_X1 U1204 ( .A(n2879), .B(DATAIN[13]), .S(n47), .Z(n3540) );
  MUX2_X1 U1205 ( .A(n2900), .B(DATAIN[12]), .S(n47), .Z(n3539) );
  MUX2_X1 U1206 ( .A(n2921), .B(DATAIN[11]), .S(n46), .Z(n3538) );
  MUX2_X1 U1207 ( .A(n2942), .B(DATAIN[10]), .S(n46), .Z(n3537) );
  MUX2_X1 U1208 ( .A(n2963), .B(DATAIN[9]), .S(n46), .Z(n3536) );
  MUX2_X1 U1209 ( .A(n3560), .B(DATAIN[8]), .S(n46), .Z(n3535) );
  MUX2_X1 U1210 ( .A(n3581), .B(DATAIN[7]), .S(n46), .Z(n3534) );
  MUX2_X1 U1211 ( .A(n3602), .B(DATAIN[6]), .S(n46), .Z(n3533) );
  MUX2_X1 U1212 ( .A(n3623), .B(DATAIN[5]), .S(n46), .Z(n3532) );
  MUX2_X1 U1213 ( .A(n3644), .B(DATAIN[4]), .S(n46), .Z(n3531) );
  MUX2_X1 U1214 ( .A(n3665), .B(DATAIN[3]), .S(n46), .Z(n3530) );
  MUX2_X1 U1215 ( .A(n3686), .B(DATAIN[2]), .S(n46), .Z(n3529) );
  MUX2_X1 U1216 ( .A(n3707), .B(DATAIN[1]), .S(n46), .Z(n3528) );
  MUX2_X1 U1217 ( .A(n3728), .B(DATAIN[0]), .S(n46), .Z(n3527) );
  AND2_X1 U1218 ( .A1(n705), .A2(n604), .ZN(n941) );
  MUX2_X1 U1219 ( .A(n2500), .B(DATAIN[31]), .S(n51), .Z(n3526) );
  MUX2_X1 U1220 ( .A(n2521), .B(DATAIN[30]), .S(n51), .Z(n3525) );
  MUX2_X1 U1221 ( .A(n2542), .B(DATAIN[29]), .S(n51), .Z(n3524) );
  MUX2_X1 U1222 ( .A(n2563), .B(DATAIN[28]), .S(n51), .Z(n3523) );
  MUX2_X1 U1223 ( .A(n2584), .B(DATAIN[27]), .S(n51), .Z(n3522) );
  MUX2_X1 U1224 ( .A(n2605), .B(DATAIN[26]), .S(n51), .Z(n3521) );
  MUX2_X1 U1225 ( .A(n2626), .B(DATAIN[25]), .S(n51), .Z(n3520) );
  MUX2_X1 U1226 ( .A(n2647), .B(DATAIN[24]), .S(n51), .Z(n3519) );
  MUX2_X1 U1227 ( .A(n2668), .B(DATAIN[23]), .S(n50), .Z(n3518) );
  MUX2_X1 U1228 ( .A(n2689), .B(DATAIN[22]), .S(n50), .Z(n3517) );
  MUX2_X1 U1229 ( .A(n2710), .B(DATAIN[21]), .S(n50), .Z(n3516) );
  MUX2_X1 U1230 ( .A(n2731), .B(DATAIN[20]), .S(n50), .Z(n3515) );
  MUX2_X1 U1231 ( .A(n2752), .B(DATAIN[19]), .S(n50), .Z(n3514) );
  MUX2_X1 U1232 ( .A(n2773), .B(DATAIN[18]), .S(n50), .Z(n3513) );
  MUX2_X1 U1233 ( .A(n2794), .B(DATAIN[17]), .S(n50), .Z(n3512) );
  MUX2_X1 U1234 ( .A(n2815), .B(DATAIN[16]), .S(n50), .Z(n3511) );
  MUX2_X1 U1235 ( .A(n2836), .B(DATAIN[15]), .S(n50), .Z(n3510) );
  MUX2_X1 U1236 ( .A(n2857), .B(DATAIN[14]), .S(n50), .Z(n3509) );
  MUX2_X1 U1237 ( .A(n2878), .B(DATAIN[13]), .S(n50), .Z(n3508) );
  MUX2_X1 U1238 ( .A(n2899), .B(DATAIN[12]), .S(n50), .Z(n3507) );
  MUX2_X1 U1239 ( .A(n2920), .B(DATAIN[11]), .S(n49), .Z(n3506) );
  MUX2_X1 U1240 ( .A(n2941), .B(DATAIN[10]), .S(n49), .Z(n3505) );
  MUX2_X1 U1241 ( .A(n2962), .B(DATAIN[9]), .S(n49), .Z(n3504) );
  MUX2_X1 U1242 ( .A(n3559), .B(DATAIN[8]), .S(n49), .Z(n3503) );
  MUX2_X1 U1243 ( .A(n3580), .B(DATAIN[7]), .S(n49), .Z(n3502) );
  MUX2_X1 U1244 ( .A(n3601), .B(DATAIN[6]), .S(n49), .Z(n3501) );
  MUX2_X1 U1245 ( .A(n3622), .B(DATAIN[5]), .S(n49), .Z(n3500) );
  MUX2_X1 U1246 ( .A(n3643), .B(DATAIN[4]), .S(n49), .Z(n3499) );
  MUX2_X1 U1247 ( .A(n3664), .B(DATAIN[3]), .S(n49), .Z(n3498) );
  MUX2_X1 U1248 ( .A(n3685), .B(DATAIN[2]), .S(n49), .Z(n3497) );
  MUX2_X1 U1249 ( .A(n3706), .B(DATAIN[1]), .S(n49), .Z(n3496) );
  MUX2_X1 U1250 ( .A(n3727), .B(DATAIN[0]), .S(n49), .Z(n3495) );
  AND2_X1 U1251 ( .A1(n739), .A2(n604), .ZN(n942) );
  MUX2_X1 U1252 ( .A(n2499), .B(DATAIN[31]), .S(n54), .Z(n3494) );
  MUX2_X1 U1253 ( .A(n2520), .B(DATAIN[30]), .S(n54), .Z(n3493) );
  MUX2_X1 U1254 ( .A(n2541), .B(DATAIN[29]), .S(n54), .Z(n3492) );
  MUX2_X1 U1255 ( .A(n2562), .B(DATAIN[28]), .S(n54), .Z(n3491) );
  MUX2_X1 U1256 ( .A(n2583), .B(DATAIN[27]), .S(n54), .Z(n3490) );
  MUX2_X1 U1257 ( .A(n2604), .B(DATAIN[26]), .S(n54), .Z(n3489) );
  MUX2_X1 U1258 ( .A(n2625), .B(DATAIN[25]), .S(n54), .Z(n3488) );
  MUX2_X1 U1259 ( .A(n2646), .B(DATAIN[24]), .S(n54), .Z(n3487) );
  MUX2_X1 U1260 ( .A(n2667), .B(DATAIN[23]), .S(n53), .Z(n3486) );
  MUX2_X1 U1261 ( .A(n2688), .B(DATAIN[22]), .S(n53), .Z(n3485) );
  MUX2_X1 U1262 ( .A(n2709), .B(DATAIN[21]), .S(n53), .Z(n3484) );
  MUX2_X1 U1263 ( .A(n2730), .B(DATAIN[20]), .S(n53), .Z(n3483) );
  MUX2_X1 U1264 ( .A(n2751), .B(DATAIN[19]), .S(n53), .Z(n3482) );
  MUX2_X1 U1265 ( .A(n2772), .B(DATAIN[18]), .S(n53), .Z(n3481) );
  MUX2_X1 U1266 ( .A(n2793), .B(DATAIN[17]), .S(n53), .Z(n3480) );
  MUX2_X1 U1267 ( .A(n2814), .B(DATAIN[16]), .S(n53), .Z(n3479) );
  MUX2_X1 U1268 ( .A(n2835), .B(DATAIN[15]), .S(n53), .Z(n3478) );
  MUX2_X1 U1269 ( .A(n2856), .B(DATAIN[14]), .S(n53), .Z(n3477) );
  MUX2_X1 U1270 ( .A(n2877), .B(DATAIN[13]), .S(n53), .Z(n3476) );
  MUX2_X1 U1271 ( .A(n2898), .B(DATAIN[12]), .S(n53), .Z(n3475) );
  MUX2_X1 U1272 ( .A(n2919), .B(DATAIN[11]), .S(n52), .Z(n3474) );
  MUX2_X1 U1273 ( .A(n2940), .B(DATAIN[10]), .S(n52), .Z(n3473) );
  MUX2_X1 U1274 ( .A(n2961), .B(DATAIN[9]), .S(n52), .Z(n3472) );
  MUX2_X1 U1275 ( .A(n2982), .B(DATAIN[8]), .S(n52), .Z(n3471) );
  MUX2_X1 U1276 ( .A(n3579), .B(DATAIN[7]), .S(n52), .Z(n3470) );
  MUX2_X1 U1277 ( .A(n3600), .B(DATAIN[6]), .S(n52), .Z(n3469) );
  MUX2_X1 U1278 ( .A(n3621), .B(DATAIN[5]), .S(n52), .Z(n3468) );
  MUX2_X1 U1279 ( .A(n3642), .B(DATAIN[4]), .S(n52), .Z(n3467) );
  MUX2_X1 U1280 ( .A(n3663), .B(DATAIN[3]), .S(n52), .Z(n3466) );
  MUX2_X1 U1281 ( .A(n3684), .B(DATAIN[2]), .S(n52), .Z(n3465) );
  MUX2_X1 U1282 ( .A(n3705), .B(DATAIN[1]), .S(n52), .Z(n3464) );
  MUX2_X1 U1283 ( .A(n3726), .B(DATAIN[0]), .S(n52), .Z(n3463) );
  AND2_X1 U1284 ( .A1(n773), .A2(n604), .ZN(n943) );
  MUX2_X1 U1285 ( .A(n2498), .B(DATAIN[31]), .S(n57), .Z(n3462) );
  MUX2_X1 U1286 ( .A(n2519), .B(DATAIN[30]), .S(n57), .Z(n3461) );
  MUX2_X1 U1287 ( .A(n2540), .B(DATAIN[29]), .S(n57), .Z(n3460) );
  MUX2_X1 U1288 ( .A(n2561), .B(DATAIN[28]), .S(n57), .Z(n3459) );
  MUX2_X1 U1289 ( .A(n2582), .B(DATAIN[27]), .S(n57), .Z(n3458) );
  MUX2_X1 U1290 ( .A(n2603), .B(DATAIN[26]), .S(n57), .Z(n3457) );
  MUX2_X1 U1291 ( .A(n2624), .B(DATAIN[25]), .S(n57), .Z(n3456) );
  MUX2_X1 U1292 ( .A(n2645), .B(DATAIN[24]), .S(n57), .Z(n3455) );
  MUX2_X1 U1293 ( .A(n2666), .B(DATAIN[23]), .S(n56), .Z(n3454) );
  MUX2_X1 U1294 ( .A(n2687), .B(DATAIN[22]), .S(n56), .Z(n3453) );
  MUX2_X1 U1295 ( .A(n2708), .B(DATAIN[21]), .S(n56), .Z(n3452) );
  MUX2_X1 U1296 ( .A(n2729), .B(DATAIN[20]), .S(n56), .Z(n3451) );
  MUX2_X1 U1297 ( .A(n2750), .B(DATAIN[19]), .S(n56), .Z(n3450) );
  MUX2_X1 U1298 ( .A(n2771), .B(DATAIN[18]), .S(n56), .Z(n3449) );
  MUX2_X1 U1299 ( .A(n2792), .B(DATAIN[17]), .S(n56), .Z(n3448) );
  MUX2_X1 U1300 ( .A(n2813), .B(DATAIN[16]), .S(n56), .Z(n3447) );
  MUX2_X1 U1301 ( .A(n2834), .B(DATAIN[15]), .S(n56), .Z(n3446) );
  MUX2_X1 U1302 ( .A(n2855), .B(DATAIN[14]), .S(n56), .Z(n3445) );
  MUX2_X1 U1303 ( .A(n2876), .B(DATAIN[13]), .S(n56), .Z(n3444) );
  MUX2_X1 U1304 ( .A(n2897), .B(DATAIN[12]), .S(n56), .Z(n3443) );
  MUX2_X1 U1305 ( .A(n2918), .B(DATAIN[11]), .S(n55), .Z(n3442) );
  MUX2_X1 U1306 ( .A(n2939), .B(DATAIN[10]), .S(n55), .Z(n3441) );
  MUX2_X1 U1307 ( .A(n2960), .B(DATAIN[9]), .S(n55), .Z(n3440) );
  MUX2_X1 U1308 ( .A(n2981), .B(DATAIN[8]), .S(n55), .Z(n3439) );
  MUX2_X1 U1309 ( .A(n3578), .B(DATAIN[7]), .S(n55), .Z(n3438) );
  MUX2_X1 U1310 ( .A(n3599), .B(DATAIN[6]), .S(n55), .Z(n3437) );
  MUX2_X1 U1311 ( .A(n3620), .B(DATAIN[5]), .S(n55), .Z(n3436) );
  MUX2_X1 U1312 ( .A(n3641), .B(DATAIN[4]), .S(n55), .Z(n3435) );
  MUX2_X1 U1313 ( .A(n3662), .B(DATAIN[3]), .S(n55), .Z(n3434) );
  MUX2_X1 U1314 ( .A(n3683), .B(DATAIN[2]), .S(n55), .Z(n3433) );
  MUX2_X1 U1315 ( .A(n3704), .B(DATAIN[1]), .S(n55), .Z(n3432) );
  MUX2_X1 U1316 ( .A(n3725), .B(DATAIN[0]), .S(n55), .Z(n3431) );
  AND2_X1 U1317 ( .A1(n807), .A2(n604), .ZN(n944) );
  AND3_X1 U1318 ( .A1(n945), .A2(n946), .A3(n947), .ZN(n604) );
  MUX2_X1 U1319 ( .A(n2497), .B(DATAIN[31]), .S(n60), .Z(n3430) );
  MUX2_X1 U1320 ( .A(n2518), .B(DATAIN[30]), .S(n60), .Z(n3429) );
  MUX2_X1 U1321 ( .A(n2539), .B(DATAIN[29]), .S(n60), .Z(n3428) );
  MUX2_X1 U1322 ( .A(n2560), .B(DATAIN[28]), .S(n60), .Z(n3427) );
  MUX2_X1 U1323 ( .A(n2581), .B(DATAIN[27]), .S(n60), .Z(n3426) );
  MUX2_X1 U1324 ( .A(n2602), .B(DATAIN[26]), .S(n60), .Z(n3425) );
  MUX2_X1 U1325 ( .A(n2623), .B(DATAIN[25]), .S(n60), .Z(n3424) );
  MUX2_X1 U1326 ( .A(n2644), .B(DATAIN[24]), .S(n60), .Z(n3423) );
  MUX2_X1 U1327 ( .A(n2665), .B(DATAIN[23]), .S(n59), .Z(n3422) );
  MUX2_X1 U1328 ( .A(n2686), .B(DATAIN[22]), .S(n59), .Z(n3421) );
  MUX2_X1 U1329 ( .A(n2707), .B(DATAIN[21]), .S(n59), .Z(n3420) );
  MUX2_X1 U1330 ( .A(n2728), .B(DATAIN[20]), .S(n59), .Z(n3419) );
  MUX2_X1 U1331 ( .A(n2749), .B(DATAIN[19]), .S(n59), .Z(n3418) );
  MUX2_X1 U1332 ( .A(n2770), .B(DATAIN[18]), .S(n59), .Z(n3417) );
  MUX2_X1 U1333 ( .A(n2791), .B(DATAIN[17]), .S(n59), .Z(n3416) );
  MUX2_X1 U1334 ( .A(n2812), .B(DATAIN[16]), .S(n59), .Z(n3415) );
  MUX2_X1 U1335 ( .A(n2833), .B(DATAIN[15]), .S(n59), .Z(n3414) );
  MUX2_X1 U1336 ( .A(n2854), .B(DATAIN[14]), .S(n59), .Z(n3413) );
  MUX2_X1 U1337 ( .A(n2875), .B(DATAIN[13]), .S(n59), .Z(n3412) );
  MUX2_X1 U1338 ( .A(n2896), .B(DATAIN[12]), .S(n59), .Z(n3411) );
  MUX2_X1 U1339 ( .A(n2917), .B(DATAIN[11]), .S(n58), .Z(n3410) );
  MUX2_X1 U1340 ( .A(n2938), .B(DATAIN[10]), .S(n58), .Z(n3409) );
  MUX2_X1 U1341 ( .A(n2959), .B(DATAIN[9]), .S(n58), .Z(n3408) );
  MUX2_X1 U1342 ( .A(n2980), .B(DATAIN[8]), .S(n58), .Z(n3407) );
  MUX2_X1 U1343 ( .A(n3577), .B(DATAIN[7]), .S(n58), .Z(n3406) );
  MUX2_X1 U1344 ( .A(n3598), .B(DATAIN[6]), .S(n58), .Z(n3405) );
  MUX2_X1 U1345 ( .A(n3619), .B(DATAIN[5]), .S(n58), .Z(n3404) );
  MUX2_X1 U1346 ( .A(n3640), .B(DATAIN[4]), .S(n58), .Z(n3403) );
  MUX2_X1 U1347 ( .A(n3661), .B(DATAIN[3]), .S(n58), .Z(n3402) );
  MUX2_X1 U1348 ( .A(n3682), .B(DATAIN[2]), .S(n58), .Z(n3401) );
  MUX2_X1 U1349 ( .A(n3703), .B(DATAIN[1]), .S(n58), .Z(n3400) );
  MUX2_X1 U1350 ( .A(n3724), .B(DATAIN[0]), .S(n58), .Z(n3399) );
  AND2_X1 U1351 ( .A1(n705), .A2(n467), .ZN(n948) );
  MUX2_X1 U1352 ( .A(n2496), .B(DATAIN[31]), .S(n63), .Z(n3398) );
  MUX2_X1 U1353 ( .A(n2517), .B(DATAIN[30]), .S(n63), .Z(n3397) );
  MUX2_X1 U1354 ( .A(n2538), .B(DATAIN[29]), .S(n63), .Z(n3396) );
  MUX2_X1 U1355 ( .A(n2559), .B(DATAIN[28]), .S(n63), .Z(n3395) );
  MUX2_X1 U1356 ( .A(n2580), .B(DATAIN[27]), .S(n63), .Z(n3394) );
  MUX2_X1 U1357 ( .A(n2601), .B(DATAIN[26]), .S(n63), .Z(n3393) );
  MUX2_X1 U1358 ( .A(n2622), .B(DATAIN[25]), .S(n63), .Z(n3392) );
  MUX2_X1 U1359 ( .A(n2643), .B(DATAIN[24]), .S(n63), .Z(n3391) );
  MUX2_X1 U1360 ( .A(n2664), .B(DATAIN[23]), .S(n62), .Z(n3390) );
  MUX2_X1 U1361 ( .A(n2685), .B(DATAIN[22]), .S(n62), .Z(n3389) );
  MUX2_X1 U1362 ( .A(n2706), .B(DATAIN[21]), .S(n62), .Z(n3388) );
  MUX2_X1 U1363 ( .A(n2727), .B(DATAIN[20]), .S(n62), .Z(n3387) );
  MUX2_X1 U1364 ( .A(n2748), .B(DATAIN[19]), .S(n62), .Z(n3386) );
  MUX2_X1 U1365 ( .A(n2769), .B(DATAIN[18]), .S(n62), .Z(n3385) );
  MUX2_X1 U1366 ( .A(n2790), .B(DATAIN[17]), .S(n62), .Z(n3384) );
  MUX2_X1 U1367 ( .A(n2811), .B(DATAIN[16]), .S(n62), .Z(n3383) );
  MUX2_X1 U1368 ( .A(n2832), .B(DATAIN[15]), .S(n62), .Z(n3382) );
  MUX2_X1 U1369 ( .A(n2853), .B(DATAIN[14]), .S(n62), .Z(n3381) );
  MUX2_X1 U1370 ( .A(n2874), .B(DATAIN[13]), .S(n62), .Z(n3380) );
  MUX2_X1 U1371 ( .A(n2895), .B(DATAIN[12]), .S(n62), .Z(n3379) );
  MUX2_X1 U1372 ( .A(n2916), .B(DATAIN[11]), .S(n61), .Z(n3378) );
  MUX2_X1 U1373 ( .A(n2937), .B(DATAIN[10]), .S(n61), .Z(n3377) );
  MUX2_X1 U1374 ( .A(n2958), .B(DATAIN[9]), .S(n61), .Z(n3376) );
  MUX2_X1 U1375 ( .A(n2979), .B(DATAIN[8]), .S(n61), .Z(n3375) );
  MUX2_X1 U1376 ( .A(n3576), .B(DATAIN[7]), .S(n61), .Z(n3374) );
  MUX2_X1 U1377 ( .A(n3597), .B(DATAIN[6]), .S(n61), .Z(n3373) );
  MUX2_X1 U1378 ( .A(n3618), .B(DATAIN[5]), .S(n61), .Z(n3372) );
  MUX2_X1 U1379 ( .A(n3639), .B(DATAIN[4]), .S(n61), .Z(n3371) );
  MUX2_X1 U1380 ( .A(n3660), .B(DATAIN[3]), .S(n61), .Z(n3370) );
  MUX2_X1 U1381 ( .A(n3681), .B(DATAIN[2]), .S(n61), .Z(n3369) );
  MUX2_X1 U1382 ( .A(n3702), .B(DATAIN[1]), .S(n61), .Z(n3368) );
  MUX2_X1 U1383 ( .A(n3723), .B(DATAIN[0]), .S(n61), .Z(n3367) );
  AND2_X1 U1384 ( .A1(n739), .A2(n467), .ZN(n949) );
  MUX2_X1 U1385 ( .A(n2493), .B(DATAIN[31]), .S(n66), .Z(n3366) );
  MUX2_X1 U1386 ( .A(n2514), .B(DATAIN[30]), .S(n66), .Z(n3365) );
  MUX2_X1 U1387 ( .A(n2535), .B(DATAIN[29]), .S(n66), .Z(n3364) );
  MUX2_X1 U1388 ( .A(n2556), .B(DATAIN[28]), .S(n66), .Z(n3363) );
  MUX2_X1 U1389 ( .A(n2577), .B(DATAIN[27]), .S(n66), .Z(n3362) );
  MUX2_X1 U1390 ( .A(n2598), .B(DATAIN[26]), .S(n66), .Z(n3361) );
  MUX2_X1 U1391 ( .A(n2619), .B(DATAIN[25]), .S(n66), .Z(n3360) );
  MUX2_X1 U1392 ( .A(n2640), .B(DATAIN[24]), .S(n66), .Z(n3359) );
  MUX2_X1 U1393 ( .A(n2661), .B(DATAIN[23]), .S(n65), .Z(n3358) );
  MUX2_X1 U1394 ( .A(n2682), .B(DATAIN[22]), .S(n65), .Z(n3357) );
  MUX2_X1 U1395 ( .A(n2703), .B(DATAIN[21]), .S(n65), .Z(n3356) );
  MUX2_X1 U1396 ( .A(n2724), .B(DATAIN[20]), .S(n65), .Z(n3355) );
  MUX2_X1 U1397 ( .A(n2745), .B(DATAIN[19]), .S(n65), .Z(n3354) );
  MUX2_X1 U1398 ( .A(n2766), .B(DATAIN[18]), .S(n65), .Z(n3353) );
  MUX2_X1 U1399 ( .A(n2787), .B(DATAIN[17]), .S(n65), .Z(n3352) );
  MUX2_X1 U1400 ( .A(n2808), .B(DATAIN[16]), .S(n65), .Z(n3351) );
  MUX2_X1 U1401 ( .A(n2829), .B(DATAIN[15]), .S(n65), .Z(n3350) );
  MUX2_X1 U1402 ( .A(n2850), .B(DATAIN[14]), .S(n65), .Z(n3349) );
  MUX2_X1 U1403 ( .A(n2871), .B(DATAIN[13]), .S(n65), .Z(n3348) );
  MUX2_X1 U1404 ( .A(n2892), .B(DATAIN[12]), .S(n65), .Z(n3347) );
  MUX2_X1 U1405 ( .A(n2913), .B(DATAIN[11]), .S(n64), .Z(n3346) );
  MUX2_X1 U1406 ( .A(n2934), .B(DATAIN[10]), .S(n64), .Z(n3345) );
  MUX2_X1 U1407 ( .A(n2955), .B(DATAIN[9]), .S(n64), .Z(n3344) );
  MUX2_X1 U1408 ( .A(n2976), .B(DATAIN[8]), .S(n64), .Z(n3343) );
  MUX2_X1 U1409 ( .A(n3573), .B(DATAIN[7]), .S(n64), .Z(n3342) );
  MUX2_X1 U1410 ( .A(n3594), .B(DATAIN[6]), .S(n64), .Z(n3341) );
  MUX2_X1 U1411 ( .A(n3615), .B(DATAIN[5]), .S(n64), .Z(n3340) );
  MUX2_X1 U1412 ( .A(n3636), .B(DATAIN[4]), .S(n64), .Z(n3339) );
  MUX2_X1 U1413 ( .A(n3657), .B(DATAIN[3]), .S(n64), .Z(n3338) );
  MUX2_X1 U1414 ( .A(n3678), .B(DATAIN[2]), .S(n64), .Z(n3337) );
  MUX2_X1 U1415 ( .A(n3699), .B(DATAIN[1]), .S(n64), .Z(n3336) );
  MUX2_X1 U1416 ( .A(n3720), .B(DATAIN[0]), .S(n64), .Z(n3335) );
  AND2_X1 U1417 ( .A1(n773), .A2(n467), .ZN(n950) );
  MUX2_X1 U1418 ( .A(n2492), .B(DATAIN[31]), .S(n69), .Z(n3334) );
  MUX2_X1 U1419 ( .A(n2513), .B(DATAIN[30]), .S(n69), .Z(n3333) );
  MUX2_X1 U1420 ( .A(n2534), .B(DATAIN[29]), .S(n69), .Z(n3332) );
  MUX2_X1 U1421 ( .A(n2555), .B(DATAIN[28]), .S(n69), .Z(n3331) );
  MUX2_X1 U1422 ( .A(n2576), .B(DATAIN[27]), .S(n69), .Z(n3330) );
  MUX2_X1 U1423 ( .A(n2597), .B(DATAIN[26]), .S(n69), .Z(n3329) );
  MUX2_X1 U1424 ( .A(n2618), .B(DATAIN[25]), .S(n69), .Z(n3328) );
  MUX2_X1 U1425 ( .A(n2639), .B(DATAIN[24]), .S(n69), .Z(n3327) );
  MUX2_X1 U1426 ( .A(n2660), .B(DATAIN[23]), .S(n68), .Z(n3326) );
  MUX2_X1 U1427 ( .A(n2681), .B(DATAIN[22]), .S(n68), .Z(n3325) );
  MUX2_X1 U1428 ( .A(n2702), .B(DATAIN[21]), .S(n68), .Z(n3324) );
  MUX2_X1 U1429 ( .A(n2723), .B(DATAIN[20]), .S(n68), .Z(n3323) );
  MUX2_X1 U1430 ( .A(n2744), .B(DATAIN[19]), .S(n68), .Z(n3322) );
  MUX2_X1 U1431 ( .A(n2765), .B(DATAIN[18]), .S(n68), .Z(n3321) );
  MUX2_X1 U1432 ( .A(n2786), .B(DATAIN[17]), .S(n68), .Z(n3320) );
  MUX2_X1 U1433 ( .A(n2807), .B(DATAIN[16]), .S(n68), .Z(n3319) );
  MUX2_X1 U1434 ( .A(n2828), .B(DATAIN[15]), .S(n68), .Z(n3318) );
  MUX2_X1 U1435 ( .A(n2849), .B(DATAIN[14]), .S(n68), .Z(n3317) );
  MUX2_X1 U1436 ( .A(n2870), .B(DATAIN[13]), .S(n68), .Z(n3316) );
  MUX2_X1 U1437 ( .A(n2891), .B(DATAIN[12]), .S(n68), .Z(n3315) );
  MUX2_X1 U1438 ( .A(n2912), .B(DATAIN[11]), .S(n67), .Z(n3314) );
  MUX2_X1 U1439 ( .A(n2933), .B(DATAIN[10]), .S(n67), .Z(n3313) );
  MUX2_X1 U1440 ( .A(n2954), .B(DATAIN[9]), .S(n67), .Z(n3312) );
  MUX2_X1 U1441 ( .A(n2975), .B(DATAIN[8]), .S(n67), .Z(n3311) );
  MUX2_X1 U1442 ( .A(n3572), .B(DATAIN[7]), .S(n67), .Z(n3310) );
  MUX2_X1 U1443 ( .A(n3593), .B(DATAIN[6]), .S(n67), .Z(n3309) );
  MUX2_X1 U1444 ( .A(n3614), .B(DATAIN[5]), .S(n67), .Z(n3308) );
  MUX2_X1 U1445 ( .A(n3635), .B(DATAIN[4]), .S(n67), .Z(n3307) );
  MUX2_X1 U1446 ( .A(n3656), .B(DATAIN[3]), .S(n67), .Z(n3306) );
  MUX2_X1 U1447 ( .A(n3677), .B(DATAIN[2]), .S(n67), .Z(n3305) );
  MUX2_X1 U1448 ( .A(n3698), .B(DATAIN[1]), .S(n67), .Z(n3304) );
  MUX2_X1 U1449 ( .A(n3719), .B(DATAIN[0]), .S(n67), .Z(n3303) );
  AND2_X1 U1450 ( .A1(n807), .A2(n467), .ZN(n951) );
  AND3_X1 U1451 ( .A1(n947), .A2(n946), .A3(ADD_WR[3]), .ZN(n467) );
  INV_X1 U1452 ( .A(ADD_WR[4]), .ZN(n946) );
  MUX2_X1 U1453 ( .A(n2509), .B(DATAIN[31]), .S(n72), .Z(n3302) );
  MUX2_X1 U1454 ( .A(n2530), .B(DATAIN[30]), .S(n72), .Z(n3301) );
  MUX2_X1 U1455 ( .A(n2551), .B(DATAIN[29]), .S(n72), .Z(n3300) );
  MUX2_X1 U1456 ( .A(n2572), .B(DATAIN[28]), .S(n72), .Z(n3299) );
  MUX2_X1 U1457 ( .A(n2593), .B(DATAIN[27]), .S(n72), .Z(n3298) );
  MUX2_X1 U1458 ( .A(n2614), .B(DATAIN[26]), .S(n72), .Z(n3297) );
  MUX2_X1 U1459 ( .A(n2635), .B(DATAIN[25]), .S(n72), .Z(n3296) );
  MUX2_X1 U1460 ( .A(n2656), .B(DATAIN[24]), .S(n72), .Z(n3295) );
  MUX2_X1 U1461 ( .A(n2677), .B(DATAIN[23]), .S(n71), .Z(n3294) );
  MUX2_X1 U1462 ( .A(n2698), .B(DATAIN[22]), .S(n71), .Z(n3293) );
  MUX2_X1 U1463 ( .A(n2719), .B(DATAIN[21]), .S(n71), .Z(n3292) );
  MUX2_X1 U1464 ( .A(n2740), .B(DATAIN[20]), .S(n71), .Z(n3291) );
  MUX2_X1 U1465 ( .A(n2761), .B(DATAIN[19]), .S(n71), .Z(n3290) );
  MUX2_X1 U1466 ( .A(n2782), .B(DATAIN[18]), .S(n71), .Z(n3289) );
  MUX2_X1 U1467 ( .A(n2803), .B(DATAIN[17]), .S(n71), .Z(n3288) );
  MUX2_X1 U1468 ( .A(n2824), .B(DATAIN[16]), .S(n71), .Z(n3287) );
  MUX2_X1 U1469 ( .A(n2845), .B(DATAIN[15]), .S(n71), .Z(n3286) );
  MUX2_X1 U1470 ( .A(n2866), .B(DATAIN[14]), .S(n71), .Z(n3285) );
  MUX2_X1 U1471 ( .A(n2887), .B(DATAIN[13]), .S(n71), .Z(n3284) );
  MUX2_X1 U1472 ( .A(n2908), .B(DATAIN[12]), .S(n71), .Z(n3283) );
  MUX2_X1 U1473 ( .A(n2929), .B(DATAIN[11]), .S(n70), .Z(n3282) );
  MUX2_X1 U1474 ( .A(n2950), .B(DATAIN[10]), .S(n70), .Z(n3281) );
  MUX2_X1 U1475 ( .A(n2971), .B(DATAIN[9]), .S(n70), .Z(n3280) );
  MUX2_X1 U1476 ( .A(n3568), .B(DATAIN[8]), .S(n70), .Z(n3279) );
  MUX2_X1 U1477 ( .A(n3589), .B(DATAIN[7]), .S(n70), .Z(n3278) );
  MUX2_X1 U1478 ( .A(n3610), .B(DATAIN[6]), .S(n70), .Z(n3277) );
  MUX2_X1 U1479 ( .A(n3631), .B(DATAIN[5]), .S(n70), .Z(n3276) );
  MUX2_X1 U1480 ( .A(n3652), .B(DATAIN[4]), .S(n70), .Z(n3275) );
  MUX2_X1 U1481 ( .A(n3673), .B(DATAIN[3]), .S(n70), .Z(n3274) );
  MUX2_X1 U1482 ( .A(n3694), .B(DATAIN[2]), .S(n70), .Z(n3273) );
  MUX2_X1 U1483 ( .A(n3715), .B(DATAIN[1]), .S(n70), .Z(n3272) );
  MUX2_X1 U1484 ( .A(n3736), .B(DATAIN[0]), .S(n70), .Z(n3271) );
  AND2_X1 U1485 ( .A1(n841), .A2(n705), .ZN(n952) );
  AND3_X1 U1486 ( .A1(n953), .A2(n954), .A3(ADD_WR[1]), .ZN(n705) );
  MUX2_X1 U1487 ( .A(n2508), .B(DATAIN[31]), .S(n75), .Z(n3270) );
  MUX2_X1 U1488 ( .A(n2529), .B(DATAIN[30]), .S(n75), .Z(n3269) );
  MUX2_X1 U1489 ( .A(n2550), .B(DATAIN[29]), .S(n75), .Z(n3268) );
  MUX2_X1 U1490 ( .A(n2571), .B(DATAIN[28]), .S(n75), .Z(n3267) );
  MUX2_X1 U1491 ( .A(n2592), .B(DATAIN[27]), .S(n75), .Z(n3266) );
  MUX2_X1 U1492 ( .A(n2613), .B(DATAIN[26]), .S(n75), .Z(n3265) );
  MUX2_X1 U1493 ( .A(n2634), .B(DATAIN[25]), .S(n75), .Z(n3264) );
  MUX2_X1 U1494 ( .A(n2655), .B(DATAIN[24]), .S(n75), .Z(n3263) );
  MUX2_X1 U1495 ( .A(n2676), .B(DATAIN[23]), .S(n74), .Z(n3262) );
  MUX2_X1 U1496 ( .A(n2697), .B(DATAIN[22]), .S(n74), .Z(n3261) );
  MUX2_X1 U1497 ( .A(n2718), .B(DATAIN[21]), .S(n74), .Z(n3260) );
  MUX2_X1 U1498 ( .A(n2739), .B(DATAIN[20]), .S(n74), .Z(n3259) );
  MUX2_X1 U1499 ( .A(n2760), .B(DATAIN[19]), .S(n74), .Z(n3258) );
  MUX2_X1 U1500 ( .A(n2781), .B(DATAIN[18]), .S(n74), .Z(n3257) );
  MUX2_X1 U1501 ( .A(n2802), .B(DATAIN[17]), .S(n74), .Z(n3256) );
  MUX2_X1 U1502 ( .A(n2823), .B(DATAIN[16]), .S(n74), .Z(n3255) );
  MUX2_X1 U1503 ( .A(n2844), .B(DATAIN[15]), .S(n74), .Z(n3254) );
  MUX2_X1 U1504 ( .A(n2865), .B(DATAIN[14]), .S(n74), .Z(n3253) );
  MUX2_X1 U1505 ( .A(n2886), .B(DATAIN[13]), .S(n74), .Z(n3252) );
  MUX2_X1 U1506 ( .A(n2907), .B(DATAIN[12]), .S(n74), .Z(n3251) );
  MUX2_X1 U1507 ( .A(n2928), .B(DATAIN[11]), .S(n73), .Z(n3250) );
  MUX2_X1 U1508 ( .A(n2949), .B(DATAIN[10]), .S(n73), .Z(n3249) );
  MUX2_X1 U1509 ( .A(n2970), .B(DATAIN[9]), .S(n73), .Z(n3248) );
  MUX2_X1 U1510 ( .A(n3567), .B(DATAIN[8]), .S(n73), .Z(n3247) );
  MUX2_X1 U1511 ( .A(n3588), .B(DATAIN[7]), .S(n73), .Z(n3246) );
  MUX2_X1 U1512 ( .A(n3609), .B(DATAIN[6]), .S(n73), .Z(n3245) );
  MUX2_X1 U1513 ( .A(n3630), .B(DATAIN[5]), .S(n73), .Z(n3244) );
  MUX2_X1 U1514 ( .A(n3651), .B(DATAIN[4]), .S(n73), .Z(n3243) );
  MUX2_X1 U1515 ( .A(n3672), .B(DATAIN[3]), .S(n73), .Z(n3242) );
  MUX2_X1 U1516 ( .A(n3693), .B(DATAIN[2]), .S(n73), .Z(n3241) );
  MUX2_X1 U1517 ( .A(n3714), .B(DATAIN[1]), .S(n73), .Z(n3240) );
  MUX2_X1 U1518 ( .A(n3735), .B(DATAIN[0]), .S(n73), .Z(n3239) );
  AND2_X1 U1519 ( .A1(n841), .A2(n739), .ZN(n955) );
  AND3_X1 U1520 ( .A1(ADD_WR[0]), .A2(n954), .A3(ADD_WR[1]), .ZN(n739) );
  MUX2_X1 U1521 ( .A(n2506), .B(DATAIN[31]), .S(n78), .Z(n3238) );
  MUX2_X1 U1522 ( .A(n2527), .B(DATAIN[30]), .S(n78), .Z(n3237) );
  MUX2_X1 U1523 ( .A(n2548), .B(DATAIN[29]), .S(n78), .Z(n3236) );
  MUX2_X1 U1524 ( .A(n2569), .B(DATAIN[28]), .S(n78), .Z(n3235) );
  MUX2_X1 U1525 ( .A(n2590), .B(DATAIN[27]), .S(n78), .Z(n3234) );
  MUX2_X1 U1526 ( .A(n2611), .B(DATAIN[26]), .S(n78), .Z(n3233) );
  MUX2_X1 U1527 ( .A(n2632), .B(DATAIN[25]), .S(n78), .Z(n3232) );
  MUX2_X1 U1528 ( .A(n2653), .B(DATAIN[24]), .S(n78), .Z(n3231) );
  MUX2_X1 U1529 ( .A(n2674), .B(DATAIN[23]), .S(n77), .Z(n3230) );
  MUX2_X1 U1530 ( .A(n2695), .B(DATAIN[22]), .S(n77), .Z(n3229) );
  MUX2_X1 U1531 ( .A(n2716), .B(DATAIN[21]), .S(n77), .Z(n3228) );
  MUX2_X1 U1532 ( .A(n2737), .B(DATAIN[20]), .S(n77), .Z(n3227) );
  MUX2_X1 U1533 ( .A(n2758), .B(DATAIN[19]), .S(n77), .Z(n3226) );
  MUX2_X1 U1534 ( .A(n2779), .B(DATAIN[18]), .S(n77), .Z(n3225) );
  MUX2_X1 U1535 ( .A(n2800), .B(DATAIN[17]), .S(n77), .Z(n3224) );
  MUX2_X1 U1536 ( .A(n2821), .B(DATAIN[16]), .S(n77), .Z(n3223) );
  MUX2_X1 U1537 ( .A(n2842), .B(DATAIN[15]), .S(n77), .Z(n3222) );
  MUX2_X1 U1538 ( .A(n2863), .B(DATAIN[14]), .S(n77), .Z(n3221) );
  MUX2_X1 U1539 ( .A(n2884), .B(DATAIN[13]), .S(n77), .Z(n3220) );
  MUX2_X1 U1540 ( .A(n2905), .B(DATAIN[12]), .S(n77), .Z(n3219) );
  MUX2_X1 U1541 ( .A(n2926), .B(DATAIN[11]), .S(n76), .Z(n3218) );
  MUX2_X1 U1542 ( .A(n2947), .B(DATAIN[10]), .S(n76), .Z(n3217) );
  MUX2_X1 U1543 ( .A(n2968), .B(DATAIN[9]), .S(n76), .Z(n3216) );
  MUX2_X1 U1544 ( .A(n3565), .B(DATAIN[8]), .S(n76), .Z(n3215) );
  MUX2_X1 U1545 ( .A(n3586), .B(DATAIN[7]), .S(n76), .Z(n3214) );
  MUX2_X1 U1546 ( .A(n3607), .B(DATAIN[6]), .S(n76), .Z(n3213) );
  MUX2_X1 U1547 ( .A(n3628), .B(DATAIN[5]), .S(n76), .Z(n3212) );
  MUX2_X1 U1548 ( .A(n3649), .B(DATAIN[4]), .S(n76), .Z(n3211) );
  MUX2_X1 U1549 ( .A(n3670), .B(DATAIN[3]), .S(n76), .Z(n3210) );
  MUX2_X1 U1550 ( .A(n3691), .B(DATAIN[2]), .S(n76), .Z(n3209) );
  MUX2_X1 U1551 ( .A(n3712), .B(DATAIN[1]), .S(n76), .Z(n3208) );
  MUX2_X1 U1552 ( .A(n3733), .B(DATAIN[0]), .S(n76), .Z(n3207) );
  AND2_X1 U1553 ( .A1(n841), .A2(n773), .ZN(n956) );
  AND3_X1 U1554 ( .A1(ADD_WR[2]), .A2(n953), .A3(ADD_WR[1]), .ZN(n773) );
  MUX2_X1 U1555 ( .A(n2505), .B(DATAIN[31]), .S(n81), .Z(n3206) );
  MUX2_X1 U1556 ( .A(n2526), .B(DATAIN[30]), .S(n81), .Z(n3205) );
  MUX2_X1 U1557 ( .A(n2547), .B(DATAIN[29]), .S(n81), .Z(n3204) );
  MUX2_X1 U1558 ( .A(n2568), .B(DATAIN[28]), .S(n81), .Z(n3203) );
  MUX2_X1 U1559 ( .A(n2589), .B(DATAIN[27]), .S(n81), .Z(n3202) );
  MUX2_X1 U1560 ( .A(n2610), .B(DATAIN[26]), .S(n81), .Z(n3201) );
  MUX2_X1 U1561 ( .A(n2631), .B(DATAIN[25]), .S(n81), .Z(n3200) );
  MUX2_X1 U1562 ( .A(n2652), .B(DATAIN[24]), .S(n81), .Z(n3199) );
  MUX2_X1 U1563 ( .A(n2673), .B(DATAIN[23]), .S(n80), .Z(n3198) );
  MUX2_X1 U1564 ( .A(n2694), .B(DATAIN[22]), .S(n80), .Z(n3197) );
  MUX2_X1 U1565 ( .A(n2715), .B(DATAIN[21]), .S(n80), .Z(n3196) );
  MUX2_X1 U1566 ( .A(n2736), .B(DATAIN[20]), .S(n80), .Z(n3195) );
  MUX2_X1 U1567 ( .A(n2757), .B(DATAIN[19]), .S(n80), .Z(n3194) );
  MUX2_X1 U1568 ( .A(n2778), .B(DATAIN[18]), .S(n80), .Z(n3193) );
  MUX2_X1 U1569 ( .A(n2799), .B(DATAIN[17]), .S(n80), .Z(n3192) );
  MUX2_X1 U1570 ( .A(n2820), .B(DATAIN[16]), .S(n80), .Z(n3191) );
  MUX2_X1 U1571 ( .A(n2841), .B(DATAIN[15]), .S(n80), .Z(n3190) );
  MUX2_X1 U1572 ( .A(n2862), .B(DATAIN[14]), .S(n80), .Z(n3189) );
  MUX2_X1 U1573 ( .A(n2883), .B(DATAIN[13]), .S(n80), .Z(n3188) );
  MUX2_X1 U1574 ( .A(n2904), .B(DATAIN[12]), .S(n80), .Z(n3187) );
  MUX2_X1 U1575 ( .A(n2925), .B(DATAIN[11]), .S(n79), .Z(n3186) );
  MUX2_X1 U1576 ( .A(n2946), .B(DATAIN[10]), .S(n79), .Z(n3185) );
  MUX2_X1 U1577 ( .A(n2967), .B(DATAIN[9]), .S(n79), .Z(n3184) );
  MUX2_X1 U1578 ( .A(n3564), .B(DATAIN[8]), .S(n79), .Z(n3183) );
  MUX2_X1 U1579 ( .A(n3585), .B(DATAIN[7]), .S(n79), .Z(n3182) );
  MUX2_X1 U1580 ( .A(n3606), .B(DATAIN[6]), .S(n79), .Z(n3181) );
  MUX2_X1 U1581 ( .A(n3627), .B(DATAIN[5]), .S(n79), .Z(n3180) );
  MUX2_X1 U1582 ( .A(n3648), .B(DATAIN[4]), .S(n79), .Z(n3179) );
  MUX2_X1 U1583 ( .A(n3669), .B(DATAIN[3]), .S(n79), .Z(n3178) );
  MUX2_X1 U1584 ( .A(n3690), .B(DATAIN[2]), .S(n79), .Z(n3177) );
  MUX2_X1 U1585 ( .A(n3711), .B(DATAIN[1]), .S(n79), .Z(n3176) );
  MUX2_X1 U1586 ( .A(n3732), .B(DATAIN[0]), .S(n79), .Z(n3175) );
  AND2_X1 U1587 ( .A1(n841), .A2(n807), .ZN(n957) );
  AND3_X1 U1588 ( .A1(ADD_WR[2]), .A2(ADD_WR[0]), .A3(ADD_WR[1]), .ZN(n807) );
  AND3_X1 U1589 ( .A1(n947), .A2(n945), .A3(ADD_WR[4]), .ZN(n841) );
  INV_X1 U1590 ( .A(ADD_WR[3]), .ZN(n945) );
  MUX2_X1 U1591 ( .A(n2503), .B(DATAIN[31]), .S(n84), .Z(n3174) );
  MUX2_X1 U1592 ( .A(n2524), .B(DATAIN[30]), .S(n84), .Z(n3173) );
  MUX2_X1 U1593 ( .A(n2545), .B(DATAIN[29]), .S(n84), .Z(n3172) );
  MUX2_X1 U1594 ( .A(n2566), .B(DATAIN[28]), .S(n84), .Z(n3171) );
  MUX2_X1 U1595 ( .A(n2587), .B(DATAIN[27]), .S(n84), .Z(n3170) );
  MUX2_X1 U1596 ( .A(n2608), .B(DATAIN[26]), .S(n84), .Z(n3169) );
  MUX2_X1 U1597 ( .A(n2629), .B(DATAIN[25]), .S(n84), .Z(n3168) );
  MUX2_X1 U1598 ( .A(n2650), .B(DATAIN[24]), .S(n84), .Z(n3167) );
  MUX2_X1 U1599 ( .A(n2671), .B(DATAIN[23]), .S(n83), .Z(n3166) );
  MUX2_X1 U1600 ( .A(n2692), .B(DATAIN[22]), .S(n83), .Z(n3165) );
  MUX2_X1 U1601 ( .A(n2713), .B(DATAIN[21]), .S(n83), .Z(n3164) );
  MUX2_X1 U1602 ( .A(n2734), .B(DATAIN[20]), .S(n83), .Z(n3163) );
  MUX2_X1 U1603 ( .A(n2755), .B(DATAIN[19]), .S(n83), .Z(n3162) );
  MUX2_X1 U1604 ( .A(n2776), .B(DATAIN[18]), .S(n83), .Z(n3161) );
  MUX2_X1 U1605 ( .A(n2797), .B(DATAIN[17]), .S(n83), .Z(n3160) );
  MUX2_X1 U1606 ( .A(n2818), .B(DATAIN[16]), .S(n83), .Z(n3159) );
  MUX2_X1 U1607 ( .A(n2839), .B(DATAIN[15]), .S(n83), .Z(n3158) );
  MUX2_X1 U1608 ( .A(n2860), .B(DATAIN[14]), .S(n83), .Z(n3157) );
  MUX2_X1 U1609 ( .A(n2881), .B(DATAIN[13]), .S(n83), .Z(n3156) );
  MUX2_X1 U1610 ( .A(n2902), .B(DATAIN[12]), .S(n83), .Z(n3155) );
  MUX2_X1 U1611 ( .A(n2923), .B(DATAIN[11]), .S(n82), .Z(n3154) );
  MUX2_X1 U1612 ( .A(n2944), .B(DATAIN[10]), .S(n82), .Z(n3153) );
  MUX2_X1 U1613 ( .A(n2965), .B(DATAIN[9]), .S(n82), .Z(n3152) );
  MUX2_X1 U1614 ( .A(n3562), .B(DATAIN[8]), .S(n82), .Z(n3151) );
  MUX2_X1 U1615 ( .A(n3583), .B(DATAIN[7]), .S(n82), .Z(n3150) );
  MUX2_X1 U1616 ( .A(n3604), .B(DATAIN[6]), .S(n82), .Z(n3149) );
  MUX2_X1 U1617 ( .A(n3625), .B(DATAIN[5]), .S(n82), .Z(n3148) );
  MUX2_X1 U1618 ( .A(n3646), .B(DATAIN[4]), .S(n82), .Z(n3147) );
  MUX2_X1 U1619 ( .A(n3667), .B(DATAIN[3]), .S(n82), .Z(n3146) );
  MUX2_X1 U1620 ( .A(n3688), .B(DATAIN[2]), .S(n82), .Z(n3145) );
  MUX2_X1 U1621 ( .A(n3709), .B(DATAIN[1]), .S(n82), .Z(n3144) );
  MUX2_X1 U1622 ( .A(n3730), .B(DATAIN[0]), .S(n82), .Z(n3143) );
  AND2_X1 U1623 ( .A1(n704), .A2(n468), .ZN(n958) );
  NOR3_X1 U1624 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(ADD_WR[0]), .ZN(n468) );
  MUX2_X1 U1625 ( .A(n2502), .B(DATAIN[31]), .S(n87), .Z(n3142) );
  MUX2_X1 U1626 ( .A(n2523), .B(DATAIN[30]), .S(n87), .Z(n3141) );
  MUX2_X1 U1627 ( .A(n2544), .B(DATAIN[29]), .S(n87), .Z(n3140) );
  MUX2_X1 U1628 ( .A(n2565), .B(DATAIN[28]), .S(n87), .Z(n3139) );
  MUX2_X1 U1629 ( .A(n2586), .B(DATAIN[27]), .S(n87), .Z(n3138) );
  MUX2_X1 U1630 ( .A(n2607), .B(DATAIN[26]), .S(n87), .Z(n3137) );
  MUX2_X1 U1631 ( .A(n2628), .B(DATAIN[25]), .S(n87), .Z(n3136) );
  MUX2_X1 U1632 ( .A(n2649), .B(DATAIN[24]), .S(n87), .Z(n3135) );
  MUX2_X1 U1633 ( .A(n2670), .B(DATAIN[23]), .S(n86), .Z(n3134) );
  MUX2_X1 U1634 ( .A(n2691), .B(DATAIN[22]), .S(n86), .Z(n3133) );
  MUX2_X1 U1635 ( .A(n2712), .B(DATAIN[21]), .S(n86), .Z(n3132) );
  MUX2_X1 U1636 ( .A(n2733), .B(DATAIN[20]), .S(n86), .Z(n3131) );
  MUX2_X1 U1637 ( .A(n2754), .B(DATAIN[19]), .S(n86), .Z(n3130) );
  MUX2_X1 U1638 ( .A(n2775), .B(DATAIN[18]), .S(n86), .Z(n3129) );
  MUX2_X1 U1639 ( .A(n2796), .B(DATAIN[17]), .S(n86), .Z(n3128) );
  MUX2_X1 U1640 ( .A(n2817), .B(DATAIN[16]), .S(n86), .Z(n3127) );
  MUX2_X1 U1641 ( .A(n2838), .B(DATAIN[15]), .S(n86), .Z(n3126) );
  MUX2_X1 U1642 ( .A(n2859), .B(DATAIN[14]), .S(n86), .Z(n3125) );
  MUX2_X1 U1643 ( .A(n2880), .B(DATAIN[13]), .S(n86), .Z(n3124) );
  MUX2_X1 U1644 ( .A(n2901), .B(DATAIN[12]), .S(n86), .Z(n3123) );
  MUX2_X1 U1645 ( .A(n2922), .B(DATAIN[11]), .S(n85), .Z(n3122) );
  MUX2_X1 U1646 ( .A(n2943), .B(DATAIN[10]), .S(n85), .Z(n3121) );
  MUX2_X1 U1647 ( .A(n2964), .B(DATAIN[9]), .S(n85), .Z(n3120) );
  MUX2_X1 U1648 ( .A(n3561), .B(DATAIN[8]), .S(n85), .Z(n3119) );
  MUX2_X1 U1649 ( .A(n3582), .B(DATAIN[7]), .S(n85), .Z(n3118) );
  MUX2_X1 U1650 ( .A(n3603), .B(DATAIN[6]), .S(n85), .Z(n3117) );
  MUX2_X1 U1651 ( .A(n3624), .B(DATAIN[5]), .S(n85), .Z(n3116) );
  MUX2_X1 U1652 ( .A(n3645), .B(DATAIN[4]), .S(n85), .Z(n3115) );
  MUX2_X1 U1653 ( .A(n3666), .B(DATAIN[3]), .S(n85), .Z(n3114) );
  MUX2_X1 U1654 ( .A(n3687), .B(DATAIN[2]), .S(n85), .Z(n3113) );
  MUX2_X1 U1655 ( .A(n3708), .B(DATAIN[1]), .S(n85), .Z(n3112) );
  MUX2_X1 U1656 ( .A(n3729), .B(DATAIN[0]), .S(n85), .Z(n3111) );
  AND2_X1 U1657 ( .A1(n704), .A2(n502), .ZN(n959) );
  NOR3_X1 U1658 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(n953), .ZN(n502) );
  MUX2_X1 U1659 ( .A(n3832), .B(DATAIN[31]), .S(n90), .Z(n3110) );
  MUX2_X1 U1660 ( .A(n3831), .B(DATAIN[30]), .S(n90), .Z(n3109) );
  MUX2_X1 U1661 ( .A(n3830), .B(DATAIN[29]), .S(n90), .Z(n3108) );
  MUX2_X1 U1662 ( .A(n3829), .B(DATAIN[28]), .S(n90), .Z(n3107) );
  MUX2_X1 U1663 ( .A(n3828), .B(DATAIN[27]), .S(n90), .Z(n3106) );
  MUX2_X1 U1664 ( .A(n3827), .B(DATAIN[26]), .S(n90), .Z(n3105) );
  MUX2_X1 U1665 ( .A(n3826), .B(DATAIN[25]), .S(n90), .Z(n3104) );
  MUX2_X1 U1666 ( .A(n3825), .B(DATAIN[24]), .S(n90), .Z(n3103) );
  MUX2_X1 U1667 ( .A(n3824), .B(DATAIN[23]), .S(n89), .Z(n3102) );
  MUX2_X1 U1668 ( .A(n3823), .B(DATAIN[22]), .S(n89), .Z(n3101) );
  MUX2_X1 U1669 ( .A(n3822), .B(DATAIN[21]), .S(n89), .Z(n3100) );
  MUX2_X1 U1670 ( .A(n3821), .B(DATAIN[20]), .S(n89), .Z(n3099) );
  MUX2_X1 U1671 ( .A(n3820), .B(DATAIN[19]), .S(n89), .Z(n3098) );
  MUX2_X1 U1672 ( .A(n3819), .B(DATAIN[18]), .S(n89), .Z(n3097) );
  MUX2_X1 U1673 ( .A(n3818), .B(DATAIN[17]), .S(n89), .Z(n3096) );
  MUX2_X1 U1674 ( .A(n3817), .B(DATAIN[16]), .S(n89), .Z(n3095) );
  MUX2_X1 U1675 ( .A(n3816), .B(DATAIN[15]), .S(n89), .Z(n3094) );
  MUX2_X1 U1676 ( .A(n3815), .B(DATAIN[14]), .S(n89), .Z(n3093) );
  MUX2_X1 U1677 ( .A(n3814), .B(DATAIN[13]), .S(n89), .Z(n3092) );
  MUX2_X1 U1678 ( .A(n3813), .B(DATAIN[12]), .S(n89), .Z(n3091) );
  MUX2_X1 U1679 ( .A(n3812), .B(DATAIN[11]), .S(n88), .Z(n3090) );
  MUX2_X1 U1680 ( .A(n3811), .B(DATAIN[10]), .S(n88), .Z(n3089) );
  MUX2_X1 U1681 ( .A(n3810), .B(DATAIN[9]), .S(n88), .Z(n3088) );
  MUX2_X1 U1682 ( .A(n3809), .B(DATAIN[8]), .S(n88), .Z(n3087) );
  MUX2_X1 U1683 ( .A(n3808), .B(DATAIN[7]), .S(n88), .Z(n3086) );
  MUX2_X1 U1684 ( .A(n3807), .B(DATAIN[6]), .S(n88), .Z(n3085) );
  MUX2_X1 U1685 ( .A(n3806), .B(DATAIN[5]), .S(n88), .Z(n3084) );
  MUX2_X1 U1686 ( .A(n3805), .B(DATAIN[4]), .S(n88), .Z(n3083) );
  MUX2_X1 U1687 ( .A(n3804), .B(DATAIN[3]), .S(n88), .Z(n3082) );
  MUX2_X1 U1688 ( .A(n3803), .B(DATAIN[2]), .S(n88), .Z(n3081) );
  MUX2_X1 U1689 ( .A(n3802), .B(DATAIN[1]), .S(n88), .Z(n3080) );
  MUX2_X1 U1690 ( .A(n3801), .B(DATAIN[0]), .S(n88), .Z(n3079) );
  AND2_X1 U1691 ( .A1(n704), .A2(n536), .ZN(n960) );
  NOR3_X1 U1692 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(n954), .ZN(n536) );
  MUX2_X1 U1693 ( .A(n3800), .B(DATAIN[31]), .S(n93), .Z(n3078) );
  MUX2_X1 U1694 ( .A(n3799), .B(DATAIN[30]), .S(n93), .Z(n3077) );
  MUX2_X1 U1695 ( .A(n3798), .B(DATAIN[29]), .S(n93), .Z(n3076) );
  MUX2_X1 U1696 ( .A(n3797), .B(DATAIN[28]), .S(n93), .Z(n3075) );
  MUX2_X1 U1697 ( .A(n3796), .B(DATAIN[27]), .S(n93), .Z(n3074) );
  MUX2_X1 U1698 ( .A(n3795), .B(DATAIN[26]), .S(n93), .Z(n3073) );
  MUX2_X1 U1699 ( .A(n3794), .B(DATAIN[25]), .S(n93), .Z(n3072) );
  MUX2_X1 U1700 ( .A(n3793), .B(DATAIN[24]), .S(n93), .Z(n3071) );
  MUX2_X1 U1701 ( .A(n3792), .B(DATAIN[23]), .S(n92), .Z(n3070) );
  MUX2_X1 U1702 ( .A(n3791), .B(DATAIN[22]), .S(n92), .Z(n3069) );
  MUX2_X1 U1703 ( .A(n3790), .B(DATAIN[21]), .S(n92), .Z(n3068) );
  MUX2_X1 U1704 ( .A(n3789), .B(DATAIN[20]), .S(n92), .Z(n3067) );
  MUX2_X1 U1705 ( .A(n3788), .B(DATAIN[19]), .S(n92), .Z(n3066) );
  MUX2_X1 U1706 ( .A(n3787), .B(DATAIN[18]), .S(n92), .Z(n3065) );
  MUX2_X1 U1707 ( .A(n3786), .B(DATAIN[17]), .S(n92), .Z(n3064) );
  MUX2_X1 U1708 ( .A(n3785), .B(DATAIN[16]), .S(n92), .Z(n3063) );
  MUX2_X1 U1709 ( .A(n3784), .B(DATAIN[15]), .S(n92), .Z(n3062) );
  MUX2_X1 U1710 ( .A(n3783), .B(DATAIN[14]), .S(n92), .Z(n3061) );
  MUX2_X1 U1711 ( .A(n3782), .B(DATAIN[13]), .S(n92), .Z(n3060) );
  MUX2_X1 U1712 ( .A(n3781), .B(DATAIN[12]), .S(n92), .Z(n3059) );
  MUX2_X1 U1713 ( .A(n3780), .B(DATAIN[11]), .S(n91), .Z(n3058) );
  MUX2_X1 U1714 ( .A(n3779), .B(DATAIN[10]), .S(n91), .Z(n3057) );
  MUX2_X1 U1715 ( .A(n3778), .B(DATAIN[9]), .S(n91), .Z(n3056) );
  MUX2_X1 U1716 ( .A(n3777), .B(DATAIN[8]), .S(n91), .Z(n3055) );
  MUX2_X1 U1717 ( .A(n3776), .B(DATAIN[7]), .S(n91), .Z(n3054) );
  MUX2_X1 U1718 ( .A(n3775), .B(DATAIN[6]), .S(n91), .Z(n3053) );
  MUX2_X1 U1719 ( .A(n3774), .B(DATAIN[5]), .S(n91), .Z(n3052) );
  MUX2_X1 U1720 ( .A(n3773), .B(DATAIN[4]), .S(n91), .Z(n3051) );
  MUX2_X1 U1721 ( .A(n3772), .B(DATAIN[3]), .S(n91), .Z(n3050) );
  MUX2_X1 U1722 ( .A(n3771), .B(DATAIN[2]), .S(n91), .Z(n3049) );
  MUX2_X1 U1723 ( .A(n3770), .B(DATAIN[1]), .S(n91), .Z(n3048) );
  MUX2_X1 U1724 ( .A(n3769), .B(DATAIN[0]), .S(n91), .Z(n3047) );
  AND2_X1 U1725 ( .A1(n704), .A2(n570), .ZN(n961) );
  NOR3_X1 U1726 ( .A1(n953), .A2(ADD_WR[1]), .A3(n954), .ZN(n570) );
  INV_X1 U1727 ( .A(ADD_WR[2]), .ZN(n954) );
  AND3_X1 U1728 ( .A1(ADD_WR[3]), .A2(n947), .A3(ADD_WR[4]), .ZN(n704) );
  AND2_X1 U1729 ( .A1(WR), .A2(ENABLE), .ZN(n947) );
  OAI222_X1 U1730 ( .A1(n298), .A2(n96), .B1(n963), .B2(n99), .C1(n3716), .C2(
        n102), .ZN(n3046) );
  NOR4_X1 U1731 ( .A1(n966), .A2(n967), .A3(n968), .A4(n969), .ZN(n963) );
  OAI221_X1 U1732 ( .B1(n3833), .B2(n105), .C1(n971), .C2(n108), .A(n973), 
        .ZN(n969) );
  AOI22_X1 U1733 ( .A1(n111), .A2(n3730), .B1(n114), .B2(n673), .ZN(n973) );
  OAI221_X1 U1734 ( .B1(n976), .B2(n117), .C1(n3737), .C2(n120), .A(n979), 
        .ZN(n968) );
  AOI22_X1 U1735 ( .A1(n123), .A2(n774), .B1(n126), .B2(n3729), .ZN(n979) );
  OAI211_X1 U1736 ( .C1(n3734), .C2(n129), .A(n983), .B(n984), .ZN(n967) );
  AOI221_X1 U1737 ( .B1(n132), .B2(n908), .C1(n135), .C2(n3735), .A(n987), 
        .ZN(n984) );
  OAI22_X1 U1738 ( .A1(n3731), .A2(n138), .B1(n989), .B2(n141), .ZN(n987) );
  AOI22_X1 U1739 ( .A1(n144), .A2(n3736), .B1(n147), .B2(n808), .ZN(n983) );
  NAND4_X1 U1740 ( .A1(n993), .A2(n994), .A3(n995), .A4(n996), .ZN(n966) );
  AOI221_X1 U1741 ( .B1(n150), .B2(n3719), .C1(n153), .C2(n3720), .A(n999), 
        .ZN(n996) );
  OAI22_X1 U1742 ( .A1(n3718), .A2(n156), .B1(n3717), .B2(n159), .ZN(n999) );
  AOI221_X1 U1743 ( .B1(n162), .B2(n3723), .C1(n165), .C2(n3724), .A(n1004), 
        .ZN(n995) );
  OAI22_X1 U1744 ( .A1(n3722), .A2(n168), .B1(n3721), .B2(n171), .ZN(n1004) );
  AOI221_X1 U1745 ( .B1(n174), .B2(n605), .C1(n177), .C2(n638), .A(n1009), 
        .ZN(n994) );
  OAI22_X1 U1746 ( .A1(n1010), .A2(n180), .B1(n1012), .B2(n183), .ZN(n1009) );
  AOI221_X1 U1747 ( .B1(n186), .B2(n571), .C1(n189), .C2(n3769), .A(n1016), 
        .ZN(n993) );
  OAI22_X1 U1748 ( .A1(n1017), .A2(n192), .B1(n1019), .B2(n195), .ZN(n1016) );
  OAI222_X1 U1749 ( .A1(n299), .A2(n96), .B1(n1021), .B2(n99), .C1(n3695), 
        .C2(n102), .ZN(n3045) );
  NOR4_X1 U1750 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1021)
         );
  OAI221_X1 U1751 ( .B1(n3834), .B2(n105), .C1(n1026), .C2(n108), .A(n1027), 
        .ZN(n1025) );
  AOI22_X1 U1752 ( .A1(n111), .A2(n3709), .B1(n114), .B2(n674), .ZN(n1027) );
  OAI221_X1 U1753 ( .B1(n1028), .B2(n117), .C1(n3738), .C2(n120), .A(n1029), 
        .ZN(n1024) );
  AOI22_X1 U1754 ( .A1(n123), .A2(n776), .B1(n126), .B2(n3708), .ZN(n1029) );
  OAI211_X1 U1755 ( .C1(n3713), .C2(n129), .A(n1030), .B(n1031), .ZN(n1023) );
  AOI221_X1 U1756 ( .B1(n132), .B2(n910), .C1(n135), .C2(n3714), .A(n1032), 
        .ZN(n1031) );
  OAI22_X1 U1757 ( .A1(n3710), .A2(n138), .B1(n1033), .B2(n141), .ZN(n1032) );
  AOI22_X1 U1758 ( .A1(n144), .A2(n3715), .B1(n147), .B2(n810), .ZN(n1030) );
  NAND4_X1 U1759 ( .A1(n1034), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1022)
         );
  AOI221_X1 U1760 ( .B1(n150), .B2(n3698), .C1(n153), .C2(n3699), .A(n1038), 
        .ZN(n1037) );
  OAI22_X1 U1761 ( .A1(n3697), .A2(n156), .B1(n3696), .B2(n159), .ZN(n1038) );
  AOI221_X1 U1762 ( .B1(n162), .B2(n3702), .C1(n165), .C2(n3703), .A(n1039), 
        .ZN(n1036) );
  OAI22_X1 U1763 ( .A1(n3701), .A2(n168), .B1(n3700), .B2(n171), .ZN(n1039) );
  AOI221_X1 U1764 ( .B1(n174), .B2(n607), .C1(n177), .C2(n640), .A(n1040), 
        .ZN(n1035) );
  OAI22_X1 U1765 ( .A1(n1041), .A2(n180), .B1(n1042), .B2(n183), .ZN(n1040) );
  AOI221_X1 U1766 ( .B1(n186), .B2(n573), .C1(n189), .C2(n3770), .A(n1043), 
        .ZN(n1034) );
  OAI22_X1 U1767 ( .A1(n1044), .A2(n192), .B1(n1045), .B2(n195), .ZN(n1043) );
  OAI222_X1 U1768 ( .A1(n300), .A2(n96), .B1(n1046), .B2(n99), .C1(n3674), 
        .C2(n102), .ZN(n3044) );
  NOR4_X1 U1769 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046)
         );
  OAI221_X1 U1770 ( .B1(n3835), .B2(n105), .C1(n1051), .C2(n108), .A(n1052), 
        .ZN(n1050) );
  AOI22_X1 U1771 ( .A1(n111), .A2(n3688), .B1(n114), .B2(n675), .ZN(n1052) );
  OAI221_X1 U1772 ( .B1(n1053), .B2(n117), .C1(n3739), .C2(n120), .A(n1054), 
        .ZN(n1049) );
  AOI22_X1 U1773 ( .A1(n123), .A2(n777), .B1(n126), .B2(n3687), .ZN(n1054) );
  OAI211_X1 U1774 ( .C1(n3692), .C2(n129), .A(n1055), .B(n1056), .ZN(n1048) );
  AOI221_X1 U1775 ( .B1(n132), .B2(n911), .C1(n135), .C2(n3693), .A(n1057), 
        .ZN(n1056) );
  OAI22_X1 U1776 ( .A1(n3689), .A2(n138), .B1(n1058), .B2(n141), .ZN(n1057) );
  AOI22_X1 U1777 ( .A1(n144), .A2(n3694), .B1(n147), .B2(n811), .ZN(n1055) );
  NAND4_X1 U1778 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1047)
         );
  AOI221_X1 U1779 ( .B1(n150), .B2(n3677), .C1(n153), .C2(n3678), .A(n1063), 
        .ZN(n1062) );
  OAI22_X1 U1780 ( .A1(n3676), .A2(n156), .B1(n3675), .B2(n159), .ZN(n1063) );
  AOI221_X1 U1781 ( .B1(n162), .B2(n3681), .C1(n165), .C2(n3682), .A(n1064), 
        .ZN(n1061) );
  OAI22_X1 U1782 ( .A1(n3680), .A2(n168), .B1(n3679), .B2(n171), .ZN(n1064) );
  AOI221_X1 U1783 ( .B1(n174), .B2(n608), .C1(n177), .C2(n641), .A(n1065), 
        .ZN(n1060) );
  OAI22_X1 U1784 ( .A1(n1066), .A2(n180), .B1(n1067), .B2(n183), .ZN(n1065) );
  AOI221_X1 U1785 ( .B1(n186), .B2(n574), .C1(n189), .C2(n3771), .A(n1068), 
        .ZN(n1059) );
  OAI22_X1 U1786 ( .A1(n1069), .A2(n192), .B1(n1070), .B2(n195), .ZN(n1068) );
  OAI222_X1 U1787 ( .A1(n301), .A2(n96), .B1(n1071), .B2(n99), .C1(n3653), 
        .C2(n102), .ZN(n3043) );
  NOR4_X1 U1788 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1071)
         );
  OAI221_X1 U1789 ( .B1(n3836), .B2(n105), .C1(n1076), .C2(n108), .A(n1077), 
        .ZN(n1075) );
  AOI22_X1 U1790 ( .A1(n111), .A2(n3667), .B1(n114), .B2(n676), .ZN(n1077) );
  OAI221_X1 U1791 ( .B1(n1078), .B2(n117), .C1(n3740), .C2(n120), .A(n1079), 
        .ZN(n1074) );
  AOI22_X1 U1792 ( .A1(n123), .A2(n778), .B1(n126), .B2(n3666), .ZN(n1079) );
  OAI211_X1 U1793 ( .C1(n3671), .C2(n129), .A(n1080), .B(n1081), .ZN(n1073) );
  AOI221_X1 U1794 ( .B1(n132), .B2(n912), .C1(n135), .C2(n3672), .A(n1082), 
        .ZN(n1081) );
  OAI22_X1 U1795 ( .A1(n3668), .A2(n138), .B1(n1083), .B2(n141), .ZN(n1082) );
  AOI22_X1 U1796 ( .A1(n144), .A2(n3673), .B1(n147), .B2(n812), .ZN(n1080) );
  NAND4_X1 U1797 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1072)
         );
  AOI221_X1 U1798 ( .B1(n150), .B2(n3656), .C1(n153), .C2(n3657), .A(n1088), 
        .ZN(n1087) );
  OAI22_X1 U1799 ( .A1(n3655), .A2(n156), .B1(n3654), .B2(n159), .ZN(n1088) );
  AOI221_X1 U1800 ( .B1(n162), .B2(n3660), .C1(n165), .C2(n3661), .A(n1089), 
        .ZN(n1086) );
  OAI22_X1 U1801 ( .A1(n3659), .A2(n168), .B1(n3658), .B2(n171), .ZN(n1089) );
  AOI221_X1 U1802 ( .B1(n174), .B2(n609), .C1(n177), .C2(n642), .A(n1090), 
        .ZN(n1085) );
  OAI22_X1 U1803 ( .A1(n1091), .A2(n180), .B1(n1092), .B2(n183), .ZN(n1090) );
  AOI221_X1 U1804 ( .B1(n186), .B2(n575), .C1(n189), .C2(n3772), .A(n1093), 
        .ZN(n1084) );
  OAI22_X1 U1805 ( .A1(n1094), .A2(n192), .B1(n1095), .B2(n195), .ZN(n1093) );
  OAI222_X1 U1806 ( .A1(n302), .A2(n96), .B1(n1096), .B2(n99), .C1(n3632), 
        .C2(n102), .ZN(n3042) );
  NOR4_X1 U1807 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1096)
         );
  OAI221_X1 U1808 ( .B1(n3837), .B2(n105), .C1(n1101), .C2(n108), .A(n1102), 
        .ZN(n1100) );
  AOI22_X1 U1809 ( .A1(n111), .A2(n3646), .B1(n114), .B2(n677), .ZN(n1102) );
  OAI221_X1 U1810 ( .B1(n1103), .B2(n117), .C1(n3741), .C2(n120), .A(n1104), 
        .ZN(n1099) );
  AOI22_X1 U1811 ( .A1(n123), .A2(n779), .B1(n126), .B2(n3645), .ZN(n1104) );
  OAI211_X1 U1812 ( .C1(n3650), .C2(n129), .A(n1105), .B(n1106), .ZN(n1098) );
  AOI221_X1 U1813 ( .B1(n132), .B2(n913), .C1(n135), .C2(n3651), .A(n1107), 
        .ZN(n1106) );
  OAI22_X1 U1814 ( .A1(n3647), .A2(n138), .B1(n1108), .B2(n141), .ZN(n1107) );
  AOI22_X1 U1815 ( .A1(n144), .A2(n3652), .B1(n147), .B2(n813), .ZN(n1105) );
  NAND4_X1 U1816 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1097)
         );
  AOI221_X1 U1817 ( .B1(n150), .B2(n3635), .C1(n153), .C2(n3636), .A(n1113), 
        .ZN(n1112) );
  OAI22_X1 U1818 ( .A1(n3634), .A2(n156), .B1(n3633), .B2(n159), .ZN(n1113) );
  AOI221_X1 U1819 ( .B1(n162), .B2(n3639), .C1(n165), .C2(n3640), .A(n1114), 
        .ZN(n1111) );
  OAI22_X1 U1820 ( .A1(n3638), .A2(n168), .B1(n3637), .B2(n171), .ZN(n1114) );
  AOI221_X1 U1821 ( .B1(n174), .B2(n610), .C1(n177), .C2(n643), .A(n1115), 
        .ZN(n1110) );
  OAI22_X1 U1822 ( .A1(n1116), .A2(n180), .B1(n1117), .B2(n183), .ZN(n1115) );
  AOI221_X1 U1823 ( .B1(n186), .B2(n576), .C1(n189), .C2(n3773), .A(n1118), 
        .ZN(n1109) );
  OAI22_X1 U1824 ( .A1(n1119), .A2(n192), .B1(n1120), .B2(n195), .ZN(n1118) );
  OAI222_X1 U1825 ( .A1(n303), .A2(n96), .B1(n1121), .B2(n99), .C1(n3611), 
        .C2(n102), .ZN(n3041) );
  NOR4_X1 U1826 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1121)
         );
  OAI221_X1 U1827 ( .B1(n3838), .B2(n105), .C1(n1126), .C2(n108), .A(n1127), 
        .ZN(n1125) );
  AOI22_X1 U1828 ( .A1(n111), .A2(n3625), .B1(n114), .B2(n678), .ZN(n1127) );
  OAI221_X1 U1829 ( .B1(n1128), .B2(n117), .C1(n3742), .C2(n120), .A(n1129), 
        .ZN(n1124) );
  AOI22_X1 U1830 ( .A1(n123), .A2(n780), .B1(n126), .B2(n3624), .ZN(n1129) );
  OAI211_X1 U1831 ( .C1(n3629), .C2(n129), .A(n1130), .B(n1131), .ZN(n1123) );
  AOI221_X1 U1832 ( .B1(n132), .B2(n914), .C1(n135), .C2(n3630), .A(n1132), 
        .ZN(n1131) );
  OAI22_X1 U1833 ( .A1(n3626), .A2(n138), .B1(n1133), .B2(n141), .ZN(n1132) );
  AOI22_X1 U1834 ( .A1(n144), .A2(n3631), .B1(n147), .B2(n814), .ZN(n1130) );
  NAND4_X1 U1835 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1122)
         );
  AOI221_X1 U1836 ( .B1(n150), .B2(n3614), .C1(n153), .C2(n3615), .A(n1138), 
        .ZN(n1137) );
  OAI22_X1 U1837 ( .A1(n3613), .A2(n156), .B1(n3612), .B2(n159), .ZN(n1138) );
  AOI221_X1 U1838 ( .B1(n162), .B2(n3618), .C1(n165), .C2(n3619), .A(n1139), 
        .ZN(n1136) );
  OAI22_X1 U1839 ( .A1(n3617), .A2(n168), .B1(n3616), .B2(n171), .ZN(n1139) );
  AOI221_X1 U1840 ( .B1(n174), .B2(n611), .C1(n177), .C2(n644), .A(n1140), 
        .ZN(n1135) );
  OAI22_X1 U1841 ( .A1(n1141), .A2(n180), .B1(n1142), .B2(n183), .ZN(n1140) );
  AOI221_X1 U1842 ( .B1(n186), .B2(n577), .C1(n189), .C2(n3774), .A(n1143), 
        .ZN(n1134) );
  OAI22_X1 U1843 ( .A1(n1144), .A2(n192), .B1(n1145), .B2(n195), .ZN(n1143) );
  OAI222_X1 U1844 ( .A1(n304), .A2(n96), .B1(n1146), .B2(n99), .C1(n3590), 
        .C2(n102), .ZN(n3040) );
  NOR4_X1 U1845 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1146)
         );
  OAI221_X1 U1846 ( .B1(n3839), .B2(n105), .C1(n1151), .C2(n108), .A(n1152), 
        .ZN(n1150) );
  AOI22_X1 U1847 ( .A1(n111), .A2(n3604), .B1(n114), .B2(n679), .ZN(n1152) );
  OAI221_X1 U1848 ( .B1(n1153), .B2(n117), .C1(n3743), .C2(n120), .A(n1154), 
        .ZN(n1149) );
  AOI22_X1 U1849 ( .A1(n123), .A2(n781), .B1(n126), .B2(n3603), .ZN(n1154) );
  OAI211_X1 U1850 ( .C1(n3608), .C2(n129), .A(n1155), .B(n1156), .ZN(n1148) );
  AOI221_X1 U1851 ( .B1(n132), .B2(n915), .C1(n135), .C2(n3609), .A(n1157), 
        .ZN(n1156) );
  OAI22_X1 U1852 ( .A1(n3605), .A2(n138), .B1(n1158), .B2(n141), .ZN(n1157) );
  AOI22_X1 U1853 ( .A1(n144), .A2(n3610), .B1(n147), .B2(n815), .ZN(n1155) );
  NAND4_X1 U1854 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1147)
         );
  AOI221_X1 U1855 ( .B1(n150), .B2(n3593), .C1(n153), .C2(n3594), .A(n1163), 
        .ZN(n1162) );
  OAI22_X1 U1856 ( .A1(n3592), .A2(n156), .B1(n3591), .B2(n159), .ZN(n1163) );
  AOI221_X1 U1857 ( .B1(n162), .B2(n3597), .C1(n165), .C2(n3598), .A(n1164), 
        .ZN(n1161) );
  OAI22_X1 U1858 ( .A1(n3596), .A2(n168), .B1(n3595), .B2(n171), .ZN(n1164) );
  AOI221_X1 U1859 ( .B1(n174), .B2(n612), .C1(n177), .C2(n645), .A(n1165), 
        .ZN(n1160) );
  OAI22_X1 U1860 ( .A1(n1166), .A2(n180), .B1(n1167), .B2(n183), .ZN(n1165) );
  AOI221_X1 U1861 ( .B1(n186), .B2(n578), .C1(n189), .C2(n3775), .A(n1168), 
        .ZN(n1159) );
  OAI22_X1 U1862 ( .A1(n1169), .A2(n192), .B1(n1170), .B2(n195), .ZN(n1168) );
  OAI222_X1 U1863 ( .A1(n305), .A2(n96), .B1(n1171), .B2(n99), .C1(n3569), 
        .C2(n102), .ZN(n3039) );
  NOR4_X1 U1864 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1171)
         );
  OAI221_X1 U1865 ( .B1(n3840), .B2(n105), .C1(n1176), .C2(n108), .A(n1177), 
        .ZN(n1175) );
  AOI22_X1 U1866 ( .A1(n111), .A2(n3583), .B1(n114), .B2(n680), .ZN(n1177) );
  OAI221_X1 U1867 ( .B1(n1178), .B2(n117), .C1(n3744), .C2(n120), .A(n1179), 
        .ZN(n1174) );
  AOI22_X1 U1868 ( .A1(n123), .A2(n782), .B1(n126), .B2(n3582), .ZN(n1179) );
  OAI211_X1 U1869 ( .C1(n3587), .C2(n129), .A(n1180), .B(n1181), .ZN(n1173) );
  AOI221_X1 U1870 ( .B1(n132), .B2(n916), .C1(n135), .C2(n3588), .A(n1182), 
        .ZN(n1181) );
  OAI22_X1 U1871 ( .A1(n3584), .A2(n138), .B1(n1183), .B2(n141), .ZN(n1182) );
  AOI22_X1 U1872 ( .A1(n144), .A2(n3589), .B1(n147), .B2(n816), .ZN(n1180) );
  NAND4_X1 U1873 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1172)
         );
  AOI221_X1 U1874 ( .B1(n150), .B2(n3572), .C1(n153), .C2(n3573), .A(n1188), 
        .ZN(n1187) );
  OAI22_X1 U1875 ( .A1(n3571), .A2(n156), .B1(n3570), .B2(n159), .ZN(n1188) );
  AOI221_X1 U1876 ( .B1(n162), .B2(n3576), .C1(n165), .C2(n3577), .A(n1189), 
        .ZN(n1186) );
  OAI22_X1 U1877 ( .A1(n3575), .A2(n168), .B1(n3574), .B2(n171), .ZN(n1189) );
  AOI221_X1 U1878 ( .B1(n174), .B2(n613), .C1(n177), .C2(n646), .A(n1190), 
        .ZN(n1185) );
  OAI22_X1 U1879 ( .A1(n1191), .A2(n180), .B1(n1192), .B2(n183), .ZN(n1190) );
  AOI221_X1 U1880 ( .B1(n186), .B2(n579), .C1(n189), .C2(n3776), .A(n1193), 
        .ZN(n1184) );
  OAI22_X1 U1881 ( .A1(n1194), .A2(n192), .B1(n1195), .B2(n195), .ZN(n1193) );
  OAI222_X1 U1882 ( .A1(n306), .A2(n95), .B1(n1196), .B2(n98), .C1(n2972), 
        .C2(n102), .ZN(n3038) );
  NOR4_X1 U1883 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1196)
         );
  OAI221_X1 U1884 ( .B1(n3841), .B2(n104), .C1(n1201), .C2(n107), .A(n1202), 
        .ZN(n1200) );
  AOI22_X1 U1885 ( .A1(n110), .A2(n3562), .B1(n113), .B2(n681), .ZN(n1202) );
  OAI221_X1 U1886 ( .B1(n1203), .B2(n116), .C1(n3745), .C2(n119), .A(n1204), 
        .ZN(n1199) );
  AOI22_X1 U1887 ( .A1(n122), .A2(n783), .B1(n125), .B2(n3561), .ZN(n1204) );
  OAI211_X1 U1888 ( .C1(n3566), .C2(n128), .A(n1205), .B(n1206), .ZN(n1198) );
  AOI221_X1 U1889 ( .B1(n131), .B2(n917), .C1(n134), .C2(n3567), .A(n1207), 
        .ZN(n1206) );
  OAI22_X1 U1890 ( .A1(n3563), .A2(n137), .B1(n1208), .B2(n140), .ZN(n1207) );
  AOI22_X1 U1891 ( .A1(n143), .A2(n3568), .B1(n146), .B2(n817), .ZN(n1205) );
  NAND4_X1 U1892 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1197)
         );
  AOI221_X1 U1893 ( .B1(n149), .B2(n2975), .C1(n152), .C2(n2976), .A(n1213), 
        .ZN(n1212) );
  OAI22_X1 U1894 ( .A1(n2974), .A2(n155), .B1(n2973), .B2(n158), .ZN(n1213) );
  AOI221_X1 U1895 ( .B1(n161), .B2(n2979), .C1(n164), .C2(n2980), .A(n1214), 
        .ZN(n1211) );
  OAI22_X1 U1896 ( .A1(n2978), .A2(n167), .B1(n2977), .B2(n170), .ZN(n1214) );
  AOI221_X1 U1897 ( .B1(n173), .B2(n614), .C1(n176), .C2(n647), .A(n1215), 
        .ZN(n1210) );
  OAI22_X1 U1898 ( .A1(n1216), .A2(n179), .B1(n1217), .B2(n182), .ZN(n1215) );
  AOI221_X1 U1899 ( .B1(n185), .B2(n580), .C1(n188), .C2(n3777), .A(n1218), 
        .ZN(n1209) );
  OAI22_X1 U1900 ( .A1(n1219), .A2(n191), .B1(n1220), .B2(n194), .ZN(n1218) );
  OAI222_X1 U1901 ( .A1(n307), .A2(n95), .B1(n1221), .B2(n98), .C1(n2951), 
        .C2(n102), .ZN(n3037) );
  NOR4_X1 U1902 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1221)
         );
  OAI221_X1 U1903 ( .B1(n3842), .B2(n104), .C1(n1226), .C2(n107), .A(n1227), 
        .ZN(n1225) );
  AOI22_X1 U1904 ( .A1(n110), .A2(n2965), .B1(n113), .B2(n682), .ZN(n1227) );
  OAI221_X1 U1905 ( .B1(n1228), .B2(n116), .C1(n3746), .C2(n119), .A(n1229), 
        .ZN(n1224) );
  AOI22_X1 U1906 ( .A1(n122), .A2(n784), .B1(n125), .B2(n2964), .ZN(n1229) );
  OAI211_X1 U1907 ( .C1(n2969), .C2(n128), .A(n1230), .B(n1231), .ZN(n1223) );
  AOI221_X1 U1908 ( .B1(n131), .B2(n918), .C1(n134), .C2(n2970), .A(n1232), 
        .ZN(n1231) );
  OAI22_X1 U1909 ( .A1(n2966), .A2(n137), .B1(n1233), .B2(n140), .ZN(n1232) );
  AOI22_X1 U1910 ( .A1(n143), .A2(n2971), .B1(n146), .B2(n818), .ZN(n1230) );
  NAND4_X1 U1911 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1222)
         );
  AOI221_X1 U1912 ( .B1(n149), .B2(n2954), .C1(n152), .C2(n2955), .A(n1238), 
        .ZN(n1237) );
  OAI22_X1 U1913 ( .A1(n2953), .A2(n155), .B1(n2952), .B2(n158), .ZN(n1238) );
  AOI221_X1 U1914 ( .B1(n161), .B2(n2958), .C1(n164), .C2(n2959), .A(n1239), 
        .ZN(n1236) );
  OAI22_X1 U1915 ( .A1(n2957), .A2(n167), .B1(n2956), .B2(n170), .ZN(n1239) );
  AOI221_X1 U1916 ( .B1(n173), .B2(n615), .C1(n176), .C2(n648), .A(n1240), 
        .ZN(n1235) );
  OAI22_X1 U1917 ( .A1(n1241), .A2(n179), .B1(n1242), .B2(n182), .ZN(n1240) );
  AOI221_X1 U1918 ( .B1(n185), .B2(n581), .C1(n188), .C2(n3778), .A(n1243), 
        .ZN(n1234) );
  OAI22_X1 U1919 ( .A1(n1244), .A2(n191), .B1(n1245), .B2(n194), .ZN(n1243) );
  OAI222_X1 U1920 ( .A1(n308), .A2(n95), .B1(n1246), .B2(n98), .C1(n2930), 
        .C2(n101), .ZN(n3036) );
  NOR4_X1 U1921 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1246)
         );
  OAI221_X1 U1922 ( .B1(n3843), .B2(n104), .C1(n1251), .C2(n107), .A(n1252), 
        .ZN(n1250) );
  AOI22_X1 U1923 ( .A1(n110), .A2(n2944), .B1(n113), .B2(n683), .ZN(n1252) );
  OAI221_X1 U1924 ( .B1(n1253), .B2(n116), .C1(n3747), .C2(n119), .A(n1254), 
        .ZN(n1249) );
  AOI22_X1 U1925 ( .A1(n122), .A2(n785), .B1(n125), .B2(n2943), .ZN(n1254) );
  OAI211_X1 U1926 ( .C1(n2948), .C2(n128), .A(n1255), .B(n1256), .ZN(n1248) );
  AOI221_X1 U1927 ( .B1(n131), .B2(n919), .C1(n134), .C2(n2949), .A(n1257), 
        .ZN(n1256) );
  OAI22_X1 U1928 ( .A1(n2945), .A2(n137), .B1(n1258), .B2(n140), .ZN(n1257) );
  AOI22_X1 U1929 ( .A1(n143), .A2(n2950), .B1(n146), .B2(n819), .ZN(n1255) );
  NAND4_X1 U1930 ( .A1(n1259), .A2(n1260), .A3(n1261), .A4(n1262), .ZN(n1247)
         );
  AOI221_X1 U1931 ( .B1(n149), .B2(n2933), .C1(n152), .C2(n2934), .A(n1263), 
        .ZN(n1262) );
  OAI22_X1 U1932 ( .A1(n2932), .A2(n155), .B1(n2931), .B2(n158), .ZN(n1263) );
  AOI221_X1 U1933 ( .B1(n161), .B2(n2937), .C1(n164), .C2(n2938), .A(n1264), 
        .ZN(n1261) );
  OAI22_X1 U1934 ( .A1(n2936), .A2(n167), .B1(n2935), .B2(n170), .ZN(n1264) );
  AOI221_X1 U1935 ( .B1(n173), .B2(n616), .C1(n176), .C2(n649), .A(n1265), 
        .ZN(n1260) );
  OAI22_X1 U1936 ( .A1(n1266), .A2(n179), .B1(n1267), .B2(n182), .ZN(n1265) );
  AOI221_X1 U1937 ( .B1(n185), .B2(n582), .C1(n188), .C2(n3779), .A(n1268), 
        .ZN(n1259) );
  OAI22_X1 U1938 ( .A1(n1269), .A2(n191), .B1(n1270), .B2(n194), .ZN(n1268) );
  OAI222_X1 U1939 ( .A1(n309), .A2(n95), .B1(n1271), .B2(n98), .C1(n2909), 
        .C2(n101), .ZN(n3035) );
  NOR4_X1 U1940 ( .A1(n1272), .A2(n1273), .A3(n1274), .A4(n1275), .ZN(n1271)
         );
  OAI221_X1 U1941 ( .B1(n3844), .B2(n104), .C1(n1276), .C2(n107), .A(n1277), 
        .ZN(n1275) );
  AOI22_X1 U1942 ( .A1(n110), .A2(n2923), .B1(n113), .B2(n684), .ZN(n1277) );
  OAI221_X1 U1943 ( .B1(n1278), .B2(n116), .C1(n3748), .C2(n119), .A(n1279), 
        .ZN(n1274) );
  AOI22_X1 U1944 ( .A1(n122), .A2(n786), .B1(n125), .B2(n2922), .ZN(n1279) );
  OAI211_X1 U1945 ( .C1(n2927), .C2(n128), .A(n1280), .B(n1281), .ZN(n1273) );
  AOI221_X1 U1946 ( .B1(n131), .B2(n920), .C1(n134), .C2(n2928), .A(n1282), 
        .ZN(n1281) );
  OAI22_X1 U1947 ( .A1(n2924), .A2(n137), .B1(n1283), .B2(n140), .ZN(n1282) );
  AOI22_X1 U1948 ( .A1(n143), .A2(n2929), .B1(n146), .B2(n820), .ZN(n1280) );
  NAND4_X1 U1949 ( .A1(n1284), .A2(n1285), .A3(n1286), .A4(n1287), .ZN(n1272)
         );
  AOI221_X1 U1950 ( .B1(n149), .B2(n2912), .C1(n152), .C2(n2913), .A(n1288), 
        .ZN(n1287) );
  OAI22_X1 U1951 ( .A1(n2911), .A2(n155), .B1(n2910), .B2(n158), .ZN(n1288) );
  AOI221_X1 U1952 ( .B1(n161), .B2(n2916), .C1(n164), .C2(n2917), .A(n1289), 
        .ZN(n1286) );
  OAI22_X1 U1953 ( .A1(n2915), .A2(n167), .B1(n2914), .B2(n170), .ZN(n1289) );
  AOI221_X1 U1954 ( .B1(n173), .B2(n617), .C1(n176), .C2(n650), .A(n1290), 
        .ZN(n1285) );
  OAI22_X1 U1955 ( .A1(n1291), .A2(n179), .B1(n1292), .B2(n182), .ZN(n1290) );
  AOI221_X1 U1956 ( .B1(n185), .B2(n583), .C1(n188), .C2(n3780), .A(n1293), 
        .ZN(n1284) );
  OAI22_X1 U1957 ( .A1(n1294), .A2(n191), .B1(n1295), .B2(n194), .ZN(n1293) );
  OAI222_X1 U1958 ( .A1(n310), .A2(n95), .B1(n1296), .B2(n98), .C1(n2888), 
        .C2(n101), .ZN(n3034) );
  NOR4_X1 U1959 ( .A1(n1297), .A2(n1298), .A3(n1299), .A4(n1300), .ZN(n1296)
         );
  OAI221_X1 U1960 ( .B1(n3845), .B2(n104), .C1(n1301), .C2(n107), .A(n1302), 
        .ZN(n1300) );
  AOI22_X1 U1961 ( .A1(n110), .A2(n2902), .B1(n113), .B2(n685), .ZN(n1302) );
  OAI221_X1 U1962 ( .B1(n1303), .B2(n116), .C1(n3749), .C2(n119), .A(n1304), 
        .ZN(n1299) );
  AOI22_X1 U1963 ( .A1(n122), .A2(n787), .B1(n125), .B2(n2901), .ZN(n1304) );
  OAI211_X1 U1964 ( .C1(n2906), .C2(n128), .A(n1305), .B(n1306), .ZN(n1298) );
  AOI221_X1 U1965 ( .B1(n131), .B2(n921), .C1(n134), .C2(n2907), .A(n1307), 
        .ZN(n1306) );
  OAI22_X1 U1966 ( .A1(n2903), .A2(n137), .B1(n1308), .B2(n140), .ZN(n1307) );
  AOI22_X1 U1967 ( .A1(n143), .A2(n2908), .B1(n146), .B2(n821), .ZN(n1305) );
  NAND4_X1 U1968 ( .A1(n1309), .A2(n1310), .A3(n1311), .A4(n1312), .ZN(n1297)
         );
  AOI221_X1 U1969 ( .B1(n149), .B2(n2891), .C1(n152), .C2(n2892), .A(n1313), 
        .ZN(n1312) );
  OAI22_X1 U1970 ( .A1(n2890), .A2(n155), .B1(n2889), .B2(n158), .ZN(n1313) );
  AOI221_X1 U1971 ( .B1(n161), .B2(n2895), .C1(n164), .C2(n2896), .A(n1314), 
        .ZN(n1311) );
  OAI22_X1 U1972 ( .A1(n2894), .A2(n167), .B1(n2893), .B2(n170), .ZN(n1314) );
  AOI221_X1 U1973 ( .B1(n173), .B2(n618), .C1(n176), .C2(n651), .A(n1315), 
        .ZN(n1310) );
  OAI22_X1 U1974 ( .A1(n1316), .A2(n179), .B1(n1317), .B2(n182), .ZN(n1315) );
  AOI221_X1 U1975 ( .B1(n185), .B2(n584), .C1(n188), .C2(n3781), .A(n1318), 
        .ZN(n1309) );
  OAI22_X1 U1976 ( .A1(n1319), .A2(n191), .B1(n1320), .B2(n194), .ZN(n1318) );
  OAI222_X1 U1977 ( .A1(n311), .A2(n95), .B1(n1321), .B2(n98), .C1(n2867), 
        .C2(n101), .ZN(n3033) );
  NOR4_X1 U1978 ( .A1(n1322), .A2(n1323), .A3(n1324), .A4(n1325), .ZN(n1321)
         );
  OAI221_X1 U1979 ( .B1(n3846), .B2(n104), .C1(n1326), .C2(n107), .A(n1327), 
        .ZN(n1325) );
  AOI22_X1 U1980 ( .A1(n110), .A2(n2881), .B1(n113), .B2(n686), .ZN(n1327) );
  OAI221_X1 U1981 ( .B1(n1328), .B2(n116), .C1(n3750), .C2(n119), .A(n1329), 
        .ZN(n1324) );
  AOI22_X1 U1982 ( .A1(n122), .A2(n788), .B1(n125), .B2(n2880), .ZN(n1329) );
  OAI211_X1 U1983 ( .C1(n2885), .C2(n128), .A(n1330), .B(n1331), .ZN(n1323) );
  AOI221_X1 U1984 ( .B1(n131), .B2(n922), .C1(n134), .C2(n2886), .A(n1332), 
        .ZN(n1331) );
  OAI22_X1 U1985 ( .A1(n2882), .A2(n137), .B1(n1333), .B2(n140), .ZN(n1332) );
  AOI22_X1 U1986 ( .A1(n143), .A2(n2887), .B1(n146), .B2(n822), .ZN(n1330) );
  NAND4_X1 U1987 ( .A1(n1334), .A2(n1335), .A3(n1336), .A4(n1337), .ZN(n1322)
         );
  AOI221_X1 U1988 ( .B1(n149), .B2(n2870), .C1(n152), .C2(n2871), .A(n1338), 
        .ZN(n1337) );
  OAI22_X1 U1989 ( .A1(n2869), .A2(n155), .B1(n2868), .B2(n158), .ZN(n1338) );
  AOI221_X1 U1990 ( .B1(n161), .B2(n2874), .C1(n164), .C2(n2875), .A(n1339), 
        .ZN(n1336) );
  OAI22_X1 U1991 ( .A1(n2873), .A2(n167), .B1(n2872), .B2(n170), .ZN(n1339) );
  AOI221_X1 U1992 ( .B1(n173), .B2(n619), .C1(n176), .C2(n652), .A(n1340), 
        .ZN(n1335) );
  OAI22_X1 U1993 ( .A1(n1341), .A2(n179), .B1(n1342), .B2(n182), .ZN(n1340) );
  AOI221_X1 U1994 ( .B1(n185), .B2(n585), .C1(n188), .C2(n3782), .A(n1343), 
        .ZN(n1334) );
  OAI22_X1 U1995 ( .A1(n1344), .A2(n191), .B1(n1345), .B2(n194), .ZN(n1343) );
  OAI222_X1 U1996 ( .A1(n312), .A2(n95), .B1(n1346), .B2(n98), .C1(n2846), 
        .C2(n101), .ZN(n3032) );
  NOR4_X1 U1997 ( .A1(n1347), .A2(n1348), .A3(n1349), .A4(n1350), .ZN(n1346)
         );
  OAI221_X1 U1998 ( .B1(n3847), .B2(n104), .C1(n1351), .C2(n107), .A(n1352), 
        .ZN(n1350) );
  AOI22_X1 U1999 ( .A1(n110), .A2(n2860), .B1(n113), .B2(n687), .ZN(n1352) );
  OAI221_X1 U2000 ( .B1(n1353), .B2(n116), .C1(n3751), .C2(n119), .A(n1354), 
        .ZN(n1349) );
  AOI22_X1 U2001 ( .A1(n122), .A2(n789), .B1(n125), .B2(n2859), .ZN(n1354) );
  OAI211_X1 U2002 ( .C1(n2864), .C2(n128), .A(n1355), .B(n1356), .ZN(n1348) );
  AOI221_X1 U2003 ( .B1(n131), .B2(n923), .C1(n134), .C2(n2865), .A(n1357), 
        .ZN(n1356) );
  OAI22_X1 U2004 ( .A1(n2861), .A2(n137), .B1(n1358), .B2(n140), .ZN(n1357) );
  AOI22_X1 U2005 ( .A1(n143), .A2(n2866), .B1(n146), .B2(n823), .ZN(n1355) );
  NAND4_X1 U2006 ( .A1(n1359), .A2(n1360), .A3(n1361), .A4(n1362), .ZN(n1347)
         );
  AOI221_X1 U2007 ( .B1(n149), .B2(n2849), .C1(n152), .C2(n2850), .A(n1363), 
        .ZN(n1362) );
  OAI22_X1 U2008 ( .A1(n2848), .A2(n155), .B1(n2847), .B2(n158), .ZN(n1363) );
  AOI221_X1 U2009 ( .B1(n161), .B2(n2853), .C1(n164), .C2(n2854), .A(n1364), 
        .ZN(n1361) );
  OAI22_X1 U2010 ( .A1(n2852), .A2(n167), .B1(n2851), .B2(n170), .ZN(n1364) );
  AOI221_X1 U2011 ( .B1(n173), .B2(n620), .C1(n176), .C2(n653), .A(n1365), 
        .ZN(n1360) );
  OAI22_X1 U2012 ( .A1(n1366), .A2(n179), .B1(n1367), .B2(n182), .ZN(n1365) );
  AOI221_X1 U2013 ( .B1(n185), .B2(n586), .C1(n188), .C2(n3783), .A(n1368), 
        .ZN(n1359) );
  OAI22_X1 U2014 ( .A1(n1369), .A2(n191), .B1(n1370), .B2(n194), .ZN(n1368) );
  OAI222_X1 U2015 ( .A1(n313), .A2(n95), .B1(n1371), .B2(n98), .C1(n2825), 
        .C2(n101), .ZN(n3031) );
  NOR4_X1 U2016 ( .A1(n1372), .A2(n1373), .A3(n1374), .A4(n1375), .ZN(n1371)
         );
  OAI221_X1 U2017 ( .B1(n3848), .B2(n104), .C1(n1376), .C2(n107), .A(n1377), 
        .ZN(n1375) );
  AOI22_X1 U2018 ( .A1(n110), .A2(n2839), .B1(n113), .B2(n688), .ZN(n1377) );
  OAI221_X1 U2019 ( .B1(n1378), .B2(n116), .C1(n3752), .C2(n119), .A(n1379), 
        .ZN(n1374) );
  AOI22_X1 U2020 ( .A1(n122), .A2(n790), .B1(n125), .B2(n2838), .ZN(n1379) );
  OAI211_X1 U2021 ( .C1(n2843), .C2(n128), .A(n1380), .B(n1381), .ZN(n1373) );
  AOI221_X1 U2022 ( .B1(n131), .B2(n924), .C1(n134), .C2(n2844), .A(n1382), 
        .ZN(n1381) );
  OAI22_X1 U2023 ( .A1(n2840), .A2(n137), .B1(n1383), .B2(n140), .ZN(n1382) );
  AOI22_X1 U2024 ( .A1(n143), .A2(n2845), .B1(n146), .B2(n824), .ZN(n1380) );
  NAND4_X1 U2025 ( .A1(n1384), .A2(n1385), .A3(n1386), .A4(n1387), .ZN(n1372)
         );
  AOI221_X1 U2026 ( .B1(n149), .B2(n2828), .C1(n152), .C2(n2829), .A(n1388), 
        .ZN(n1387) );
  OAI22_X1 U2027 ( .A1(n2827), .A2(n155), .B1(n2826), .B2(n158), .ZN(n1388) );
  AOI221_X1 U2028 ( .B1(n161), .B2(n2832), .C1(n164), .C2(n2833), .A(n1389), 
        .ZN(n1386) );
  OAI22_X1 U2029 ( .A1(n2831), .A2(n167), .B1(n2830), .B2(n170), .ZN(n1389) );
  AOI221_X1 U2030 ( .B1(n173), .B2(n621), .C1(n176), .C2(n654), .A(n1390), 
        .ZN(n1385) );
  OAI22_X1 U2031 ( .A1(n1391), .A2(n179), .B1(n1392), .B2(n182), .ZN(n1390) );
  AOI221_X1 U2032 ( .B1(n185), .B2(n587), .C1(n188), .C2(n3784), .A(n1393), 
        .ZN(n1384) );
  OAI22_X1 U2033 ( .A1(n1394), .A2(n191), .B1(n1395), .B2(n194), .ZN(n1393) );
  OAI222_X1 U2034 ( .A1(n314), .A2(n95), .B1(n1396), .B2(n98), .C1(n2804), 
        .C2(n101), .ZN(n3030) );
  NOR4_X1 U2035 ( .A1(n1397), .A2(n1398), .A3(n1399), .A4(n1400), .ZN(n1396)
         );
  OAI221_X1 U2036 ( .B1(n3849), .B2(n104), .C1(n1401), .C2(n107), .A(n1402), 
        .ZN(n1400) );
  AOI22_X1 U2037 ( .A1(n110), .A2(n2818), .B1(n113), .B2(n689), .ZN(n1402) );
  OAI221_X1 U2038 ( .B1(n1403), .B2(n116), .C1(n3753), .C2(n119), .A(n1404), 
        .ZN(n1399) );
  AOI22_X1 U2039 ( .A1(n122), .A2(n791), .B1(n125), .B2(n2817), .ZN(n1404) );
  OAI211_X1 U2040 ( .C1(n2822), .C2(n128), .A(n1405), .B(n1406), .ZN(n1398) );
  AOI221_X1 U2041 ( .B1(n131), .B2(n925), .C1(n134), .C2(n2823), .A(n1407), 
        .ZN(n1406) );
  OAI22_X1 U2042 ( .A1(n2819), .A2(n137), .B1(n1408), .B2(n140), .ZN(n1407) );
  AOI22_X1 U2043 ( .A1(n143), .A2(n2824), .B1(n146), .B2(n825), .ZN(n1405) );
  NAND4_X1 U2044 ( .A1(n1409), .A2(n1410), .A3(n1411), .A4(n1412), .ZN(n1397)
         );
  AOI221_X1 U2045 ( .B1(n149), .B2(n2807), .C1(n152), .C2(n2808), .A(n1413), 
        .ZN(n1412) );
  OAI22_X1 U2046 ( .A1(n2806), .A2(n155), .B1(n2805), .B2(n158), .ZN(n1413) );
  AOI221_X1 U2047 ( .B1(n161), .B2(n2811), .C1(n164), .C2(n2812), .A(n1414), 
        .ZN(n1411) );
  OAI22_X1 U2048 ( .A1(n2810), .A2(n167), .B1(n2809), .B2(n170), .ZN(n1414) );
  AOI221_X1 U2049 ( .B1(n173), .B2(n622), .C1(n176), .C2(n655), .A(n1415), 
        .ZN(n1410) );
  OAI22_X1 U2050 ( .A1(n1416), .A2(n179), .B1(n1417), .B2(n182), .ZN(n1415) );
  AOI221_X1 U2051 ( .B1(n185), .B2(n588), .C1(n188), .C2(n3785), .A(n1418), 
        .ZN(n1409) );
  OAI22_X1 U2052 ( .A1(n1419), .A2(n191), .B1(n1420), .B2(n194), .ZN(n1418) );
  OAI222_X1 U2053 ( .A1(n315), .A2(n95), .B1(n1421), .B2(n98), .C1(n2783), 
        .C2(n101), .ZN(n3029) );
  NOR4_X1 U2054 ( .A1(n1422), .A2(n1423), .A3(n1424), .A4(n1425), .ZN(n1421)
         );
  OAI221_X1 U2055 ( .B1(n3850), .B2(n104), .C1(n1426), .C2(n107), .A(n1427), 
        .ZN(n1425) );
  AOI22_X1 U2056 ( .A1(n110), .A2(n2797), .B1(n113), .B2(n690), .ZN(n1427) );
  OAI221_X1 U2057 ( .B1(n1428), .B2(n116), .C1(n3754), .C2(n119), .A(n1429), 
        .ZN(n1424) );
  AOI22_X1 U2058 ( .A1(n122), .A2(n792), .B1(n125), .B2(n2796), .ZN(n1429) );
  OAI211_X1 U2059 ( .C1(n2801), .C2(n128), .A(n1430), .B(n1431), .ZN(n1423) );
  AOI221_X1 U2060 ( .B1(n131), .B2(n926), .C1(n134), .C2(n2802), .A(n1432), 
        .ZN(n1431) );
  OAI22_X1 U2061 ( .A1(n2798), .A2(n137), .B1(n1433), .B2(n140), .ZN(n1432) );
  AOI22_X1 U2062 ( .A1(n143), .A2(n2803), .B1(n146), .B2(n826), .ZN(n1430) );
  NAND4_X1 U2063 ( .A1(n1434), .A2(n1435), .A3(n1436), .A4(n1437), .ZN(n1422)
         );
  AOI221_X1 U2064 ( .B1(n149), .B2(n2786), .C1(n152), .C2(n2787), .A(n1438), 
        .ZN(n1437) );
  OAI22_X1 U2065 ( .A1(n2785), .A2(n155), .B1(n2784), .B2(n158), .ZN(n1438) );
  AOI221_X1 U2066 ( .B1(n161), .B2(n2790), .C1(n164), .C2(n2791), .A(n1439), 
        .ZN(n1436) );
  OAI22_X1 U2067 ( .A1(n2789), .A2(n167), .B1(n2788), .B2(n170), .ZN(n1439) );
  AOI221_X1 U2068 ( .B1(n173), .B2(n623), .C1(n176), .C2(n656), .A(n1440), 
        .ZN(n1435) );
  OAI22_X1 U2069 ( .A1(n1441), .A2(n179), .B1(n1442), .B2(n182), .ZN(n1440) );
  AOI221_X1 U2070 ( .B1(n185), .B2(n589), .C1(n188), .C2(n3786), .A(n1443), 
        .ZN(n1434) );
  OAI22_X1 U2071 ( .A1(n1444), .A2(n191), .B1(n1445), .B2(n194), .ZN(n1443) );
  OAI222_X1 U2072 ( .A1(n316), .A2(n95), .B1(n1446), .B2(n98), .C1(n2762), 
        .C2(n101), .ZN(n3028) );
  NOR4_X1 U2073 ( .A1(n1447), .A2(n1448), .A3(n1449), .A4(n1450), .ZN(n1446)
         );
  OAI221_X1 U2074 ( .B1(n3851), .B2(n104), .C1(n1451), .C2(n107), .A(n1452), 
        .ZN(n1450) );
  AOI22_X1 U2075 ( .A1(n110), .A2(n2776), .B1(n113), .B2(n691), .ZN(n1452) );
  OAI221_X1 U2076 ( .B1(n1453), .B2(n116), .C1(n3755), .C2(n119), .A(n1454), 
        .ZN(n1449) );
  AOI22_X1 U2077 ( .A1(n122), .A2(n793), .B1(n125), .B2(n2775), .ZN(n1454) );
  OAI211_X1 U2078 ( .C1(n2780), .C2(n128), .A(n1455), .B(n1456), .ZN(n1448) );
  AOI221_X1 U2079 ( .B1(n131), .B2(n927), .C1(n134), .C2(n2781), .A(n1457), 
        .ZN(n1456) );
  OAI22_X1 U2080 ( .A1(n2777), .A2(n137), .B1(n1458), .B2(n140), .ZN(n1457) );
  AOI22_X1 U2081 ( .A1(n143), .A2(n2782), .B1(n146), .B2(n827), .ZN(n1455) );
  NAND4_X1 U2082 ( .A1(n1459), .A2(n1460), .A3(n1461), .A4(n1462), .ZN(n1447)
         );
  AOI221_X1 U2083 ( .B1(n149), .B2(n2765), .C1(n152), .C2(n2766), .A(n1463), 
        .ZN(n1462) );
  OAI22_X1 U2084 ( .A1(n2764), .A2(n155), .B1(n2763), .B2(n158), .ZN(n1463) );
  AOI221_X1 U2085 ( .B1(n161), .B2(n2769), .C1(n164), .C2(n2770), .A(n1464), 
        .ZN(n1461) );
  OAI22_X1 U2086 ( .A1(n2768), .A2(n167), .B1(n2767), .B2(n170), .ZN(n1464) );
  AOI221_X1 U2087 ( .B1(n173), .B2(n624), .C1(n176), .C2(n657), .A(n1465), 
        .ZN(n1460) );
  OAI22_X1 U2088 ( .A1(n1466), .A2(n179), .B1(n1467), .B2(n182), .ZN(n1465) );
  AOI221_X1 U2089 ( .B1(n185), .B2(n590), .C1(n188), .C2(n3787), .A(n1468), 
        .ZN(n1459) );
  OAI22_X1 U2090 ( .A1(n1469), .A2(n191), .B1(n1470), .B2(n194), .ZN(n1468) );
  OAI222_X1 U2091 ( .A1(n317), .A2(n95), .B1(n1471), .B2(n98), .C1(n2741), 
        .C2(n101), .ZN(n3027) );
  NOR4_X1 U2092 ( .A1(n1472), .A2(n1473), .A3(n1474), .A4(n1475), .ZN(n1471)
         );
  OAI221_X1 U2093 ( .B1(n3852), .B2(n104), .C1(n1476), .C2(n107), .A(n1477), 
        .ZN(n1475) );
  AOI22_X1 U2094 ( .A1(n110), .A2(n2755), .B1(n113), .B2(n692), .ZN(n1477) );
  OAI221_X1 U2095 ( .B1(n1478), .B2(n116), .C1(n3756), .C2(n119), .A(n1479), 
        .ZN(n1474) );
  AOI22_X1 U2096 ( .A1(n122), .A2(n794), .B1(n125), .B2(n2754), .ZN(n1479) );
  OAI211_X1 U2097 ( .C1(n2759), .C2(n128), .A(n1480), .B(n1481), .ZN(n1473) );
  AOI221_X1 U2098 ( .B1(n131), .B2(n928), .C1(n134), .C2(n2760), .A(n1482), 
        .ZN(n1481) );
  OAI22_X1 U2099 ( .A1(n2756), .A2(n137), .B1(n1483), .B2(n140), .ZN(n1482) );
  AOI22_X1 U2100 ( .A1(n143), .A2(n2761), .B1(n146), .B2(n828), .ZN(n1480) );
  NAND4_X1 U2101 ( .A1(n1484), .A2(n1485), .A3(n1486), .A4(n1487), .ZN(n1472)
         );
  AOI221_X1 U2102 ( .B1(n149), .B2(n2744), .C1(n152), .C2(n2745), .A(n1488), 
        .ZN(n1487) );
  OAI22_X1 U2103 ( .A1(n2743), .A2(n155), .B1(n2742), .B2(n158), .ZN(n1488) );
  AOI221_X1 U2104 ( .B1(n161), .B2(n2748), .C1(n164), .C2(n2749), .A(n1489), 
        .ZN(n1486) );
  OAI22_X1 U2105 ( .A1(n2747), .A2(n167), .B1(n2746), .B2(n170), .ZN(n1489) );
  AOI221_X1 U2106 ( .B1(n173), .B2(n625), .C1(n176), .C2(n658), .A(n1490), 
        .ZN(n1485) );
  OAI22_X1 U2107 ( .A1(n1491), .A2(n179), .B1(n1492), .B2(n182), .ZN(n1490) );
  AOI221_X1 U2108 ( .B1(n185), .B2(n591), .C1(n188), .C2(n3788), .A(n1493), 
        .ZN(n1484) );
  OAI22_X1 U2109 ( .A1(n1494), .A2(n191), .B1(n1495), .B2(n194), .ZN(n1493) );
  OAI222_X1 U2110 ( .A1(n318), .A2(n94), .B1(n1496), .B2(n97), .C1(n2720), 
        .C2(n101), .ZN(n3026) );
  NOR4_X1 U2111 ( .A1(n1497), .A2(n1498), .A3(n1499), .A4(n1500), .ZN(n1496)
         );
  OAI221_X1 U2112 ( .B1(n3853), .B2(n103), .C1(n1501), .C2(n106), .A(n1502), 
        .ZN(n1500) );
  AOI22_X1 U2113 ( .A1(n109), .A2(n2734), .B1(n112), .B2(n693), .ZN(n1502) );
  OAI221_X1 U2114 ( .B1(n1503), .B2(n115), .C1(n3757), .C2(n118), .A(n1504), 
        .ZN(n1499) );
  AOI22_X1 U2115 ( .A1(n121), .A2(n795), .B1(n124), .B2(n2733), .ZN(n1504) );
  OAI211_X1 U2116 ( .C1(n2738), .C2(n127), .A(n1505), .B(n1506), .ZN(n1498) );
  AOI221_X1 U2117 ( .B1(n130), .B2(n929), .C1(n133), .C2(n2739), .A(n1507), 
        .ZN(n1506) );
  OAI22_X1 U2118 ( .A1(n2735), .A2(n136), .B1(n1508), .B2(n139), .ZN(n1507) );
  AOI22_X1 U2119 ( .A1(n142), .A2(n2740), .B1(n145), .B2(n829), .ZN(n1505) );
  NAND4_X1 U2120 ( .A1(n1509), .A2(n1510), .A3(n1511), .A4(n1512), .ZN(n1497)
         );
  AOI221_X1 U2121 ( .B1(n148), .B2(n2723), .C1(n151), .C2(n2724), .A(n1513), 
        .ZN(n1512) );
  OAI22_X1 U2122 ( .A1(n2722), .A2(n154), .B1(n2721), .B2(n157), .ZN(n1513) );
  AOI221_X1 U2123 ( .B1(n160), .B2(n2727), .C1(n163), .C2(n2728), .A(n1514), 
        .ZN(n1511) );
  OAI22_X1 U2124 ( .A1(n2726), .A2(n166), .B1(n2725), .B2(n169), .ZN(n1514) );
  AOI221_X1 U2125 ( .B1(n172), .B2(n626), .C1(n175), .C2(n659), .A(n1515), 
        .ZN(n1510) );
  OAI22_X1 U2126 ( .A1(n1516), .A2(n178), .B1(n1517), .B2(n181), .ZN(n1515) );
  AOI221_X1 U2127 ( .B1(n184), .B2(n592), .C1(n187), .C2(n3789), .A(n1518), 
        .ZN(n1509) );
  OAI22_X1 U2128 ( .A1(n1519), .A2(n190), .B1(n1520), .B2(n193), .ZN(n1518) );
  OAI222_X1 U2129 ( .A1(n319), .A2(n94), .B1(n1521), .B2(n97), .C1(n2699), 
        .C2(n101), .ZN(n3025) );
  NOR4_X1 U2130 ( .A1(n1522), .A2(n1523), .A3(n1524), .A4(n1525), .ZN(n1521)
         );
  OAI221_X1 U2131 ( .B1(n3854), .B2(n103), .C1(n1526), .C2(n106), .A(n1527), 
        .ZN(n1525) );
  AOI22_X1 U2132 ( .A1(n109), .A2(n2713), .B1(n112), .B2(n694), .ZN(n1527) );
  OAI221_X1 U2133 ( .B1(n1528), .B2(n115), .C1(n3758), .C2(n118), .A(n1529), 
        .ZN(n1524) );
  AOI22_X1 U2134 ( .A1(n121), .A2(n796), .B1(n124), .B2(n2712), .ZN(n1529) );
  OAI211_X1 U2135 ( .C1(n2717), .C2(n127), .A(n1530), .B(n1531), .ZN(n1523) );
  AOI221_X1 U2136 ( .B1(n130), .B2(n930), .C1(n133), .C2(n2718), .A(n1532), 
        .ZN(n1531) );
  OAI22_X1 U2137 ( .A1(n2714), .A2(n136), .B1(n1533), .B2(n139), .ZN(n1532) );
  AOI22_X1 U2138 ( .A1(n142), .A2(n2719), .B1(n145), .B2(n830), .ZN(n1530) );
  NAND4_X1 U2139 ( .A1(n1534), .A2(n1535), .A3(n1536), .A4(n1537), .ZN(n1522)
         );
  AOI221_X1 U2140 ( .B1(n148), .B2(n2702), .C1(n151), .C2(n2703), .A(n1538), 
        .ZN(n1537) );
  OAI22_X1 U2141 ( .A1(n2701), .A2(n154), .B1(n2700), .B2(n157), .ZN(n1538) );
  AOI221_X1 U2142 ( .B1(n160), .B2(n2706), .C1(n163), .C2(n2707), .A(n1539), 
        .ZN(n1536) );
  OAI22_X1 U2143 ( .A1(n2705), .A2(n166), .B1(n2704), .B2(n169), .ZN(n1539) );
  AOI221_X1 U2144 ( .B1(n172), .B2(n627), .C1(n175), .C2(n660), .A(n1540), 
        .ZN(n1535) );
  OAI22_X1 U2145 ( .A1(n1541), .A2(n178), .B1(n1542), .B2(n181), .ZN(n1540) );
  AOI221_X1 U2146 ( .B1(n184), .B2(n593), .C1(n187), .C2(n3790), .A(n1543), 
        .ZN(n1534) );
  OAI22_X1 U2147 ( .A1(n1544), .A2(n190), .B1(n1545), .B2(n193), .ZN(n1543) );
  OAI222_X1 U2148 ( .A1(n320), .A2(n94), .B1(n1546), .B2(n97), .C1(n2678), 
        .C2(n100), .ZN(n3024) );
  NOR4_X1 U2149 ( .A1(n1547), .A2(n1548), .A3(n1549), .A4(n1550), .ZN(n1546)
         );
  OAI221_X1 U2150 ( .B1(n3855), .B2(n103), .C1(n1551), .C2(n106), .A(n1552), 
        .ZN(n1550) );
  AOI22_X1 U2151 ( .A1(n109), .A2(n2692), .B1(n112), .B2(n695), .ZN(n1552) );
  OAI221_X1 U2152 ( .B1(n1553), .B2(n115), .C1(n3759), .C2(n118), .A(n1554), 
        .ZN(n1549) );
  AOI22_X1 U2153 ( .A1(n121), .A2(n797), .B1(n124), .B2(n2691), .ZN(n1554) );
  OAI211_X1 U2154 ( .C1(n2696), .C2(n127), .A(n1555), .B(n1556), .ZN(n1548) );
  AOI221_X1 U2155 ( .B1(n130), .B2(n931), .C1(n133), .C2(n2697), .A(n1557), 
        .ZN(n1556) );
  OAI22_X1 U2156 ( .A1(n2693), .A2(n136), .B1(n1558), .B2(n139), .ZN(n1557) );
  AOI22_X1 U2157 ( .A1(n142), .A2(n2698), .B1(n145), .B2(n831), .ZN(n1555) );
  NAND4_X1 U2158 ( .A1(n1559), .A2(n1560), .A3(n1561), .A4(n1562), .ZN(n1547)
         );
  AOI221_X1 U2159 ( .B1(n148), .B2(n2681), .C1(n151), .C2(n2682), .A(n1563), 
        .ZN(n1562) );
  OAI22_X1 U2160 ( .A1(n2680), .A2(n154), .B1(n2679), .B2(n157), .ZN(n1563) );
  AOI221_X1 U2161 ( .B1(n160), .B2(n2685), .C1(n163), .C2(n2686), .A(n1564), 
        .ZN(n1561) );
  OAI22_X1 U2162 ( .A1(n2684), .A2(n166), .B1(n2683), .B2(n169), .ZN(n1564) );
  AOI221_X1 U2163 ( .B1(n172), .B2(n628), .C1(n175), .C2(n661), .A(n1565), 
        .ZN(n1560) );
  OAI22_X1 U2164 ( .A1(n1566), .A2(n178), .B1(n1567), .B2(n181), .ZN(n1565) );
  AOI221_X1 U2165 ( .B1(n184), .B2(n594), .C1(n187), .C2(n3791), .A(n1568), 
        .ZN(n1559) );
  OAI22_X1 U2166 ( .A1(n1569), .A2(n190), .B1(n1570), .B2(n193), .ZN(n1568) );
  OAI222_X1 U2167 ( .A1(n321), .A2(n94), .B1(n1571), .B2(n97), .C1(n2657), 
        .C2(n100), .ZN(n3023) );
  NOR4_X1 U2168 ( .A1(n1572), .A2(n1573), .A3(n1574), .A4(n1575), .ZN(n1571)
         );
  OAI221_X1 U2169 ( .B1(n3856), .B2(n103), .C1(n1576), .C2(n106), .A(n1577), 
        .ZN(n1575) );
  AOI22_X1 U2170 ( .A1(n109), .A2(n2671), .B1(n112), .B2(n696), .ZN(n1577) );
  OAI221_X1 U2171 ( .B1(n1578), .B2(n115), .C1(n3760), .C2(n118), .A(n1579), 
        .ZN(n1574) );
  AOI22_X1 U2172 ( .A1(n121), .A2(n798), .B1(n124), .B2(n2670), .ZN(n1579) );
  OAI211_X1 U2173 ( .C1(n2675), .C2(n127), .A(n1580), .B(n1581), .ZN(n1573) );
  AOI221_X1 U2174 ( .B1(n130), .B2(n932), .C1(n133), .C2(n2676), .A(n1582), 
        .ZN(n1581) );
  OAI22_X1 U2175 ( .A1(n2672), .A2(n136), .B1(n1583), .B2(n139), .ZN(n1582) );
  AOI22_X1 U2176 ( .A1(n142), .A2(n2677), .B1(n145), .B2(n832), .ZN(n1580) );
  NAND4_X1 U2177 ( .A1(n1584), .A2(n1585), .A3(n1586), .A4(n1587), .ZN(n1572)
         );
  AOI221_X1 U2178 ( .B1(n148), .B2(n2660), .C1(n151), .C2(n2661), .A(n1588), 
        .ZN(n1587) );
  OAI22_X1 U2179 ( .A1(n2659), .A2(n154), .B1(n2658), .B2(n157), .ZN(n1588) );
  AOI221_X1 U2180 ( .B1(n160), .B2(n2664), .C1(n163), .C2(n2665), .A(n1589), 
        .ZN(n1586) );
  OAI22_X1 U2181 ( .A1(n2663), .A2(n166), .B1(n2662), .B2(n169), .ZN(n1589) );
  AOI221_X1 U2182 ( .B1(n172), .B2(n629), .C1(n175), .C2(n662), .A(n1590), 
        .ZN(n1585) );
  OAI22_X1 U2183 ( .A1(n1591), .A2(n178), .B1(n1592), .B2(n181), .ZN(n1590) );
  AOI221_X1 U2184 ( .B1(n184), .B2(n595), .C1(n187), .C2(n3792), .A(n1593), 
        .ZN(n1584) );
  OAI22_X1 U2185 ( .A1(n1594), .A2(n190), .B1(n1595), .B2(n193), .ZN(n1593) );
  OAI222_X1 U2186 ( .A1(n322), .A2(n94), .B1(n1596), .B2(n97), .C1(n2636), 
        .C2(n100), .ZN(n3022) );
  NOR4_X1 U2187 ( .A1(n1597), .A2(n1598), .A3(n1599), .A4(n1600), .ZN(n1596)
         );
  OAI221_X1 U2188 ( .B1(n3857), .B2(n103), .C1(n1601), .C2(n106), .A(n1602), 
        .ZN(n1600) );
  AOI22_X1 U2189 ( .A1(n109), .A2(n2650), .B1(n112), .B2(n697), .ZN(n1602) );
  OAI221_X1 U2190 ( .B1(n1603), .B2(n115), .C1(n3761), .C2(n118), .A(n1604), 
        .ZN(n1599) );
  AOI22_X1 U2191 ( .A1(n121), .A2(n799), .B1(n124), .B2(n2649), .ZN(n1604) );
  OAI211_X1 U2192 ( .C1(n2654), .C2(n127), .A(n1605), .B(n1606), .ZN(n1598) );
  AOI221_X1 U2193 ( .B1(n130), .B2(n933), .C1(n133), .C2(n2655), .A(n1607), 
        .ZN(n1606) );
  OAI22_X1 U2194 ( .A1(n2651), .A2(n136), .B1(n1608), .B2(n139), .ZN(n1607) );
  AOI22_X1 U2195 ( .A1(n142), .A2(n2656), .B1(n145), .B2(n833), .ZN(n1605) );
  NAND4_X1 U2196 ( .A1(n1609), .A2(n1610), .A3(n1611), .A4(n1612), .ZN(n1597)
         );
  AOI221_X1 U2197 ( .B1(n148), .B2(n2639), .C1(n151), .C2(n2640), .A(n1613), 
        .ZN(n1612) );
  OAI22_X1 U2198 ( .A1(n2638), .A2(n154), .B1(n2637), .B2(n157), .ZN(n1613) );
  AOI221_X1 U2199 ( .B1(n160), .B2(n2643), .C1(n163), .C2(n2644), .A(n1614), 
        .ZN(n1611) );
  OAI22_X1 U2200 ( .A1(n2642), .A2(n166), .B1(n2641), .B2(n169), .ZN(n1614) );
  AOI221_X1 U2201 ( .B1(n172), .B2(n630), .C1(n175), .C2(n663), .A(n1615), 
        .ZN(n1610) );
  OAI22_X1 U2202 ( .A1(n1616), .A2(n178), .B1(n1617), .B2(n181), .ZN(n1615) );
  AOI221_X1 U2203 ( .B1(n184), .B2(n596), .C1(n187), .C2(n3793), .A(n1618), 
        .ZN(n1609) );
  OAI22_X1 U2204 ( .A1(n1619), .A2(n190), .B1(n1620), .B2(n193), .ZN(n1618) );
  OAI222_X1 U2205 ( .A1(n323), .A2(n94), .B1(n1621), .B2(n97), .C1(n2615), 
        .C2(n100), .ZN(n3021) );
  NOR4_X1 U2206 ( .A1(n1622), .A2(n1623), .A3(n1624), .A4(n1625), .ZN(n1621)
         );
  OAI221_X1 U2207 ( .B1(n3858), .B2(n103), .C1(n1626), .C2(n106), .A(n1627), 
        .ZN(n1625) );
  AOI22_X1 U2208 ( .A1(n109), .A2(n2629), .B1(n112), .B2(n698), .ZN(n1627) );
  OAI221_X1 U2209 ( .B1(n1628), .B2(n115), .C1(n3762), .C2(n118), .A(n1629), 
        .ZN(n1624) );
  AOI22_X1 U2210 ( .A1(n121), .A2(n800), .B1(n124), .B2(n2628), .ZN(n1629) );
  OAI211_X1 U2211 ( .C1(n2633), .C2(n127), .A(n1630), .B(n1631), .ZN(n1623) );
  AOI221_X1 U2212 ( .B1(n130), .B2(n934), .C1(n133), .C2(n2634), .A(n1632), 
        .ZN(n1631) );
  OAI22_X1 U2213 ( .A1(n2630), .A2(n136), .B1(n1633), .B2(n139), .ZN(n1632) );
  AOI22_X1 U2214 ( .A1(n142), .A2(n2635), .B1(n145), .B2(n834), .ZN(n1630) );
  NAND4_X1 U2215 ( .A1(n1634), .A2(n1635), .A3(n1636), .A4(n1637), .ZN(n1622)
         );
  AOI221_X1 U2216 ( .B1(n148), .B2(n2618), .C1(n151), .C2(n2619), .A(n1638), 
        .ZN(n1637) );
  OAI22_X1 U2217 ( .A1(n2617), .A2(n154), .B1(n2616), .B2(n157), .ZN(n1638) );
  AOI221_X1 U2218 ( .B1(n160), .B2(n2622), .C1(n163), .C2(n2623), .A(n1639), 
        .ZN(n1636) );
  OAI22_X1 U2219 ( .A1(n2621), .A2(n166), .B1(n2620), .B2(n169), .ZN(n1639) );
  AOI221_X1 U2220 ( .B1(n172), .B2(n631), .C1(n175), .C2(n664), .A(n1640), 
        .ZN(n1635) );
  OAI22_X1 U2221 ( .A1(n1641), .A2(n178), .B1(n1642), .B2(n181), .ZN(n1640) );
  AOI221_X1 U2222 ( .B1(n184), .B2(n597), .C1(n187), .C2(n3794), .A(n1643), 
        .ZN(n1634) );
  OAI22_X1 U2223 ( .A1(n1644), .A2(n190), .B1(n1645), .B2(n193), .ZN(n1643) );
  OAI222_X1 U2224 ( .A1(n324), .A2(n94), .B1(n1646), .B2(n97), .C1(n2594), 
        .C2(n100), .ZN(n3020) );
  NOR4_X1 U2225 ( .A1(n1647), .A2(n1648), .A3(n1649), .A4(n1650), .ZN(n1646)
         );
  OAI221_X1 U2226 ( .B1(n3859), .B2(n103), .C1(n1651), .C2(n106), .A(n1652), 
        .ZN(n1650) );
  AOI22_X1 U2227 ( .A1(n109), .A2(n2608), .B1(n112), .B2(n699), .ZN(n1652) );
  OAI221_X1 U2228 ( .B1(n1653), .B2(n115), .C1(n3763), .C2(n118), .A(n1654), 
        .ZN(n1649) );
  AOI22_X1 U2229 ( .A1(n121), .A2(n801), .B1(n124), .B2(n2607), .ZN(n1654) );
  OAI211_X1 U2230 ( .C1(n2612), .C2(n127), .A(n1655), .B(n1656), .ZN(n1648) );
  AOI221_X1 U2231 ( .B1(n130), .B2(n935), .C1(n133), .C2(n2613), .A(n1657), 
        .ZN(n1656) );
  OAI22_X1 U2232 ( .A1(n2609), .A2(n136), .B1(n1658), .B2(n139), .ZN(n1657) );
  AOI22_X1 U2233 ( .A1(n142), .A2(n2614), .B1(n145), .B2(n835), .ZN(n1655) );
  NAND4_X1 U2234 ( .A1(n1659), .A2(n1660), .A3(n1661), .A4(n1662), .ZN(n1647)
         );
  AOI221_X1 U2235 ( .B1(n148), .B2(n2597), .C1(n151), .C2(n2598), .A(n1663), 
        .ZN(n1662) );
  OAI22_X1 U2236 ( .A1(n2596), .A2(n154), .B1(n2595), .B2(n157), .ZN(n1663) );
  AOI221_X1 U2237 ( .B1(n160), .B2(n2601), .C1(n163), .C2(n2602), .A(n1664), 
        .ZN(n1661) );
  OAI22_X1 U2238 ( .A1(n2600), .A2(n166), .B1(n2599), .B2(n169), .ZN(n1664) );
  AOI221_X1 U2239 ( .B1(n172), .B2(n632), .C1(n175), .C2(n665), .A(n1665), 
        .ZN(n1660) );
  OAI22_X1 U2240 ( .A1(n1666), .A2(n178), .B1(n1667), .B2(n181), .ZN(n1665) );
  AOI221_X1 U2241 ( .B1(n184), .B2(n598), .C1(n187), .C2(n3795), .A(n1668), 
        .ZN(n1659) );
  OAI22_X1 U2242 ( .A1(n1669), .A2(n190), .B1(n1670), .B2(n193), .ZN(n1668) );
  OAI222_X1 U2243 ( .A1(n325), .A2(n94), .B1(n1671), .B2(n97), .C1(n2573), 
        .C2(n100), .ZN(n3019) );
  NOR4_X1 U2244 ( .A1(n1672), .A2(n1673), .A3(n1674), .A4(n1675), .ZN(n1671)
         );
  OAI221_X1 U2245 ( .B1(n3860), .B2(n103), .C1(n1676), .C2(n106), .A(n1677), 
        .ZN(n1675) );
  AOI22_X1 U2246 ( .A1(n109), .A2(n2587), .B1(n112), .B2(n700), .ZN(n1677) );
  OAI221_X1 U2247 ( .B1(n1678), .B2(n115), .C1(n3764), .C2(n118), .A(n1679), 
        .ZN(n1674) );
  AOI22_X1 U2248 ( .A1(n121), .A2(n802), .B1(n124), .B2(n2586), .ZN(n1679) );
  OAI211_X1 U2249 ( .C1(n2591), .C2(n127), .A(n1680), .B(n1681), .ZN(n1673) );
  AOI221_X1 U2250 ( .B1(n130), .B2(n936), .C1(n133), .C2(n2592), .A(n1682), 
        .ZN(n1681) );
  OAI22_X1 U2251 ( .A1(n2588), .A2(n136), .B1(n1683), .B2(n139), .ZN(n1682) );
  AOI22_X1 U2252 ( .A1(n142), .A2(n2593), .B1(n145), .B2(n836), .ZN(n1680) );
  NAND4_X1 U2253 ( .A1(n1684), .A2(n1685), .A3(n1686), .A4(n1687), .ZN(n1672)
         );
  AOI221_X1 U2254 ( .B1(n148), .B2(n2576), .C1(n151), .C2(n2577), .A(n1688), 
        .ZN(n1687) );
  OAI22_X1 U2255 ( .A1(n2575), .A2(n154), .B1(n2574), .B2(n157), .ZN(n1688) );
  AOI221_X1 U2256 ( .B1(n160), .B2(n2580), .C1(n163), .C2(n2581), .A(n1689), 
        .ZN(n1686) );
  OAI22_X1 U2257 ( .A1(n2579), .A2(n166), .B1(n2578), .B2(n169), .ZN(n1689) );
  AOI221_X1 U2258 ( .B1(n172), .B2(n633), .C1(n175), .C2(n666), .A(n1690), 
        .ZN(n1685) );
  OAI22_X1 U2259 ( .A1(n1691), .A2(n178), .B1(n1692), .B2(n181), .ZN(n1690) );
  AOI221_X1 U2260 ( .B1(n184), .B2(n599), .C1(n187), .C2(n3796), .A(n1693), 
        .ZN(n1684) );
  OAI22_X1 U2261 ( .A1(n1694), .A2(n190), .B1(n1695), .B2(n193), .ZN(n1693) );
  OAI222_X1 U2262 ( .A1(n326), .A2(n94), .B1(n1696), .B2(n97), .C1(n2552), 
        .C2(n100), .ZN(n3018) );
  NOR4_X1 U2263 ( .A1(n1697), .A2(n1698), .A3(n1699), .A4(n1700), .ZN(n1696)
         );
  OAI221_X1 U2264 ( .B1(n3861), .B2(n103), .C1(n1701), .C2(n106), .A(n1702), 
        .ZN(n1700) );
  AOI22_X1 U2265 ( .A1(n109), .A2(n2566), .B1(n112), .B2(n701), .ZN(n1702) );
  OAI221_X1 U2266 ( .B1(n1703), .B2(n115), .C1(n3765), .C2(n118), .A(n1704), 
        .ZN(n1699) );
  AOI22_X1 U2267 ( .A1(n121), .A2(n803), .B1(n124), .B2(n2565), .ZN(n1704) );
  OAI211_X1 U2268 ( .C1(n2570), .C2(n127), .A(n1705), .B(n1706), .ZN(n1698) );
  AOI221_X1 U2269 ( .B1(n130), .B2(n937), .C1(n133), .C2(n2571), .A(n1707), 
        .ZN(n1706) );
  OAI22_X1 U2270 ( .A1(n2567), .A2(n136), .B1(n1708), .B2(n139), .ZN(n1707) );
  AOI22_X1 U2271 ( .A1(n142), .A2(n2572), .B1(n145), .B2(n837), .ZN(n1705) );
  NAND4_X1 U2272 ( .A1(n1709), .A2(n1710), .A3(n1711), .A4(n1712), .ZN(n1697)
         );
  AOI221_X1 U2273 ( .B1(n148), .B2(n2555), .C1(n151), .C2(n2556), .A(n1713), 
        .ZN(n1712) );
  OAI22_X1 U2274 ( .A1(n2554), .A2(n154), .B1(n2553), .B2(n157), .ZN(n1713) );
  AOI221_X1 U2275 ( .B1(n160), .B2(n2559), .C1(n163), .C2(n2560), .A(n1714), 
        .ZN(n1711) );
  OAI22_X1 U2276 ( .A1(n2558), .A2(n166), .B1(n2557), .B2(n169), .ZN(n1714) );
  AOI221_X1 U2277 ( .B1(n172), .B2(n634), .C1(n175), .C2(n667), .A(n1715), 
        .ZN(n1710) );
  OAI22_X1 U2278 ( .A1(n1716), .A2(n178), .B1(n1717), .B2(n181), .ZN(n1715) );
  AOI221_X1 U2279 ( .B1(n184), .B2(n600), .C1(n187), .C2(n3797), .A(n1718), 
        .ZN(n1709) );
  OAI22_X1 U2280 ( .A1(n1719), .A2(n190), .B1(n1720), .B2(n193), .ZN(n1718) );
  OAI222_X1 U2281 ( .A1(n327), .A2(n94), .B1(n1721), .B2(n97), .C1(n2531), 
        .C2(n100), .ZN(n3017) );
  NOR4_X1 U2282 ( .A1(n1722), .A2(n1723), .A3(n1724), .A4(n1725), .ZN(n1721)
         );
  OAI221_X1 U2283 ( .B1(n3862), .B2(n103), .C1(n1726), .C2(n106), .A(n1727), 
        .ZN(n1725) );
  AOI22_X1 U2284 ( .A1(n109), .A2(n2545), .B1(n112), .B2(n702), .ZN(n1727) );
  OAI221_X1 U2285 ( .B1(n1728), .B2(n115), .C1(n3766), .C2(n118), .A(n1729), 
        .ZN(n1724) );
  AOI22_X1 U2286 ( .A1(n121), .A2(n804), .B1(n124), .B2(n2544), .ZN(n1729) );
  OAI211_X1 U2287 ( .C1(n2549), .C2(n127), .A(n1730), .B(n1731), .ZN(n1723) );
  AOI221_X1 U2288 ( .B1(n130), .B2(n938), .C1(n133), .C2(n2550), .A(n1732), 
        .ZN(n1731) );
  OAI22_X1 U2289 ( .A1(n2546), .A2(n136), .B1(n1733), .B2(n139), .ZN(n1732) );
  AOI22_X1 U2290 ( .A1(n142), .A2(n2551), .B1(n145), .B2(n838), .ZN(n1730) );
  NAND4_X1 U2291 ( .A1(n1734), .A2(n1735), .A3(n1736), .A4(n1737), .ZN(n1722)
         );
  AOI221_X1 U2292 ( .B1(n148), .B2(n2534), .C1(n151), .C2(n2535), .A(n1738), 
        .ZN(n1737) );
  OAI22_X1 U2293 ( .A1(n2533), .A2(n154), .B1(n2532), .B2(n157), .ZN(n1738) );
  AOI221_X1 U2294 ( .B1(n160), .B2(n2538), .C1(n163), .C2(n2539), .A(n1739), 
        .ZN(n1736) );
  OAI22_X1 U2295 ( .A1(n2537), .A2(n166), .B1(n2536), .B2(n169), .ZN(n1739) );
  AOI221_X1 U2296 ( .B1(n172), .B2(n635), .C1(n175), .C2(n668), .A(n1740), 
        .ZN(n1735) );
  OAI22_X1 U2297 ( .A1(n1741), .A2(n178), .B1(n1742), .B2(n181), .ZN(n1740) );
  AOI221_X1 U2298 ( .B1(n184), .B2(n601), .C1(n187), .C2(n3798), .A(n1743), 
        .ZN(n1734) );
  OAI22_X1 U2299 ( .A1(n1744), .A2(n190), .B1(n1745), .B2(n193), .ZN(n1743) );
  OAI222_X1 U2300 ( .A1(n328), .A2(n94), .B1(n1746), .B2(n97), .C1(n2510), 
        .C2(n100), .ZN(n3016) );
  NOR4_X1 U2301 ( .A1(n1747), .A2(n1748), .A3(n1749), .A4(n1750), .ZN(n1746)
         );
  OAI221_X1 U2302 ( .B1(n3863), .B2(n103), .C1(n1751), .C2(n106), .A(n1752), 
        .ZN(n1750) );
  AOI22_X1 U2303 ( .A1(n109), .A2(n2524), .B1(n112), .B2(n703), .ZN(n1752) );
  OAI221_X1 U2304 ( .B1(n1753), .B2(n115), .C1(n3767), .C2(n118), .A(n1754), 
        .ZN(n1749) );
  AOI22_X1 U2305 ( .A1(n121), .A2(n805), .B1(n124), .B2(n2523), .ZN(n1754) );
  OAI211_X1 U2306 ( .C1(n2528), .C2(n127), .A(n1755), .B(n1756), .ZN(n1748) );
  AOI221_X1 U2307 ( .B1(n130), .B2(n939), .C1(n133), .C2(n2529), .A(n1757), 
        .ZN(n1756) );
  OAI22_X1 U2308 ( .A1(n2525), .A2(n136), .B1(n1758), .B2(n139), .ZN(n1757) );
  AOI22_X1 U2309 ( .A1(n142), .A2(n2530), .B1(n145), .B2(n839), .ZN(n1755) );
  NAND4_X1 U2310 ( .A1(n1759), .A2(n1760), .A3(n1761), .A4(n1762), .ZN(n1747)
         );
  AOI221_X1 U2311 ( .B1(n148), .B2(n2513), .C1(n151), .C2(n2514), .A(n1763), 
        .ZN(n1762) );
  OAI22_X1 U2312 ( .A1(n2512), .A2(n154), .B1(n2511), .B2(n157), .ZN(n1763) );
  AOI221_X1 U2313 ( .B1(n160), .B2(n2517), .C1(n163), .C2(n2518), .A(n1764), 
        .ZN(n1761) );
  OAI22_X1 U2314 ( .A1(n2516), .A2(n166), .B1(n2515), .B2(n169), .ZN(n1764) );
  AOI221_X1 U2315 ( .B1(n172), .B2(n636), .C1(n175), .C2(n669), .A(n1765), 
        .ZN(n1760) );
  OAI22_X1 U2316 ( .A1(n1766), .A2(n178), .B1(n1767), .B2(n181), .ZN(n1765) );
  AOI221_X1 U2317 ( .B1(n184), .B2(n602), .C1(n187), .C2(n3799), .A(n1768), 
        .ZN(n1759) );
  OAI22_X1 U2318 ( .A1(n1769), .A2(n190), .B1(n1770), .B2(n193), .ZN(n1768) );
  OAI222_X1 U2319 ( .A1(n329), .A2(n94), .B1(n1771), .B2(n97), .C1(n2489), 
        .C2(n100), .ZN(n3015) );
  NAND2_X1 U2320 ( .A1(n100), .A2(n1772), .ZN(n964) );
  NOR4_X1 U2321 ( .A1(n1773), .A2(n1774), .A3(n1775), .A4(n1776), .ZN(n1771)
         );
  OAI221_X1 U2322 ( .B1(n3864), .B2(n103), .C1(n1777), .C2(n106), .A(n1778), 
        .ZN(n1776) );
  AOI22_X1 U2323 ( .A1(n109), .A2(n2503), .B1(n112), .B2(n671), .ZN(n1778) );
  AND2_X1 U2324 ( .A1(n1779), .A2(n1780), .ZN(n975) );
  AND2_X1 U2325 ( .A1(n1779), .A2(n1781), .ZN(n974) );
  NAND2_X1 U2326 ( .A1(n1782), .A2(n1783), .ZN(n972) );
  NAND2_X1 U2327 ( .A1(n1784), .A2(n1780), .ZN(n970) );
  OAI221_X1 U2328 ( .B1(n1785), .B2(n115), .C1(n3768), .C2(n118), .A(n1786), 
        .ZN(n1775) );
  AOI22_X1 U2329 ( .A1(n121), .A2(n806), .B1(n124), .B2(n2502), .ZN(n1786) );
  AND2_X1 U2330 ( .A1(n1784), .A2(n1781), .ZN(n981) );
  AND2_X1 U2331 ( .A1(n1784), .A2(n1783), .ZN(n980) );
  NAND2_X1 U2332 ( .A1(n1779), .A2(n1783), .ZN(n978) );
  NAND2_X1 U2333 ( .A1(n1779), .A2(n1787), .ZN(n977) );
  NOR3_X1 U2334 ( .A1(n1788), .A2(ADD_RS2[0]), .A3(n1789), .ZN(n1779) );
  OAI211_X1 U2335 ( .C1(n2507), .C2(n127), .A(n1790), .B(n1791), .ZN(n1774) );
  AOI221_X1 U2336 ( .B1(n130), .B2(n940), .C1(n133), .C2(n2508), .A(n1792), 
        .ZN(n1791) );
  OAI22_X1 U2337 ( .A1(n2504), .A2(n136), .B1(n1793), .B2(n139), .ZN(n1792) );
  NAND2_X1 U2338 ( .A1(n1794), .A2(n1783), .ZN(n990) );
  NAND2_X1 U2339 ( .A1(n1794), .A2(n1787), .ZN(n988) );
  AND2_X1 U2340 ( .A1(n1782), .A2(n1780), .ZN(n986) );
  AND2_X1 U2341 ( .A1(n1782), .A2(n1787), .ZN(n985) );
  AOI22_X1 U2342 ( .A1(n142), .A2(n2509), .B1(n145), .B2(n840), .ZN(n1790) );
  AND2_X1 U2343 ( .A1(n1794), .A2(n1781), .ZN(n992) );
  AND2_X1 U2344 ( .A1(n1794), .A2(n1780), .ZN(n991) );
  NOR3_X1 U2345 ( .A1(ADD_RS2[0]), .A2(ADD_RS2[3]), .A3(n1788), .ZN(n1794) );
  NAND2_X1 U2346 ( .A1(n1782), .A2(n1781), .ZN(n982) );
  NOR3_X1 U2347 ( .A1(n1795), .A2(ADD_RS2[3]), .A3(n1788), .ZN(n1782) );
  NAND4_X1 U2348 ( .A1(n1796), .A2(n1797), .A3(n1798), .A4(n1799), .ZN(n1773)
         );
  AOI221_X1 U2349 ( .B1(n148), .B2(n2492), .C1(n151), .C2(n2493), .A(n1800), 
        .ZN(n1799) );
  OAI22_X1 U2350 ( .A1(n2491), .A2(n154), .B1(n2490), .B2(n157), .ZN(n1800) );
  NAND2_X1 U2351 ( .A1(n1787), .A2(n1801), .ZN(n1001) );
  NAND2_X1 U2352 ( .A1(n1787), .A2(n1802), .ZN(n1000) );
  AND2_X1 U2353 ( .A1(n1801), .A2(n1783), .ZN(n998) );
  AND2_X1 U2354 ( .A1(n1783), .A2(n1802), .ZN(n997) );
  AOI221_X1 U2355 ( .B1(n160), .B2(n2496), .C1(n163), .C2(n2497), .A(n1803), 
        .ZN(n1798) );
  OAI22_X1 U2356 ( .A1(n2495), .A2(n166), .B1(n2494), .B2(n169), .ZN(n1803) );
  NAND2_X1 U2357 ( .A1(n1781), .A2(n1801), .ZN(n1006) );
  NAND2_X1 U2358 ( .A1(n1781), .A2(n1802), .ZN(n1005) );
  AND2_X1 U2359 ( .A1(n1780), .A2(n1801), .ZN(n1003) );
  NOR3_X1 U2360 ( .A1(ADD_RS2[0]), .A2(ADD_RS2[4]), .A3(n1789), .ZN(n1801) );
  AND2_X1 U2361 ( .A1(n1780), .A2(n1802), .ZN(n1002) );
  NOR3_X1 U2362 ( .A1(n1795), .A2(ADD_RS2[4]), .A3(n1789), .ZN(n1802) );
  AOI221_X1 U2363 ( .B1(n172), .B2(n637), .C1(n175), .C2(n670), .A(n1804), 
        .ZN(n1797) );
  OAI22_X1 U2364 ( .A1(n1805), .A2(n178), .B1(n1806), .B2(n181), .ZN(n1804) );
  NAND2_X1 U2365 ( .A1(n1807), .A2(n1783), .ZN(n1013) );
  NAND2_X1 U2366 ( .A1(n1808), .A2(n1783), .ZN(n1011) );
  NOR2_X1 U2367 ( .A1(n1809), .A2(n1810), .ZN(n1783) );
  AND2_X1 U2368 ( .A1(n1807), .A2(n1787), .ZN(n1008) );
  AND2_X1 U2369 ( .A1(n1808), .A2(n1787), .ZN(n1007) );
  AOI221_X1 U2370 ( .B1(n184), .B2(n603), .C1(n187), .C2(n3800), .A(n1811), 
        .ZN(n1796) );
  OAI22_X1 U2371 ( .A1(n1812), .A2(n190), .B1(n1813), .B2(n193), .ZN(n1811) );
  NAND2_X1 U2372 ( .A1(n1807), .A2(n1780), .ZN(n1020) );
  NAND2_X1 U2373 ( .A1(n1808), .A2(n1780), .ZN(n1018) );
  NOR2_X1 U2374 ( .A1(n1810), .A2(ADD_RS2[2]), .ZN(n1780) );
  NOR3_X1 U2375 ( .A1(ADD_RS2[3]), .A2(ADD_RS2[4]), .A3(ADD_RS2[0]), .ZN(n1808) );
  AND2_X1 U2376 ( .A1(n1784), .A2(n1787), .ZN(n1015) );
  NOR2_X1 U2377 ( .A1(n1809), .A2(ADD_RS2[1]), .ZN(n1787) );
  INV_X1 U2378 ( .A(ADD_RS2[2]), .ZN(n1809) );
  NOR3_X1 U2379 ( .A1(n1788), .A2(n1795), .A3(n1789), .ZN(n1784) );
  INV_X1 U2380 ( .A(ADD_RS2[3]), .ZN(n1789) );
  INV_X1 U2381 ( .A(ADD_RS2[4]), .ZN(n1788) );
  AND2_X1 U2382 ( .A1(n1807), .A2(n1781), .ZN(n1014) );
  NOR2_X1 U2383 ( .A1(ADD_RS2[1]), .A2(ADD_RS2[2]), .ZN(n1781) );
  NOR3_X1 U2384 ( .A1(ADD_RS2[3]), .A2(ADD_RS2[4]), .A3(n1795), .ZN(n1807) );
  INV_X1 U2385 ( .A(ADD_RS2[0]), .ZN(n1795) );
  NAND2_X1 U2386 ( .A1(n1814), .A2(n100), .ZN(n962) );
  AND3_X1 U2387 ( .A1(RD2), .A2(ENABLE), .A3(n419), .ZN(n965) );
  INV_X1 U2388 ( .A(n1772), .ZN(n1814) );
  NAND4_X1 U2389 ( .A1(n1815), .A2(n1816), .A3(n1817), .A4(n1818), .ZN(n1772)
         );
  NOR3_X1 U2390 ( .A1(n1819), .A2(n1820), .A3(n1821), .ZN(n1818) );
  XNOR2_X1 U2391 ( .A(ADD_WR[1]), .B(n1810), .ZN(n1821) );
  INV_X1 U2392 ( .A(ADD_RS2[1]), .ZN(n1810) );
  XNOR2_X1 U2393 ( .A(n953), .B(ADD_RS2[0]), .ZN(n1819) );
  XNOR2_X1 U2394 ( .A(ADD_WR[3]), .B(ADD_RS2[3]), .ZN(n1817) );
  XNOR2_X1 U2395 ( .A(ADD_WR[4]), .B(ADD_RS2[4]), .ZN(n1816) );
  XNOR2_X1 U2396 ( .A(ADD_RS2[2]), .B(ADD_WR[2]), .ZN(n1815) );
  OAI222_X1 U2397 ( .A1(n329), .A2(n198), .B1(n1823), .B2(n201), .C1(n2488), 
        .C2(n204), .ZN(n3014) );
  NOR4_X1 U2398 ( .A1(n1826), .A2(n1827), .A3(n1828), .A4(n1829), .ZN(n1823)
         );
  OAI221_X1 U2399 ( .B1(n3864), .B2(n207), .C1(n1777), .C2(n210), .A(n1832), 
        .ZN(n1829) );
  AOI22_X1 U2400 ( .A1(n213), .A2(n2503), .B1(n216), .B2(n671), .ZN(n1832) );
  OAI221_X1 U2401 ( .B1(n1785), .B2(n219), .C1(n3768), .C2(n222), .A(n1837), 
        .ZN(n1828) );
  AOI22_X1 U2402 ( .A1(n225), .A2(n806), .B1(n228), .B2(n2502), .ZN(n1837) );
  OAI211_X1 U2403 ( .C1(n2507), .C2(n231), .A(n1841), .B(n1842), .ZN(n1827) );
  AOI221_X1 U2404 ( .B1(n234), .B2(n940), .C1(n237), .C2(n2508), .A(n1845), 
        .ZN(n1842) );
  OAI22_X1 U2405 ( .A1(n2504), .A2(n240), .B1(n1793), .B2(n243), .ZN(n1845) );
  AOI22_X1 U2406 ( .A1(n246), .A2(n2509), .B1(n249), .B2(n840), .ZN(n1841) );
  NAND4_X1 U2407 ( .A1(n1850), .A2(n1851), .A3(n1852), .A4(n1853), .ZN(n1826)
         );
  AOI221_X1 U2408 ( .B1(n252), .B2(n2492), .C1(n255), .C2(n2493), .A(n1856), 
        .ZN(n1853) );
  OAI22_X1 U2409 ( .A1(n2491), .A2(n258), .B1(n2490), .B2(n261), .ZN(n1856) );
  AOI221_X1 U2410 ( .B1(n264), .B2(n2496), .C1(n267), .C2(n2497), .A(n1861), 
        .ZN(n1852) );
  OAI22_X1 U2411 ( .A1(n2495), .A2(n270), .B1(n2494), .B2(n273), .ZN(n1861) );
  AOI221_X1 U2412 ( .B1(n276), .B2(n637), .C1(n279), .C2(n670), .A(n1866), 
        .ZN(n1851) );
  OAI22_X1 U2413 ( .A1(n1805), .A2(n282), .B1(n1806), .B2(n285), .ZN(n1866) );
  AOI221_X1 U2414 ( .B1(n288), .B2(n603), .C1(n291), .C2(n3800), .A(n1871), 
        .ZN(n1850) );
  OAI22_X1 U2415 ( .A1(n1812), .A2(n294), .B1(n1813), .B2(n297), .ZN(n1871) );
  OAI222_X1 U2416 ( .A1(n328), .A2(n198), .B1(n1874), .B2(n201), .C1(n2487), 
        .C2(n204), .ZN(n3013) );
  NOR4_X1 U2417 ( .A1(n1875), .A2(n1876), .A3(n1877), .A4(n1878), .ZN(n1874)
         );
  OAI221_X1 U2418 ( .B1(n3863), .B2(n207), .C1(n1751), .C2(n210), .A(n1879), 
        .ZN(n1878) );
  AOI22_X1 U2419 ( .A1(n213), .A2(n2524), .B1(n216), .B2(n703), .ZN(n1879) );
  OAI221_X1 U2420 ( .B1(n1753), .B2(n219), .C1(n3767), .C2(n222), .A(n1880), 
        .ZN(n1877) );
  AOI22_X1 U2421 ( .A1(n225), .A2(n805), .B1(n228), .B2(n2523), .ZN(n1880) );
  OAI211_X1 U2422 ( .C1(n2528), .C2(n231), .A(n1881), .B(n1882), .ZN(n1876) );
  AOI221_X1 U2423 ( .B1(n234), .B2(n939), .C1(n237), .C2(n2529), .A(n1883), 
        .ZN(n1882) );
  OAI22_X1 U2424 ( .A1(n2525), .A2(n240), .B1(n1758), .B2(n243), .ZN(n1883) );
  AOI22_X1 U2425 ( .A1(n246), .A2(n2530), .B1(n249), .B2(n839), .ZN(n1881) );
  NAND4_X1 U2426 ( .A1(n1884), .A2(n1885), .A3(n1886), .A4(n1887), .ZN(n1875)
         );
  AOI221_X1 U2427 ( .B1(n252), .B2(n2513), .C1(n255), .C2(n2514), .A(n1888), 
        .ZN(n1887) );
  OAI22_X1 U2428 ( .A1(n2512), .A2(n258), .B1(n2511), .B2(n261), .ZN(n1888) );
  AOI221_X1 U2429 ( .B1(n264), .B2(n2517), .C1(n267), .C2(n2518), .A(n1889), 
        .ZN(n1886) );
  OAI22_X1 U2430 ( .A1(n2516), .A2(n270), .B1(n2515), .B2(n273), .ZN(n1889) );
  AOI221_X1 U2431 ( .B1(n276), .B2(n636), .C1(n279), .C2(n669), .A(n1890), 
        .ZN(n1885) );
  OAI22_X1 U2432 ( .A1(n1766), .A2(n282), .B1(n1767), .B2(n285), .ZN(n1890) );
  AOI221_X1 U2433 ( .B1(n288), .B2(n602), .C1(n291), .C2(n3799), .A(n1891), 
        .ZN(n1884) );
  OAI22_X1 U2434 ( .A1(n1769), .A2(n294), .B1(n1770), .B2(n297), .ZN(n1891) );
  OAI222_X1 U2435 ( .A1(n327), .A2(n198), .B1(n1892), .B2(n201), .C1(n2486), 
        .C2(n204), .ZN(n3012) );
  NOR4_X1 U2436 ( .A1(n1893), .A2(n1894), .A3(n1895), .A4(n1896), .ZN(n1892)
         );
  OAI221_X1 U2437 ( .B1(n3862), .B2(n207), .C1(n1726), .C2(n210), .A(n1897), 
        .ZN(n1896) );
  AOI22_X1 U2438 ( .A1(n213), .A2(n2545), .B1(n216), .B2(n702), .ZN(n1897) );
  OAI221_X1 U2439 ( .B1(n1728), .B2(n219), .C1(n3766), .C2(n222), .A(n1898), 
        .ZN(n1895) );
  AOI22_X1 U2440 ( .A1(n225), .A2(n804), .B1(n228), .B2(n2544), .ZN(n1898) );
  OAI211_X1 U2441 ( .C1(n2549), .C2(n231), .A(n1899), .B(n1900), .ZN(n1894) );
  AOI221_X1 U2442 ( .B1(n234), .B2(n938), .C1(n237), .C2(n2550), .A(n1901), 
        .ZN(n1900) );
  OAI22_X1 U2443 ( .A1(n2546), .A2(n240), .B1(n1733), .B2(n243), .ZN(n1901) );
  AOI22_X1 U2444 ( .A1(n246), .A2(n2551), .B1(n249), .B2(n838), .ZN(n1899) );
  NAND4_X1 U2445 ( .A1(n1902), .A2(n1903), .A3(n1904), .A4(n1905), .ZN(n1893)
         );
  AOI221_X1 U2446 ( .B1(n252), .B2(n2534), .C1(n255), .C2(n2535), .A(n1906), 
        .ZN(n1905) );
  OAI22_X1 U2447 ( .A1(n2533), .A2(n258), .B1(n2532), .B2(n261), .ZN(n1906) );
  AOI221_X1 U2448 ( .B1(n264), .B2(n2538), .C1(n267), .C2(n2539), .A(n1907), 
        .ZN(n1904) );
  OAI22_X1 U2449 ( .A1(n2537), .A2(n270), .B1(n2536), .B2(n273), .ZN(n1907) );
  AOI221_X1 U2450 ( .B1(n276), .B2(n635), .C1(n279), .C2(n668), .A(n1908), 
        .ZN(n1903) );
  OAI22_X1 U2451 ( .A1(n1741), .A2(n282), .B1(n1742), .B2(n285), .ZN(n1908) );
  AOI221_X1 U2452 ( .B1(n288), .B2(n601), .C1(n291), .C2(n3798), .A(n1909), 
        .ZN(n1902) );
  OAI22_X1 U2453 ( .A1(n1744), .A2(n294), .B1(n1745), .B2(n297), .ZN(n1909) );
  OAI222_X1 U2454 ( .A1(n326), .A2(n198), .B1(n1910), .B2(n201), .C1(n2485), 
        .C2(n204), .ZN(n3011) );
  NOR4_X1 U2455 ( .A1(n1911), .A2(n1912), .A3(n1913), .A4(n1914), .ZN(n1910)
         );
  OAI221_X1 U2456 ( .B1(n3861), .B2(n207), .C1(n1701), .C2(n210), .A(n1915), 
        .ZN(n1914) );
  AOI22_X1 U2457 ( .A1(n213), .A2(n2566), .B1(n216), .B2(n701), .ZN(n1915) );
  OAI221_X1 U2458 ( .B1(n1703), .B2(n219), .C1(n3765), .C2(n222), .A(n1916), 
        .ZN(n1913) );
  AOI22_X1 U2459 ( .A1(n225), .A2(n803), .B1(n228), .B2(n2565), .ZN(n1916) );
  OAI211_X1 U2460 ( .C1(n2570), .C2(n231), .A(n1917), .B(n1918), .ZN(n1912) );
  AOI221_X1 U2461 ( .B1(n234), .B2(n937), .C1(n237), .C2(n2571), .A(n1919), 
        .ZN(n1918) );
  OAI22_X1 U2462 ( .A1(n2567), .A2(n240), .B1(n1708), .B2(n243), .ZN(n1919) );
  AOI22_X1 U2463 ( .A1(n246), .A2(n2572), .B1(n249), .B2(n837), .ZN(n1917) );
  NAND4_X1 U2464 ( .A1(n1920), .A2(n1921), .A3(n1922), .A4(n1923), .ZN(n1911)
         );
  AOI221_X1 U2465 ( .B1(n252), .B2(n2555), .C1(n255), .C2(n2556), .A(n1924), 
        .ZN(n1923) );
  OAI22_X1 U2466 ( .A1(n2554), .A2(n258), .B1(n2553), .B2(n261), .ZN(n1924) );
  AOI221_X1 U2467 ( .B1(n264), .B2(n2559), .C1(n267), .C2(n2560), .A(n1925), 
        .ZN(n1922) );
  OAI22_X1 U2468 ( .A1(n2558), .A2(n270), .B1(n2557), .B2(n273), .ZN(n1925) );
  AOI221_X1 U2469 ( .B1(n276), .B2(n634), .C1(n279), .C2(n667), .A(n1926), 
        .ZN(n1921) );
  OAI22_X1 U2470 ( .A1(n1716), .A2(n282), .B1(n1717), .B2(n285), .ZN(n1926) );
  AOI221_X1 U2471 ( .B1(n288), .B2(n600), .C1(n291), .C2(n3797), .A(n1927), 
        .ZN(n1920) );
  OAI22_X1 U2472 ( .A1(n1719), .A2(n294), .B1(n1720), .B2(n297), .ZN(n1927) );
  OAI222_X1 U2473 ( .A1(n325), .A2(n198), .B1(n1928), .B2(n201), .C1(n2484), 
        .C2(n204), .ZN(n3010) );
  NOR4_X1 U2474 ( .A1(n1929), .A2(n1930), .A3(n1931), .A4(n1932), .ZN(n1928)
         );
  OAI221_X1 U2475 ( .B1(n3860), .B2(n207), .C1(n1676), .C2(n210), .A(n1933), 
        .ZN(n1932) );
  AOI22_X1 U2476 ( .A1(n213), .A2(n2587), .B1(n216), .B2(n700), .ZN(n1933) );
  OAI221_X1 U2477 ( .B1(n1678), .B2(n219), .C1(n3764), .C2(n222), .A(n1934), 
        .ZN(n1931) );
  AOI22_X1 U2478 ( .A1(n225), .A2(n802), .B1(n228), .B2(n2586), .ZN(n1934) );
  OAI211_X1 U2479 ( .C1(n2591), .C2(n231), .A(n1935), .B(n1936), .ZN(n1930) );
  AOI221_X1 U2480 ( .B1(n234), .B2(n936), .C1(n237), .C2(n2592), .A(n1937), 
        .ZN(n1936) );
  OAI22_X1 U2481 ( .A1(n2588), .A2(n240), .B1(n1683), .B2(n243), .ZN(n1937) );
  AOI22_X1 U2482 ( .A1(n246), .A2(n2593), .B1(n249), .B2(n836), .ZN(n1935) );
  NAND4_X1 U2483 ( .A1(n1938), .A2(n1939), .A3(n1940), .A4(n1941), .ZN(n1929)
         );
  AOI221_X1 U2484 ( .B1(n252), .B2(n2576), .C1(n255), .C2(n2577), .A(n1942), 
        .ZN(n1941) );
  OAI22_X1 U2485 ( .A1(n2575), .A2(n258), .B1(n2574), .B2(n261), .ZN(n1942) );
  AOI221_X1 U2486 ( .B1(n264), .B2(n2580), .C1(n267), .C2(n2581), .A(n1943), 
        .ZN(n1940) );
  OAI22_X1 U2487 ( .A1(n2579), .A2(n270), .B1(n2578), .B2(n273), .ZN(n1943) );
  AOI221_X1 U2488 ( .B1(n276), .B2(n633), .C1(n279), .C2(n666), .A(n1944), 
        .ZN(n1939) );
  OAI22_X1 U2489 ( .A1(n1691), .A2(n282), .B1(n1692), .B2(n285), .ZN(n1944) );
  AOI221_X1 U2490 ( .B1(n288), .B2(n599), .C1(n291), .C2(n3796), .A(n1945), 
        .ZN(n1938) );
  OAI22_X1 U2491 ( .A1(n1694), .A2(n294), .B1(n1695), .B2(n297), .ZN(n1945) );
  OAI222_X1 U2492 ( .A1(n324), .A2(n198), .B1(n1946), .B2(n201), .C1(n2483), 
        .C2(n204), .ZN(n3009) );
  NOR4_X1 U2493 ( .A1(n1947), .A2(n1948), .A3(n1949), .A4(n1950), .ZN(n1946)
         );
  OAI221_X1 U2494 ( .B1(n3859), .B2(n207), .C1(n1651), .C2(n210), .A(n1951), 
        .ZN(n1950) );
  AOI22_X1 U2495 ( .A1(n213), .A2(n2608), .B1(n216), .B2(n699), .ZN(n1951) );
  OAI221_X1 U2496 ( .B1(n1653), .B2(n219), .C1(n3763), .C2(n222), .A(n1952), 
        .ZN(n1949) );
  AOI22_X1 U2497 ( .A1(n225), .A2(n801), .B1(n228), .B2(n2607), .ZN(n1952) );
  OAI211_X1 U2498 ( .C1(n2612), .C2(n231), .A(n1953), .B(n1954), .ZN(n1948) );
  AOI221_X1 U2499 ( .B1(n234), .B2(n935), .C1(n237), .C2(n2613), .A(n1955), 
        .ZN(n1954) );
  OAI22_X1 U2500 ( .A1(n2609), .A2(n240), .B1(n1658), .B2(n243), .ZN(n1955) );
  AOI22_X1 U2501 ( .A1(n246), .A2(n2614), .B1(n249), .B2(n835), .ZN(n1953) );
  NAND4_X1 U2502 ( .A1(n1956), .A2(n1957), .A3(n1958), .A4(n1959), .ZN(n1947)
         );
  AOI221_X1 U2503 ( .B1(n252), .B2(n2597), .C1(n255), .C2(n2598), .A(n1960), 
        .ZN(n1959) );
  OAI22_X1 U2504 ( .A1(n2596), .A2(n258), .B1(n2595), .B2(n261), .ZN(n1960) );
  AOI221_X1 U2505 ( .B1(n264), .B2(n2601), .C1(n267), .C2(n2602), .A(n1961), 
        .ZN(n1958) );
  OAI22_X1 U2506 ( .A1(n2600), .A2(n270), .B1(n2599), .B2(n273), .ZN(n1961) );
  AOI221_X1 U2507 ( .B1(n276), .B2(n632), .C1(n279), .C2(n665), .A(n1962), 
        .ZN(n1957) );
  OAI22_X1 U2508 ( .A1(n1666), .A2(n282), .B1(n1667), .B2(n285), .ZN(n1962) );
  AOI221_X1 U2509 ( .B1(n288), .B2(n598), .C1(n291), .C2(n3795), .A(n1963), 
        .ZN(n1956) );
  OAI22_X1 U2510 ( .A1(n1669), .A2(n294), .B1(n1670), .B2(n297), .ZN(n1963) );
  OAI222_X1 U2511 ( .A1(n323), .A2(n198), .B1(n1964), .B2(n201), .C1(n2482), 
        .C2(n204), .ZN(n3008) );
  NOR4_X1 U2512 ( .A1(n1965), .A2(n1966), .A3(n1967), .A4(n1968), .ZN(n1964)
         );
  OAI221_X1 U2513 ( .B1(n3858), .B2(n207), .C1(n1626), .C2(n210), .A(n1969), 
        .ZN(n1968) );
  AOI22_X1 U2514 ( .A1(n213), .A2(n2629), .B1(n216), .B2(n698), .ZN(n1969) );
  OAI221_X1 U2515 ( .B1(n1628), .B2(n219), .C1(n3762), .C2(n222), .A(n1970), 
        .ZN(n1967) );
  AOI22_X1 U2516 ( .A1(n225), .A2(n800), .B1(n228), .B2(n2628), .ZN(n1970) );
  OAI211_X1 U2517 ( .C1(n2633), .C2(n231), .A(n1971), .B(n1972), .ZN(n1966) );
  AOI221_X1 U2518 ( .B1(n234), .B2(n934), .C1(n237), .C2(n2634), .A(n1973), 
        .ZN(n1972) );
  OAI22_X1 U2519 ( .A1(n2630), .A2(n240), .B1(n1633), .B2(n243), .ZN(n1973) );
  AOI22_X1 U2520 ( .A1(n246), .A2(n2635), .B1(n249), .B2(n834), .ZN(n1971) );
  NAND4_X1 U2521 ( .A1(n1974), .A2(n1975), .A3(n1976), .A4(n1977), .ZN(n1965)
         );
  AOI221_X1 U2522 ( .B1(n252), .B2(n2618), .C1(n255), .C2(n2619), .A(n1978), 
        .ZN(n1977) );
  OAI22_X1 U2523 ( .A1(n2617), .A2(n258), .B1(n2616), .B2(n261), .ZN(n1978) );
  AOI221_X1 U2524 ( .B1(n264), .B2(n2622), .C1(n267), .C2(n2623), .A(n1979), 
        .ZN(n1976) );
  OAI22_X1 U2525 ( .A1(n2621), .A2(n270), .B1(n2620), .B2(n273), .ZN(n1979) );
  AOI221_X1 U2526 ( .B1(n276), .B2(n631), .C1(n279), .C2(n664), .A(n1980), 
        .ZN(n1975) );
  OAI22_X1 U2527 ( .A1(n1641), .A2(n282), .B1(n1642), .B2(n285), .ZN(n1980) );
  AOI221_X1 U2528 ( .B1(n288), .B2(n597), .C1(n291), .C2(n3794), .A(n1981), 
        .ZN(n1974) );
  OAI22_X1 U2529 ( .A1(n1644), .A2(n294), .B1(n1645), .B2(n297), .ZN(n1981) );
  OAI222_X1 U2530 ( .A1(n322), .A2(n198), .B1(n1982), .B2(n201), .C1(n2481), 
        .C2(n204), .ZN(n3007) );
  NOR4_X1 U2531 ( .A1(n1983), .A2(n1984), .A3(n1985), .A4(n1986), .ZN(n1982)
         );
  OAI221_X1 U2532 ( .B1(n3857), .B2(n207), .C1(n1601), .C2(n210), .A(n1987), 
        .ZN(n1986) );
  AOI22_X1 U2533 ( .A1(n213), .A2(n2650), .B1(n216), .B2(n697), .ZN(n1987) );
  OAI221_X1 U2534 ( .B1(n1603), .B2(n219), .C1(n3761), .C2(n222), .A(n1988), 
        .ZN(n1985) );
  AOI22_X1 U2535 ( .A1(n225), .A2(n799), .B1(n228), .B2(n2649), .ZN(n1988) );
  OAI211_X1 U2536 ( .C1(n2654), .C2(n231), .A(n1989), .B(n1990), .ZN(n1984) );
  AOI221_X1 U2537 ( .B1(n234), .B2(n933), .C1(n237), .C2(n2655), .A(n1991), 
        .ZN(n1990) );
  OAI22_X1 U2538 ( .A1(n2651), .A2(n240), .B1(n1608), .B2(n243), .ZN(n1991) );
  AOI22_X1 U2539 ( .A1(n246), .A2(n2656), .B1(n249), .B2(n833), .ZN(n1989) );
  NAND4_X1 U2540 ( .A1(n1992), .A2(n1993), .A3(n1994), .A4(n1995), .ZN(n1983)
         );
  AOI221_X1 U2541 ( .B1(n252), .B2(n2639), .C1(n255), .C2(n2640), .A(n1996), 
        .ZN(n1995) );
  OAI22_X1 U2542 ( .A1(n2638), .A2(n258), .B1(n2637), .B2(n261), .ZN(n1996) );
  AOI221_X1 U2543 ( .B1(n264), .B2(n2643), .C1(n267), .C2(n2644), .A(n1997), 
        .ZN(n1994) );
  OAI22_X1 U2544 ( .A1(n2642), .A2(n270), .B1(n2641), .B2(n273), .ZN(n1997) );
  AOI221_X1 U2545 ( .B1(n276), .B2(n630), .C1(n279), .C2(n663), .A(n1998), 
        .ZN(n1993) );
  OAI22_X1 U2546 ( .A1(n1616), .A2(n282), .B1(n1617), .B2(n285), .ZN(n1998) );
  AOI221_X1 U2547 ( .B1(n288), .B2(n596), .C1(n291), .C2(n3793), .A(n1999), 
        .ZN(n1992) );
  OAI22_X1 U2548 ( .A1(n1619), .A2(n294), .B1(n1620), .B2(n297), .ZN(n1999) );
  OAI222_X1 U2549 ( .A1(n321), .A2(n197), .B1(n2000), .B2(n200), .C1(n2480), 
        .C2(n204), .ZN(n3006) );
  NOR4_X1 U2550 ( .A1(n2001), .A2(n2002), .A3(n2003), .A4(n2004), .ZN(n2000)
         );
  OAI221_X1 U2551 ( .B1(n3856), .B2(n206), .C1(n1576), .C2(n209), .A(n2005), 
        .ZN(n2004) );
  AOI22_X1 U2552 ( .A1(n212), .A2(n2671), .B1(n215), .B2(n696), .ZN(n2005) );
  OAI221_X1 U2553 ( .B1(n1578), .B2(n218), .C1(n3760), .C2(n221), .A(n2006), 
        .ZN(n2003) );
  AOI22_X1 U2554 ( .A1(n224), .A2(n798), .B1(n227), .B2(n2670), .ZN(n2006) );
  OAI211_X1 U2555 ( .C1(n2675), .C2(n230), .A(n2007), .B(n2008), .ZN(n2002) );
  AOI221_X1 U2556 ( .B1(n233), .B2(n932), .C1(n236), .C2(n2676), .A(n2009), 
        .ZN(n2008) );
  OAI22_X1 U2557 ( .A1(n2672), .A2(n239), .B1(n1583), .B2(n242), .ZN(n2009) );
  AOI22_X1 U2558 ( .A1(n245), .A2(n2677), .B1(n248), .B2(n832), .ZN(n2007) );
  NAND4_X1 U2559 ( .A1(n2010), .A2(n2011), .A3(n2012), .A4(n2013), .ZN(n2001)
         );
  AOI221_X1 U2560 ( .B1(n251), .B2(n2660), .C1(n254), .C2(n2661), .A(n2014), 
        .ZN(n2013) );
  OAI22_X1 U2561 ( .A1(n2659), .A2(n257), .B1(n2658), .B2(n260), .ZN(n2014) );
  AOI221_X1 U2562 ( .B1(n263), .B2(n2664), .C1(n266), .C2(n2665), .A(n2015), 
        .ZN(n2012) );
  OAI22_X1 U2563 ( .A1(n2663), .A2(n269), .B1(n2662), .B2(n272), .ZN(n2015) );
  AOI221_X1 U2564 ( .B1(n275), .B2(n629), .C1(n278), .C2(n662), .A(n2016), 
        .ZN(n2011) );
  OAI22_X1 U2565 ( .A1(n1591), .A2(n281), .B1(n1592), .B2(n284), .ZN(n2016) );
  AOI221_X1 U2566 ( .B1(n287), .B2(n595), .C1(n290), .C2(n3792), .A(n2017), 
        .ZN(n2010) );
  OAI22_X1 U2567 ( .A1(n1594), .A2(n293), .B1(n1595), .B2(n296), .ZN(n2017) );
  OAI222_X1 U2568 ( .A1(n320), .A2(n197), .B1(n2018), .B2(n200), .C1(n2479), 
        .C2(n204), .ZN(n3005) );
  NOR4_X1 U2569 ( .A1(n2019), .A2(n2020), .A3(n2021), .A4(n2022), .ZN(n2018)
         );
  OAI221_X1 U2570 ( .B1(n3855), .B2(n206), .C1(n1551), .C2(n209), .A(n2023), 
        .ZN(n2022) );
  AOI22_X1 U2571 ( .A1(n212), .A2(n2692), .B1(n215), .B2(n695), .ZN(n2023) );
  OAI221_X1 U2572 ( .B1(n1553), .B2(n218), .C1(n3759), .C2(n221), .A(n2024), 
        .ZN(n2021) );
  AOI22_X1 U2573 ( .A1(n224), .A2(n797), .B1(n227), .B2(n2691), .ZN(n2024) );
  OAI211_X1 U2574 ( .C1(n2696), .C2(n230), .A(n2025), .B(n2026), .ZN(n2020) );
  AOI221_X1 U2575 ( .B1(n233), .B2(n931), .C1(n236), .C2(n2697), .A(n2027), 
        .ZN(n2026) );
  OAI22_X1 U2576 ( .A1(n2693), .A2(n239), .B1(n1558), .B2(n242), .ZN(n2027) );
  AOI22_X1 U2577 ( .A1(n245), .A2(n2698), .B1(n248), .B2(n831), .ZN(n2025) );
  NAND4_X1 U2578 ( .A1(n2028), .A2(n2029), .A3(n2030), .A4(n2031), .ZN(n2019)
         );
  AOI221_X1 U2579 ( .B1(n251), .B2(n2681), .C1(n254), .C2(n2682), .A(n2032), 
        .ZN(n2031) );
  OAI22_X1 U2580 ( .A1(n2680), .A2(n257), .B1(n2679), .B2(n260), .ZN(n2032) );
  AOI221_X1 U2581 ( .B1(n263), .B2(n2685), .C1(n266), .C2(n2686), .A(n2033), 
        .ZN(n2030) );
  OAI22_X1 U2582 ( .A1(n2684), .A2(n269), .B1(n2683), .B2(n272), .ZN(n2033) );
  AOI221_X1 U2583 ( .B1(n275), .B2(n628), .C1(n278), .C2(n661), .A(n2034), 
        .ZN(n2029) );
  OAI22_X1 U2584 ( .A1(n1566), .A2(n281), .B1(n1567), .B2(n284), .ZN(n2034) );
  AOI221_X1 U2585 ( .B1(n287), .B2(n594), .C1(n290), .C2(n3791), .A(n2035), 
        .ZN(n2028) );
  OAI22_X1 U2586 ( .A1(n1569), .A2(n293), .B1(n1570), .B2(n296), .ZN(n2035) );
  OAI222_X1 U2587 ( .A1(n319), .A2(n197), .B1(n2036), .B2(n200), .C1(n2478), 
        .C2(n203), .ZN(n3004) );
  NOR4_X1 U2588 ( .A1(n2037), .A2(n2038), .A3(n2039), .A4(n2040), .ZN(n2036)
         );
  OAI221_X1 U2589 ( .B1(n3854), .B2(n206), .C1(n1526), .C2(n209), .A(n2041), 
        .ZN(n2040) );
  AOI22_X1 U2590 ( .A1(n212), .A2(n2713), .B1(n215), .B2(n694), .ZN(n2041) );
  OAI221_X1 U2591 ( .B1(n1528), .B2(n218), .C1(n3758), .C2(n221), .A(n2042), 
        .ZN(n2039) );
  AOI22_X1 U2592 ( .A1(n224), .A2(n796), .B1(n227), .B2(n2712), .ZN(n2042) );
  OAI211_X1 U2593 ( .C1(n2717), .C2(n230), .A(n2043), .B(n2044), .ZN(n2038) );
  AOI221_X1 U2594 ( .B1(n233), .B2(n930), .C1(n236), .C2(n2718), .A(n2045), 
        .ZN(n2044) );
  OAI22_X1 U2595 ( .A1(n2714), .A2(n239), .B1(n1533), .B2(n242), .ZN(n2045) );
  AOI22_X1 U2596 ( .A1(n245), .A2(n2719), .B1(n248), .B2(n830), .ZN(n2043) );
  NAND4_X1 U2597 ( .A1(n2046), .A2(n2047), .A3(n2048), .A4(n2049), .ZN(n2037)
         );
  AOI221_X1 U2598 ( .B1(n251), .B2(n2702), .C1(n254), .C2(n2703), .A(n2050), 
        .ZN(n2049) );
  OAI22_X1 U2599 ( .A1(n2701), .A2(n257), .B1(n2700), .B2(n260), .ZN(n2050) );
  AOI221_X1 U2600 ( .B1(n263), .B2(n2706), .C1(n266), .C2(n2707), .A(n2051), 
        .ZN(n2048) );
  OAI22_X1 U2601 ( .A1(n2705), .A2(n269), .B1(n2704), .B2(n272), .ZN(n2051) );
  AOI221_X1 U2602 ( .B1(n275), .B2(n627), .C1(n278), .C2(n660), .A(n2052), 
        .ZN(n2047) );
  OAI22_X1 U2603 ( .A1(n1541), .A2(n281), .B1(n1542), .B2(n284), .ZN(n2052) );
  AOI221_X1 U2604 ( .B1(n287), .B2(n593), .C1(n290), .C2(n3790), .A(n2053), 
        .ZN(n2046) );
  OAI22_X1 U2605 ( .A1(n1544), .A2(n293), .B1(n1545), .B2(n296), .ZN(n2053) );
  OAI222_X1 U2606 ( .A1(n318), .A2(n197), .B1(n2054), .B2(n200), .C1(n2477), 
        .C2(n203), .ZN(n3003) );
  NOR4_X1 U2607 ( .A1(n2055), .A2(n2056), .A3(n2057), .A4(n2058), .ZN(n2054)
         );
  OAI221_X1 U2608 ( .B1(n3853), .B2(n206), .C1(n1501), .C2(n209), .A(n2059), 
        .ZN(n2058) );
  AOI22_X1 U2609 ( .A1(n212), .A2(n2734), .B1(n215), .B2(n693), .ZN(n2059) );
  OAI221_X1 U2610 ( .B1(n1503), .B2(n218), .C1(n3757), .C2(n221), .A(n2060), 
        .ZN(n2057) );
  AOI22_X1 U2611 ( .A1(n224), .A2(n795), .B1(n227), .B2(n2733), .ZN(n2060) );
  OAI211_X1 U2612 ( .C1(n2738), .C2(n230), .A(n2061), .B(n2062), .ZN(n2056) );
  AOI221_X1 U2613 ( .B1(n233), .B2(n929), .C1(n236), .C2(n2739), .A(n2063), 
        .ZN(n2062) );
  OAI22_X1 U2614 ( .A1(n2735), .A2(n239), .B1(n1508), .B2(n242), .ZN(n2063) );
  AOI22_X1 U2615 ( .A1(n245), .A2(n2740), .B1(n248), .B2(n829), .ZN(n2061) );
  NAND4_X1 U2616 ( .A1(n2064), .A2(n2065), .A3(n2066), .A4(n2067), .ZN(n2055)
         );
  AOI221_X1 U2617 ( .B1(n251), .B2(n2723), .C1(n254), .C2(n2724), .A(n2068), 
        .ZN(n2067) );
  OAI22_X1 U2618 ( .A1(n2722), .A2(n257), .B1(n2721), .B2(n260), .ZN(n2068) );
  AOI221_X1 U2619 ( .B1(n263), .B2(n2727), .C1(n266), .C2(n2728), .A(n2069), 
        .ZN(n2066) );
  OAI22_X1 U2620 ( .A1(n2726), .A2(n269), .B1(n2725), .B2(n272), .ZN(n2069) );
  AOI221_X1 U2621 ( .B1(n275), .B2(n626), .C1(n278), .C2(n659), .A(n2070), 
        .ZN(n2065) );
  OAI22_X1 U2622 ( .A1(n1516), .A2(n281), .B1(n1517), .B2(n284), .ZN(n2070) );
  AOI221_X1 U2623 ( .B1(n287), .B2(n592), .C1(n290), .C2(n3789), .A(n2071), 
        .ZN(n2064) );
  OAI22_X1 U2624 ( .A1(n1519), .A2(n293), .B1(n1520), .B2(n296), .ZN(n2071) );
  OAI222_X1 U2625 ( .A1(n317), .A2(n197), .B1(n2072), .B2(n200), .C1(n2476), 
        .C2(n203), .ZN(n3002) );
  NOR4_X1 U2626 ( .A1(n2073), .A2(n2074), .A3(n2075), .A4(n2076), .ZN(n2072)
         );
  OAI221_X1 U2627 ( .B1(n3852), .B2(n206), .C1(n1476), .C2(n209), .A(n2077), 
        .ZN(n2076) );
  AOI22_X1 U2628 ( .A1(n212), .A2(n2755), .B1(n215), .B2(n692), .ZN(n2077) );
  OAI221_X1 U2629 ( .B1(n1478), .B2(n218), .C1(n3756), .C2(n221), .A(n2078), 
        .ZN(n2075) );
  AOI22_X1 U2630 ( .A1(n224), .A2(n794), .B1(n227), .B2(n2754), .ZN(n2078) );
  OAI211_X1 U2631 ( .C1(n2759), .C2(n230), .A(n2079), .B(n2080), .ZN(n2074) );
  AOI221_X1 U2632 ( .B1(n233), .B2(n928), .C1(n236), .C2(n2760), .A(n2081), 
        .ZN(n2080) );
  OAI22_X1 U2633 ( .A1(n2756), .A2(n239), .B1(n1483), .B2(n242), .ZN(n2081) );
  AOI22_X1 U2634 ( .A1(n245), .A2(n2761), .B1(n248), .B2(n828), .ZN(n2079) );
  NAND4_X1 U2635 ( .A1(n2082), .A2(n2083), .A3(n2084), .A4(n2085), .ZN(n2073)
         );
  AOI221_X1 U2636 ( .B1(n251), .B2(n2744), .C1(n254), .C2(n2745), .A(n2086), 
        .ZN(n2085) );
  OAI22_X1 U2637 ( .A1(n2743), .A2(n257), .B1(n2742), .B2(n260), .ZN(n2086) );
  AOI221_X1 U2638 ( .B1(n263), .B2(n2748), .C1(n266), .C2(n2749), .A(n2087), 
        .ZN(n2084) );
  OAI22_X1 U2639 ( .A1(n2747), .A2(n269), .B1(n2746), .B2(n272), .ZN(n2087) );
  AOI221_X1 U2640 ( .B1(n275), .B2(n625), .C1(n278), .C2(n658), .A(n2088), 
        .ZN(n2083) );
  OAI22_X1 U2641 ( .A1(n1491), .A2(n281), .B1(n1492), .B2(n284), .ZN(n2088) );
  AOI221_X1 U2642 ( .B1(n287), .B2(n591), .C1(n290), .C2(n3788), .A(n2089), 
        .ZN(n2082) );
  OAI22_X1 U2643 ( .A1(n1494), .A2(n293), .B1(n1495), .B2(n296), .ZN(n2089) );
  OAI222_X1 U2644 ( .A1(n316), .A2(n197), .B1(n2090), .B2(n200), .C1(n2475), 
        .C2(n203), .ZN(n3001) );
  NOR4_X1 U2645 ( .A1(n2091), .A2(n2092), .A3(n2093), .A4(n2094), .ZN(n2090)
         );
  OAI221_X1 U2646 ( .B1(n3851), .B2(n206), .C1(n1451), .C2(n209), .A(n2095), 
        .ZN(n2094) );
  AOI22_X1 U2647 ( .A1(n212), .A2(n2776), .B1(n215), .B2(n691), .ZN(n2095) );
  OAI221_X1 U2648 ( .B1(n1453), .B2(n218), .C1(n3755), .C2(n221), .A(n2096), 
        .ZN(n2093) );
  AOI22_X1 U2649 ( .A1(n224), .A2(n793), .B1(n227), .B2(n2775), .ZN(n2096) );
  OAI211_X1 U2650 ( .C1(n2780), .C2(n230), .A(n2097), .B(n2098), .ZN(n2092) );
  AOI221_X1 U2651 ( .B1(n233), .B2(n927), .C1(n236), .C2(n2781), .A(n2099), 
        .ZN(n2098) );
  OAI22_X1 U2652 ( .A1(n2777), .A2(n239), .B1(n1458), .B2(n242), .ZN(n2099) );
  AOI22_X1 U2653 ( .A1(n245), .A2(n2782), .B1(n248), .B2(n827), .ZN(n2097) );
  NAND4_X1 U2654 ( .A1(n2100), .A2(n2101), .A3(n2102), .A4(n2103), .ZN(n2091)
         );
  AOI221_X1 U2655 ( .B1(n251), .B2(n2765), .C1(n254), .C2(n2766), .A(n2104), 
        .ZN(n2103) );
  OAI22_X1 U2656 ( .A1(n2764), .A2(n257), .B1(n2763), .B2(n260), .ZN(n2104) );
  AOI221_X1 U2657 ( .B1(n263), .B2(n2769), .C1(n266), .C2(n2770), .A(n2105), 
        .ZN(n2102) );
  OAI22_X1 U2658 ( .A1(n2768), .A2(n269), .B1(n2767), .B2(n272), .ZN(n2105) );
  AOI221_X1 U2659 ( .B1(n275), .B2(n624), .C1(n278), .C2(n657), .A(n2106), 
        .ZN(n2101) );
  OAI22_X1 U2660 ( .A1(n1466), .A2(n281), .B1(n1467), .B2(n284), .ZN(n2106) );
  AOI221_X1 U2661 ( .B1(n287), .B2(n590), .C1(n290), .C2(n3787), .A(n2107), 
        .ZN(n2100) );
  OAI22_X1 U2662 ( .A1(n1469), .A2(n293), .B1(n1470), .B2(n296), .ZN(n2107) );
  OAI222_X1 U2663 ( .A1(n315), .A2(n197), .B1(n2108), .B2(n200), .C1(n2474), 
        .C2(n203), .ZN(n3000) );
  NOR4_X1 U2664 ( .A1(n2109), .A2(n2110), .A3(n2111), .A4(n2112), .ZN(n2108)
         );
  OAI221_X1 U2665 ( .B1(n3850), .B2(n206), .C1(n1426), .C2(n209), .A(n2113), 
        .ZN(n2112) );
  AOI22_X1 U2666 ( .A1(n212), .A2(n2797), .B1(n215), .B2(n690), .ZN(n2113) );
  OAI221_X1 U2667 ( .B1(n1428), .B2(n218), .C1(n3754), .C2(n221), .A(n2114), 
        .ZN(n2111) );
  AOI22_X1 U2668 ( .A1(n224), .A2(n792), .B1(n227), .B2(n2796), .ZN(n2114) );
  OAI211_X1 U2669 ( .C1(n2801), .C2(n230), .A(n2115), .B(n2116), .ZN(n2110) );
  AOI221_X1 U2670 ( .B1(n233), .B2(n926), .C1(n236), .C2(n2802), .A(n2117), 
        .ZN(n2116) );
  OAI22_X1 U2671 ( .A1(n2798), .A2(n239), .B1(n1433), .B2(n242), .ZN(n2117) );
  AOI22_X1 U2672 ( .A1(n245), .A2(n2803), .B1(n248), .B2(n826), .ZN(n2115) );
  NAND4_X1 U2673 ( .A1(n2118), .A2(n2119), .A3(n2120), .A4(n2121), .ZN(n2109)
         );
  AOI221_X1 U2674 ( .B1(n251), .B2(n2786), .C1(n254), .C2(n2787), .A(n2122), 
        .ZN(n2121) );
  OAI22_X1 U2675 ( .A1(n2785), .A2(n257), .B1(n2784), .B2(n260), .ZN(n2122) );
  AOI221_X1 U2676 ( .B1(n263), .B2(n2790), .C1(n266), .C2(n2791), .A(n2123), 
        .ZN(n2120) );
  OAI22_X1 U2677 ( .A1(n2789), .A2(n269), .B1(n2788), .B2(n272), .ZN(n2123) );
  AOI221_X1 U2678 ( .B1(n275), .B2(n623), .C1(n278), .C2(n656), .A(n2124), 
        .ZN(n2119) );
  OAI22_X1 U2679 ( .A1(n1441), .A2(n281), .B1(n1442), .B2(n284), .ZN(n2124) );
  AOI221_X1 U2680 ( .B1(n287), .B2(n589), .C1(n290), .C2(n3786), .A(n2125), 
        .ZN(n2118) );
  OAI22_X1 U2681 ( .A1(n1444), .A2(n293), .B1(n1445), .B2(n296), .ZN(n2125) );
  OAI222_X1 U2682 ( .A1(n314), .A2(n197), .B1(n2126), .B2(n200), .C1(n2473), 
        .C2(n203), .ZN(n2999) );
  NOR4_X1 U2683 ( .A1(n2127), .A2(n2128), .A3(n2129), .A4(n2130), .ZN(n2126)
         );
  OAI221_X1 U2684 ( .B1(n3849), .B2(n206), .C1(n1401), .C2(n209), .A(n2131), 
        .ZN(n2130) );
  AOI22_X1 U2685 ( .A1(n212), .A2(n2818), .B1(n215), .B2(n689), .ZN(n2131) );
  OAI221_X1 U2686 ( .B1(n1403), .B2(n218), .C1(n3753), .C2(n221), .A(n2132), 
        .ZN(n2129) );
  AOI22_X1 U2687 ( .A1(n224), .A2(n791), .B1(n227), .B2(n2817), .ZN(n2132) );
  OAI211_X1 U2688 ( .C1(n2822), .C2(n230), .A(n2133), .B(n2134), .ZN(n2128) );
  AOI221_X1 U2689 ( .B1(n233), .B2(n925), .C1(n236), .C2(n2823), .A(n2135), 
        .ZN(n2134) );
  OAI22_X1 U2690 ( .A1(n2819), .A2(n239), .B1(n1408), .B2(n242), .ZN(n2135) );
  AOI22_X1 U2691 ( .A1(n245), .A2(n2824), .B1(n248), .B2(n825), .ZN(n2133) );
  NAND4_X1 U2692 ( .A1(n2136), .A2(n2137), .A3(n2138), .A4(n2139), .ZN(n2127)
         );
  AOI221_X1 U2693 ( .B1(n251), .B2(n2807), .C1(n254), .C2(n2808), .A(n2140), 
        .ZN(n2139) );
  OAI22_X1 U2694 ( .A1(n2806), .A2(n257), .B1(n2805), .B2(n260), .ZN(n2140) );
  AOI221_X1 U2695 ( .B1(n263), .B2(n2811), .C1(n266), .C2(n2812), .A(n2141), 
        .ZN(n2138) );
  OAI22_X1 U2696 ( .A1(n2810), .A2(n269), .B1(n2809), .B2(n272), .ZN(n2141) );
  AOI221_X1 U2697 ( .B1(n275), .B2(n622), .C1(n278), .C2(n655), .A(n2142), 
        .ZN(n2137) );
  OAI22_X1 U2698 ( .A1(n1416), .A2(n281), .B1(n1417), .B2(n284), .ZN(n2142) );
  AOI221_X1 U2699 ( .B1(n287), .B2(n588), .C1(n290), .C2(n3785), .A(n2143), 
        .ZN(n2136) );
  OAI22_X1 U2700 ( .A1(n1419), .A2(n293), .B1(n1420), .B2(n296), .ZN(n2143) );
  OAI222_X1 U2701 ( .A1(n313), .A2(n197), .B1(n2144), .B2(n200), .C1(n2472), 
        .C2(n203), .ZN(n2998) );
  NOR4_X1 U2702 ( .A1(n2145), .A2(n2146), .A3(n2147), .A4(n2148), .ZN(n2144)
         );
  OAI221_X1 U2703 ( .B1(n3848), .B2(n206), .C1(n1376), .C2(n209), .A(n2149), 
        .ZN(n2148) );
  AOI22_X1 U2704 ( .A1(n212), .A2(n2839), .B1(n215), .B2(n688), .ZN(n2149) );
  OAI221_X1 U2705 ( .B1(n1378), .B2(n218), .C1(n3752), .C2(n221), .A(n2150), 
        .ZN(n2147) );
  AOI22_X1 U2706 ( .A1(n224), .A2(n790), .B1(n227), .B2(n2838), .ZN(n2150) );
  OAI211_X1 U2707 ( .C1(n2843), .C2(n230), .A(n2151), .B(n2152), .ZN(n2146) );
  AOI221_X1 U2708 ( .B1(n233), .B2(n924), .C1(n236), .C2(n2844), .A(n2153), 
        .ZN(n2152) );
  OAI22_X1 U2709 ( .A1(n2840), .A2(n239), .B1(n1383), .B2(n242), .ZN(n2153) );
  AOI22_X1 U2710 ( .A1(n245), .A2(n2845), .B1(n248), .B2(n824), .ZN(n2151) );
  NAND4_X1 U2711 ( .A1(n2154), .A2(n2155), .A3(n2156), .A4(n2157), .ZN(n2145)
         );
  AOI221_X1 U2712 ( .B1(n251), .B2(n2828), .C1(n254), .C2(n2829), .A(n2158), 
        .ZN(n2157) );
  OAI22_X1 U2713 ( .A1(n2827), .A2(n257), .B1(n2826), .B2(n260), .ZN(n2158) );
  AOI221_X1 U2714 ( .B1(n263), .B2(n2832), .C1(n266), .C2(n2833), .A(n2159), 
        .ZN(n2156) );
  OAI22_X1 U2715 ( .A1(n2831), .A2(n269), .B1(n2830), .B2(n272), .ZN(n2159) );
  AOI221_X1 U2716 ( .B1(n275), .B2(n621), .C1(n278), .C2(n654), .A(n2160), 
        .ZN(n2155) );
  OAI22_X1 U2717 ( .A1(n1391), .A2(n281), .B1(n1392), .B2(n284), .ZN(n2160) );
  AOI221_X1 U2718 ( .B1(n287), .B2(n587), .C1(n290), .C2(n3784), .A(n2161), 
        .ZN(n2154) );
  OAI22_X1 U2719 ( .A1(n1394), .A2(n293), .B1(n1395), .B2(n296), .ZN(n2161) );
  OAI222_X1 U2720 ( .A1(n312), .A2(n197), .B1(n2162), .B2(n200), .C1(n2471), 
        .C2(n203), .ZN(n2997) );
  NOR4_X1 U2721 ( .A1(n2163), .A2(n2164), .A3(n2165), .A4(n2166), .ZN(n2162)
         );
  OAI221_X1 U2722 ( .B1(n3847), .B2(n206), .C1(n1351), .C2(n209), .A(n2167), 
        .ZN(n2166) );
  AOI22_X1 U2723 ( .A1(n212), .A2(n2860), .B1(n215), .B2(n687), .ZN(n2167) );
  OAI221_X1 U2724 ( .B1(n1353), .B2(n218), .C1(n3751), .C2(n221), .A(n2168), 
        .ZN(n2165) );
  AOI22_X1 U2725 ( .A1(n224), .A2(n789), .B1(n227), .B2(n2859), .ZN(n2168) );
  OAI211_X1 U2726 ( .C1(n2864), .C2(n230), .A(n2169), .B(n2170), .ZN(n2164) );
  AOI221_X1 U2727 ( .B1(n233), .B2(n923), .C1(n236), .C2(n2865), .A(n2171), 
        .ZN(n2170) );
  OAI22_X1 U2728 ( .A1(n2861), .A2(n239), .B1(n1358), .B2(n242), .ZN(n2171) );
  AOI22_X1 U2729 ( .A1(n245), .A2(n2866), .B1(n248), .B2(n823), .ZN(n2169) );
  NAND4_X1 U2730 ( .A1(n2172), .A2(n2173), .A3(n2174), .A4(n2175), .ZN(n2163)
         );
  AOI221_X1 U2731 ( .B1(n251), .B2(n2849), .C1(n254), .C2(n2850), .A(n2176), 
        .ZN(n2175) );
  OAI22_X1 U2732 ( .A1(n2848), .A2(n257), .B1(n2847), .B2(n260), .ZN(n2176) );
  AOI221_X1 U2733 ( .B1(n263), .B2(n2853), .C1(n266), .C2(n2854), .A(n2177), 
        .ZN(n2174) );
  OAI22_X1 U2734 ( .A1(n2852), .A2(n269), .B1(n2851), .B2(n272), .ZN(n2177) );
  AOI221_X1 U2735 ( .B1(n275), .B2(n620), .C1(n278), .C2(n653), .A(n2178), 
        .ZN(n2173) );
  OAI22_X1 U2736 ( .A1(n1366), .A2(n281), .B1(n1367), .B2(n284), .ZN(n2178) );
  AOI221_X1 U2737 ( .B1(n287), .B2(n586), .C1(n290), .C2(n3783), .A(n2179), 
        .ZN(n2172) );
  OAI22_X1 U2738 ( .A1(n1369), .A2(n293), .B1(n1370), .B2(n296), .ZN(n2179) );
  OAI222_X1 U2739 ( .A1(n311), .A2(n197), .B1(n2180), .B2(n200), .C1(n2470), 
        .C2(n203), .ZN(n2996) );
  NOR4_X1 U2740 ( .A1(n2181), .A2(n2182), .A3(n2183), .A4(n2184), .ZN(n2180)
         );
  OAI221_X1 U2741 ( .B1(n3846), .B2(n206), .C1(n1326), .C2(n209), .A(n2185), 
        .ZN(n2184) );
  AOI22_X1 U2742 ( .A1(n212), .A2(n2881), .B1(n215), .B2(n686), .ZN(n2185) );
  OAI221_X1 U2743 ( .B1(n1328), .B2(n218), .C1(n3750), .C2(n221), .A(n2186), 
        .ZN(n2183) );
  AOI22_X1 U2744 ( .A1(n224), .A2(n788), .B1(n227), .B2(n2880), .ZN(n2186) );
  OAI211_X1 U2745 ( .C1(n2885), .C2(n230), .A(n2187), .B(n2188), .ZN(n2182) );
  AOI221_X1 U2746 ( .B1(n233), .B2(n922), .C1(n236), .C2(n2886), .A(n2189), 
        .ZN(n2188) );
  OAI22_X1 U2747 ( .A1(n2882), .A2(n239), .B1(n1333), .B2(n242), .ZN(n2189) );
  AOI22_X1 U2748 ( .A1(n245), .A2(n2887), .B1(n248), .B2(n822), .ZN(n2187) );
  NAND4_X1 U2749 ( .A1(n2190), .A2(n2191), .A3(n2192), .A4(n2193), .ZN(n2181)
         );
  AOI221_X1 U2750 ( .B1(n251), .B2(n2870), .C1(n254), .C2(n2871), .A(n2194), 
        .ZN(n2193) );
  OAI22_X1 U2751 ( .A1(n2869), .A2(n257), .B1(n2868), .B2(n260), .ZN(n2194) );
  AOI221_X1 U2752 ( .B1(n263), .B2(n2874), .C1(n266), .C2(n2875), .A(n2195), 
        .ZN(n2192) );
  OAI22_X1 U2753 ( .A1(n2873), .A2(n269), .B1(n2872), .B2(n272), .ZN(n2195) );
  AOI221_X1 U2754 ( .B1(n275), .B2(n619), .C1(n278), .C2(n652), .A(n2196), 
        .ZN(n2191) );
  OAI22_X1 U2755 ( .A1(n1341), .A2(n281), .B1(n1342), .B2(n284), .ZN(n2196) );
  AOI221_X1 U2756 ( .B1(n287), .B2(n585), .C1(n290), .C2(n3782), .A(n2197), 
        .ZN(n2190) );
  OAI22_X1 U2757 ( .A1(n1344), .A2(n293), .B1(n1345), .B2(n296), .ZN(n2197) );
  OAI222_X1 U2758 ( .A1(n310), .A2(n197), .B1(n2198), .B2(n200), .C1(n2469), 
        .C2(n203), .ZN(n2995) );
  NOR4_X1 U2759 ( .A1(n2199), .A2(n2200), .A3(n2201), .A4(n2202), .ZN(n2198)
         );
  OAI221_X1 U2760 ( .B1(n3845), .B2(n206), .C1(n1301), .C2(n209), .A(n2203), 
        .ZN(n2202) );
  AOI22_X1 U2761 ( .A1(n212), .A2(n2902), .B1(n215), .B2(n685), .ZN(n2203) );
  OAI221_X1 U2762 ( .B1(n1303), .B2(n218), .C1(n3749), .C2(n221), .A(n2204), 
        .ZN(n2201) );
  AOI22_X1 U2763 ( .A1(n224), .A2(n787), .B1(n227), .B2(n2901), .ZN(n2204) );
  OAI211_X1 U2764 ( .C1(n2906), .C2(n230), .A(n2205), .B(n2206), .ZN(n2200) );
  AOI221_X1 U2765 ( .B1(n233), .B2(n921), .C1(n236), .C2(n2907), .A(n2207), 
        .ZN(n2206) );
  OAI22_X1 U2766 ( .A1(n2903), .A2(n239), .B1(n1308), .B2(n242), .ZN(n2207) );
  AOI22_X1 U2767 ( .A1(n245), .A2(n2908), .B1(n248), .B2(n821), .ZN(n2205) );
  NAND4_X1 U2768 ( .A1(n2208), .A2(n2209), .A3(n2210), .A4(n2211), .ZN(n2199)
         );
  AOI221_X1 U2769 ( .B1(n251), .B2(n2891), .C1(n254), .C2(n2892), .A(n2212), 
        .ZN(n2211) );
  OAI22_X1 U2770 ( .A1(n2890), .A2(n257), .B1(n2889), .B2(n260), .ZN(n2212) );
  AOI221_X1 U2771 ( .B1(n263), .B2(n2895), .C1(n266), .C2(n2896), .A(n2213), 
        .ZN(n2210) );
  OAI22_X1 U2772 ( .A1(n2894), .A2(n269), .B1(n2893), .B2(n272), .ZN(n2213) );
  AOI221_X1 U2773 ( .B1(n275), .B2(n618), .C1(n278), .C2(n651), .A(n2214), 
        .ZN(n2209) );
  OAI22_X1 U2774 ( .A1(n1316), .A2(n281), .B1(n1317), .B2(n284), .ZN(n2214) );
  AOI221_X1 U2775 ( .B1(n287), .B2(n584), .C1(n290), .C2(n3781), .A(n2215), 
        .ZN(n2208) );
  OAI22_X1 U2776 ( .A1(n1319), .A2(n293), .B1(n1320), .B2(n296), .ZN(n2215) );
  OAI222_X1 U2777 ( .A1(n309), .A2(n196), .B1(n2216), .B2(n199), .C1(n2468), 
        .C2(n203), .ZN(n2994) );
  NOR4_X1 U2778 ( .A1(n2217), .A2(n2218), .A3(n2219), .A4(n2220), .ZN(n2216)
         );
  OAI221_X1 U2779 ( .B1(n3844), .B2(n205), .C1(n1276), .C2(n208), .A(n2221), 
        .ZN(n2220) );
  AOI22_X1 U2780 ( .A1(n211), .A2(n2923), .B1(n214), .B2(n684), .ZN(n2221) );
  OAI221_X1 U2781 ( .B1(n1278), .B2(n217), .C1(n3748), .C2(n220), .A(n2222), 
        .ZN(n2219) );
  AOI22_X1 U2782 ( .A1(n223), .A2(n786), .B1(n226), .B2(n2922), .ZN(n2222) );
  OAI211_X1 U2783 ( .C1(n2927), .C2(n229), .A(n2223), .B(n2224), .ZN(n2218) );
  AOI221_X1 U2784 ( .B1(n232), .B2(n920), .C1(n235), .C2(n2928), .A(n2225), 
        .ZN(n2224) );
  OAI22_X1 U2785 ( .A1(n2924), .A2(n238), .B1(n1283), .B2(n241), .ZN(n2225) );
  AOI22_X1 U2786 ( .A1(n244), .A2(n2929), .B1(n247), .B2(n820), .ZN(n2223) );
  NAND4_X1 U2787 ( .A1(n2226), .A2(n2227), .A3(n2228), .A4(n2229), .ZN(n2217)
         );
  AOI221_X1 U2788 ( .B1(n250), .B2(n2912), .C1(n253), .C2(n2913), .A(n2230), 
        .ZN(n2229) );
  OAI22_X1 U2789 ( .A1(n2911), .A2(n256), .B1(n2910), .B2(n259), .ZN(n2230) );
  AOI221_X1 U2790 ( .B1(n262), .B2(n2916), .C1(n265), .C2(n2917), .A(n2231), 
        .ZN(n2228) );
  OAI22_X1 U2791 ( .A1(n2915), .A2(n268), .B1(n2914), .B2(n271), .ZN(n2231) );
  AOI221_X1 U2792 ( .B1(n274), .B2(n617), .C1(n277), .C2(n650), .A(n2232), 
        .ZN(n2227) );
  OAI22_X1 U2793 ( .A1(n1291), .A2(n280), .B1(n1292), .B2(n283), .ZN(n2232) );
  AOI221_X1 U2794 ( .B1(n286), .B2(n583), .C1(n289), .C2(n3780), .A(n2233), 
        .ZN(n2226) );
  OAI22_X1 U2795 ( .A1(n1294), .A2(n292), .B1(n1295), .B2(n295), .ZN(n2233) );
  OAI222_X1 U2796 ( .A1(n308), .A2(n196), .B1(n2234), .B2(n199), .C1(n2467), 
        .C2(n203), .ZN(n2993) );
  NOR4_X1 U2797 ( .A1(n2235), .A2(n2236), .A3(n2237), .A4(n2238), .ZN(n2234)
         );
  OAI221_X1 U2798 ( .B1(n3843), .B2(n205), .C1(n1251), .C2(n208), .A(n2239), 
        .ZN(n2238) );
  AOI22_X1 U2799 ( .A1(n211), .A2(n2944), .B1(n214), .B2(n683), .ZN(n2239) );
  OAI221_X1 U2800 ( .B1(n1253), .B2(n217), .C1(n3747), .C2(n220), .A(n2240), 
        .ZN(n2237) );
  AOI22_X1 U2801 ( .A1(n223), .A2(n785), .B1(n226), .B2(n2943), .ZN(n2240) );
  OAI211_X1 U2802 ( .C1(n2948), .C2(n229), .A(n2241), .B(n2242), .ZN(n2236) );
  AOI221_X1 U2803 ( .B1(n232), .B2(n919), .C1(n235), .C2(n2949), .A(n2243), 
        .ZN(n2242) );
  OAI22_X1 U2804 ( .A1(n2945), .A2(n238), .B1(n1258), .B2(n241), .ZN(n2243) );
  AOI22_X1 U2805 ( .A1(n244), .A2(n2950), .B1(n247), .B2(n819), .ZN(n2241) );
  NAND4_X1 U2806 ( .A1(n2244), .A2(n2245), .A3(n2246), .A4(n2247), .ZN(n2235)
         );
  AOI221_X1 U2807 ( .B1(n250), .B2(n2933), .C1(n253), .C2(n2934), .A(n2248), 
        .ZN(n2247) );
  OAI22_X1 U2808 ( .A1(n2932), .A2(n256), .B1(n2931), .B2(n259), .ZN(n2248) );
  AOI221_X1 U2809 ( .B1(n262), .B2(n2937), .C1(n265), .C2(n2938), .A(n2249), 
        .ZN(n2246) );
  OAI22_X1 U2810 ( .A1(n2936), .A2(n268), .B1(n2935), .B2(n271), .ZN(n2249) );
  AOI221_X1 U2811 ( .B1(n274), .B2(n616), .C1(n277), .C2(n649), .A(n2250), 
        .ZN(n2245) );
  OAI22_X1 U2812 ( .A1(n1266), .A2(n280), .B1(n1267), .B2(n283), .ZN(n2250) );
  AOI221_X1 U2813 ( .B1(n286), .B2(n582), .C1(n289), .C2(n3779), .A(n2251), 
        .ZN(n2244) );
  OAI22_X1 U2814 ( .A1(n1269), .A2(n292), .B1(n1270), .B2(n295), .ZN(n2251) );
  OAI222_X1 U2815 ( .A1(n307), .A2(n196), .B1(n2252), .B2(n199), .C1(n2466), 
        .C2(n202), .ZN(n2992) );
  NOR4_X1 U2816 ( .A1(n2253), .A2(n2254), .A3(n2255), .A4(n2256), .ZN(n2252)
         );
  OAI221_X1 U2817 ( .B1(n3842), .B2(n205), .C1(n1226), .C2(n208), .A(n2257), 
        .ZN(n2256) );
  AOI22_X1 U2818 ( .A1(n211), .A2(n2965), .B1(n214), .B2(n682), .ZN(n2257) );
  OAI221_X1 U2819 ( .B1(n1228), .B2(n217), .C1(n3746), .C2(n220), .A(n2258), 
        .ZN(n2255) );
  AOI22_X1 U2820 ( .A1(n223), .A2(n784), .B1(n226), .B2(n2964), .ZN(n2258) );
  OAI211_X1 U2821 ( .C1(n2969), .C2(n229), .A(n2259), .B(n2260), .ZN(n2254) );
  AOI221_X1 U2822 ( .B1(n232), .B2(n918), .C1(n235), .C2(n2970), .A(n2261), 
        .ZN(n2260) );
  OAI22_X1 U2823 ( .A1(n2966), .A2(n238), .B1(n1233), .B2(n241), .ZN(n2261) );
  AOI22_X1 U2824 ( .A1(n244), .A2(n2971), .B1(n247), .B2(n818), .ZN(n2259) );
  NAND4_X1 U2825 ( .A1(n2262), .A2(n2263), .A3(n2264), .A4(n2265), .ZN(n2253)
         );
  AOI221_X1 U2826 ( .B1(n250), .B2(n2954), .C1(n253), .C2(n2955), .A(n2266), 
        .ZN(n2265) );
  OAI22_X1 U2827 ( .A1(n2953), .A2(n256), .B1(n2952), .B2(n259), .ZN(n2266) );
  AOI221_X1 U2828 ( .B1(n262), .B2(n2958), .C1(n265), .C2(n2959), .A(n2267), 
        .ZN(n2264) );
  OAI22_X1 U2829 ( .A1(n2957), .A2(n268), .B1(n2956), .B2(n271), .ZN(n2267) );
  AOI221_X1 U2830 ( .B1(n274), .B2(n615), .C1(n277), .C2(n648), .A(n2268), 
        .ZN(n2263) );
  OAI22_X1 U2831 ( .A1(n1241), .A2(n280), .B1(n1242), .B2(n283), .ZN(n2268) );
  AOI221_X1 U2832 ( .B1(n286), .B2(n581), .C1(n289), .C2(n3778), .A(n2269), 
        .ZN(n2262) );
  OAI22_X1 U2833 ( .A1(n1244), .A2(n292), .B1(n1245), .B2(n295), .ZN(n2269) );
  OAI222_X1 U2834 ( .A1(n306), .A2(n196), .B1(n2270), .B2(n199), .C1(n2465), 
        .C2(n202), .ZN(n2991) );
  NOR4_X1 U2835 ( .A1(n2271), .A2(n2272), .A3(n2273), .A4(n2274), .ZN(n2270)
         );
  OAI221_X1 U2836 ( .B1(n3841), .B2(n205), .C1(n1201), .C2(n208), .A(n2275), 
        .ZN(n2274) );
  AOI22_X1 U2837 ( .A1(n211), .A2(n3562), .B1(n214), .B2(n681), .ZN(n2275) );
  OAI221_X1 U2838 ( .B1(n1203), .B2(n217), .C1(n3745), .C2(n220), .A(n2276), 
        .ZN(n2273) );
  AOI22_X1 U2839 ( .A1(n223), .A2(n783), .B1(n226), .B2(n3561), .ZN(n2276) );
  OAI211_X1 U2840 ( .C1(n3566), .C2(n229), .A(n2277), .B(n2278), .ZN(n2272) );
  AOI221_X1 U2841 ( .B1(n232), .B2(n917), .C1(n235), .C2(n3567), .A(n2279), 
        .ZN(n2278) );
  OAI22_X1 U2842 ( .A1(n3563), .A2(n238), .B1(n1208), .B2(n241), .ZN(n2279) );
  AOI22_X1 U2843 ( .A1(n244), .A2(n3568), .B1(n247), .B2(n817), .ZN(n2277) );
  NAND4_X1 U2844 ( .A1(n2280), .A2(n2281), .A3(n2282), .A4(n2283), .ZN(n2271)
         );
  AOI221_X1 U2845 ( .B1(n250), .B2(n2975), .C1(n253), .C2(n2976), .A(n2284), 
        .ZN(n2283) );
  OAI22_X1 U2846 ( .A1(n2974), .A2(n256), .B1(n2973), .B2(n259), .ZN(n2284) );
  AOI221_X1 U2847 ( .B1(n262), .B2(n2979), .C1(n265), .C2(n2980), .A(n2285), 
        .ZN(n2282) );
  OAI22_X1 U2848 ( .A1(n2978), .A2(n268), .B1(n2977), .B2(n271), .ZN(n2285) );
  AOI221_X1 U2849 ( .B1(n274), .B2(n614), .C1(n277), .C2(n647), .A(n2286), 
        .ZN(n2281) );
  OAI22_X1 U2850 ( .A1(n1216), .A2(n280), .B1(n1217), .B2(n283), .ZN(n2286) );
  AOI221_X1 U2851 ( .B1(n286), .B2(n580), .C1(n289), .C2(n3777), .A(n2287), 
        .ZN(n2280) );
  OAI22_X1 U2852 ( .A1(n1219), .A2(n292), .B1(n1220), .B2(n295), .ZN(n2287) );
  OAI222_X1 U2853 ( .A1(n305), .A2(n196), .B1(n2288), .B2(n199), .C1(n2464), 
        .C2(n202), .ZN(n2990) );
  NOR4_X1 U2854 ( .A1(n2289), .A2(n2290), .A3(n2291), .A4(n2292), .ZN(n2288)
         );
  OAI221_X1 U2855 ( .B1(n3840), .B2(n205), .C1(n1176), .C2(n208), .A(n2293), 
        .ZN(n2292) );
  AOI22_X1 U2856 ( .A1(n211), .A2(n3583), .B1(n214), .B2(n680), .ZN(n2293) );
  OAI221_X1 U2857 ( .B1(n1178), .B2(n217), .C1(n3744), .C2(n220), .A(n2294), 
        .ZN(n2291) );
  AOI22_X1 U2858 ( .A1(n223), .A2(n782), .B1(n226), .B2(n3582), .ZN(n2294) );
  OAI211_X1 U2859 ( .C1(n3587), .C2(n229), .A(n2295), .B(n2296), .ZN(n2290) );
  AOI221_X1 U2860 ( .B1(n232), .B2(n916), .C1(n235), .C2(n3588), .A(n2297), 
        .ZN(n2296) );
  OAI22_X1 U2861 ( .A1(n3584), .A2(n238), .B1(n1183), .B2(n241), .ZN(n2297) );
  AOI22_X1 U2862 ( .A1(n244), .A2(n3589), .B1(n247), .B2(n816), .ZN(n2295) );
  NAND4_X1 U2863 ( .A1(n2298), .A2(n2299), .A3(n2300), .A4(n2301), .ZN(n2289)
         );
  AOI221_X1 U2864 ( .B1(n250), .B2(n3572), .C1(n253), .C2(n3573), .A(n2302), 
        .ZN(n2301) );
  OAI22_X1 U2865 ( .A1(n3571), .A2(n256), .B1(n3570), .B2(n259), .ZN(n2302) );
  AOI221_X1 U2866 ( .B1(n262), .B2(n3576), .C1(n265), .C2(n3577), .A(n2303), 
        .ZN(n2300) );
  OAI22_X1 U2867 ( .A1(n3575), .A2(n268), .B1(n3574), .B2(n271), .ZN(n2303) );
  AOI221_X1 U2868 ( .B1(n274), .B2(n613), .C1(n277), .C2(n646), .A(n2304), 
        .ZN(n2299) );
  OAI22_X1 U2869 ( .A1(n1191), .A2(n280), .B1(n1192), .B2(n283), .ZN(n2304) );
  AOI221_X1 U2870 ( .B1(n286), .B2(n579), .C1(n289), .C2(n3776), .A(n2305), 
        .ZN(n2298) );
  OAI22_X1 U2871 ( .A1(n1194), .A2(n292), .B1(n1195), .B2(n295), .ZN(n2305) );
  OAI222_X1 U2872 ( .A1(n304), .A2(n196), .B1(n2306), .B2(n199), .C1(n2463), 
        .C2(n202), .ZN(n2989) );
  NOR4_X1 U2873 ( .A1(n2307), .A2(n2308), .A3(n2309), .A4(n2310), .ZN(n2306)
         );
  OAI221_X1 U2874 ( .B1(n3839), .B2(n205), .C1(n1151), .C2(n208), .A(n2311), 
        .ZN(n2310) );
  AOI22_X1 U2875 ( .A1(n211), .A2(n3604), .B1(n214), .B2(n679), .ZN(n2311) );
  OAI221_X1 U2876 ( .B1(n1153), .B2(n217), .C1(n3743), .C2(n220), .A(n2312), 
        .ZN(n2309) );
  AOI22_X1 U2877 ( .A1(n223), .A2(n781), .B1(n226), .B2(n3603), .ZN(n2312) );
  OAI211_X1 U2878 ( .C1(n3608), .C2(n229), .A(n2313), .B(n2314), .ZN(n2308) );
  AOI221_X1 U2879 ( .B1(n232), .B2(n915), .C1(n235), .C2(n3609), .A(n2315), 
        .ZN(n2314) );
  OAI22_X1 U2880 ( .A1(n3605), .A2(n238), .B1(n1158), .B2(n241), .ZN(n2315) );
  AOI22_X1 U2881 ( .A1(n244), .A2(n3610), .B1(n247), .B2(n815), .ZN(n2313) );
  NAND4_X1 U2882 ( .A1(n2316), .A2(n2317), .A3(n2318), .A4(n2319), .ZN(n2307)
         );
  AOI221_X1 U2883 ( .B1(n250), .B2(n3593), .C1(n253), .C2(n3594), .A(n2320), 
        .ZN(n2319) );
  OAI22_X1 U2884 ( .A1(n3592), .A2(n256), .B1(n3591), .B2(n259), .ZN(n2320) );
  AOI221_X1 U2885 ( .B1(n262), .B2(n3597), .C1(n265), .C2(n3598), .A(n2321), 
        .ZN(n2318) );
  OAI22_X1 U2886 ( .A1(n3596), .A2(n268), .B1(n3595), .B2(n271), .ZN(n2321) );
  AOI221_X1 U2887 ( .B1(n274), .B2(n612), .C1(n277), .C2(n645), .A(n2322), 
        .ZN(n2317) );
  OAI22_X1 U2888 ( .A1(n1166), .A2(n280), .B1(n1167), .B2(n283), .ZN(n2322) );
  AOI221_X1 U2889 ( .B1(n286), .B2(n578), .C1(n289), .C2(n3775), .A(n2323), 
        .ZN(n2316) );
  OAI22_X1 U2890 ( .A1(n1169), .A2(n292), .B1(n1170), .B2(n295), .ZN(n2323) );
  OAI222_X1 U2891 ( .A1(n303), .A2(n196), .B1(n2324), .B2(n199), .C1(n2462), 
        .C2(n202), .ZN(n2988) );
  NOR4_X1 U2892 ( .A1(n2325), .A2(n2326), .A3(n2327), .A4(n2328), .ZN(n2324)
         );
  OAI221_X1 U2893 ( .B1(n3838), .B2(n205), .C1(n1126), .C2(n208), .A(n2329), 
        .ZN(n2328) );
  AOI22_X1 U2894 ( .A1(n211), .A2(n3625), .B1(n214), .B2(n678), .ZN(n2329) );
  OAI221_X1 U2895 ( .B1(n1128), .B2(n217), .C1(n3742), .C2(n220), .A(n2330), 
        .ZN(n2327) );
  AOI22_X1 U2896 ( .A1(n223), .A2(n780), .B1(n226), .B2(n3624), .ZN(n2330) );
  OAI211_X1 U2897 ( .C1(n3629), .C2(n229), .A(n2331), .B(n2332), .ZN(n2326) );
  AOI221_X1 U2898 ( .B1(n232), .B2(n914), .C1(n235), .C2(n3630), .A(n2333), 
        .ZN(n2332) );
  OAI22_X1 U2899 ( .A1(n3626), .A2(n238), .B1(n1133), .B2(n241), .ZN(n2333) );
  AOI22_X1 U2900 ( .A1(n244), .A2(n3631), .B1(n247), .B2(n814), .ZN(n2331) );
  NAND4_X1 U2901 ( .A1(n2334), .A2(n2335), .A3(n2336), .A4(n2337), .ZN(n2325)
         );
  AOI221_X1 U2902 ( .B1(n250), .B2(n3614), .C1(n253), .C2(n3615), .A(n2338), 
        .ZN(n2337) );
  OAI22_X1 U2903 ( .A1(n3613), .A2(n256), .B1(n3612), .B2(n259), .ZN(n2338) );
  AOI221_X1 U2904 ( .B1(n262), .B2(n3618), .C1(n265), .C2(n3619), .A(n2339), 
        .ZN(n2336) );
  OAI22_X1 U2905 ( .A1(n3617), .A2(n268), .B1(n3616), .B2(n271), .ZN(n2339) );
  AOI221_X1 U2906 ( .B1(n274), .B2(n611), .C1(n277), .C2(n644), .A(n2340), 
        .ZN(n2335) );
  OAI22_X1 U2907 ( .A1(n1141), .A2(n280), .B1(n1142), .B2(n283), .ZN(n2340) );
  AOI221_X1 U2908 ( .B1(n286), .B2(n577), .C1(n289), .C2(n3774), .A(n2341), 
        .ZN(n2334) );
  OAI22_X1 U2909 ( .A1(n1144), .A2(n292), .B1(n1145), .B2(n295), .ZN(n2341) );
  OAI222_X1 U2910 ( .A1(n302), .A2(n196), .B1(n2342), .B2(n199), .C1(n2461), 
        .C2(n202), .ZN(n2987) );
  NOR4_X1 U2911 ( .A1(n2343), .A2(n2344), .A3(n2345), .A4(n2346), .ZN(n2342)
         );
  OAI221_X1 U2912 ( .B1(n3837), .B2(n205), .C1(n1101), .C2(n208), .A(n2347), 
        .ZN(n2346) );
  AOI22_X1 U2913 ( .A1(n211), .A2(n3646), .B1(n214), .B2(n677), .ZN(n2347) );
  OAI221_X1 U2914 ( .B1(n1103), .B2(n217), .C1(n3741), .C2(n220), .A(n2348), 
        .ZN(n2345) );
  AOI22_X1 U2915 ( .A1(n223), .A2(n779), .B1(n226), .B2(n3645), .ZN(n2348) );
  OAI211_X1 U2916 ( .C1(n3650), .C2(n229), .A(n2349), .B(n2350), .ZN(n2344) );
  AOI221_X1 U2917 ( .B1(n232), .B2(n913), .C1(n235), .C2(n3651), .A(n2351), 
        .ZN(n2350) );
  OAI22_X1 U2918 ( .A1(n3647), .A2(n238), .B1(n1108), .B2(n241), .ZN(n2351) );
  AOI22_X1 U2919 ( .A1(n244), .A2(n3652), .B1(n247), .B2(n813), .ZN(n2349) );
  NAND4_X1 U2920 ( .A1(n2352), .A2(n2353), .A3(n2354), .A4(n2355), .ZN(n2343)
         );
  AOI221_X1 U2921 ( .B1(n250), .B2(n3635), .C1(n253), .C2(n3636), .A(n2356), 
        .ZN(n2355) );
  OAI22_X1 U2922 ( .A1(n3634), .A2(n256), .B1(n3633), .B2(n259), .ZN(n2356) );
  AOI221_X1 U2923 ( .B1(n262), .B2(n3639), .C1(n265), .C2(n3640), .A(n2357), 
        .ZN(n2354) );
  OAI22_X1 U2924 ( .A1(n3638), .A2(n268), .B1(n3637), .B2(n271), .ZN(n2357) );
  AOI221_X1 U2925 ( .B1(n274), .B2(n610), .C1(n277), .C2(n643), .A(n2358), 
        .ZN(n2353) );
  OAI22_X1 U2926 ( .A1(n1116), .A2(n280), .B1(n1117), .B2(n283), .ZN(n2358) );
  AOI221_X1 U2927 ( .B1(n286), .B2(n576), .C1(n289), .C2(n3773), .A(n2359), 
        .ZN(n2352) );
  OAI22_X1 U2928 ( .A1(n1119), .A2(n292), .B1(n1120), .B2(n295), .ZN(n2359) );
  OAI222_X1 U2929 ( .A1(n301), .A2(n196), .B1(n2360), .B2(n199), .C1(n2460), 
        .C2(n202), .ZN(n2986) );
  NOR4_X1 U2930 ( .A1(n2361), .A2(n2362), .A3(n2363), .A4(n2364), .ZN(n2360)
         );
  OAI221_X1 U2931 ( .B1(n3836), .B2(n205), .C1(n1076), .C2(n208), .A(n2365), 
        .ZN(n2364) );
  AOI22_X1 U2932 ( .A1(n211), .A2(n3667), .B1(n214), .B2(n676), .ZN(n2365) );
  OAI221_X1 U2933 ( .B1(n1078), .B2(n217), .C1(n3740), .C2(n220), .A(n2366), 
        .ZN(n2363) );
  AOI22_X1 U2934 ( .A1(n223), .A2(n778), .B1(n226), .B2(n3666), .ZN(n2366) );
  OAI211_X1 U2935 ( .C1(n3671), .C2(n229), .A(n2367), .B(n2368), .ZN(n2362) );
  AOI221_X1 U2936 ( .B1(n232), .B2(n912), .C1(n235), .C2(n3672), .A(n2369), 
        .ZN(n2368) );
  OAI22_X1 U2937 ( .A1(n3668), .A2(n238), .B1(n1083), .B2(n241), .ZN(n2369) );
  AOI22_X1 U2938 ( .A1(n244), .A2(n3673), .B1(n247), .B2(n812), .ZN(n2367) );
  NAND4_X1 U2939 ( .A1(n2370), .A2(n2371), .A3(n2372), .A4(n2373), .ZN(n2361)
         );
  AOI221_X1 U2940 ( .B1(n250), .B2(n3656), .C1(n253), .C2(n3657), .A(n2374), 
        .ZN(n2373) );
  OAI22_X1 U2941 ( .A1(n3655), .A2(n256), .B1(n3654), .B2(n259), .ZN(n2374) );
  AOI221_X1 U2942 ( .B1(n262), .B2(n3660), .C1(n265), .C2(n3661), .A(n2375), 
        .ZN(n2372) );
  OAI22_X1 U2943 ( .A1(n3659), .A2(n268), .B1(n3658), .B2(n271), .ZN(n2375) );
  AOI221_X1 U2944 ( .B1(n274), .B2(n609), .C1(n277), .C2(n642), .A(n2376), 
        .ZN(n2371) );
  OAI22_X1 U2945 ( .A1(n1091), .A2(n280), .B1(n1092), .B2(n283), .ZN(n2376) );
  AOI221_X1 U2946 ( .B1(n286), .B2(n575), .C1(n289), .C2(n3772), .A(n2377), 
        .ZN(n2370) );
  OAI22_X1 U2947 ( .A1(n1094), .A2(n292), .B1(n1095), .B2(n295), .ZN(n2377) );
  OAI222_X1 U2948 ( .A1(n300), .A2(n196), .B1(n2378), .B2(n199), .C1(n2459), 
        .C2(n202), .ZN(n2985) );
  NOR4_X1 U2949 ( .A1(n2379), .A2(n2380), .A3(n2381), .A4(n2382), .ZN(n2378)
         );
  OAI221_X1 U2950 ( .B1(n3835), .B2(n205), .C1(n1051), .C2(n208), .A(n2383), 
        .ZN(n2382) );
  AOI22_X1 U2951 ( .A1(n211), .A2(n3688), .B1(n214), .B2(n675), .ZN(n2383) );
  OAI221_X1 U2952 ( .B1(n1053), .B2(n217), .C1(n3739), .C2(n220), .A(n2384), 
        .ZN(n2381) );
  AOI22_X1 U2953 ( .A1(n223), .A2(n777), .B1(n226), .B2(n3687), .ZN(n2384) );
  OAI211_X1 U2954 ( .C1(n3692), .C2(n229), .A(n2385), .B(n2386), .ZN(n2380) );
  AOI221_X1 U2955 ( .B1(n232), .B2(n911), .C1(n235), .C2(n3693), .A(n2387), 
        .ZN(n2386) );
  OAI22_X1 U2956 ( .A1(n3689), .A2(n238), .B1(n1058), .B2(n241), .ZN(n2387) );
  AOI22_X1 U2957 ( .A1(n244), .A2(n3694), .B1(n247), .B2(n811), .ZN(n2385) );
  NAND4_X1 U2958 ( .A1(n2388), .A2(n2389), .A3(n2390), .A4(n2391), .ZN(n2379)
         );
  AOI221_X1 U2959 ( .B1(n250), .B2(n3677), .C1(n253), .C2(n3678), .A(n2392), 
        .ZN(n2391) );
  OAI22_X1 U2960 ( .A1(n3676), .A2(n256), .B1(n3675), .B2(n259), .ZN(n2392) );
  AOI221_X1 U2961 ( .B1(n262), .B2(n3681), .C1(n265), .C2(n3682), .A(n2393), 
        .ZN(n2390) );
  OAI22_X1 U2962 ( .A1(n3680), .A2(n268), .B1(n3679), .B2(n271), .ZN(n2393) );
  AOI221_X1 U2963 ( .B1(n274), .B2(n608), .C1(n277), .C2(n641), .A(n2394), 
        .ZN(n2389) );
  OAI22_X1 U2964 ( .A1(n1066), .A2(n280), .B1(n1067), .B2(n283), .ZN(n2394) );
  AOI221_X1 U2965 ( .B1(n286), .B2(n574), .C1(n289), .C2(n3771), .A(n2395), 
        .ZN(n2388) );
  OAI22_X1 U2966 ( .A1(n1069), .A2(n292), .B1(n1070), .B2(n295), .ZN(n2395) );
  OAI222_X1 U2967 ( .A1(n299), .A2(n196), .B1(n2396), .B2(n199), .C1(n2458), 
        .C2(n202), .ZN(n2984) );
  NOR4_X1 U2968 ( .A1(n2397), .A2(n2398), .A3(n2399), .A4(n2400), .ZN(n2396)
         );
  OAI221_X1 U2969 ( .B1(n3834), .B2(n205), .C1(n1026), .C2(n208), .A(n2401), 
        .ZN(n2400) );
  AOI22_X1 U2970 ( .A1(n211), .A2(n3709), .B1(n214), .B2(n674), .ZN(n2401) );
  OAI221_X1 U2971 ( .B1(n1028), .B2(n217), .C1(n3738), .C2(n220), .A(n2402), 
        .ZN(n2399) );
  AOI22_X1 U2972 ( .A1(n223), .A2(n776), .B1(n226), .B2(n3708), .ZN(n2402) );
  OAI211_X1 U2973 ( .C1(n3713), .C2(n229), .A(n2403), .B(n2404), .ZN(n2398) );
  AOI221_X1 U2974 ( .B1(n232), .B2(n910), .C1(n235), .C2(n3714), .A(n2405), 
        .ZN(n2404) );
  OAI22_X1 U2975 ( .A1(n3710), .A2(n238), .B1(n1033), .B2(n241), .ZN(n2405) );
  AOI22_X1 U2976 ( .A1(n244), .A2(n3715), .B1(n247), .B2(n810), .ZN(n2403) );
  NAND4_X1 U2977 ( .A1(n2406), .A2(n2407), .A3(n2408), .A4(n2409), .ZN(n2397)
         );
  AOI221_X1 U2978 ( .B1(n250), .B2(n3698), .C1(n253), .C2(n3699), .A(n2410), 
        .ZN(n2409) );
  OAI22_X1 U2979 ( .A1(n3697), .A2(n256), .B1(n3696), .B2(n259), .ZN(n2410) );
  AOI221_X1 U2980 ( .B1(n262), .B2(n3702), .C1(n265), .C2(n3703), .A(n2411), 
        .ZN(n2408) );
  OAI22_X1 U2981 ( .A1(n3701), .A2(n268), .B1(n3700), .B2(n271), .ZN(n2411) );
  AOI221_X1 U2982 ( .B1(n274), .B2(n607), .C1(n277), .C2(n640), .A(n2412), 
        .ZN(n2407) );
  OAI22_X1 U2983 ( .A1(n1041), .A2(n280), .B1(n1042), .B2(n283), .ZN(n2412) );
  AOI221_X1 U2984 ( .B1(n286), .B2(n573), .C1(n289), .C2(n3770), .A(n2413), 
        .ZN(n2406) );
  OAI22_X1 U2985 ( .A1(n1044), .A2(n292), .B1(n1045), .B2(n295), .ZN(n2413) );
  OAI222_X1 U2986 ( .A1(n298), .A2(n196), .B1(n2414), .B2(n199), .C1(n2457), 
        .C2(n202), .ZN(n2983) );
  NAND2_X1 U2987 ( .A1(n202), .A2(n2415), .ZN(n1824) );
  NOR4_X1 U2988 ( .A1(n2416), .A2(n2417), .A3(n2418), .A4(n2419), .ZN(n2414)
         );
  OAI221_X1 U2989 ( .B1(n3833), .B2(n205), .C1(n971), .C2(n208), .A(n2420), 
        .ZN(n2419) );
  AOI22_X1 U2990 ( .A1(n211), .A2(n3730), .B1(n214), .B2(n673), .ZN(n2420) );
  AND2_X1 U2991 ( .A1(n2421), .A2(n2422), .ZN(n1834) );
  AND2_X1 U2992 ( .A1(n2421), .A2(n2423), .ZN(n1833) );
  NAND2_X1 U2993 ( .A1(n2424), .A2(n2425), .ZN(n1831) );
  NAND2_X1 U2994 ( .A1(n2426), .A2(n2422), .ZN(n1830) );
  OAI221_X1 U2995 ( .B1(n976), .B2(n217), .C1(n3737), .C2(n220), .A(n2427), 
        .ZN(n2418) );
  AOI22_X1 U2996 ( .A1(n223), .A2(n774), .B1(n226), .B2(n3729), .ZN(n2427) );
  AND2_X1 U2997 ( .A1(n2426), .A2(n2423), .ZN(n1839) );
  AND2_X1 U2998 ( .A1(n2426), .A2(n2425), .ZN(n1838) );
  NAND2_X1 U2999 ( .A1(n2421), .A2(n2425), .ZN(n1836) );
  NAND2_X1 U3000 ( .A1(n2421), .A2(n2428), .ZN(n1835) );
  NOR3_X1 U3001 ( .A1(n2429), .A2(ADD_RS1[0]), .A3(n2430), .ZN(n2421) );
  OAI211_X1 U3002 ( .C1(n3734), .C2(n229), .A(n2431), .B(n2432), .ZN(n2417) );
  AOI221_X1 U3003 ( .B1(n232), .B2(n908), .C1(n235), .C2(n3735), .A(n2433), 
        .ZN(n2432) );
  OAI22_X1 U3004 ( .A1(n3731), .A2(n238), .B1(n989), .B2(n241), .ZN(n2433) );
  NAND2_X1 U3005 ( .A1(n2434), .A2(n2425), .ZN(n1847) );
  NAND2_X1 U3006 ( .A1(n2434), .A2(n2428), .ZN(n1846) );
  AND2_X1 U3007 ( .A1(n2424), .A2(n2422), .ZN(n1844) );
  AND2_X1 U3008 ( .A1(n2424), .A2(n2428), .ZN(n1843) );
  AOI22_X1 U3009 ( .A1(n244), .A2(n3736), .B1(n247), .B2(n808), .ZN(n2431) );
  AND2_X1 U3010 ( .A1(n2434), .A2(n2423), .ZN(n1849) );
  AND2_X1 U3011 ( .A1(n2434), .A2(n2422), .ZN(n1848) );
  NOR3_X1 U3012 ( .A1(ADD_RS1[0]), .A2(ADD_RS1[3]), .A3(n2429), .ZN(n2434) );
  NAND2_X1 U3013 ( .A1(n2424), .A2(n2423), .ZN(n1840) );
  NOR3_X1 U3014 ( .A1(n2435), .A2(ADD_RS1[3]), .A3(n2429), .ZN(n2424) );
  NAND4_X1 U3015 ( .A1(n2436), .A2(n2437), .A3(n2438), .A4(n2439), .ZN(n2416)
         );
  AOI221_X1 U3016 ( .B1(n250), .B2(n3719), .C1(n253), .C2(n3720), .A(n2440), 
        .ZN(n2439) );
  OAI22_X1 U3017 ( .A1(n3718), .A2(n256), .B1(n3717), .B2(n259), .ZN(n2440) );
  NAND2_X1 U3018 ( .A1(n2428), .A2(n2441), .ZN(n1858) );
  NAND2_X1 U3019 ( .A1(n2428), .A2(n2442), .ZN(n1857) );
  AND2_X1 U3020 ( .A1(n2441), .A2(n2425), .ZN(n1855) );
  AND2_X1 U3021 ( .A1(n2425), .A2(n2442), .ZN(n1854) );
  AOI221_X1 U3022 ( .B1(n262), .B2(n3723), .C1(n265), .C2(n3724), .A(n2443), 
        .ZN(n2438) );
  OAI22_X1 U3023 ( .A1(n3722), .A2(n268), .B1(n3721), .B2(n271), .ZN(n2443) );
  NAND2_X1 U3024 ( .A1(n2423), .A2(n2441), .ZN(n1863) );
  NAND2_X1 U3025 ( .A1(n2423), .A2(n2442), .ZN(n1862) );
  AND2_X1 U3026 ( .A1(n2422), .A2(n2441), .ZN(n1860) );
  NOR3_X1 U3027 ( .A1(ADD_RS1[0]), .A2(ADD_RS1[4]), .A3(n2430), .ZN(n2441) );
  AND2_X1 U3028 ( .A1(n2422), .A2(n2442), .ZN(n1859) );
  NOR3_X1 U3029 ( .A1(n2435), .A2(ADD_RS1[4]), .A3(n2430), .ZN(n2442) );
  AOI221_X1 U3030 ( .B1(n274), .B2(n605), .C1(n277), .C2(n638), .A(n2444), 
        .ZN(n2437) );
  OAI22_X1 U3031 ( .A1(n1010), .A2(n280), .B1(n1012), .B2(n283), .ZN(n2444) );
  NAND2_X1 U3032 ( .A1(n2445), .A2(n2425), .ZN(n1868) );
  NAND2_X1 U3033 ( .A1(n2446), .A2(n2425), .ZN(n1867) );
  NOR2_X1 U3034 ( .A1(n2447), .A2(n2448), .ZN(n2425) );
  AND2_X1 U3035 ( .A1(n2445), .A2(n2428), .ZN(n1865) );
  AND2_X1 U3036 ( .A1(n2446), .A2(n2428), .ZN(n1864) );
  AOI221_X1 U3037 ( .B1(n286), .B2(n571), .C1(n289), .C2(n3769), .A(n2449), 
        .ZN(n2436) );
  OAI22_X1 U3038 ( .A1(n1017), .A2(n292), .B1(n1019), .B2(n295), .ZN(n2449) );
  NAND2_X1 U3039 ( .A1(n2445), .A2(n2422), .ZN(n1873) );
  NAND2_X1 U3040 ( .A1(n2446), .A2(n2422), .ZN(n1872) );
  NOR2_X1 U3041 ( .A1(n2448), .A2(ADD_RS1[2]), .ZN(n2422) );
  NOR3_X1 U3042 ( .A1(ADD_RS1[3]), .A2(ADD_RS1[4]), .A3(ADD_RS1[0]), .ZN(n2446) );
  AND2_X1 U3043 ( .A1(n2426), .A2(n2428), .ZN(n1870) );
  NOR2_X1 U3044 ( .A1(n2447), .A2(ADD_RS1[1]), .ZN(n2428) );
  INV_X1 U3045 ( .A(ADD_RS1[2]), .ZN(n2447) );
  NOR3_X1 U3046 ( .A1(n2429), .A2(n2435), .A3(n2430), .ZN(n2426) );
  INV_X1 U3047 ( .A(ADD_RS1[3]), .ZN(n2430) );
  INV_X1 U3048 ( .A(ADD_RS1[4]), .ZN(n2429) );
  AND2_X1 U3049 ( .A1(n2445), .A2(n2423), .ZN(n1869) );
  NOR2_X1 U3050 ( .A1(ADD_RS1[1]), .A2(ADD_RS1[2]), .ZN(n2423) );
  NOR3_X1 U3051 ( .A1(ADD_RS1[3]), .A2(ADD_RS1[4]), .A3(n2435), .ZN(n2445) );
  INV_X1 U3052 ( .A(ADD_RS1[0]), .ZN(n2435) );
  NAND2_X1 U3053 ( .A1(n2450), .A2(n202), .ZN(n1822) );
  AND3_X1 U3054 ( .A1(n419), .A2(ENABLE), .A3(RD1), .ZN(n1825) );
  INV_X1 U3055 ( .A(n2415), .ZN(n2450) );
  NAND4_X1 U3056 ( .A1(n2451), .A2(n2452), .A3(n2453), .A4(n2454), .ZN(n2415)
         );
  NOR3_X1 U3057 ( .A1(n2455), .A2(n1820), .A3(n2456), .ZN(n2454) );
  XNOR2_X1 U3058 ( .A(ADD_WR[1]), .B(n2448), .ZN(n2456) );
  INV_X1 U3059 ( .A(ADD_RS1[1]), .ZN(n2448) );
  INV_X1 U3060 ( .A(WR), .ZN(n1820) );
  XNOR2_X1 U3061 ( .A(n953), .B(ADD_RS1[0]), .ZN(n2455) );
  INV_X1 U3062 ( .A(ADD_WR[0]), .ZN(n953) );
  XNOR2_X1 U3063 ( .A(ADD_WR[3]), .B(ADD_RS1[3]), .ZN(n2453) );
  XNOR2_X1 U3064 ( .A(ADD_WR[4]), .B(ADD_RS1[4]), .ZN(n2452) );
  XNOR2_X1 U3065 ( .A(ADD_RS1[2]), .B(ADD_WR[2]), .ZN(n2451) );
endmodule


module Decode ( CLK, RST, REG_LATCH_EN, RD1, RD2, RF_WE, ZERO_FLAG, PC_IN, 
        INS_IN, ADD_WR, DATA_WR_IN, PC_OUT, A_OUT, B_OUT, IMM_OUT, ADD_RS1_HDU, 
        ADD_RS2_HDU, ADD_WR_OUT, ADD_RS1_OUT, ADD_RS2_OUT );
  input [31:0] PC_IN;
  input [31:0] INS_IN;
  input [4:0] ADD_WR;
  input [31:0] DATA_WR_IN;
  output [31:0] PC_OUT;
  output [31:0] A_OUT;
  output [31:0] B_OUT;
  output [31:0] IMM_OUT;
  output [4:0] ADD_RS1_HDU;
  output [4:0] ADD_RS2_HDU;
  output [4:0] ADD_WR_OUT;
  output [4:0] ADD_RS1_OUT;
  output [4:0] ADD_RS2_OUT;
  input CLK, RST, REG_LATCH_EN, RD1, RD2, RF_WE, ZERO_FLAG;
  wire   sig_RST, sig_Rtype, sig_Itype, sig_Jtype, n1;
  wire   [4:0] sig_ADD_WR;
  wire   [31:0] sig_IMM;

  NOR2_X2 U2 ( .A1(ZERO_FLAG), .A2(n1), .ZN(sig_RST) );
  instruction_type ins_type ( .INST_IN(INS_IN), .Rtype(sig_Rtype), .Itype(
        sig_Itype), .Jtype(sig_Jtype) );
  instruction_decomposition ins_dec ( .INST_IN(INS_IN), .Rtype(sig_Rtype), 
        .Itype(sig_Itype), .Jtype(sig_Jtype), .ADD_RS1(ADD_RS1_HDU), .ADD_RS2(
        ADD_RS2_HDU), .ADD_WR(sig_ADD_WR), .IMM(sig_IMM) );
  regn_N32_8 regPC ( .DIN(PC_IN), .CLK(CLK), .EN(1'b1), .RST(sig_RST), .DOUT(
        PC_OUT) );
  regn_N32_7 regIMM ( .DIN(sig_IMM), .CLK(CLK), .EN(REG_LATCH_EN), .RST(
        sig_RST), .DOUT(IMM_OUT) );
  regn_N5_0 regWR ( .DIN(sig_ADD_WR), .CLK(CLK), .EN(REG_LATCH_EN), .RST(
        sig_RST), .DOUT(ADD_WR_OUT) );
  regn_N5_4 regRS1 ( .DIN(ADD_RS1_HDU), .CLK(CLK), .EN(REG_LATCH_EN), .RST(
        sig_RST), .DOUT(ADD_RS1_OUT) );
  regn_N5_3 regRS2 ( .DIN(ADD_RS2_HDU), .CLK(CLK), .EN(REG_LATCH_EN), .RST(
        sig_RST), .DOUT(ADD_RS2_OUT) );
  register_file_NBIT_ADD5_NBIT_DATA32 rf ( .CLK(CLK), .RST(RST), .ENABLE(
        REG_LATCH_EN), .RD1(RD1), .RD2(RD2), .WR(RF_WE), .ADD_WR(ADD_WR), 
        .ADD_RS1(ADD_RS1_HDU), .ADD_RS2(ADD_RS2_HDU), .DATAIN(DATA_WR_IN), 
        .OUT1(A_OUT), .OUT2(B_OUT) );
  INV_X1 U3 ( .A(RST), .ZN(n1) );
endmodule


module Branch_Cond_Unit_NBIT32 ( RST, A, .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , 
        \ALU_OPC[1] , \ALU_OPC[0] }), JUMP_TYPE, PC_SEL, ZERO );
  input [31:0] A;
  input [1:0] JUMP_TYPE;
  output [1:0] PC_SEL;
  input RST, \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] ;
  output ZERO;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n1, n2;
  wire   [3:0] ALU_OPC;

  NOR4_X1 U3 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n15) );
  NOR4_X1 U4 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n19) );
  NAND4_X1 U5 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .ZN(n11) );
  NOR4_X1 U6 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n12) );
  NOR4_X1 U7 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n13) );
  NOR4_X1 U8 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n14) );
  NAND4_X1 U9 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .ZN(n10) );
  NOR4_X1 U10 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n16) );
  NOR4_X1 U11 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n17) );
  NOR4_X1 U12 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n18) );
  NOR4_X1 U13 ( .A1(ALU_OPC[0]), .A2(n1), .A3(ALU_OPC[2]), .A4(ALU_OPC[1]), 
        .ZN(n7) );
  OAI211_X1 U14 ( .C1(n5), .C2(n6), .A(JUMP_TYPE[0]), .B(RST), .ZN(n4) );
  AND2_X1 U15 ( .A1(n7), .A2(n8), .ZN(n6) );
  NOR4_X1 U16 ( .A1(n8), .A2(n9), .A3(n7), .A4(n1), .ZN(n5) );
  NOR2_X1 U17 ( .A1(n10), .A2(n11), .ZN(n8) );
  NAND2_X1 U18 ( .A1(JUMP_TYPE[1]), .A2(RST), .ZN(n3) );
  INV_X1 U19 ( .A(ALU_OPC[3]), .ZN(n1) );
  NAND2_X1 U20 ( .A1(n3), .A2(n4), .ZN(ZERO) );
  OAI22_X1 U21 ( .A1(JUMP_TYPE[0]), .A2(n3), .B1(JUMP_TYPE[1]), .B2(n4), .ZN(
        PC_SEL[0]) );
  NOR2_X1 U22 ( .A1(n2), .A2(n3), .ZN(PC_SEL[1]) );
  INV_X1 U23 ( .A(JUMP_TYPE[0]), .ZN(n2) );
  OR2_X1 U24 ( .A1(ALU_OPC[1]), .A2(ALU_OPC[2]), .ZN(n9) );
endmodule


module ff_1 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n4, n5, n6;

  DFFR_X1 Q_reg ( .D(n4), .CK(CLK), .RN(RST), .Q(Q), .QN(n5) );
  OAI21_X1 U2 ( .B1(n5), .B2(EN), .A(n6), .ZN(n4) );
  NAND2_X1 U3 ( .A1(EN), .A2(D), .ZN(n6) );
endmodule


module regn_N2 ( DIN, CLK, EN, RST, DOUT );
  input [1:0] DIN;
  output [1:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n4, n5, n6;

  DFFR_X1 \DOUT_reg[1]  ( .D(n6), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n4) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n5), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n3) );
  OAI21_X1 U2 ( .B1(n3), .B2(EN), .A(n1), .ZN(n5) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n1) );
  OAI21_X1 U4 ( .B1(n4), .B2(EN), .A(n2), .ZN(n6) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n2) );
endmodule


module FWD_Unit ( RST, ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB, RF_WE_MEM, 
        RF_WE_WB, FWDA, FWDB );
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [4:0] ADD_WR_MEM;
  input [4:0] ADD_WR_WB;
  output [1:0] FWDA;
  output [1:0] FWDB;
  input RST, RF_WE_MEM, RF_WE_WB;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42;

  NOR2_X1 U3 ( .A1(n1), .A2(n2), .ZN(FWDB[1]) );
  AOI21_X1 U4 ( .B1(n3), .B2(n4), .A(n5), .ZN(n1) );
  INV_X1 U5 ( .A(n6), .ZN(n3) );
  NOR2_X1 U6 ( .A1(n2), .A2(n7), .ZN(FWDB[0]) );
  MUX2_X1 U7 ( .A(n6), .B(n8), .S(n5), .Z(n7) );
  AND4_X1 U8 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n5) );
  NOR2_X1 U9 ( .A1(n13), .A2(n14), .ZN(n12) );
  XOR2_X1 U10 ( .A(ADD_WR_MEM[4]), .B(ADD_RS2[4]), .Z(n14) );
  XOR2_X1 U11 ( .A(ADD_WR_MEM[3]), .B(ADD_RS2[3]), .Z(n13) );
  XNOR2_X1 U12 ( .A(ADD_RS2[1]), .B(ADD_WR_MEM[1]), .ZN(n11) );
  XNOR2_X1 U13 ( .A(ADD_RS2[2]), .B(ADD_WR_MEM[2]), .ZN(n10) );
  XNOR2_X1 U14 ( .A(ADD_RS2[0]), .B(ADD_WR_MEM[0]), .ZN(n9) );
  NAND4_X1 U15 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(n6) );
  NOR2_X1 U16 ( .A1(n19), .A2(n20), .ZN(n18) );
  XOR2_X1 U17 ( .A(ADD_WR_WB[3]), .B(ADD_RS2[3]), .Z(n20) );
  XOR2_X1 U18 ( .A(ADD_WR_WB[2]), .B(ADD_RS2[2]), .Z(n19) );
  XNOR2_X1 U19 ( .A(ADD_RS2[4]), .B(ADD_WR_WB[4]), .ZN(n17) );
  XNOR2_X1 U20 ( .A(ADD_RS2[1]), .B(ADD_WR_WB[1]), .ZN(n16) );
  XNOR2_X1 U21 ( .A(ADD_RS2[0]), .B(ADD_WR_WB[0]), .ZN(n15) );
  NOR2_X1 U22 ( .A1(n21), .A2(n2), .ZN(FWDA[1]) );
  AOI21_X1 U23 ( .B1(n22), .B2(n4), .A(n23), .ZN(n21) );
  OAI21_X1 U24 ( .B1(n24), .B2(n25), .A(RF_WE_WB), .ZN(n4) );
  OR2_X1 U25 ( .A1(ADD_WR_WB[0]), .A2(ADD_WR_WB[1]), .ZN(n25) );
  OR3_X1 U26 ( .A1(ADD_WR_WB[3]), .A2(ADD_WR_WB[4]), .A3(ADD_WR_WB[2]), .ZN(
        n24) );
  INV_X1 U27 ( .A(n26), .ZN(n22) );
  NOR2_X1 U28 ( .A1(n2), .A2(n27), .ZN(FWDA[0]) );
  MUX2_X1 U29 ( .A(n26), .B(n8), .S(n23), .Z(n27) );
  AND4_X1 U30 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n23) );
  NOR2_X1 U31 ( .A1(n32), .A2(n33), .ZN(n31) );
  XOR2_X1 U32 ( .A(ADD_WR_MEM[4]), .B(ADD_RS1[4]), .Z(n33) );
  XOR2_X1 U33 ( .A(ADD_WR_MEM[3]), .B(ADD_RS1[3]), .Z(n32) );
  XNOR2_X1 U34 ( .A(ADD_RS1[1]), .B(ADD_WR_MEM[1]), .ZN(n30) );
  XNOR2_X1 U35 ( .A(ADD_RS1[2]), .B(ADD_WR_MEM[2]), .ZN(n29) );
  XNOR2_X1 U36 ( .A(ADD_RS1[0]), .B(ADD_WR_MEM[0]), .ZN(n28) );
  INV_X1 U37 ( .A(n34), .ZN(n8) );
  OAI21_X1 U38 ( .B1(n35), .B2(n36), .A(RF_WE_MEM), .ZN(n34) );
  OR2_X1 U39 ( .A1(ADD_WR_MEM[0]), .A2(ADD_WR_MEM[1]), .ZN(n36) );
  OR3_X1 U40 ( .A1(ADD_WR_MEM[3]), .A2(ADD_WR_MEM[4]), .A3(ADD_WR_MEM[2]), 
        .ZN(n35) );
  NAND4_X1 U41 ( .A1(n37), .A2(n38), .A3(n39), .A4(n40), .ZN(n26) );
  NOR2_X1 U42 ( .A1(n41), .A2(n42), .ZN(n40) );
  XOR2_X1 U43 ( .A(ADD_WR_WB[3]), .B(ADD_RS1[3]), .Z(n42) );
  XOR2_X1 U44 ( .A(ADD_WR_WB[2]), .B(ADD_RS1[2]), .Z(n41) );
  XNOR2_X1 U45 ( .A(ADD_RS1[4]), .B(ADD_WR_WB[4]), .ZN(n39) );
  XNOR2_X1 U46 ( .A(ADD_RS1[1]), .B(ADD_WR_WB[1]), .ZN(n38) );
  XNOR2_X1 U47 ( .A(ADD_RS1[0]), .B(ADD_WR_WB[0]), .ZN(n37) );
  INV_X1 U48 ( .A(RST), .ZN(n2) );
endmodule


module mux41_NBIT32_0 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n1, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  BUF_X1 U1 ( .A(n6), .Z(n72) );
  BUF_X1 U2 ( .A(n6), .Z(n73) );
  BUF_X1 U3 ( .A(n4), .Z(n78) );
  BUF_X1 U4 ( .A(n4), .Z(n79) );
  BUF_X1 U5 ( .A(n7), .Z(n1) );
  BUF_X1 U6 ( .A(n7), .Z(n70) );
  BUF_X1 U7 ( .A(n5), .Z(n75) );
  BUF_X1 U8 ( .A(n5), .Z(n76) );
  BUF_X1 U9 ( .A(n6), .Z(n74) );
  BUF_X1 U10 ( .A(n4), .Z(n80) );
  BUF_X1 U11 ( .A(n7), .Z(n71) );
  BUF_X1 U12 ( .A(n5), .Z(n77) );
  NOR2_X1 U13 ( .A1(n81), .A2(S[1]), .ZN(n6) );
  NOR2_X1 U14 ( .A1(S[0]), .A2(S[1]), .ZN(n7) );
  AND2_X1 U15 ( .A1(S[1]), .A2(S[0]), .ZN(n4) );
  AND2_X1 U16 ( .A1(S[1]), .A2(n81), .ZN(n5) );
  INV_X1 U17 ( .A(S[0]), .ZN(n81) );
  NAND2_X1 U18 ( .A1(n68), .A2(n69), .ZN(Z[0]) );
  AOI22_X1 U19 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n69) );
  AOI22_X1 U20 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n68) );
  NAND2_X1 U21 ( .A1(n44), .A2(n45), .ZN(Z[20]) );
  AOI22_X1 U22 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n45) );
  AOI22_X1 U23 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n44) );
  NAND2_X1 U24 ( .A1(n52), .A2(n53), .ZN(Z[17]) );
  AOI22_X1 U25 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n53) );
  AOI22_X1 U26 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n52) );
  NAND2_X1 U27 ( .A1(n60), .A2(n61), .ZN(Z[13]) );
  AOI22_X1 U28 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n61) );
  AOI22_X1 U29 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n60) );
  NAND2_X1 U30 ( .A1(n12), .A2(n13), .ZN(Z[6]) );
  AOI22_X1 U31 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n13) );
  AOI22_X1 U32 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n12) );
  NAND2_X1 U33 ( .A1(n20), .A2(n21), .ZN(Z[31]) );
  AOI22_X1 U34 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n21) );
  AOI22_X1 U35 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n20) );
  NAND2_X1 U36 ( .A1(n28), .A2(n29), .ZN(Z[28]) );
  AOI22_X1 U37 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n29) );
  AOI22_X1 U38 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n28) );
  NAND2_X1 U39 ( .A1(n36), .A2(n37), .ZN(Z[24]) );
  AOI22_X1 U40 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n37) );
  AOI22_X1 U41 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n36) );
  NAND2_X1 U42 ( .A1(n42), .A2(n43), .ZN(Z[21]) );
  AOI22_X1 U43 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n43) );
  AOI22_X1 U44 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n42) );
  NAND2_X1 U45 ( .A1(n50), .A2(n51), .ZN(Z[18]) );
  AOI22_X1 U46 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n51) );
  AOI22_X1 U47 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n50) );
  NAND2_X1 U48 ( .A1(n58), .A2(n59), .ZN(Z[14]) );
  AOI22_X1 U49 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n59) );
  AOI22_X1 U50 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n58) );
  NAND2_X1 U51 ( .A1(n66), .A2(n67), .ZN(Z[10]) );
  AOI22_X1 U52 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n67) );
  AOI22_X1 U53 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n66) );
  NAND2_X1 U54 ( .A1(n10), .A2(n11), .ZN(Z[7]) );
  AOI22_X1 U55 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n11) );
  AOI22_X1 U56 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n10) );
  NAND2_X1 U57 ( .A1(n18), .A2(n19), .ZN(Z[3]) );
  AOI22_X1 U58 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n19) );
  AOI22_X1 U59 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n18) );
  NAND2_X1 U60 ( .A1(n26), .A2(n27), .ZN(Z[29]) );
  AOI22_X1 U61 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n27) );
  AOI22_X1 U62 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n26) );
  NAND2_X1 U63 ( .A1(n34), .A2(n35), .ZN(Z[25]) );
  AOI22_X1 U64 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n35) );
  AOI22_X1 U65 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n34) );
  NAND2_X1 U66 ( .A1(n40), .A2(n41), .ZN(Z[22]) );
  AOI22_X1 U67 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n41) );
  AOI22_X1 U68 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n40) );
  NAND2_X1 U69 ( .A1(n48), .A2(n49), .ZN(Z[19]) );
  AOI22_X1 U70 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n49) );
  AOI22_X1 U71 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n48) );
  NAND2_X1 U72 ( .A1(n56), .A2(n57), .ZN(Z[15]) );
  AOI22_X1 U73 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n57) );
  AOI22_X1 U74 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n56) );
  NAND2_X1 U75 ( .A1(n64), .A2(n65), .ZN(Z[11]) );
  AOI22_X1 U76 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n65) );
  AOI22_X1 U77 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n64) );
  NAND2_X1 U78 ( .A1(n8), .A2(n9), .ZN(Z[8]) );
  AOI22_X1 U79 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n9) );
  AOI22_X1 U80 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n8) );
  NAND2_X1 U81 ( .A1(n16), .A2(n17), .ZN(Z[4]) );
  AOI22_X1 U82 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n17) );
  AOI22_X1 U83 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n16) );
  NAND2_X1 U84 ( .A1(n24), .A2(n25), .ZN(Z[2]) );
  AOI22_X1 U85 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n25) );
  AOI22_X1 U86 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n24) );
  NAND2_X1 U87 ( .A1(n32), .A2(n33), .ZN(Z[26]) );
  AOI22_X1 U88 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n33) );
  AOI22_X1 U89 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n32) );
  NAND2_X1 U90 ( .A1(n38), .A2(n39), .ZN(Z[23]) );
  AOI22_X1 U91 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n39) );
  AOI22_X1 U92 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n38) );
  NAND2_X1 U93 ( .A1(n46), .A2(n47), .ZN(Z[1]) );
  AOI22_X1 U94 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n47) );
  AOI22_X1 U95 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n46) );
  NAND2_X1 U96 ( .A1(n54), .A2(n55), .ZN(Z[16]) );
  AOI22_X1 U97 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n55) );
  AOI22_X1 U98 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n54) );
  NAND2_X1 U99 ( .A1(n62), .A2(n63), .ZN(Z[12]) );
  AOI22_X1 U100 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n63) );
  AOI22_X1 U101 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n62) );
  NAND2_X1 U102 ( .A1(n2), .A2(n3), .ZN(Z[9]) );
  AOI22_X1 U103 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n3) );
  AOI22_X1 U104 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n2) );
  NAND2_X1 U105 ( .A1(n14), .A2(n15), .ZN(Z[5]) );
  AOI22_X1 U106 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n15) );
  AOI22_X1 U107 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n14) );
  NAND2_X1 U108 ( .A1(n22), .A2(n23), .ZN(Z[30]) );
  AOI22_X1 U109 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n23) );
  AOI22_X1 U110 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n22) );
  NAND2_X1 U111 ( .A1(n30), .A2(n31), .ZN(Z[27]) );
  AOI22_X1 U112 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n31) );
  AOI22_X1 U113 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n30) );
endmodule


module mux41_NBIT32_4 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149;

  BUF_X1 U1 ( .A(n145), .Z(n72) );
  BUF_X1 U2 ( .A(n145), .Z(n73) );
  BUF_X1 U3 ( .A(n147), .Z(n78) );
  BUF_X1 U4 ( .A(n147), .Z(n79) );
  BUF_X1 U5 ( .A(n144), .Z(n1) );
  BUF_X1 U6 ( .A(n144), .Z(n70) );
  BUF_X1 U7 ( .A(n146), .Z(n75) );
  BUF_X1 U8 ( .A(n146), .Z(n76) );
  BUF_X1 U9 ( .A(n145), .Z(n74) );
  BUF_X1 U10 ( .A(n147), .Z(n80) );
  BUF_X1 U11 ( .A(n144), .Z(n71) );
  BUF_X1 U12 ( .A(n146), .Z(n77) );
  NOR2_X1 U13 ( .A1(n81), .A2(S[1]), .ZN(n145) );
  NOR2_X1 U14 ( .A1(S[0]), .A2(S[1]), .ZN(n144) );
  AND2_X1 U15 ( .A1(S[1]), .A2(S[0]), .ZN(n147) );
  AND2_X1 U16 ( .A1(S[1]), .A2(n81), .ZN(n146) );
  INV_X1 U17 ( .A(S[0]), .ZN(n81) );
  NAND2_X1 U18 ( .A1(n83), .A2(n82), .ZN(Z[0]) );
  AOI22_X1 U19 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n82) );
  AOI22_X1 U20 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n83) );
  NAND2_X1 U21 ( .A1(n105), .A2(n104), .ZN(Z[1]) );
  AOI22_X1 U22 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n104) );
  AOI22_X1 U23 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n105) );
  NAND2_X1 U24 ( .A1(n127), .A2(n126), .ZN(Z[2]) );
  AOI22_X1 U25 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n126) );
  AOI22_X1 U26 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n127) );
  NAND2_X1 U27 ( .A1(n139), .A2(n138), .ZN(Z[6]) );
  AOI22_X1 U28 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n138) );
  AOI22_X1 U29 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n139) );
  NAND2_X1 U30 ( .A1(n137), .A2(n136), .ZN(Z[5]) );
  AOI22_X1 U31 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n136) );
  AOI22_X1 U32 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n137) );
  NAND2_X1 U33 ( .A1(n135), .A2(n134), .ZN(Z[4]) );
  AOI22_X1 U34 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n134) );
  AOI22_X1 U35 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n135) );
  NAND2_X1 U36 ( .A1(n91), .A2(n90), .ZN(Z[13]) );
  AOI22_X1 U37 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n90) );
  AOI22_X1 U38 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n91) );
  NAND2_X1 U39 ( .A1(n93), .A2(n92), .ZN(Z[14]) );
  AOI22_X1 U40 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n92) );
  AOI22_X1 U41 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n93) );
  NAND2_X1 U42 ( .A1(n89), .A2(n88), .ZN(Z[12]) );
  AOI22_X1 U43 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n88) );
  AOI22_X1 U44 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n89) );
  NAND2_X1 U45 ( .A1(n97), .A2(n96), .ZN(Z[16]) );
  AOI22_X1 U46 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n96) );
  AOI22_X1 U47 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n97) );
  NAND2_X1 U48 ( .A1(n99), .A2(n98), .ZN(Z[17]) );
  AOI22_X1 U49 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n98) );
  AOI22_X1 U50 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n99) );
  NAND2_X1 U51 ( .A1(n143), .A2(n142), .ZN(Z[8]) );
  AOI22_X1 U52 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n142) );
  AOI22_X1 U53 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n143) );
  NAND2_X1 U54 ( .A1(n149), .A2(n148), .ZN(Z[9]) );
  AOI22_X1 U55 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n148) );
  AOI22_X1 U56 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n149) );
  NAND2_X1 U57 ( .A1(n85), .A2(n84), .ZN(Z[10]) );
  AOI22_X1 U58 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n84) );
  AOI22_X1 U59 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n85) );
  NAND2_X1 U60 ( .A1(n101), .A2(n100), .ZN(Z[18]) );
  AOI22_X1 U61 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n100) );
  AOI22_X1 U62 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n101) );
  NAND2_X1 U63 ( .A1(n109), .A2(n108), .ZN(Z[21]) );
  AOI22_X1 U64 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n108) );
  AOI22_X1 U65 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n109) );
  NAND2_X1 U66 ( .A1(n107), .A2(n106), .ZN(Z[20]) );
  AOI22_X1 U67 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n106) );
  AOI22_X1 U68 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n107) );
  NAND2_X1 U69 ( .A1(n129), .A2(n128), .ZN(Z[30]) );
  AOI22_X1 U70 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n128) );
  AOI22_X1 U71 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n129) );
  NAND2_X1 U72 ( .A1(n125), .A2(n124), .ZN(Z[29]) );
  AOI22_X1 U73 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n124) );
  AOI22_X1 U74 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n125) );
  NAND2_X1 U75 ( .A1(n115), .A2(n114), .ZN(Z[24]) );
  AOI22_X1 U76 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n114) );
  AOI22_X1 U77 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n115) );
  NAND2_X1 U78 ( .A1(n111), .A2(n110), .ZN(Z[22]) );
  AOI22_X1 U79 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n110) );
  AOI22_X1 U80 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n111) );
  NAND2_X1 U81 ( .A1(n117), .A2(n116), .ZN(Z[25]) );
  AOI22_X1 U82 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n116) );
  AOI22_X1 U83 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n117) );
  NAND2_X1 U84 ( .A1(n119), .A2(n118), .ZN(Z[26]) );
  AOI22_X1 U85 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n118) );
  AOI22_X1 U86 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n119) );
  NAND2_X1 U87 ( .A1(n123), .A2(n122), .ZN(Z[28]) );
  AOI22_X1 U88 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n122) );
  AOI22_X1 U89 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n123) );
  NAND2_X1 U90 ( .A1(n133), .A2(n132), .ZN(Z[3]) );
  AOI22_X1 U91 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n132) );
  AOI22_X1 U92 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n133) );
  NAND2_X1 U93 ( .A1(n141), .A2(n140), .ZN(Z[7]) );
  AOI22_X1 U94 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n140) );
  AOI22_X1 U95 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n141) );
  NAND2_X1 U96 ( .A1(n87), .A2(n86), .ZN(Z[11]) );
  AOI22_X1 U97 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n86) );
  AOI22_X1 U98 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n87) );
  NAND2_X1 U99 ( .A1(n95), .A2(n94), .ZN(Z[15]) );
  AOI22_X1 U100 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n94) );
  AOI22_X1 U101 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n95) );
  NAND2_X1 U102 ( .A1(n103), .A2(n102), .ZN(Z[19]) );
  AOI22_X1 U103 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n102) );
  AOI22_X1 U104 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n103) );
  NAND2_X1 U105 ( .A1(n113), .A2(n112), .ZN(Z[23]) );
  AOI22_X1 U106 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n112) );
  AOI22_X1 U107 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n113) );
  NAND2_X1 U108 ( .A1(n121), .A2(n120), .ZN(Z[27]) );
  AOI22_X1 U109 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n120) );
  AOI22_X1 U110 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n121) );
  NAND2_X1 U111 ( .A1(n131), .A2(n130), .ZN(Z[31]) );
  AOI22_X1 U112 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n130) );
  AOI22_X1 U113 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n131) );
endmodule


module mux21_NBIT32_3 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100;

  BUF_X1 U1 ( .A(n68), .Z(n1) );
  BUF_X1 U2 ( .A(n68), .Z(n2) );
  BUF_X1 U3 ( .A(n68), .Z(n3) );
  INV_X1 U4 ( .A(n69), .ZN(Z[0]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n1), .B1(B[0]), .B2(S), .ZN(n69) );
  INV_X1 U6 ( .A(n81), .ZN(Z[20]) );
  AOI22_X1 U7 ( .A1(A[20]), .A2(n2), .B1(B[20]), .B2(S), .ZN(n81) );
  INV_X1 U8 ( .A(n73), .ZN(Z[13]) );
  AOI22_X1 U9 ( .A1(A[13]), .A2(n1), .B1(B[13]), .B2(S), .ZN(n73) );
  INV_X1 U10 ( .A(n77), .ZN(Z[17]) );
  AOI22_X1 U11 ( .A1(A[17]), .A2(n1), .B1(B[17]), .B2(S), .ZN(n77) );
  INV_X1 U12 ( .A(n97), .ZN(Z[6]) );
  AOI22_X1 U13 ( .A1(A[6]), .A2(n3), .B1(B[6]), .B2(S), .ZN(n97) );
  INV_X1 U14 ( .A(n85), .ZN(Z[24]) );
  AOI22_X1 U15 ( .A1(A[24]), .A2(n2), .B1(B[24]), .B2(S), .ZN(n85) );
  INV_X1 U16 ( .A(n89), .ZN(Z[28]) );
  AOI22_X1 U17 ( .A1(A[28]), .A2(n2), .B1(B[28]), .B2(S), .ZN(n89) );
  INV_X1 U18 ( .A(n93), .ZN(Z[31]) );
  AOI22_X1 U19 ( .A1(A[31]), .A2(n3), .B1(B[31]), .B2(S), .ZN(n93) );
  INV_X1 U20 ( .A(n70), .ZN(Z[10]) );
  AOI22_X1 U21 ( .A1(A[10]), .A2(n1), .B1(B[10]), .B2(S), .ZN(n70) );
  INV_X1 U22 ( .A(n82), .ZN(Z[21]) );
  AOI22_X1 U23 ( .A1(A[21]), .A2(n2), .B1(B[21]), .B2(S), .ZN(n82) );
  INV_X1 U24 ( .A(n74), .ZN(Z[14]) );
  AOI22_X1 U25 ( .A1(A[14]), .A2(n1), .B1(B[14]), .B2(S), .ZN(n74) );
  INV_X1 U26 ( .A(n78), .ZN(Z[18]) );
  AOI22_X1 U27 ( .A1(A[18]), .A2(n1), .B1(B[18]), .B2(S), .ZN(n78) );
  INV_X1 U28 ( .A(n86), .ZN(Z[25]) );
  AOI22_X1 U29 ( .A1(A[25]), .A2(n2), .B1(B[25]), .B2(S), .ZN(n86) );
  INV_X1 U30 ( .A(n90), .ZN(Z[29]) );
  AOI22_X1 U31 ( .A1(A[29]), .A2(n2), .B1(B[29]), .B2(S), .ZN(n90) );
  INV_X1 U32 ( .A(n94), .ZN(Z[3]) );
  AOI22_X1 U33 ( .A1(A[3]), .A2(n3), .B1(B[3]), .B2(S), .ZN(n94) );
  INV_X1 U34 ( .A(n98), .ZN(Z[7]) );
  AOI22_X1 U35 ( .A1(A[7]), .A2(n3), .B1(B[7]), .B2(S), .ZN(n98) );
  INV_X1 U36 ( .A(n95), .ZN(Z[4]) );
  AOI22_X1 U37 ( .A1(A[4]), .A2(n3), .B1(B[4]), .B2(S), .ZN(n95) );
  INV_X1 U38 ( .A(n83), .ZN(Z[22]) );
  AOI22_X1 U39 ( .A1(A[22]), .A2(n2), .B1(B[22]), .B2(S), .ZN(n83) );
  INV_X1 U40 ( .A(n91), .ZN(Z[2]) );
  AOI22_X1 U41 ( .A1(A[2]), .A2(n2), .B1(B[2]), .B2(S), .ZN(n91) );
  INV_X1 U42 ( .A(n99), .ZN(Z[8]) );
  AOI22_X1 U43 ( .A1(A[8]), .A2(n3), .B1(B[8]), .B2(S), .ZN(n99) );
  INV_X1 U44 ( .A(n87), .ZN(Z[26]) );
  AOI22_X1 U45 ( .A1(A[26]), .A2(n2), .B1(B[26]), .B2(S), .ZN(n87) );
  INV_X1 U46 ( .A(n71), .ZN(Z[11]) );
  AOI22_X1 U47 ( .A1(A[11]), .A2(n1), .B1(B[11]), .B2(S), .ZN(n71) );
  INV_X1 U48 ( .A(n75), .ZN(Z[15]) );
  AOI22_X1 U49 ( .A1(A[15]), .A2(n1), .B1(B[15]), .B2(S), .ZN(n75) );
  INV_X1 U50 ( .A(n79), .ZN(Z[19]) );
  AOI22_X1 U51 ( .A1(A[19]), .A2(n1), .B1(B[19]), .B2(S), .ZN(n79) );
  INV_X1 U52 ( .A(n76), .ZN(Z[16]) );
  AOI22_X1 U53 ( .A1(A[16]), .A2(n1), .B1(B[16]), .B2(S), .ZN(n76) );
  INV_X1 U54 ( .A(n72), .ZN(Z[12]) );
  AOI22_X1 U55 ( .A1(A[12]), .A2(n1), .B1(B[12]), .B2(S), .ZN(n72) );
  INV_X1 U56 ( .A(n80), .ZN(Z[1]) );
  AOI22_X1 U57 ( .A1(A[1]), .A2(n1), .B1(B[1]), .B2(S), .ZN(n80) );
  INV_X1 U58 ( .A(n96), .ZN(Z[5]) );
  AOI22_X1 U59 ( .A1(A[5]), .A2(n3), .B1(B[5]), .B2(S), .ZN(n96) );
  INV_X1 U60 ( .A(n92), .ZN(Z[30]) );
  AOI22_X1 U61 ( .A1(A[30]), .A2(n2), .B1(B[30]), .B2(S), .ZN(n92) );
  INV_X1 U62 ( .A(n84), .ZN(Z[23]) );
  AOI22_X1 U63 ( .A1(A[23]), .A2(n2), .B1(B[23]), .B2(S), .ZN(n84) );
  INV_X1 U64 ( .A(n88), .ZN(Z[27]) );
  AOI22_X1 U65 ( .A1(A[27]), .A2(n2), .B1(B[27]), .B2(S), .ZN(n88) );
  INV_X1 U66 ( .A(n100), .ZN(Z[9]) );
  AOI22_X1 U67 ( .A1(A[9]), .A2(n3), .B1(S), .B2(B[9]), .ZN(n100) );
  INV_X1 U68 ( .A(S), .ZN(n68) );
endmodule


module mux41_NBIT32_3 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149;

  BUF_X1 U1 ( .A(n145), .Z(n72) );
  BUF_X1 U2 ( .A(n147), .Z(n78) );
  BUF_X1 U3 ( .A(n145), .Z(n73) );
  BUF_X1 U4 ( .A(n147), .Z(n79) );
  BUF_X1 U5 ( .A(n144), .Z(n1) );
  BUF_X1 U6 ( .A(n146), .Z(n75) );
  BUF_X1 U7 ( .A(n144), .Z(n70) );
  BUF_X1 U8 ( .A(n146), .Z(n76) );
  BUF_X1 U9 ( .A(n145), .Z(n74) );
  BUF_X1 U10 ( .A(n147), .Z(n80) );
  BUF_X1 U11 ( .A(n144), .Z(n71) );
  BUF_X1 U12 ( .A(n146), .Z(n77) );
  NAND2_X1 U13 ( .A1(n83), .A2(n82), .ZN(Z[0]) );
  AOI22_X1 U14 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n82) );
  AOI22_X1 U15 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n83) );
  NAND2_X1 U16 ( .A1(n105), .A2(n104), .ZN(Z[1]) );
  AOI22_X1 U17 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n104) );
  AOI22_X1 U18 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n105) );
  NAND2_X1 U19 ( .A1(n127), .A2(n126), .ZN(Z[2]) );
  AOI22_X1 U20 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n126) );
  AOI22_X1 U21 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n127) );
  NAND2_X1 U22 ( .A1(n139), .A2(n138), .ZN(Z[6]) );
  AOI22_X1 U23 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n138) );
  AOI22_X1 U24 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n139) );
  NAND2_X1 U25 ( .A1(n137), .A2(n136), .ZN(Z[5]) );
  AOI22_X1 U26 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n136) );
  AOI22_X1 U27 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n137) );
  NAND2_X1 U28 ( .A1(n135), .A2(n134), .ZN(Z[4]) );
  AOI22_X1 U29 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n134) );
  AOI22_X1 U30 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n135) );
  NAND2_X1 U31 ( .A1(n91), .A2(n90), .ZN(Z[13]) );
  AOI22_X1 U32 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n90) );
  AOI22_X1 U33 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n91) );
  NAND2_X1 U34 ( .A1(n93), .A2(n92), .ZN(Z[14]) );
  AOI22_X1 U35 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n92) );
  AOI22_X1 U36 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n93) );
  NAND2_X1 U37 ( .A1(n89), .A2(n88), .ZN(Z[12]) );
  AOI22_X1 U38 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n88) );
  AOI22_X1 U39 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n89) );
  NAND2_X1 U40 ( .A1(n97), .A2(n96), .ZN(Z[16]) );
  AOI22_X1 U41 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n96) );
  AOI22_X1 U42 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n97) );
  NAND2_X1 U43 ( .A1(n99), .A2(n98), .ZN(Z[17]) );
  AOI22_X1 U44 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n98) );
  AOI22_X1 U45 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n99) );
  NAND2_X1 U46 ( .A1(n143), .A2(n142), .ZN(Z[8]) );
  AOI22_X1 U47 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n142) );
  AOI22_X1 U48 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n143) );
  NAND2_X1 U49 ( .A1(n149), .A2(n148), .ZN(Z[9]) );
  AOI22_X1 U50 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n148) );
  AOI22_X1 U51 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n149) );
  NAND2_X1 U52 ( .A1(n85), .A2(n84), .ZN(Z[10]) );
  AOI22_X1 U53 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n84) );
  AOI22_X1 U54 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n85) );
  NAND2_X1 U55 ( .A1(n101), .A2(n100), .ZN(Z[18]) );
  AOI22_X1 U56 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n100) );
  AOI22_X1 U57 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n101) );
  NAND2_X1 U58 ( .A1(n109), .A2(n108), .ZN(Z[21]) );
  AOI22_X1 U59 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n108) );
  AOI22_X1 U60 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n109) );
  NAND2_X1 U61 ( .A1(n107), .A2(n106), .ZN(Z[20]) );
  AOI22_X1 U62 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n106) );
  AOI22_X1 U63 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n107) );
  NAND2_X1 U64 ( .A1(n129), .A2(n128), .ZN(Z[30]) );
  AOI22_X1 U65 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n128) );
  AOI22_X1 U66 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n129) );
  NAND2_X1 U67 ( .A1(n125), .A2(n124), .ZN(Z[29]) );
  AOI22_X1 U68 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n124) );
  AOI22_X1 U69 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n125) );
  NAND2_X1 U70 ( .A1(n115), .A2(n114), .ZN(Z[24]) );
  AOI22_X1 U71 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n114) );
  AOI22_X1 U72 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n115) );
  NAND2_X1 U73 ( .A1(n111), .A2(n110), .ZN(Z[22]) );
  AOI22_X1 U74 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n110) );
  AOI22_X1 U75 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n111) );
  NAND2_X1 U76 ( .A1(n117), .A2(n116), .ZN(Z[25]) );
  AOI22_X1 U77 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n116) );
  AOI22_X1 U78 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n117) );
  NAND2_X1 U79 ( .A1(n119), .A2(n118), .ZN(Z[26]) );
  AOI22_X1 U80 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n118) );
  AOI22_X1 U81 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n119) );
  NAND2_X1 U82 ( .A1(n123), .A2(n122), .ZN(Z[28]) );
  AOI22_X1 U83 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n122) );
  AOI22_X1 U84 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n123) );
  NAND2_X1 U85 ( .A1(n133), .A2(n132), .ZN(Z[3]) );
  AOI22_X1 U86 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n132) );
  AOI22_X1 U87 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n133) );
  NAND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(Z[7]) );
  AOI22_X1 U89 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n140) );
  AOI22_X1 U90 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n141) );
  NAND2_X1 U91 ( .A1(n87), .A2(n86), .ZN(Z[11]) );
  AOI22_X1 U92 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n86) );
  AOI22_X1 U93 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n87) );
  NAND2_X1 U94 ( .A1(n95), .A2(n94), .ZN(Z[15]) );
  AOI22_X1 U95 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n94) );
  AOI22_X1 U96 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n95) );
  NAND2_X1 U97 ( .A1(n103), .A2(n102), .ZN(Z[19]) );
  AOI22_X1 U98 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n102) );
  AOI22_X1 U99 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n103) );
  NAND2_X1 U100 ( .A1(n113), .A2(n112), .ZN(Z[23]) );
  AOI22_X1 U101 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n112) );
  AOI22_X1 U102 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n113) );
  NAND2_X1 U103 ( .A1(n121), .A2(n120), .ZN(Z[27]) );
  AOI22_X1 U104 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n120) );
  AOI22_X1 U105 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n121) );
  NAND2_X1 U106 ( .A1(n131), .A2(n130), .ZN(Z[31]) );
  AOI22_X1 U107 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n130) );
  AOI22_X1 U108 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n131) );
  NOR2_X1 U109 ( .A1(n81), .A2(S[1]), .ZN(n145) );
  NOR2_X1 U110 ( .A1(S[0]), .A2(S[1]), .ZN(n144) );
  AND2_X1 U111 ( .A1(S[1]), .A2(S[0]), .ZN(n147) );
  AND2_X1 U112 ( .A1(S[1]), .A2(n81), .ZN(n146) );
  INV_X1 U113 ( .A(S[0]), .ZN(n81) );
endmodule


module comparator_NBIT32_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202;

  INV_X1 U1 ( .A(n142), .ZN(n10) );
  INV_X1 U2 ( .A(n130), .ZN(n14) );
  INV_X1 U3 ( .A(n118), .ZN(n18) );
  INV_X1 U4 ( .A(n106), .ZN(n22) );
  INV_X1 U5 ( .A(n94), .ZN(n26) );
  INV_X1 U6 ( .A(n82), .ZN(n30) );
  INV_X1 U7 ( .A(GE), .ZN(LT) );
  INV_X1 U8 ( .A(NE), .ZN(EQ) );
  INV_X1 U9 ( .A(n139), .ZN(n12) );
  INV_X1 U10 ( .A(n127), .ZN(n16) );
  INV_X1 U11 ( .A(n115), .ZN(n20) );
  INV_X1 U12 ( .A(n103), .ZN(n24) );
  INV_X1 U13 ( .A(n91), .ZN(n28) );
  INV_X1 U14 ( .A(n79), .ZN(n32) );
  INV_X1 U15 ( .A(GT), .ZN(LE) );
  INV_X1 U16 ( .A(n144), .ZN(n9) );
  INV_X1 U17 ( .A(n132), .ZN(n13) );
  INV_X1 U18 ( .A(n120), .ZN(n17) );
  INV_X1 U19 ( .A(n108), .ZN(n21) );
  INV_X1 U20 ( .A(n96), .ZN(n25) );
  INV_X1 U21 ( .A(n84), .ZN(n29) );
  INV_X1 U22 ( .A(n154), .ZN(n7) );
  INV_X1 U23 ( .A(n141), .ZN(n11) );
  INV_X1 U24 ( .A(n129), .ZN(n15) );
  INV_X1 U25 ( .A(n117), .ZN(n19) );
  INV_X1 U26 ( .A(n105), .ZN(n23) );
  INV_X1 U27 ( .A(n93), .ZN(n27) );
  INV_X1 U28 ( .A(n81), .ZN(n31) );
  INV_X1 U29 ( .A(n68), .ZN(n3) );
  INV_X1 U30 ( .A(A[30]), .ZN(n65) );
  INV_X1 U31 ( .A(n72), .ZN(n33) );
  INV_X1 U32 ( .A(n151), .ZN(n8) );
  INV_X1 U33 ( .A(n202), .ZN(n5) );
  INV_X1 U34 ( .A(B[30]), .ZN(n34) );
  INV_X1 U35 ( .A(A[0]), .ZN(n36) );
  INV_X1 U36 ( .A(A[3]), .ZN(n38) );
  INV_X1 U37 ( .A(A[5]), .ZN(n40) );
  INV_X1 U38 ( .A(A[7]), .ZN(n42) );
  INV_X1 U39 ( .A(A[9]), .ZN(n44) );
  INV_X1 U40 ( .A(A[11]), .ZN(n46) );
  INV_X1 U41 ( .A(A[13]), .ZN(n48) );
  INV_X1 U42 ( .A(A[15]), .ZN(n50) );
  INV_X1 U43 ( .A(A[17]), .ZN(n52) );
  INV_X1 U44 ( .A(A[19]), .ZN(n54) );
  INV_X1 U45 ( .A(A[21]), .ZN(n56) );
  INV_X1 U46 ( .A(A[23]), .ZN(n58) );
  INV_X1 U47 ( .A(A[25]), .ZN(n60) );
  INV_X1 U48 ( .A(A[27]), .ZN(n62) );
  INV_X1 U49 ( .A(A[29]), .ZN(n64) );
  INV_X1 U50 ( .A(B[31]), .ZN(n35) );
  INV_X1 U51 ( .A(B[1]), .ZN(n6) );
  INV_X1 U52 ( .A(A[4]), .ZN(n39) );
  INV_X1 U53 ( .A(A[8]), .ZN(n43) );
  INV_X1 U54 ( .A(A[12]), .ZN(n47) );
  INV_X1 U55 ( .A(A[16]), .ZN(n51) );
  INV_X1 U56 ( .A(A[20]), .ZN(n55) );
  INV_X1 U57 ( .A(A[24]), .ZN(n59) );
  INV_X1 U58 ( .A(A[28]), .ZN(n63) );
  INV_X1 U59 ( .A(A[2]), .ZN(n37) );
  INV_X1 U60 ( .A(A[6]), .ZN(n41) );
  INV_X1 U61 ( .A(A[10]), .ZN(n45) );
  INV_X1 U62 ( .A(A[14]), .ZN(n49) );
  INV_X1 U63 ( .A(A[18]), .ZN(n53) );
  INV_X1 U64 ( .A(A[22]), .ZN(n57) );
  INV_X1 U65 ( .A(A[26]), .ZN(n61) );
  NAND2_X1 U66 ( .A1(LE), .A2(GE), .ZN(NE) );
  AOI21_X1 U67 ( .B1(n66), .B2(n3), .A(n67), .ZN(GE) );
  AOI22_X1 U68 ( .A1(B[30]), .A2(n65), .B1(n69), .B2(n70), .ZN(n68) );
  AOI21_X1 U69 ( .B1(n71), .B2(n72), .A(n73), .ZN(n69) );
  AOI21_X1 U70 ( .B1(n74), .B2(n75), .A(n76), .ZN(n71) );
  AOI21_X1 U71 ( .B1(n77), .B2(n78), .A(n79), .ZN(n74) );
  AOI21_X1 U72 ( .B1(n80), .B2(n30), .A(n31), .ZN(n77) );
  AOI21_X1 U73 ( .B1(n83), .B2(n84), .A(n85), .ZN(n80) );
  AOI21_X1 U74 ( .B1(n86), .B2(n87), .A(n88), .ZN(n83) );
  AOI21_X1 U75 ( .B1(n89), .B2(n90), .A(n91), .ZN(n86) );
  AOI21_X1 U76 ( .B1(n92), .B2(n26), .A(n27), .ZN(n89) );
  AOI21_X1 U77 ( .B1(n95), .B2(n96), .A(n97), .ZN(n92) );
  AOI21_X1 U78 ( .B1(n98), .B2(n99), .A(n100), .ZN(n95) );
  AOI21_X1 U79 ( .B1(n101), .B2(n102), .A(n103), .ZN(n98) );
  AOI21_X1 U80 ( .B1(n104), .B2(n22), .A(n23), .ZN(n101) );
  AOI21_X1 U81 ( .B1(n107), .B2(n108), .A(n109), .ZN(n104) );
  AOI21_X1 U82 ( .B1(n110), .B2(n111), .A(n112), .ZN(n107) );
  AOI21_X1 U83 ( .B1(n113), .B2(n114), .A(n115), .ZN(n110) );
  AOI21_X1 U84 ( .B1(n116), .B2(n18), .A(n19), .ZN(n113) );
  AOI21_X1 U85 ( .B1(n119), .B2(n120), .A(n121), .ZN(n116) );
  AOI21_X1 U86 ( .B1(n122), .B2(n123), .A(n124), .ZN(n119) );
  AOI21_X1 U87 ( .B1(n125), .B2(n126), .A(n127), .ZN(n122) );
  AOI21_X1 U88 ( .B1(n128), .B2(n14), .A(n15), .ZN(n125) );
  AOI21_X1 U89 ( .B1(n131), .B2(n132), .A(n133), .ZN(n128) );
  AOI21_X1 U90 ( .B1(n134), .B2(n135), .A(n136), .ZN(n131) );
  AOI21_X1 U91 ( .B1(n137), .B2(n138), .A(n139), .ZN(n134) );
  AOI21_X1 U92 ( .B1(n140), .B2(n10), .A(n11), .ZN(n137) );
  AOI21_X1 U93 ( .B1(n143), .B2(n144), .A(n145), .ZN(n140) );
  AOI21_X1 U94 ( .B1(n146), .B2(n147), .A(n148), .ZN(n143) );
  AOI21_X1 U95 ( .B1(n149), .B2(n150), .A(n151), .ZN(n146) );
  AOI21_X1 U96 ( .B1(n152), .B2(n153), .A(n7), .ZN(n149) );
  AOI22_X1 U97 ( .A1(n155), .A2(n6), .B1(A[1]), .B2(n156), .ZN(n152) );
  OR2_X1 U98 ( .A1(n156), .A2(A[1]), .ZN(n155) );
  NAND2_X1 U99 ( .A1(B[0]), .A2(n36), .ZN(n156) );
  OAI21_X1 U100 ( .B1(n67), .B2(n157), .A(n66), .ZN(GT) );
  NAND2_X1 U101 ( .A1(A[31]), .A2(n35), .ZN(n66) );
  AOI22_X1 U102 ( .A1(A[30]), .A2(n34), .B1(n158), .B2(n70), .ZN(n157) );
  XOR2_X1 U103 ( .A(A[30]), .B(n34), .Z(n70) );
  AOI21_X1 U104 ( .B1(n159), .B2(n160), .A(n33), .ZN(n158) );
  NAND2_X1 U105 ( .A1(B[29]), .A2(n64), .ZN(n72) );
  OAI211_X1 U106 ( .C1(n161), .C2(n162), .A(n78), .B(n75), .ZN(n160) );
  NOR2_X1 U107 ( .A1(n163), .A2(n76), .ZN(n75) );
  AND2_X1 U108 ( .A1(B[28]), .A2(n63), .ZN(n76) );
  NAND2_X1 U109 ( .A1(B[27]), .A2(n62), .ZN(n78) );
  NAND2_X1 U110 ( .A1(n32), .A2(n164), .ZN(n162) );
  NOR2_X1 U111 ( .A1(n62), .A2(B[27]), .ZN(n79) );
  AOI211_X1 U112 ( .C1(n165), .C2(n166), .A(n82), .B(n29), .ZN(n161) );
  NAND2_X1 U113 ( .A1(B[25]), .A2(n60), .ZN(n84) );
  NAND2_X1 U114 ( .A1(n164), .A2(n81), .ZN(n82) );
  NAND2_X1 U115 ( .A1(B[26]), .A2(n61), .ZN(n81) );
  OR2_X1 U116 ( .A1(n61), .A2(B[26]), .ZN(n164) );
  OAI211_X1 U117 ( .C1(n167), .C2(n168), .A(n90), .B(n87), .ZN(n166) );
  NOR2_X1 U118 ( .A1(n169), .A2(n88), .ZN(n87) );
  AND2_X1 U119 ( .A1(B[24]), .A2(n59), .ZN(n88) );
  NAND2_X1 U120 ( .A1(B[23]), .A2(n58), .ZN(n90) );
  NAND2_X1 U121 ( .A1(n28), .A2(n170), .ZN(n168) );
  NOR2_X1 U122 ( .A1(n58), .A2(B[23]), .ZN(n91) );
  AOI211_X1 U123 ( .C1(n171), .C2(n172), .A(n94), .B(n25), .ZN(n167) );
  NAND2_X1 U124 ( .A1(B[21]), .A2(n56), .ZN(n96) );
  NAND2_X1 U125 ( .A1(n170), .A2(n93), .ZN(n94) );
  NAND2_X1 U126 ( .A1(B[22]), .A2(n57), .ZN(n93) );
  OR2_X1 U127 ( .A1(n57), .A2(B[22]), .ZN(n170) );
  OAI211_X1 U128 ( .C1(n173), .C2(n174), .A(n102), .B(n99), .ZN(n172) );
  NOR2_X1 U129 ( .A1(n175), .A2(n100), .ZN(n99) );
  AND2_X1 U130 ( .A1(B[20]), .A2(n55), .ZN(n100) );
  NAND2_X1 U131 ( .A1(B[19]), .A2(n54), .ZN(n102) );
  NAND2_X1 U132 ( .A1(n24), .A2(n176), .ZN(n174) );
  NOR2_X1 U133 ( .A1(n54), .A2(B[19]), .ZN(n103) );
  AOI211_X1 U134 ( .C1(n177), .C2(n178), .A(n106), .B(n21), .ZN(n173) );
  NAND2_X1 U135 ( .A1(B[17]), .A2(n52), .ZN(n108) );
  NAND2_X1 U136 ( .A1(n176), .A2(n105), .ZN(n106) );
  NAND2_X1 U137 ( .A1(B[18]), .A2(n53), .ZN(n105) );
  OR2_X1 U138 ( .A1(n53), .A2(B[18]), .ZN(n176) );
  OAI211_X1 U139 ( .C1(n179), .C2(n180), .A(n114), .B(n111), .ZN(n178) );
  NOR2_X1 U140 ( .A1(n181), .A2(n112), .ZN(n111) );
  AND2_X1 U141 ( .A1(B[16]), .A2(n51), .ZN(n112) );
  NAND2_X1 U142 ( .A1(B[15]), .A2(n50), .ZN(n114) );
  NAND2_X1 U143 ( .A1(n20), .A2(n182), .ZN(n180) );
  NOR2_X1 U144 ( .A1(n50), .A2(B[15]), .ZN(n115) );
  AOI211_X1 U145 ( .C1(n183), .C2(n184), .A(n118), .B(n17), .ZN(n179) );
  NAND2_X1 U146 ( .A1(B[13]), .A2(n48), .ZN(n120) );
  NAND2_X1 U147 ( .A1(n182), .A2(n117), .ZN(n118) );
  NAND2_X1 U148 ( .A1(B[14]), .A2(n49), .ZN(n117) );
  OR2_X1 U149 ( .A1(n49), .A2(B[14]), .ZN(n182) );
  OAI211_X1 U150 ( .C1(n185), .C2(n186), .A(n126), .B(n123), .ZN(n184) );
  NOR2_X1 U151 ( .A1(n187), .A2(n124), .ZN(n123) );
  AND2_X1 U152 ( .A1(B[12]), .A2(n47), .ZN(n124) );
  NAND2_X1 U153 ( .A1(B[11]), .A2(n46), .ZN(n126) );
  NAND2_X1 U154 ( .A1(n16), .A2(n188), .ZN(n186) );
  NOR2_X1 U155 ( .A1(n46), .A2(B[11]), .ZN(n127) );
  AOI211_X1 U156 ( .C1(n189), .C2(n190), .A(n130), .B(n13), .ZN(n185) );
  NAND2_X1 U157 ( .A1(B[9]), .A2(n44), .ZN(n132) );
  NAND2_X1 U158 ( .A1(n188), .A2(n129), .ZN(n130) );
  NAND2_X1 U159 ( .A1(B[10]), .A2(n45), .ZN(n129) );
  OR2_X1 U160 ( .A1(n45), .A2(B[10]), .ZN(n188) );
  OAI211_X1 U161 ( .C1(n191), .C2(n192), .A(n138), .B(n135), .ZN(n190) );
  NOR2_X1 U162 ( .A1(n193), .A2(n136), .ZN(n135) );
  AND2_X1 U163 ( .A1(B[8]), .A2(n43), .ZN(n136) );
  NAND2_X1 U164 ( .A1(B[7]), .A2(n42), .ZN(n138) );
  NAND2_X1 U165 ( .A1(n12), .A2(n194), .ZN(n192) );
  NOR2_X1 U166 ( .A1(n42), .A2(B[7]), .ZN(n139) );
  AOI211_X1 U167 ( .C1(n195), .C2(n196), .A(n142), .B(n9), .ZN(n191) );
  NAND2_X1 U168 ( .A1(B[5]), .A2(n40), .ZN(n144) );
  NAND2_X1 U169 ( .A1(n194), .A2(n141), .ZN(n142) );
  NAND2_X1 U170 ( .A1(B[6]), .A2(n41), .ZN(n141) );
  OR2_X1 U171 ( .A1(n41), .A2(B[6]), .ZN(n194) );
  NAND3_X1 U172 ( .A1(n197), .A2(n150), .A3(n147), .ZN(n196) );
  NOR2_X1 U173 ( .A1(n198), .A2(n148), .ZN(n147) );
  AND2_X1 U174 ( .A1(B[4]), .A2(n39), .ZN(n148) );
  NAND2_X1 U175 ( .A1(B[3]), .A2(n38), .ZN(n150) );
  NAND3_X1 U176 ( .A1(n8), .A2(n199), .A3(n200), .ZN(n197) );
  OAI211_X1 U177 ( .C1(A[1]), .C2(n201), .A(n5), .B(n153), .ZN(n200) );
  AND2_X1 U178 ( .A1(n199), .A2(n154), .ZN(n153) );
  NAND2_X1 U179 ( .A1(B[2]), .A2(n37), .ZN(n154) );
  AOI21_X1 U180 ( .B1(A[1]), .B2(n201), .A(n6), .ZN(n202) );
  NOR2_X1 U181 ( .A1(n36), .A2(B[0]), .ZN(n201) );
  OR2_X1 U182 ( .A1(n37), .A2(B[2]), .ZN(n199) );
  NOR2_X1 U183 ( .A1(n38), .A2(B[3]), .ZN(n151) );
  NOR2_X1 U184 ( .A1(n198), .A2(n145), .ZN(n195) );
  NOR2_X1 U185 ( .A1(n40), .A2(B[5]), .ZN(n145) );
  NOR2_X1 U186 ( .A1(n39), .A2(B[4]), .ZN(n198) );
  NOR2_X1 U187 ( .A1(n193), .A2(n133), .ZN(n189) );
  NOR2_X1 U188 ( .A1(n44), .A2(B[9]), .ZN(n133) );
  NOR2_X1 U189 ( .A1(n43), .A2(B[8]), .ZN(n193) );
  NOR2_X1 U190 ( .A1(n187), .A2(n121), .ZN(n183) );
  NOR2_X1 U191 ( .A1(n48), .A2(B[13]), .ZN(n121) );
  NOR2_X1 U192 ( .A1(n47), .A2(B[12]), .ZN(n187) );
  NOR2_X1 U193 ( .A1(n181), .A2(n109), .ZN(n177) );
  NOR2_X1 U194 ( .A1(n52), .A2(B[17]), .ZN(n109) );
  NOR2_X1 U195 ( .A1(n51), .A2(B[16]), .ZN(n181) );
  NOR2_X1 U196 ( .A1(n175), .A2(n97), .ZN(n171) );
  NOR2_X1 U197 ( .A1(n56), .A2(B[21]), .ZN(n97) );
  NOR2_X1 U198 ( .A1(n55), .A2(B[20]), .ZN(n175) );
  NOR2_X1 U199 ( .A1(n169), .A2(n85), .ZN(n165) );
  NOR2_X1 U200 ( .A1(n60), .A2(B[25]), .ZN(n85) );
  NOR2_X1 U201 ( .A1(n59), .A2(B[24]), .ZN(n169) );
  NOR2_X1 U202 ( .A1(n163), .A2(n73), .ZN(n159) );
  NOR2_X1 U203 ( .A1(n64), .A2(B[29]), .ZN(n73) );
  NOR2_X1 U204 ( .A1(n63), .A2(B[28]), .ZN(n163) );
  NOR2_X1 U205 ( .A1(n35), .A2(A[31]), .ZN(n67) );
endmodule


module comparator_NBIT32 ( A, B, .OPSel({\OPSel[2] , \OPSel[1] , \OPSel[0] }), 
        RES );
  input [31:0] A;
  input [31:0] B;
  output [31:0] RES;
  input \OPSel[2] , \OPSel[1] , \OPSel[0] ;
  wire   N26, N27, N28, N29, N30, N31, n15, n16, n17, n18, n19, n20, n2, n3,
         n4;
  wire   [2:0] OPSel;
  assign RES[1] = 1'b0;
  assign RES[2] = 1'b0;
  assign RES[3] = 1'b0;
  assign RES[4] = 1'b0;
  assign RES[5] = 1'b0;
  assign RES[6] = 1'b0;
  assign RES[7] = 1'b0;
  assign RES[8] = 1'b0;
  assign RES[9] = 1'b0;
  assign RES[10] = 1'b0;
  assign RES[11] = 1'b0;
  assign RES[12] = 1'b0;
  assign RES[13] = 1'b0;
  assign RES[14] = 1'b0;
  assign RES[15] = 1'b0;
  assign RES[16] = 1'b0;
  assign RES[17] = 1'b0;
  assign RES[18] = 1'b0;
  assign RES[19] = 1'b0;
  assign RES[20] = 1'b0;
  assign RES[21] = 1'b0;
  assign RES[22] = 1'b0;
  assign RES[23] = 1'b0;
  assign RES[24] = 1'b0;
  assign RES[25] = 1'b0;
  assign RES[26] = 1'b0;
  assign RES[27] = 1'b0;
  assign RES[28] = 1'b0;
  assign RES[29] = 1'b0;
  assign RES[30] = 1'b0;
  assign RES[31] = 1'b0;

  comparator_NBIT32_DW01_cmp6_0 r57 ( .A(A), .B(B), .TC(1'b0), .LT(N30), .GT(
        N28), .EQ(N26), .LE(N31), .GE(N29), .NE(N27) );
  INV_X1 U3 ( .A(n15), .ZN(RES[0]) );
  AOI21_X1 U4 ( .B1(n16), .B2(n4), .A(n17), .ZN(n15) );
  NOR3_X1 U5 ( .A1(n4), .A2(OPSel[1]), .A3(n18), .ZN(n17) );
  OAI22_X1 U6 ( .A1(n19), .A2(n3), .B1(OPSel[1]), .B2(n20), .ZN(n16) );
  INV_X1 U7 ( .A(OPSel[1]), .ZN(n3) );
  AOI22_X1 U8 ( .A1(N28), .A2(n2), .B1(N29), .B2(OPSel[0]), .ZN(n19) );
  INV_X1 U9 ( .A(OPSel[0]), .ZN(n2) );
  AOI22_X1 U10 ( .A1(N30), .A2(n2), .B1(OPSel[0]), .B2(N31), .ZN(n18) );
  AOI22_X1 U11 ( .A1(N26), .A2(n2), .B1(N27), .B2(OPSel[0]), .ZN(n20) );
  INV_X1 U12 ( .A(OPSel[2]), .ZN(n4) );
endmodule


module shifter_NBIT32 ( A, B, LOGIC_ARITH, LEFT_RIGHT, RES );
  input [31:0] A;
  input [31:0] B;
  output [31:0] RES;
  input LOGIC_ARITH, LEFT_RIGHT;
  wire   n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n266, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648;

  AOI21_X2 U264 ( .B1(A[31]), .B2(B[18]), .A(n483), .ZN(n282) );
  OAI21_X2 U267 ( .B1(n612), .B2(n628), .A(n486), .ZN(n285) );
  AOI21_X2 U269 ( .B1(A[31]), .B2(n38), .A(n487), .ZN(n288) );
  AOI221_X2 U388 ( .B1(n30), .B2(A[18]), .C1(n21), .C2(A[17]), .A(n568), .ZN(
        n196) );
  NOR2_X2 U428 ( .A1(n638), .A2(n38), .ZN(n165) );
  NOR2_X2 U461 ( .A1(n642), .A2(n38), .ZN(n199) );
  NAND3_X1 U637 ( .A1(n227), .A2(n646), .A3(n228), .ZN(n226) );
  NAND3_X1 U638 ( .A1(n227), .A2(n646), .A3(B[4]), .ZN(n428) );
  NAND3_X1 U639 ( .A1(n445), .A2(n199), .A3(LEFT_RIGHT), .ZN(n240) );
  NAND3_X1 U641 ( .A1(n489), .A2(n628), .A3(n579), .ZN(n255) );
  NAND3_X1 U642 ( .A1(n7), .A2(n199), .A3(n445), .ZN(n138) );
  NOR4_X1 U2 ( .A1(B[20]), .A2(B[21]), .A3(B[19]), .A4(n594), .ZN(n484) );
  NOR2_X2 U3 ( .A1(n639), .A2(B[3]), .ZN(n262) );
  AOI221_X1 U4 ( .B1(n29), .B2(A[6]), .C1(n19), .C2(A[7]), .A(n525), .ZN(n363)
         );
  AOI221_X1 U5 ( .B1(n30), .B2(A[7]), .C1(n20), .C2(A[8]), .A(n570), .ZN(n405)
         );
  AOI221_X1 U6 ( .B1(n29), .B2(A[8]), .C1(n21), .C2(A[9]), .A(n552), .ZN(n387)
         );
  OAI21_X2 U7 ( .B1(n266), .B2(n632), .A(n481), .ZN(n279) );
  AOI222_X1 U8 ( .A1(n11), .A2(A[1]), .B1(A[0]), .B2(n18), .C1(n7), .C2(A[2]), 
        .ZN(n293) );
  INV_X1 U9 ( .A(n167), .ZN(n635) );
  NOR2_X1 U10 ( .A1(n636), .A2(B[4]), .ZN(n167) );
  INV_X1 U11 ( .A(n169), .ZN(n644) );
  INV_X1 U12 ( .A(n165), .ZN(n637) );
  INV_X1 U13 ( .A(n199), .ZN(n641) );
  INV_X1 U14 ( .A(n28), .ZN(n26) );
  INV_X1 U15 ( .A(n31), .ZN(n24) );
  INV_X1 U16 ( .A(n31), .ZN(n25) );
  INV_X1 U17 ( .A(n21), .ZN(n14) );
  INV_X1 U18 ( .A(n19), .ZN(n16) );
  INV_X1 U19 ( .A(n19), .ZN(n15) );
  INV_X1 U20 ( .A(n505), .ZN(n643) );
  INV_X1 U21 ( .A(n29), .ZN(n27) );
  INV_X1 U22 ( .A(n493), .ZN(n640) );
  NOR2_X1 U23 ( .A1(n645), .A2(n38), .ZN(n169) );
  NAND2_X1 U24 ( .A1(n488), .A2(n454), .ZN(n161) );
  INV_X1 U25 ( .A(n41), .ZN(n38) );
  OAI222_X1 U26 ( .A1(n637), .A2(n70), .B1(n635), .B2(n92), .C1(n644), .C2(n80), .ZN(n224) );
  OAI222_X1 U27 ( .A1(n637), .A2(n67), .B1(n635), .B2(n96), .C1(n644), .C2(n83), .ZN(n212) );
  NOR2_X1 U28 ( .A1(n40), .A2(n642), .ZN(n493) );
  OAI22_X1 U29 ( .A1(n115), .A2(n642), .B1(n126), .B2(n638), .ZN(n383) );
  INV_X1 U30 ( .A(n454), .ZN(n636) );
  AOI21_X1 U31 ( .B1(n134), .B2(n2), .A(n519), .ZN(n286) );
  AOI21_X1 U32 ( .B1(n129), .B2(n3), .A(n519), .ZN(n312) );
  BUF_X1 U33 ( .A(n138), .Z(n33) );
  BUF_X1 U34 ( .A(n138), .Z(n32) );
  NOR2_X1 U35 ( .A1(n383), .A2(n359), .ZN(n197) );
  NOR2_X1 U36 ( .A1(n118), .A2(n359), .ZN(n181) );
  BUF_X1 U37 ( .A(n138), .Z(n34) );
  NAND2_X1 U38 ( .A1(n488), .A2(n5), .ZN(n505) );
  INV_X1 U39 ( .A(n182), .ZN(n118) );
  INV_X1 U40 ( .A(n172), .ZN(n54) );
  INV_X1 U41 ( .A(n139), .ZN(n58) );
  INV_X1 U42 ( .A(n348), .ZN(n52) );
  INV_X1 U43 ( .A(n337), .ZN(n44) );
  INV_X1 U44 ( .A(n480), .ZN(n88) );
  INV_X1 U45 ( .A(n314), .ZN(n56) );
  INV_X1 U46 ( .A(n290), .ZN(n50) );
  INV_X1 U47 ( .A(n271), .ZN(n46) );
  INV_X1 U48 ( .A(n257), .ZN(n101) );
  INV_X1 U49 ( .A(n440), .ZN(n93) );
  INV_X1 U50 ( .A(n302), .ZN(n97) );
  NOR2_X1 U51 ( .A1(n612), .A2(n148), .ZN(n150) );
  NOR2_X1 U52 ( .A1(n639), .A2(n646), .ZN(n454) );
  NAND2_X1 U53 ( .A1(n484), .A2(n630), .ZN(n281) );
  AOI222_X1 U54 ( .A1(n370), .A2(n262), .B1(n320), .B2(n260), .C1(n185), .C2(
        n3), .ZN(n238) );
  INV_X1 U55 ( .A(n356), .ZN(n642) );
  AOI222_X1 U56 ( .A1(n168), .A2(n262), .B1(n355), .B2(n260), .C1(n170), .C2(
        n3), .ZN(n471) );
  AOI222_X1 U57 ( .A1(n402), .A2(n262), .B1(n403), .B2(n260), .C1(n464), .C2(
        n2), .ZN(n461) );
  NAND2_X1 U58 ( .A1(n488), .A2(n262), .ZN(n157) );
  NAND2_X1 U59 ( .A1(n488), .A2(n260), .ZN(n158) );
  OAI222_X1 U60 ( .A1(n374), .A2(n638), .B1(n645), .B2(n375), .C1(n376), .C2(
        n642), .ZN(n172) );
  OAI222_X1 U61 ( .A1(n131), .A2(n638), .B1(n362), .B2(n645), .C1(n363), .C2(
        n642), .ZN(n139) );
  OAI222_X1 U62 ( .A1(n613), .A2(n638), .B1(n293), .B2(n645), .C1(n405), .C2(
        n642), .ZN(n348) );
  OAI222_X1 U63 ( .A1(n615), .A2(n638), .B1(n45), .B2(n645), .C1(n387), .C2(
        n642), .ZN(n337) );
  AOI221_X1 U64 ( .B1(n129), .B2(n262), .C1(n355), .C2(n2), .A(n359), .ZN(n159) );
  AOI221_X1 U65 ( .B1(n134), .B2(n262), .C1(n403), .C2(n3), .A(n359), .ZN(n347) );
  OAI221_X1 U66 ( .B1(n105), .B2(n638), .C1(n89), .C2(n642), .A(n607), .ZN(
        n480) );
  AOI22_X1 U67 ( .A1(n454), .A2(n320), .B1(n260), .B2(n370), .ZN(n607) );
  AOI222_X1 U68 ( .A1(n169), .A2(n185), .B1(n493), .B2(n320), .C1(n167), .C2(
        n370), .ZN(n550) );
  AOI222_X1 U69 ( .A1(n165), .A2(n166), .B1(n167), .B2(n168), .C1(n169), .C2(
        n170), .ZN(n164) );
  AOI222_X1 U70 ( .A1(n165), .A2(n516), .B1(n167), .B2(n402), .C1(n169), .C2(
        n464), .ZN(n581) );
  AOI222_X1 U71 ( .A1(n165), .A2(n184), .B1(n167), .B2(n185), .C1(n169), .C2(
        n186), .ZN(n183) );
  AOI222_X1 U72 ( .A1(n165), .A2(n178), .B1(n167), .B2(n186), .C1(n169), .C2(
        n184), .ZN(n239) );
  AOI222_X1 U73 ( .A1(n169), .A2(n168), .B1(n493), .B2(n128), .C1(n167), .C2(
        n355), .ZN(n534) );
  AOI222_X1 U74 ( .A1(n169), .A2(n402), .B1(n493), .B2(n133), .C1(n167), .C2(
        n403), .ZN(n520) );
  AOI222_X1 U75 ( .A1(n169), .A2(n453), .B1(n493), .B2(n382), .C1(n167), .C2(
        n506), .ZN(n507) );
  OAI222_X1 U76 ( .A1(n637), .A2(n74), .B1(n635), .B2(n100), .C1(n644), .C2(
        n196), .ZN(n200) );
  INV_X1 U77 ( .A(n260), .ZN(n645) );
  NOR2_X1 U78 ( .A1(n647), .A2(B[4]), .ZN(n488) );
  INV_X1 U79 ( .A(n262), .ZN(n638) );
  OAI222_X1 U80 ( .A1(n132), .A2(n14), .B1(n27), .B2(n614), .C1(n1), .C2(n102), 
        .ZN(n602) );
  OAI221_X1 U81 ( .B1(n363), .B2(n638), .C1(n61), .C2(n642), .A(n522), .ZN(
        n314) );
  AOI22_X1 U82 ( .A1(n454), .A2(n57), .B1(n260), .B2(n420), .ZN(n522) );
  OAI221_X1 U83 ( .B1(n405), .B2(n638), .C1(n72), .C2(n642), .A(n509), .ZN(
        n290) );
  AOI22_X1 U84 ( .A1(n454), .A2(n51), .B1(n260), .B2(n407), .ZN(n509) );
  OAI221_X1 U85 ( .B1(n387), .B2(n638), .C1(n75), .C2(n642), .A(n496), .ZN(
        n271) );
  AOI22_X1 U86 ( .A1(n454), .A2(n390), .B1(n260), .B2(n389), .ZN(n496) );
  INV_X1 U87 ( .A(n228), .ZN(n625) );
  OAI21_X1 U88 ( .B1(n612), .B2(n630), .A(n486), .ZN(n253) );
  AOI221_X1 U89 ( .B1(n199), .B2(n361), .C1(B[4]), .C2(n55), .A(n418), .ZN(
        n409) );
  INV_X1 U90 ( .A(n214), .ZN(n55) );
  OAI222_X1 U91 ( .A1(n61), .A2(n644), .B1(n363), .B2(n635), .C1(n81), .C2(
        n637), .ZN(n418) );
  AOI221_X1 U92 ( .B1(n199), .B2(n350), .C1(B[4]), .C2(n49), .A(n404), .ZN(
        n392) );
  INV_X1 U93 ( .A(n202), .ZN(n49) );
  OAI222_X1 U94 ( .A1(n72), .A2(n644), .B1(n405), .B2(n635), .C1(n84), .C2(
        n637), .ZN(n404) );
  AOI221_X1 U95 ( .B1(n199), .B2(n339), .C1(B[4]), .C2(n47), .A(n386), .ZN(
        n378) );
  INV_X1 U96 ( .A(n188), .ZN(n47) );
  OAI222_X1 U97 ( .A1(n75), .A2(n644), .B1(n387), .B2(n635), .C1(n86), .C2(
        n637), .ZN(n386) );
  AOI221_X1 U98 ( .B1(n199), .B2(n324), .C1(n38), .C2(n172), .A(n371), .ZN(
        n365) );
  OAI222_X1 U99 ( .A1(n78), .A2(n644), .B1(n62), .B2(n635), .C1(n90), .C2(n637), .ZN(n371) );
  AOI221_X1 U100 ( .B1(n199), .B2(n313), .C1(n38), .C2(n139), .A(n360), .ZN(
        n352) );
  OAI222_X1 U101 ( .A1(n81), .A2(n644), .B1(n61), .B2(n635), .C1(n94), .C2(
        n637), .ZN(n360) );
  AOI221_X1 U102 ( .B1(n199), .B2(n289), .C1(n38), .C2(n348), .A(n349), .ZN(
        n341) );
  OAI222_X1 U103 ( .A1(n84), .A2(n644), .B1(n72), .B2(n635), .C1(n98), .C2(
        n637), .ZN(n349) );
  AOI221_X1 U104 ( .B1(n199), .B2(n270), .C1(n38), .C2(n337), .A(n338), .ZN(
        n328) );
  OAI222_X1 U105 ( .A1(n86), .A2(n644), .B1(n75), .B2(n635), .C1(n103), .C2(
        n637), .ZN(n338) );
  NOR2_X1 U106 ( .A1(n612), .A2(n646), .ZN(n359) );
  AOI221_X1 U107 ( .B1(n276), .B2(n479), .C1(n627), .C2(n480), .A(n279), .ZN(
        n478) );
  OAI21_X1 U108 ( .B1(n482), .B2(n281), .A(n282), .ZN(n479) );
  AOI21_X1 U109 ( .B1(n283), .B2(n485), .A(n285), .ZN(n482) );
  OAI21_X1 U110 ( .B1(n88), .B2(n287), .A(n288), .ZN(n485) );
  AOI221_X1 U111 ( .B1(n276), .B2(n470), .C1(n627), .C2(n434), .A(n279), .ZN(
        n469) );
  OAI21_X1 U112 ( .B1(n472), .B2(n281), .A(n282), .ZN(n470) );
  AOI21_X1 U113 ( .B1(n283), .B2(n473), .A(n285), .ZN(n472) );
  OAI21_X1 U114 ( .B1(n93), .B2(n287), .A(n288), .ZN(n473) );
  AOI221_X1 U115 ( .B1(n276), .B2(n460), .C1(n627), .C2(n297), .A(n279), .ZN(
        n459) );
  OAI21_X1 U116 ( .B1(n462), .B2(n281), .A(n282), .ZN(n460) );
  AOI21_X1 U117 ( .B1(n283), .B2(n463), .A(n285), .ZN(n462) );
  OAI21_X1 U118 ( .B1(n97), .B2(n287), .A(n288), .ZN(n463) );
  AOI221_X1 U119 ( .B1(n276), .B2(n448), .C1(n627), .C2(n246), .A(n279), .ZN(
        n447) );
  OAI21_X1 U120 ( .B1(n450), .B2(n281), .A(n282), .ZN(n448) );
  AOI21_X1 U121 ( .B1(n283), .B2(n451), .A(n285), .ZN(n450) );
  OAI21_X1 U122 ( .B1(n101), .B2(n287), .A(n288), .ZN(n451) );
  AOI221_X1 U123 ( .B1(n276), .B2(n424), .C1(n627), .C2(n106), .A(n279), .ZN(
        n423) );
  INV_X1 U124 ( .A(n238), .ZN(n106) );
  OAI21_X1 U125 ( .B1(n425), .B2(n281), .A(n282), .ZN(n424) );
  AOI21_X1 U126 ( .B1(n283), .B2(n426), .A(n285), .ZN(n425) );
  AOI221_X1 U127 ( .B1(n276), .B2(n411), .C1(n627), .C2(n223), .A(n279), .ZN(
        n410) );
  OAI21_X1 U128 ( .B1(n414), .B2(n281), .A(n282), .ZN(n411) );
  AOI21_X1 U129 ( .B1(n283), .B2(n415), .A(n285), .ZN(n414) );
  OAI21_X1 U130 ( .B1(n109), .B2(n287), .A(n288), .ZN(n415) );
  AOI221_X1 U131 ( .B1(n276), .B2(n394), .C1(n627), .C2(n211), .A(n279), .ZN(
        n393) );
  OAI21_X1 U132 ( .B1(n397), .B2(n281), .A(n282), .ZN(n394) );
  AOI21_X1 U133 ( .B1(n283), .B2(n398), .A(n285), .ZN(n397) );
  OAI21_X1 U134 ( .B1(n112), .B2(n287), .A(n288), .ZN(n398) );
  AOI221_X1 U135 ( .B1(n276), .B2(n380), .C1(n627), .C2(n114), .A(n279), .ZN(
        n379) );
  OAI21_X1 U136 ( .B1(n384), .B2(n281), .A(n282), .ZN(n380) );
  AOI21_X1 U137 ( .B1(n283), .B2(n385), .A(n285), .ZN(n384) );
  OAI21_X1 U138 ( .B1(n197), .B2(n287), .A(n288), .ZN(n385) );
  AOI221_X1 U139 ( .B1(n276), .B2(n367), .C1(n627), .C2(n118), .A(n279), .ZN(
        n366) );
  OAI21_X1 U140 ( .B1(n368), .B2(n281), .A(n282), .ZN(n367) );
  AOI21_X1 U141 ( .B1(n283), .B2(n369), .A(n285), .ZN(n368) );
  OAI21_X1 U142 ( .B1(n181), .B2(n287), .A(n288), .ZN(n369) );
  AOI221_X1 U143 ( .B1(n276), .B2(n354), .C1(n627), .C2(n121), .A(n279), .ZN(
        n353) );
  INV_X1 U144 ( .A(n163), .ZN(n121) );
  OAI21_X1 U145 ( .B1(n357), .B2(n281), .A(n282), .ZN(n354) );
  AOI21_X1 U146 ( .B1(n283), .B2(n358), .A(n285), .ZN(n357) );
  AOI221_X1 U147 ( .B1(n276), .B2(n343), .C1(n627), .C2(n124), .A(n279), .ZN(
        n342) );
  INV_X1 U148 ( .A(n344), .ZN(n124) );
  OAI21_X1 U149 ( .B1(n345), .B2(n281), .A(n282), .ZN(n343) );
  AOI21_X1 U150 ( .B1(n283), .B2(n346), .A(n285), .ZN(n345) );
  NOR2_X1 U151 ( .A1(n612), .A2(n2), .ZN(n519) );
  AOI221_X1 U152 ( .B1(n165), .B2(n429), .C1(n199), .C2(n373), .A(n492), .ZN(
        n477) );
  OAI222_X1 U153 ( .A1(n374), .A2(n635), .B1(n375), .B2(n640), .C1(n376), .C2(
        n644), .ZN(n492) );
  AOI221_X1 U154 ( .B1(n165), .B2(n474), .C1(n199), .C2(n419), .A(n475), .ZN(
        n468) );
  OAI222_X1 U155 ( .A1(n131), .A2(n635), .B1(n362), .B2(n640), .C1(n363), .C2(
        n644), .ZN(n475) );
  AOI221_X1 U156 ( .B1(n165), .B2(n465), .C1(n199), .C2(n406), .A(n466), .ZN(
        n458) );
  OAI222_X1 U157 ( .A1(n613), .A2(n635), .B1(n293), .B2(n640), .C1(n405), .C2(
        n644), .ZN(n466) );
  AOI221_X1 U158 ( .B1(n165), .B2(n455), .C1(n199), .C2(n388), .A(n456), .ZN(
        n446) );
  OAI222_X1 U159 ( .A1(n615), .A2(n635), .B1(n45), .B2(n640), .C1(n387), .C2(
        n644), .ZN(n456) );
  AOI221_X1 U160 ( .B1(n165), .B2(n373), .C1(n199), .C2(n372), .A(n427), .ZN(
        n422) );
  OAI221_X1 U161 ( .B1(n376), .B2(n635), .C1(n62), .C2(n644), .A(n428), .ZN(
        n427) );
  OAI22_X1 U162 ( .A1(n8), .A2(n130), .B1(n1), .B2(n135), .ZN(n533) );
  NOR2_X1 U163 ( .A1(n612), .A2(n8), .ZN(n382) );
  OAI221_X1 U164 ( .B1(n109), .B2(n160), .C1(n92), .C2(n161), .A(n162), .ZN(
        n220) );
  OAI221_X1 U165 ( .B1(n112), .B2(n160), .C1(n96), .C2(n161), .A(n162), .ZN(
        n208) );
  OAI221_X1 U166 ( .B1(n197), .B2(n160), .C1(n100), .C2(n161), .A(n162), .ZN(
        n194) );
  AOI22_X1 U167 ( .A1(n480), .A2(n38), .B1(n42), .B2(n63), .ZN(n587) );
  INV_X1 U168 ( .A(n601), .ZN(n63) );
  AOI221_X1 U169 ( .B1(n4), .B2(n602), .C1(n454), .C2(n184), .A(n603), .ZN(
        n601) );
  OAI22_X1 U170 ( .A1(n617), .A2(n638), .B1(n64), .B2(n645), .ZN(n603) );
  AOI22_X1 U171 ( .A1(n420), .A2(n2), .B1(n57), .B2(n262), .ZN(n214) );
  AOI22_X1 U172 ( .A1(n407), .A2(n5), .B1(n51), .B2(n262), .ZN(n202) );
  AOI22_X1 U173 ( .A1(n389), .A2(n3), .B1(n390), .B2(n262), .ZN(n188) );
  AOI22_X1 U174 ( .A1(n452), .A2(n4), .B1(n453), .B2(n262), .ZN(n449) );
  AOI22_X1 U175 ( .A1(n168), .A2(n3), .B1(n355), .B2(n262), .ZN(n413) );
  AOI22_X1 U176 ( .A1(n402), .A2(n5), .B1(n403), .B2(n262), .ZN(n396) );
  AOI22_X1 U177 ( .A1(n370), .A2(n4), .B1(n320), .B2(n262), .ZN(n182) );
  AOI22_X1 U178 ( .A1(n355), .A2(n2), .B1(n128), .B2(n262), .ZN(n163) );
  AOI22_X1 U179 ( .A1(n403), .A2(n4), .B1(n133), .B2(n262), .ZN(n344) );
  AOI21_X1 U180 ( .B1(n148), .B2(n217), .A(n150), .ZN(n216) );
  OAI21_X1 U181 ( .B1(n218), .B2(n152), .A(n153), .ZN(n217) );
  AOI211_X1 U182 ( .C1(n643), .C2(n219), .A(n220), .B(n221), .ZN(n218) );
  OAI22_X1 U183 ( .A1(n70), .A2(n157), .B1(n80), .B2(n158), .ZN(n221) );
  AOI21_X1 U184 ( .B1(n148), .B2(n205), .A(n150), .ZN(n204) );
  OAI21_X1 U185 ( .B1(n206), .B2(n152), .A(n153), .ZN(n205) );
  AOI211_X1 U186 ( .C1(n643), .C2(n207), .A(n208), .B(n209), .ZN(n206) );
  OAI22_X1 U187 ( .A1(n67), .A2(n157), .B1(n83), .B2(n158), .ZN(n209) );
  AOI21_X1 U188 ( .B1(n148), .B2(n191), .A(n150), .ZN(n190) );
  OAI21_X1 U189 ( .B1(n192), .B2(n152), .A(n153), .ZN(n191) );
  AOI211_X1 U190 ( .C1(n643), .C2(n193), .A(n194), .B(n195), .ZN(n192) );
  OAI22_X1 U191 ( .A1(n74), .A2(n157), .B1(n196), .B2(n158), .ZN(n195) );
  OAI211_X1 U192 ( .C1(n126), .C2(n645), .A(n401), .B(n449), .ZN(n257) );
  AOI21_X1 U193 ( .B1(n320), .B2(n4), .A(n519), .ZN(n323) );
  AOI21_X1 U194 ( .B1(n506), .B2(n5), .A(n519), .ZN(n336) );
  NAND2_X1 U195 ( .A1(n484), .A2(n632), .ZN(n249) );
  OAI21_X1 U196 ( .B1(n417), .B2(n636), .A(n471), .ZN(n440) );
  OAI21_X1 U197 ( .B1(n400), .B2(n636), .A(n461), .ZN(n302) );
  OAI21_X1 U198 ( .B1(n412), .B2(n636), .A(n471), .ZN(n434) );
  OAI21_X1 U199 ( .B1(n395), .B2(n636), .A(n461), .ZN(n297) );
  OAI21_X1 U200 ( .B1(n412), .B2(n645), .A(n413), .ZN(n223) );
  OAI21_X1 U201 ( .B1(n395), .B2(n645), .A(n396), .ZN(n211) );
  OAI21_X1 U202 ( .B1(n333), .B2(n646), .A(n449), .ZN(n246) );
  NOR2_X1 U203 ( .A1(n612), .A2(n484), .ZN(n483) );
  OAI21_X1 U204 ( .B1(n237), .B2(n287), .A(n288), .ZN(n426) );
  OAI21_X1 U205 ( .B1(n159), .B2(n287), .A(n288), .ZN(n358) );
  OAI21_X1 U206 ( .B1(n347), .B2(n287), .A(n288), .ZN(n346) );
  OAI21_X1 U207 ( .B1(n336), .B2(n287), .A(n288), .ZN(n335) );
  BUF_X1 U208 ( .A(n137), .Z(n35) );
  BUF_X1 U209 ( .A(n137), .Z(n36) );
  OAI21_X1 U210 ( .B1(n233), .B2(n152), .A(n153), .ZN(n232) );
  AOI211_X1 U211 ( .C1(n643), .C2(n234), .A(n235), .B(n236), .ZN(n233) );
  OAI22_X1 U212 ( .A1(n64), .A2(n157), .B1(n77), .B2(n158), .ZN(n236) );
  OAI221_X1 U213 ( .B1(n237), .B2(n160), .C1(n89), .C2(n161), .A(n162), .ZN(
        n235) );
  OAI21_X1 U214 ( .B1(n177), .B2(n152), .A(n153), .ZN(n176) );
  AOI211_X1 U215 ( .C1(n643), .C2(n178), .A(n179), .B(n180), .ZN(n177) );
  OAI22_X1 U216 ( .A1(n77), .A2(n157), .B1(n89), .B2(n158), .ZN(n180) );
  OAI221_X1 U217 ( .B1(n181), .B2(n160), .C1(n105), .C2(n161), .A(n162), .ZN(
        n179) );
  OAI21_X1 U218 ( .B1(n151), .B2(n152), .A(n153), .ZN(n149) );
  AOI211_X1 U219 ( .C1(n643), .C2(n154), .A(n155), .B(n156), .ZN(n151) );
  OAI22_X1 U220 ( .A1(n80), .A2(n157), .B1(n92), .B2(n158), .ZN(n156) );
  OAI221_X1 U221 ( .B1(n159), .B2(n160), .C1(n108), .C2(n161), .A(n162), .ZN(
        n155) );
  OAI21_X1 U222 ( .B1(n576), .B2(n152), .A(n153), .ZN(n575) );
  AOI211_X1 U223 ( .C1(n643), .C2(n305), .A(n577), .B(n578), .ZN(n576) );
  OAI22_X1 U224 ( .A1(n83), .A2(n157), .B1(n96), .B2(n158), .ZN(n578) );
  OAI221_X1 U225 ( .B1(n347), .B2(n160), .C1(n111), .C2(n161), .A(n162), .ZN(
        n577) );
  OAI21_X1 U226 ( .B1(n559), .B2(n152), .A(n153), .ZN(n558) );
  AOI211_X1 U227 ( .C1(n643), .C2(n261), .A(n560), .B(n561), .ZN(n559) );
  OAI22_X1 U228 ( .A1(n196), .A2(n157), .B1(n100), .B2(n158), .ZN(n561) );
  OAI221_X1 U229 ( .B1(n336), .B2(n160), .C1(n115), .C2(n161), .A(n162), .ZN(
        n560) );
  OAI21_X1 U230 ( .B1(n547), .B2(n152), .A(n153), .ZN(n546) );
  AOI211_X1 U231 ( .C1(n643), .C2(n184), .A(n548), .B(n549), .ZN(n547) );
  OAI22_X1 U232 ( .A1(n89), .A2(n157), .B1(n105), .B2(n158), .ZN(n549) );
  OAI221_X1 U233 ( .B1(n323), .B2(n160), .C1(n117), .C2(n161), .A(n162), .ZN(
        n548) );
  OAI21_X1 U234 ( .B1(n530), .B2(n152), .A(n153), .ZN(n529) );
  AOI211_X1 U235 ( .C1(n643), .C2(n166), .A(n531), .B(n532), .ZN(n530) );
  OAI22_X1 U236 ( .A1(n92), .A2(n157), .B1(n108), .B2(n158), .ZN(n532) );
  OAI221_X1 U237 ( .B1(n312), .B2(n160), .C1(n120), .C2(n161), .A(n162), .ZN(
        n531) );
  OAI21_X1 U238 ( .B1(n515), .B2(n152), .A(n153), .ZN(n514) );
  AOI211_X1 U239 ( .C1(n643), .C2(n516), .A(n517), .B(n518), .ZN(n515) );
  OAI22_X1 U240 ( .A1(n96), .A2(n157), .B1(n111), .B2(n158), .ZN(n518) );
  OAI221_X1 U241 ( .B1(n286), .B2(n160), .C1(n123), .C2(n161), .A(n162), .ZN(
        n517) );
  INV_X1 U242 ( .A(n452), .ZN(n100) );
  INV_X1 U243 ( .A(n170), .ZN(n92) );
  INV_X1 U244 ( .A(n464), .ZN(n96) );
  INV_X1 U245 ( .A(n186), .ZN(n89) );
  INV_X1 U246 ( .A(n166), .ZN(n80) );
  INV_X1 U247 ( .A(n516), .ZN(n83) );
  NOR2_X1 U248 ( .A1(n135), .A2(n8), .ZN(n580) );
  OAI21_X1 U249 ( .B1(n587), .B2(n255), .A(n256), .ZN(n595) );
  AOI21_X1 U250 ( .B1(n251), .B2(n438), .A(n253), .ZN(n437) );
  OAI21_X1 U251 ( .B1(n439), .B2(n255), .A(n256), .ZN(n438) );
  AOI22_X1 U252 ( .A1(n435), .A2(n39), .B1(B[4]), .B2(n440), .ZN(n439) );
  AOI21_X1 U253 ( .B1(n251), .B2(n300), .A(n253), .ZN(n299) );
  OAI21_X1 U254 ( .B1(n301), .B2(n255), .A(n256), .ZN(n300) );
  AOI22_X1 U255 ( .A1(n298), .A2(n39), .B1(B[4]), .B2(n302), .ZN(n301) );
  AOI21_X1 U256 ( .B1(n251), .B2(n252), .A(n253), .ZN(n248) );
  OAI21_X1 U257 ( .B1(n254), .B2(n255), .A(n256), .ZN(n252) );
  AOI22_X1 U258 ( .A1(n247), .A2(n39), .B1(B[4]), .B2(n257), .ZN(n254) );
  BUF_X1 U259 ( .A(n356), .Z(n2) );
  BUF_X1 U260 ( .A(n356), .Z(n3) );
  INV_X1 U261 ( .A(n293), .ZN(n51) );
  INV_X1 U262 ( .A(n184), .ZN(n77) );
  INV_X1 U263 ( .A(n506), .ZN(n126) );
  INV_X1 U265 ( .A(n185), .ZN(n105) );
  INV_X1 U266 ( .A(n390), .ZN(n45) );
  BUF_X1 U268 ( .A(n356), .Z(n4) );
  BUF_X1 U270 ( .A(n356), .Z(n5) );
  INV_X1 U271 ( .A(n453), .ZN(n115) );
  INV_X1 U272 ( .A(n412), .ZN(n128) );
  INV_X1 U273 ( .A(n395), .ZN(n133) );
  INV_X1 U274 ( .A(n154), .ZN(n70) );
  INV_X1 U275 ( .A(n305), .ZN(n67) );
  INV_X1 U276 ( .A(n178), .ZN(n64) );
  INV_X1 U277 ( .A(n168), .ZN(n108) );
  INV_X1 U278 ( .A(n402), .ZN(n111) );
  INV_X1 U279 ( .A(n261), .ZN(n74) );
  INV_X1 U280 ( .A(n419), .ZN(n81) );
  INV_X1 U281 ( .A(n406), .ZN(n84) );
  INV_X1 U282 ( .A(n388), .ZN(n86) );
  BUF_X1 U283 ( .A(n43), .Z(n41) );
  INV_X1 U284 ( .A(n362), .ZN(n57) );
  INV_X1 U285 ( .A(n474), .ZN(n61) );
  INV_X1 U286 ( .A(n465), .ZN(n72) );
  INV_X1 U287 ( .A(n455), .ZN(n75) );
  INV_X1 U288 ( .A(n267), .ZN(n8) );
  INV_X1 U289 ( .A(n355), .ZN(n120) );
  INV_X1 U290 ( .A(n403), .ZN(n123) );
  BUF_X1 U291 ( .A(n43), .Z(n42) );
  BUF_X1 U292 ( .A(n43), .Z(n39) );
  BUF_X1 U293 ( .A(n43), .Z(n40) );
  INV_X1 U294 ( .A(n370), .ZN(n117) );
  INV_X1 U295 ( .A(n373), .ZN(n78) );
  INV_X1 U296 ( .A(n420), .ZN(n131) );
  INV_X1 U297 ( .A(n407), .ZN(n613) );
  INV_X1 U298 ( .A(n389), .ZN(n615) );
  INV_X1 U299 ( .A(n417), .ZN(n129) );
  INV_X1 U300 ( .A(n400), .ZN(n134) );
  INV_X1 U301 ( .A(n429), .ZN(n62) );
  INV_X1 U302 ( .A(n372), .ZN(n90) );
  INV_X1 U303 ( .A(n361), .ZN(n94) );
  INV_X1 U304 ( .A(n350), .ZN(n98) );
  INV_X1 U305 ( .A(n339), .ZN(n103) );
  AND2_X1 U306 ( .A1(n238), .A2(n401), .ZN(n237) );
  INV_X1 U307 ( .A(n234), .ZN(n617) );
  INV_X1 U308 ( .A(n416), .ZN(n109) );
  OAI211_X1 U309 ( .C1(n417), .C2(n645), .A(n401), .B(n413), .ZN(n416) );
  INV_X1 U310 ( .A(n399), .ZN(n112) );
  OAI211_X1 U311 ( .C1(n400), .C2(n645), .A(n401), .B(n396), .ZN(n399) );
  INV_X1 U312 ( .A(n381), .ZN(n114) );
  AOI21_X1 U313 ( .B1(n260), .B2(n382), .A(n383), .ZN(n381) );
  BUF_X1 U314 ( .A(n137), .Z(n37) );
  OR4_X1 U315 ( .A1(B[21]), .A2(B[20]), .A3(B[19]), .A4(B[18]), .ZN(n598) );
  OAI22_X1 U316 ( .A1(n87), .A2(n1), .B1(n85), .B2(n8), .ZN(n568) );
  OAI22_X1 U317 ( .A1(n622), .A2(n1), .B1(n623), .B2(n8), .ZN(n525) );
  OAI22_X1 U318 ( .A1(n623), .A2(n1), .B1(n65), .B2(n8), .ZN(n570) );
  OAI22_X1 U319 ( .A1(n65), .A2(n1), .B1(n73), .B2(n8), .ZN(n552) );
  AOI221_X1 U320 ( .B1(n31), .B2(A[5]), .C1(n20), .C2(A[6]), .A(n541), .ZN(
        n376) );
  OAI22_X1 U321 ( .A1(n621), .A2(n1), .B1(n622), .B2(n8), .ZN(n541) );
  OAI221_X1 U322 ( .B1(n27), .B2(n612), .C1(n17), .C2(n135), .A(n609), .ZN(
        n320) );
  AOI22_X1 U323 ( .A1(A[29]), .A2(n10), .B1(A[28]), .B2(n7), .ZN(n609) );
  OAI221_X1 U324 ( .B1(n25), .B2(n127), .C1(n15), .C2(n125), .A(n535), .ZN(
        n355) );
  AOI22_X1 U325 ( .A1(A[26]), .A2(n9), .B1(A[25]), .B2(n267), .ZN(n535) );
  OAI221_X1 U326 ( .B1(n26), .B2(n130), .C1(n16), .C2(n127), .A(n585), .ZN(
        n403) );
  AOI22_X1 U327 ( .A1(A[27]), .A2(n10), .B1(A[26]), .B2(n7), .ZN(n585) );
  OR3_X1 U328 ( .A1(B[22]), .A2(B[24]), .A3(B[23]), .ZN(n594) );
  NAND3_X1 U329 ( .A1(n489), .A2(n628), .A3(n600), .ZN(n152) );
  NOR3_X1 U330 ( .A1(B[12]), .A2(B[14]), .A3(B[13]), .ZN(n600) );
  NAND3_X1 U331 ( .A1(n592), .A2(n631), .A3(n599), .ZN(n146) );
  INV_X1 U332 ( .A(B[22]), .ZN(n631) );
  NOR3_X1 U333 ( .A1(B[23]), .A2(B[25]), .A3(B[24]), .ZN(n599) );
  OAI221_X1 U334 ( .B1(n27), .B2(n85), .C1(n17), .C2(n82), .A(n606), .ZN(n184)
         );
  AOI22_X1 U335 ( .A1(A[13]), .A2(n11), .B1(A[12]), .B2(n7), .ZN(n606) );
  OAI221_X1 U336 ( .B1(n27), .B2(n125), .C1(n17), .C2(n122), .A(n608), .ZN(
        n370) );
  AOI22_X1 U337 ( .A1(A[25]), .A2(n9), .B1(A[24]), .B2(n7), .ZN(n608) );
  NAND2_X1 U338 ( .A1(n488), .A2(n489), .ZN(n287) );
  OAI221_X1 U339 ( .B1(n25), .B2(n116), .C1(n15), .C2(n113), .A(n536), .ZN(
        n168) );
  AOI22_X1 U340 ( .A1(A[22]), .A2(n9), .B1(A[21]), .B2(n267), .ZN(n536) );
  OAI221_X1 U341 ( .B1(n26), .B2(n119), .C1(n16), .C2(n116), .A(n583), .ZN(
        n402) );
  AOI22_X1 U342 ( .A1(A[23]), .A2(n10), .B1(A[22]), .B2(n7), .ZN(n583) );
  NOR2_X2 U343 ( .A1(n490), .A2(B[11]), .ZN(n283) );
  NAND2_X1 U344 ( .A1(A[31]), .A2(n647), .ZN(n162) );
  AOI221_X1 U345 ( .B1(A[1]), .B2(n31), .C1(A[2]), .C2(n21), .A(n540), .ZN(
        n374) );
  OAI22_X1 U346 ( .A1(n614), .A2(n1), .B1(n616), .B2(n8), .ZN(n540) );
  NOR2_X2 U347 ( .A1(n266), .A2(n591), .ZN(n144) );
  NAND2_X1 U348 ( .A1(A[31]), .A2(n152), .ZN(n153) );
  NAND2_X1 U349 ( .A1(A[31]), .A2(n146), .ZN(n147) );
  OAI221_X1 U350 ( .B1(n26), .B2(n135), .C1(n16), .C2(n130), .A(n564), .ZN(
        n506) );
  AOI22_X1 U351 ( .A1(A[28]), .A2(n10), .B1(A[27]), .B2(n6), .ZN(n564) );
  OAI221_X1 U352 ( .B1(n26), .B2(n122), .C1(n16), .C2(n119), .A(n565), .ZN(
        n453) );
  AOI22_X1 U353 ( .A1(A[24]), .A2(n10), .B1(A[23]), .B2(n6), .ZN(n565) );
  NOR2_X2 U354 ( .A1(n646), .A2(B[2]), .ZN(n260) );
  OAI221_X1 U355 ( .B1(n24), .B2(n113), .C1(n14), .C2(n110), .A(n611), .ZN(
        n185) );
  AOI22_X1 U356 ( .A1(A[21]), .A2(n11), .B1(A[20]), .B2(n6), .ZN(n611) );
  AOI222_X1 U357 ( .A1(n429), .A2(n5), .B1(n619), .B2(n262), .C1(n227), .C2(
        B[3]), .ZN(n327) );
  INV_X1 U358 ( .A(n376), .ZN(n619) );
  OAI221_X1 U359 ( .B1(n24), .B2(n76), .C1(n15), .C2(n73), .A(n444), .ZN(n154)
         );
  AOI22_X1 U360 ( .A1(A[10]), .A2(n11), .B1(A[9]), .B2(n267), .ZN(n444) );
  OAI221_X1 U361 ( .B1(n27), .B2(n79), .C1(n16), .C2(n76), .A(n586), .ZN(n305)
         );
  AOI22_X1 U362 ( .A1(A[11]), .A2(n10), .B1(A[10]), .B2(n7), .ZN(n586) );
  OAI221_X1 U363 ( .B1(n26), .B2(n82), .C1(n16), .C2(n79), .A(n567), .ZN(n261)
         );
  AOI22_X1 U364 ( .A1(A[12]), .A2(n10), .B1(A[11]), .B2(n6), .ZN(n567) );
  OAI221_X1 U365 ( .B1(n24), .B2(n622), .C1(n14), .C2(n621), .A(n443), .ZN(
        n219) );
  AOI22_X1 U366 ( .A1(A[6]), .A2(n11), .B1(A[5]), .B2(n267), .ZN(n443) );
  OAI221_X1 U367 ( .B1(n24), .B2(n623), .C1(n14), .C2(n622), .A(n306), .ZN(
        n207) );
  AOI22_X1 U368 ( .A1(A[7]), .A2(n11), .B1(A[6]), .B2(n7), .ZN(n306) );
  OAI221_X1 U369 ( .B1(n25), .B2(n65), .C1(n15), .C2(n623), .A(n265), .ZN(n193) );
  AOI22_X1 U370 ( .A1(A[8]), .A2(n9), .B1(A[7]), .B2(n6), .ZN(n265) );
  OAI221_X1 U371 ( .B1(n27), .B2(n99), .C1(n17), .C2(n95), .A(n610), .ZN(n186)
         );
  AOI22_X1 U372 ( .A1(A[17]), .A2(n11), .B1(A[16]), .B2(n7), .ZN(n610) );
  OAI221_X1 U373 ( .B1(n27), .B2(n73), .C1(n17), .C2(n65), .A(n604), .ZN(n178)
         );
  AOI22_X1 U374 ( .A1(A[9]), .A2(n9), .B1(A[8]), .B2(n7), .ZN(n604) );
  OAI221_X1 U375 ( .B1(n25), .B2(n87), .C1(n15), .C2(n85), .A(n537), .ZN(n166)
         );
  AOI22_X1 U376 ( .A1(A[14]), .A2(n9), .B1(A[13]), .B2(n6), .ZN(n537) );
  OAI221_X1 U377 ( .B1(n26), .B2(n91), .C1(n16), .C2(n87), .A(n584), .ZN(n516)
         );
  AOI22_X1 U378 ( .A1(A[15]), .A2(n10), .B1(A[14]), .B2(n6), .ZN(n584) );
  OAI221_X1 U379 ( .B1(n25), .B2(n79), .C1(n15), .C2(n82), .A(n494), .ZN(n373)
         );
  AOI22_X1 U380 ( .A1(A[15]), .A2(n9), .B1(A[16]), .B2(n267), .ZN(n494) );
  OAI221_X1 U381 ( .B1(n25), .B2(n132), .C1(n15), .C2(n614), .A(n523), .ZN(
        n420) );
  AOI22_X1 U382 ( .A1(A[4]), .A2(n9), .B1(A[5]), .B2(n267), .ZN(n523) );
  OAI221_X1 U383 ( .B1(n26), .B2(n614), .C1(n16), .C2(n616), .A(n571), .ZN(
        n407) );
  AOI22_X1 U384 ( .A1(A[5]), .A2(n10), .B1(A[6]), .B2(n6), .ZN(n571) );
  OAI221_X1 U385 ( .B1(n26), .B2(n616), .C1(n16), .C2(n618), .A(n554), .ZN(
        n389) );
  AOI22_X1 U386 ( .A1(A[6]), .A2(n10), .B1(A[7]), .B2(n6), .ZN(n554) );
  OAI221_X1 U387 ( .B1(n48), .B2(n27), .C1(n102), .C2(n14), .A(n553), .ZN(n390) );
  AOI22_X1 U389 ( .A1(A[2]), .A2(n10), .B1(A[3]), .B2(n6), .ZN(n553) );
  OAI221_X1 U390 ( .B1(n26), .B2(n623), .C1(n16), .C2(n65), .A(n542), .ZN(n429) );
  AOI22_X1 U391 ( .A1(A[11]), .A2(n10), .B1(A[12]), .B2(n6), .ZN(n542) );
  OAI221_X1 U392 ( .B1(n26), .B2(n110), .C1(n16), .C2(n107), .A(n566), .ZN(
        n452) );
  AOI22_X1 U393 ( .A1(A[20]), .A2(n10), .B1(A[19]), .B2(n6), .ZN(n566) );
  OAI221_X1 U394 ( .B1(n26), .B2(n104), .C1(n16), .C2(n99), .A(n538), .ZN(n170) );
  AOI22_X1 U395 ( .A1(A[18]), .A2(n10), .B1(A[17]), .B2(n6), .ZN(n538) );
  OAI221_X1 U396 ( .B1(n26), .B2(n107), .C1(n16), .C2(n104), .A(n582), .ZN(
        n464) );
  AOI22_X1 U397 ( .A1(A[19]), .A2(n10), .B1(A[18]), .B2(n6), .ZN(n582) );
  AOI22_X1 U398 ( .A1(n7), .A2(A[1]), .B1(n11), .B2(A[0]), .ZN(n362) );
  NAND2_X1 U399 ( .A1(B[4]), .A2(n579), .ZN(n160) );
  INV_X1 U400 ( .A(A[31]), .ZN(n612) );
  INV_X1 U401 ( .A(n332), .ZN(n627) );
  AOI21_X1 U402 ( .B1(A[31]), .B2(B[11]), .A(n487), .ZN(n256) );
  AOI21_X1 U403 ( .B1(A[31]), .B2(B[25]), .A(n483), .ZN(n250) );
  OAI221_X1 U404 ( .B1(n24), .B2(n91), .C1(n14), .C2(n95), .A(n430), .ZN(n372)
         );
  AOI22_X1 U405 ( .A1(A[19]), .A2(n11), .B1(A[20]), .B2(n7), .ZN(n430) );
  OAI221_X1 U406 ( .B1(n25), .B2(n82), .C1(n15), .C2(n85), .A(n476), .ZN(n419)
         );
  AOI22_X1 U407 ( .A1(A[16]), .A2(n9), .B1(A[17]), .B2(n267), .ZN(n476) );
  OAI221_X1 U408 ( .B1(n25), .B2(n85), .C1(n15), .C2(n87), .A(n467), .ZN(n406)
         );
  AOI22_X1 U409 ( .A1(A[17]), .A2(n9), .B1(A[18]), .B2(n267), .ZN(n467) );
  OAI221_X1 U410 ( .B1(n25), .B2(n87), .C1(n15), .C2(n91), .A(n457), .ZN(n388)
         );
  AOI22_X1 U411 ( .A1(A[18]), .A2(n9), .B1(A[19]), .B2(n267), .ZN(n457) );
  OAI221_X1 U412 ( .B1(n27), .B2(n621), .C1(n17), .C2(n620), .A(n605), .ZN(
        n234) );
  AOI22_X1 U413 ( .A1(A[5]), .A2(n11), .B1(A[4]), .B2(n7), .ZN(n605) );
  OAI221_X1 U414 ( .B1(n258), .B2(n642), .C1(n196), .C2(n636), .A(n259), .ZN(
        n247) );
  AOI22_X1 U415 ( .A1(n260), .A2(n261), .B1(n262), .B2(n193), .ZN(n259) );
  AOI222_X1 U416 ( .A1(A[4]), .A2(n11), .B1(A[6]), .B2(n29), .C1(A[5]), .C2(
        n18), .ZN(n258) );
  OAI221_X1 U417 ( .B1(n303), .B2(n642), .C1(n83), .C2(n636), .A(n304), .ZN(
        n298) );
  AOI22_X1 U418 ( .A1(n260), .A2(n305), .B1(n262), .B2(n207), .ZN(n304) );
  AOI222_X1 U419 ( .A1(A[3]), .A2(n11), .B1(A[5]), .B2(n28), .C1(A[4]), .C2(
        n19), .ZN(n303) );
  OAI221_X1 U420 ( .B1(n441), .B2(n642), .C1(n80), .C2(n636), .A(n442), .ZN(
        n435) );
  AOI22_X1 U421 ( .A1(n260), .A2(n154), .B1(n262), .B2(n219), .ZN(n442) );
  AOI222_X1 U422 ( .A1(A[2]), .A2(n9), .B1(A[4]), .B2(n28), .C1(A[3]), .C2(n18), .ZN(n441) );
  OAI221_X1 U423 ( .B1(n24), .B2(n95), .C1(n14), .C2(n99), .A(n421), .ZN(n361)
         );
  AOI22_X1 U424 ( .A1(A[20]), .A2(n11), .B1(A[21]), .B2(n6), .ZN(n421) );
  OAI221_X1 U425 ( .B1(n25), .B2(n65), .C1(n15), .C2(n73), .A(n524), .ZN(n474)
         );
  AOI22_X1 U426 ( .A1(A[12]), .A2(n9), .B1(A[13]), .B2(n267), .ZN(n524) );
  OAI221_X1 U427 ( .B1(n24), .B2(n99), .C1(n14), .C2(n104), .A(n408), .ZN(n350) );
  AOI22_X1 U429 ( .A1(A[21]), .A2(n9), .B1(A[22]), .B2(n7), .ZN(n408) );
  OAI221_X1 U430 ( .B1(n25), .B2(n73), .C1(n15), .C2(n76), .A(n510), .ZN(n465)
         );
  AOI22_X1 U431 ( .A1(A[13]), .A2(n9), .B1(A[14]), .B2(n267), .ZN(n510) );
  OAI221_X1 U432 ( .B1(n24), .B2(n104), .C1(n14), .C2(n107), .A(n391), .ZN(
        n339) );
  AOI22_X1 U433 ( .A1(A[22]), .A2(n10), .B1(A[23]), .B2(n6), .ZN(n391) );
  OAI221_X1 U434 ( .B1(n25), .B2(n76), .C1(n15), .C2(n79), .A(n497), .ZN(n455)
         );
  AOI22_X1 U435 ( .A1(A[14]), .A2(n9), .B1(A[15]), .B2(n6), .ZN(n497) );
  OAI221_X1 U436 ( .B1(n24), .B2(n107), .C1(n14), .C2(n110), .A(n377), .ZN(
        n324) );
  AOI22_X1 U437 ( .A1(A[23]), .A2(n9), .B1(A[24]), .B2(n7), .ZN(n377) );
  OAI221_X1 U438 ( .B1(n24), .B2(n110), .C1(n14), .C2(n113), .A(n364), .ZN(
        n313) );
  AOI22_X1 U439 ( .A1(A[24]), .A2(n11), .B1(A[25]), .B2(n6), .ZN(n364) );
  OAI221_X1 U440 ( .B1(n24), .B2(n113), .C1(n14), .C2(n116), .A(n351), .ZN(
        n289) );
  AOI22_X1 U441 ( .A1(A[25]), .A2(n9), .B1(A[26]), .B2(n7), .ZN(n351) );
  OAI221_X1 U442 ( .B1(n24), .B2(n116), .C1(n14), .C2(n119), .A(n340), .ZN(
        n270) );
  AOI22_X1 U443 ( .A1(A[26]), .A2(n10), .B1(A[27]), .B2(n6), .ZN(n340) );
  AOI221_X1 U444 ( .B1(n169), .B2(n452), .C1(n167), .C2(n453), .A(n563), .ZN(
        n562) );
  NOR3_X1 U445 ( .A1(n40), .A2(B[3]), .A3(n333), .ZN(n563) );
  AOI221_X1 U446 ( .B1(n242), .B2(n432), .C1(n626), .C2(n71), .A(n244), .ZN(
        n431) );
  INV_X1 U447 ( .A(n433), .ZN(n71) );
  OAI21_X1 U448 ( .B1(n437), .B2(n249), .A(n250), .ZN(n432) );
  AOI22_X1 U449 ( .A1(n434), .A2(n38), .B1(n41), .B2(n435), .ZN(n433) );
  AOI221_X1 U450 ( .B1(n242), .B2(n295), .C1(n626), .C2(n68), .A(n244), .ZN(
        n294) );
  INV_X1 U451 ( .A(n296), .ZN(n68) );
  OAI21_X1 U452 ( .B1(n299), .B2(n249), .A(n250), .ZN(n295) );
  AOI22_X1 U453 ( .A1(n297), .A2(n38), .B1(n41), .B2(n298), .ZN(n296) );
  AOI221_X1 U454 ( .B1(n242), .B2(n243), .C1(n626), .C2(n59), .A(n244), .ZN(
        n241) );
  INV_X1 U455 ( .A(n245), .ZN(n59) );
  OAI21_X1 U456 ( .B1(n248), .B2(n249), .A(n250), .ZN(n243) );
  AOI22_X1 U457 ( .A1(n246), .A2(n38), .B1(n42), .B2(n247), .ZN(n245) );
  AOI22_X1 U458 ( .A1(n639), .A2(n506), .B1(B[2]), .B2(n382), .ZN(n333) );
  AOI221_X1 U459 ( .B1(n276), .B2(n319), .C1(n278), .C2(n320), .A(n279), .ZN(
        n318) );
  OAI21_X1 U460 ( .B1(n321), .B2(n281), .A(n282), .ZN(n319) );
  AOI21_X1 U462 ( .B1(n283), .B2(n322), .A(n285), .ZN(n321) );
  OAI21_X1 U463 ( .B1(n323), .B2(n287), .A(n288), .ZN(n322) );
  AOI221_X1 U464 ( .B1(n276), .B2(n309), .C1(n278), .C2(n128), .A(n279), .ZN(
        n308) );
  OAI21_X1 U465 ( .B1(n310), .B2(n281), .A(n282), .ZN(n309) );
  AOI21_X1 U466 ( .B1(n283), .B2(n311), .A(n285), .ZN(n310) );
  OAI21_X1 U467 ( .B1(n312), .B2(n287), .A(n288), .ZN(n311) );
  AOI221_X1 U468 ( .B1(n276), .B2(n277), .C1(n278), .C2(n133), .A(n279), .ZN(
        n275) );
  OAI21_X1 U469 ( .B1(n280), .B2(n281), .A(n282), .ZN(n277) );
  AOI21_X1 U470 ( .B1(n283), .B2(n284), .A(n285), .ZN(n280) );
  OAI21_X1 U471 ( .B1(n286), .B2(n287), .A(n288), .ZN(n284) );
  AOI221_X1 U472 ( .B1(n165), .B2(n324), .C1(n38), .C2(n53), .A(n325), .ZN(
        n317) );
  INV_X1 U473 ( .A(n327), .ZN(n53) );
  OAI222_X1 U474 ( .A1(n78), .A2(n635), .B1(n326), .B2(n641), .C1(n90), .C2(
        n644), .ZN(n325) );
  AOI222_X1 U475 ( .A1(A[27]), .A2(n10), .B1(A[25]), .B2(n28), .C1(A[26]), 
        .C2(n19), .ZN(n326) );
  AOI221_X1 U476 ( .B1(n165), .B2(n313), .C1(n38), .C2(n314), .A(n315), .ZN(
        n307) );
  OAI222_X1 U477 ( .A1(n81), .A2(n635), .B1(n316), .B2(n641), .C1(n94), .C2(
        n644), .ZN(n315) );
  AOI222_X1 U478 ( .A1(A[28]), .A2(n11), .B1(A[26]), .B2(n28), .C1(A[27]), 
        .C2(n18), .ZN(n316) );
  AOI221_X1 U479 ( .B1(n165), .B2(n289), .C1(n38), .C2(n290), .A(n291), .ZN(
        n274) );
  OAI222_X1 U480 ( .A1(n84), .A2(n635), .B1(n292), .B2(n641), .C1(n98), .C2(
        n644), .ZN(n291) );
  AOI222_X1 U481 ( .A1(A[29]), .A2(n11), .B1(A[27]), .B2(n31), .C1(A[28]), 
        .C2(n18), .ZN(n292) );
  AOI221_X1 U482 ( .B1(n165), .B2(n270), .C1(n38), .C2(n271), .A(n272), .ZN(
        n268) );
  OAI222_X1 U483 ( .A1(n86), .A2(n635), .B1(n273), .B2(n641), .C1(n103), .C2(
        n644), .ZN(n272) );
  AOI222_X1 U484 ( .A1(A[30]), .A2(n11), .B1(A[28]), .B2(n30), .C1(A[29]), 
        .C2(n20), .ZN(n273) );
  NOR2_X1 U485 ( .A1(n490), .A2(B[18]), .ZN(n251) );
  OAI22_X1 U486 ( .A1(B[2]), .A2(n374), .B1(n639), .B2(n375), .ZN(n227) );
  AOI21_X1 U487 ( .B1(n20), .B2(A[31]), .A(n533), .ZN(n412) );
  AOI21_X1 U488 ( .B1(n11), .B2(A[31]), .A(n580), .ZN(n395) );
  AOI21_X1 U489 ( .B1(B[1]), .B2(A[31]), .A(n533), .ZN(n417) );
  AOI21_X1 U490 ( .B1(n8), .B2(A[31]), .A(n580), .ZN(n400) );
  NOR2_X1 U491 ( .A1(B[0]), .A2(B[1]), .ZN(n267) );
  AOI211_X1 U492 ( .C1(n276), .C2(n330), .A(n279), .B(n331), .ZN(n329) );
  OAI21_X1 U493 ( .B1(n334), .B2(n281), .A(n282), .ZN(n330) );
  NOR3_X1 U494 ( .A1(n332), .A2(B[3]), .A3(n333), .ZN(n331) );
  AOI21_X1 U495 ( .B1(n283), .B2(n335), .A(n285), .ZN(n334) );
  OAI221_X1 U496 ( .B1(n587), .B2(n436), .C1(n48), .C2(n32), .A(n588), .ZN(
        RES[0]) );
  AOI21_X1 U497 ( .B1(n242), .B2(n589), .A(n244), .ZN(n588) );
  OAI21_X1 U498 ( .B1(n593), .B2(n249), .A(n250), .ZN(n589) );
  AOI21_X1 U499 ( .B1(n251), .B2(n595), .A(n253), .ZN(n593) );
  AND2_X1 U500 ( .A1(n491), .A2(n632), .ZN(n276) );
  NAND2_X1 U501 ( .A1(A[31]), .A2(n490), .ZN(n486) );
  NOR2_X1 U502 ( .A1(B[2]), .A2(B[3]), .ZN(n356) );
  INV_X1 U503 ( .A(A[10]), .ZN(n65) );
  NAND2_X1 U504 ( .A1(n454), .A2(A[31]), .ZN(n401) );
  OAI21_X1 U505 ( .B1(n489), .B2(n612), .A(n162), .ZN(n487) );
  INV_X1 U506 ( .A(B[3]), .ZN(n646) );
  INV_X1 U507 ( .A(A[11]), .ZN(n73) );
  INV_X1 U508 ( .A(A[15]), .ZN(n85) );
  INV_X1 U509 ( .A(A[16]), .ZN(n87) );
  INV_X1 U510 ( .A(A[9]), .ZN(n623) );
  OAI21_X1 U511 ( .B1(n502), .B2(n152), .A(n153), .ZN(n501) );
  AOI211_X1 U512 ( .C1(B[4]), .C2(A[31]), .A(n503), .B(n504), .ZN(n502) );
  OAI22_X1 U513 ( .A1(n196), .A2(n505), .B1(n100), .B2(n157), .ZN(n504) );
  OAI221_X1 U514 ( .B1(n126), .B2(n161), .C1(n115), .C2(n158), .A(n162), .ZN(
        n503) );
  NAND2_X1 U515 ( .A1(A[0]), .A2(n7), .ZN(n375) );
  NOR2_X1 U516 ( .A1(n269), .A2(n38), .ZN(n228) );
  INV_X1 U517 ( .A(A[30]), .ZN(n135) );
  INV_X1 U518 ( .A(A[12]), .ZN(n76) );
  INV_X1 U519 ( .A(A[13]), .ZN(n79) );
  INV_X1 U520 ( .A(A[14]), .ZN(n82) );
  INV_X1 U521 ( .A(A[19]), .ZN(n99) );
  INV_X1 U522 ( .A(A[20]), .ZN(n104) );
  INV_X1 U523 ( .A(A[21]), .ZN(n107) );
  INV_X1 U524 ( .A(A[22]), .ZN(n110) );
  INV_X1 U525 ( .A(A[23]), .ZN(n113) );
  INV_X1 U526 ( .A(A[24]), .ZN(n116) );
  OR4_X1 U527 ( .A1(B[13]), .A2(B[14]), .A3(B[12]), .A4(n596), .ZN(n490) );
  OR3_X1 U528 ( .A1(B[15]), .A2(B[17]), .A3(B[16]), .ZN(n596) );
  INV_X1 U529 ( .A(B[2]), .ZN(n639) );
  INV_X1 U530 ( .A(A[8]), .ZN(n622) );
  INV_X1 U531 ( .A(A[3]), .ZN(n614) );
  AND3_X1 U532 ( .A1(n579), .A2(n591), .A3(n597), .ZN(n445) );
  NOR3_X1 U533 ( .A1(n152), .A2(n146), .A3(n629), .ZN(n597) );
  INV_X1 U534 ( .A(n148), .ZN(n629) );
  AND2_X1 U535 ( .A1(n491), .A2(n648), .ZN(n242) );
  INV_X1 U536 ( .A(A[17]), .ZN(n91) );
  INV_X1 U537 ( .A(A[7]), .ZN(n621) );
  INV_X1 U538 ( .A(A[18]), .ZN(n95) );
  INV_X1 U539 ( .A(A[25]), .ZN(n119) );
  INV_X1 U540 ( .A(A[29]), .ZN(n130) );
  INV_X1 U541 ( .A(B[25]), .ZN(n632) );
  INV_X1 U542 ( .A(A[4]), .ZN(n616) );
  INV_X1 U543 ( .A(A[27]), .ZN(n125) );
  INV_X1 U544 ( .A(A[26]), .ZN(n122) );
  INV_X1 U545 ( .A(A[6]), .ZN(n620) );
  INV_X1 U546 ( .A(A[5]), .ZN(n618) );
  INV_X1 U547 ( .A(A[28]), .ZN(n127) );
  NAND2_X1 U548 ( .A1(n34), .A2(n648), .ZN(n137) );
  INV_X1 U549 ( .A(A[2]), .ZN(n132) );
  INV_X1 U550 ( .A(n579), .ZN(n647) );
  OR2_X1 U551 ( .A1(n624), .A2(B[1]), .ZN(n1) );
  INV_X1 U552 ( .A(n436), .ZN(n626) );
  NAND2_X1 U553 ( .A1(B[1]), .A2(B[0]), .ZN(n263) );
  NAND2_X1 U554 ( .A1(B[1]), .A2(n624), .ZN(n264) );
  INV_X1 U555 ( .A(A[1]), .ZN(n102) );
  INV_X1 U556 ( .A(B[11]), .ZN(n628) );
  INV_X1 U557 ( .A(A[0]), .ZN(n48) );
  INV_X1 U558 ( .A(B[18]), .ZN(n630) );
  INV_X1 U559 ( .A(B[0]), .ZN(n624) );
  INV_X1 U560 ( .A(B[4]), .ZN(n43) );
  NOR3_X1 U561 ( .A1(B[9]), .A2(B[8]), .A3(B[10]), .ZN(n489) );
  NOR3_X1 U562 ( .A1(B[7]), .A2(B[6]), .A3(B[5]), .ZN(n579) );
  NOR3_X1 U563 ( .A1(B[28]), .A2(B[27]), .A3(B[26]), .ZN(n592) );
  NAND3_X1 U564 ( .A1(n445), .A2(n34), .A3(LEFT_RIGHT), .ZN(n269) );
  NOR2_X1 U565 ( .A1(n481), .A2(LEFT_RIGHT), .ZN(n244) );
  AOI221_X1 U566 ( .B1(n140), .B2(n229), .C1(n142), .C2(n230), .A(n144), .ZN(
        n225) );
  OAI21_X1 U567 ( .B1(n231), .B2(n146), .A(n147), .ZN(n230) );
  OAI221_X1 U568 ( .B1(n617), .B2(n641), .C1(n238), .C2(n40), .A(n239), .ZN(
        n229) );
  AOI21_X1 U569 ( .B1(n148), .B2(n232), .A(n150), .ZN(n231) );
  AOI221_X1 U570 ( .B1(n140), .B2(n498), .C1(n142), .C2(n499), .A(n144), .ZN(
        n495) );
  OAI21_X1 U571 ( .B1(n500), .B2(n146), .A(n147), .ZN(n499) );
  OAI221_X1 U572 ( .B1(n100), .B2(n637), .C1(n196), .C2(n641), .A(n507), .ZN(
        n498) );
  AOI21_X1 U573 ( .B1(n148), .B2(n501), .A(n150), .ZN(n500) );
  AOI221_X1 U574 ( .B1(n140), .B2(n69), .C1(n142), .C2(n215), .A(n144), .ZN(
        n213) );
  INV_X1 U575 ( .A(n222), .ZN(n69) );
  OAI21_X1 U576 ( .B1(n216), .B2(n146), .A(n147), .ZN(n215) );
  AOI221_X1 U577 ( .B1(n219), .B2(n199), .C1(n223), .C2(n38), .A(n224), .ZN(
        n222) );
  AOI221_X1 U578 ( .B1(n140), .B2(n66), .C1(n142), .C2(n203), .A(n144), .ZN(
        n201) );
  INV_X1 U579 ( .A(n210), .ZN(n66) );
  OAI21_X1 U580 ( .B1(n204), .B2(n146), .A(n147), .ZN(n203) );
  AOI221_X1 U581 ( .B1(n207), .B2(n199), .C1(n211), .C2(n38), .A(n212), .ZN(
        n210) );
  AOI221_X1 U582 ( .B1(n140), .B2(n60), .C1(n142), .C2(n189), .A(n144), .ZN(
        n187) );
  INV_X1 U583 ( .A(n198), .ZN(n60) );
  OAI21_X1 U584 ( .B1(n190), .B2(n146), .A(n147), .ZN(n189) );
  AOI221_X1 U585 ( .B1(n193), .B2(n199), .C1(n114), .C2(n38), .A(n200), .ZN(
        n198) );
  AOI221_X1 U586 ( .B1(n140), .B2(n173), .C1(n142), .C2(n174), .A(n144), .ZN(
        n171) );
  OAI21_X1 U587 ( .B1(n175), .B2(n146), .A(n147), .ZN(n174) );
  OAI221_X1 U588 ( .B1(n64), .B2(n641), .C1(n182), .C2(n40), .A(n183), .ZN(
        n173) );
  AOI21_X1 U589 ( .B1(n148), .B2(n176), .A(n150), .ZN(n175) );
  AOI221_X1 U590 ( .B1(n140), .B2(n141), .C1(n142), .C2(n143), .A(n144), .ZN(
        n136) );
  OAI21_X1 U591 ( .B1(n145), .B2(n146), .A(n147), .ZN(n143) );
  OAI221_X1 U592 ( .B1(n70), .B2(n641), .C1(n163), .C2(n41), .A(n164), .ZN(
        n141) );
  AOI21_X1 U593 ( .B1(n148), .B2(n149), .A(n150), .ZN(n145) );
  AOI221_X1 U594 ( .B1(n140), .B2(n572), .C1(n142), .C2(n573), .A(n144), .ZN(
        n569) );
  OAI21_X1 U595 ( .B1(n574), .B2(n146), .A(n147), .ZN(n573) );
  OAI221_X1 U596 ( .B1(n67), .B2(n641), .C1(n344), .C2(n41), .A(n581), .ZN(
        n572) );
  AOI21_X1 U597 ( .B1(n148), .B2(n575), .A(n150), .ZN(n574) );
  AOI221_X1 U598 ( .B1(n140), .B2(n555), .C1(n142), .C2(n556), .A(n144), .ZN(
        n551) );
  OAI21_X1 U599 ( .B1(n557), .B2(n146), .A(n147), .ZN(n556) );
  OAI221_X1 U600 ( .B1(n196), .B2(n637), .C1(n74), .C2(n641), .A(n562), .ZN(
        n555) );
  AOI21_X1 U601 ( .B1(n148), .B2(n558), .A(n150), .ZN(n557) );
  AOI221_X1 U602 ( .B1(n140), .B2(n543), .C1(n142), .C2(n544), .A(n144), .ZN(
        n539) );
  OAI21_X1 U603 ( .B1(n545), .B2(n146), .A(n147), .ZN(n544) );
  OAI221_X1 U604 ( .B1(n89), .B2(n637), .C1(n77), .C2(n641), .A(n550), .ZN(
        n543) );
  AOI21_X1 U605 ( .B1(n148), .B2(n546), .A(n150), .ZN(n545) );
  AOI221_X1 U606 ( .B1(n140), .B2(n526), .C1(n142), .C2(n527), .A(n144), .ZN(
        n521) );
  OAI21_X1 U607 ( .B1(n528), .B2(n146), .A(n147), .ZN(n527) );
  OAI221_X1 U608 ( .B1(n92), .B2(n637), .C1(n80), .C2(n641), .A(n534), .ZN(
        n526) );
  AOI21_X1 U609 ( .B1(n148), .B2(n529), .A(n150), .ZN(n528) );
  AOI221_X1 U610 ( .B1(n140), .B2(n511), .C1(n142), .C2(n512), .A(n144), .ZN(
        n508) );
  OAI21_X1 U611 ( .B1(n513), .B2(n146), .A(n147), .ZN(n512) );
  OAI221_X1 U612 ( .B1(n96), .B2(n637), .C1(n83), .C2(n641), .A(n520), .ZN(
        n511) );
  AOI21_X1 U613 ( .B1(n148), .B2(n514), .A(n150), .ZN(n513) );
  AOI21_X1 U614 ( .B1(n633), .B2(n590), .A(n144), .ZN(n481) );
  INV_X1 U615 ( .A(n592), .ZN(n633) );
  NOR2_X1 U616 ( .A1(B[29]), .A2(B[30]), .ZN(n591) );
  INV_X1 U617 ( .A(n590), .ZN(n266) );
  AND2_X1 U618 ( .A1(n140), .A2(n199), .ZN(n278) );
  NAND2_X1 U619 ( .A1(n140), .A2(n39), .ZN(n332) );
  NAND2_X1 U620 ( .A1(n140), .A2(n648), .ZN(n436) );
  INV_X1 U621 ( .A(LEFT_RIGHT), .ZN(n648) );
  AND2_X1 U622 ( .A1(n142), .A2(n592), .ZN(n491) );
  NOR2_X2 U623 ( .A1(n634), .A2(LOGIC_ARITH), .ZN(n142) );
  INV_X1 U624 ( .A(n591), .ZN(n634) );
  AND2_X1 U625 ( .A1(LOGIC_ARITH), .A2(n445), .ZN(n140) );
  NOR2_X1 U626 ( .A1(n612), .A2(LOGIC_ARITH), .ZN(n590) );
  OAI222_X1 U627 ( .A1(n268), .A2(n269), .B1(LEFT_RIGHT), .B2(n266), .C1(n612), 
        .C2(n33), .ZN(RES[31]) );
  OAI222_X1 U628 ( .A1(n187), .A2(n35), .B1(n188), .B2(n625), .C1(n621), .C2(
        n32), .ZN(RES[7]) );
  OAI222_X1 U629 ( .A1(n171), .A2(n35), .B1(n54), .B2(n625), .C1(n622), .C2(
        n32), .ZN(RES[8]) );
  OAI222_X1 U630 ( .A1(n136), .A2(n35), .B1(n58), .B2(n625), .C1(n623), .C2(
        n32), .ZN(RES[9]) );
  OAI222_X1 U631 ( .A1(n539), .A2(n35), .B1(n327), .B2(n625), .C1(n76), .C2(
        n34), .ZN(RES[12]) );
  OAI222_X1 U632 ( .A1(n521), .A2(n35), .B1(n56), .B2(n625), .C1(n79), .C2(n34), .ZN(RES[13]) );
  OAI222_X1 U633 ( .A1(n508), .A2(n35), .B1(n50), .B2(n625), .C1(n82), .C2(n34), .ZN(RES[14]) );
  OAI222_X1 U634 ( .A1(n468), .A2(n269), .B1(n469), .B2(n36), .C1(n91), .C2(
        n33), .ZN(RES[17]) );
  OAI222_X1 U635 ( .A1(n495), .A2(n35), .B1(n46), .B2(n625), .C1(n85), .C2(n34), .ZN(RES[15]) );
  OAI222_X1 U636 ( .A1(n458), .A2(n269), .B1(n459), .B2(n37), .C1(n95), .C2(
        n33), .ZN(RES[18]) );
  OAI222_X1 U640 ( .A1(n477), .A2(n269), .B1(n478), .B2(n37), .C1(n87), .C2(
        n34), .ZN(RES[16]) );
  OAI222_X1 U643 ( .A1(n446), .A2(n269), .B1(n447), .B2(n36), .C1(n99), .C2(
        n33), .ZN(RES[19]) );
  OAI222_X1 U644 ( .A1(n422), .A2(n269), .B1(n423), .B2(n36), .C1(n104), .C2(
        n33), .ZN(RES[20]) );
  OAI222_X1 U645 ( .A1(n409), .A2(n269), .B1(n410), .B2(n36), .C1(n107), .C2(
        n33), .ZN(RES[21]) );
  OAI222_X1 U646 ( .A1(n392), .A2(n269), .B1(n393), .B2(n36), .C1(n110), .C2(
        n33), .ZN(RES[22]) );
  OAI222_X1 U647 ( .A1(n378), .A2(n269), .B1(n379), .B2(n36), .C1(n113), .C2(
        n33), .ZN(RES[23]) );
  OAI222_X1 U648 ( .A1(n365), .A2(n269), .B1(n366), .B2(n36), .C1(n116), .C2(
        n33), .ZN(RES[24]) );
  OAI222_X1 U649 ( .A1(n352), .A2(n269), .B1(n353), .B2(n36), .C1(n119), .C2(
        n33), .ZN(RES[25]) );
  OAI222_X1 U650 ( .A1(n201), .A2(n35), .B1(n202), .B2(n625), .C1(n620), .C2(
        n32), .ZN(RES[6]) );
  OAI222_X1 U651 ( .A1(n569), .A2(n35), .B1(n52), .B2(n625), .C1(n65), .C2(n34), .ZN(RES[10]) );
  OAI222_X1 U652 ( .A1(n551), .A2(n35), .B1(n44), .B2(n625), .C1(n73), .C2(n34), .ZN(RES[11]) );
  OAI222_X1 U653 ( .A1(n341), .A2(n269), .B1(n342), .B2(n36), .C1(n122), .C2(
        n33), .ZN(RES[26]) );
  OAI222_X1 U654 ( .A1(n328), .A2(n269), .B1(n329), .B2(n36), .C1(n125), .C2(
        n33), .ZN(RES[27]) );
  OAI222_X1 U655 ( .A1(n213), .A2(n35), .B1(n214), .B2(n625), .C1(n618), .C2(
        n32), .ZN(RES[5]) );
  OAI222_X1 U656 ( .A1(n317), .A2(n269), .B1(n318), .B2(n36), .C1(n127), .C2(
        n33), .ZN(RES[28]) );
  OAI222_X1 U657 ( .A1(n307), .A2(n269), .B1(n308), .B2(n36), .C1(n130), .C2(
        n32), .ZN(RES[29]) );
  OAI222_X1 U658 ( .A1(n274), .A2(n269), .B1(n275), .B2(n37), .C1(n135), .C2(
        n32), .ZN(RES[30]) );
  OAI221_X1 U659 ( .B1(n293), .B2(n240), .C1(n132), .C2(n32), .A(n294), .ZN(
        RES[2]) );
  OAI221_X1 U660 ( .B1(n362), .B2(n240), .C1(n102), .C2(n32), .A(n431), .ZN(
        RES[1]) );
  OAI221_X1 U661 ( .B1(n45), .B2(n240), .C1(n614), .C2(n32), .A(n241), .ZN(
        RES[3]) );
  OAI221_X1 U662 ( .B1(n225), .B2(n35), .C1(n616), .C2(n32), .A(n226), .ZN(
        RES[4]) );
  NOR4_X4 U663 ( .A1(B[16]), .A2(B[17]), .A3(B[15]), .A4(n598), .ZN(n148) );
  INV_X1 U664 ( .A(n8), .ZN(n6) );
  INV_X1 U665 ( .A(n8), .ZN(n7) );
  INV_X1 U666 ( .A(n1), .ZN(n9) );
  INV_X1 U667 ( .A(n1), .ZN(n10) );
  INV_X1 U668 ( .A(n1), .ZN(n11) );
  CLKBUF_X1 U669 ( .A(n264), .Z(n12) );
  CLKBUF_X1 U670 ( .A(n264), .Z(n13) );
  INV_X1 U671 ( .A(n20), .ZN(n17) );
  INV_X1 U672 ( .A(n12), .ZN(n18) );
  INV_X1 U673 ( .A(n12), .ZN(n19) );
  INV_X1 U674 ( .A(n12), .ZN(n20) );
  INV_X1 U675 ( .A(n13), .ZN(n21) );
  CLKBUF_X1 U676 ( .A(n263), .Z(n22) );
  CLKBUF_X1 U677 ( .A(n263), .Z(n23) );
  INV_X1 U678 ( .A(n22), .ZN(n28) );
  INV_X1 U679 ( .A(n23), .ZN(n29) );
  INV_X1 U680 ( .A(n23), .ZN(n30) );
  INV_X1 U681 ( .A(n263), .ZN(n31) );
endmodule


module PG_net_0 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_30 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_29 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_28 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_27 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_26 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_25 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_24 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_23 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_22 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_21 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_20 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_19 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_18 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_17 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_16 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_15 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_14 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_13 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_12 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_11 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_10 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_9 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_8 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_7 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_6 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_5 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_4 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_3 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_2 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_1 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module Gblock_0 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n2) );
endmodule


module Gblock_8 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_7 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_6 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_5 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_4 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_3 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_2 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_1 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module PGblock_0 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n2) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_26 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_25 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_24 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_23 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_22 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_21 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_20 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_19 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_18 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_17 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_16 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_15 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_14 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_13 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_12 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_11 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_10 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_9 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_8 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_7 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_6 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_5 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_4 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_3 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_2 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_1 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module carry_generator_NBIT32_NBIT_PER_BLOCK4 ( A, B, Cin, Co );
  input [32:1] A;
  input [32:1] B;
  output [7:0] Co;
  input Cin;
  wire   \G[16][16] , \G[16][15] , \G[16][13] , \G[16][9] , \G[15][15] ,
         \G[14][14] , \G[14][13] , \G[13][13] , \G[12][12] , \G[12][11] ,
         \G[12][9] , \G[11][11] , \G[10][10] , \G[10][9] , \G[9][9] ,
         \G[8][8] , \G[8][7] , \G[8][5] , \G[7][7] , \G[6][6] , \G[6][5] ,
         \G[5][5] , \G[4][4] , \G[4][3] , \G[3][3] , \G[2][2] , \G[2][1] ,
         \G[1][1] , \P[16][16] , \P[16][15] , \P[16][13] , \P[16][9] ,
         \P[15][15] , \P[14][14] , \P[14][13] , \P[13][13] , \P[12][12] ,
         \P[12][11] , \P[12][9] , \P[11][11] , \P[10][10] , \P[10][9] ,
         \P[9][9] , \P[8][8] , \P[8][7] , \P[8][5] , \P[7][7] , \P[6][6] ,
         \P[6][5] , \P[5][5] , \P[4][4] , \P[4][3] , \P[3][3] , \P[2][2] ,
         \G[32][32] , \G[32][31] , \G[32][29] , \G[32][25] , \G[32][17] ,
         \G[31][31] , \G[30][30] , \G[30][29] , \G[29][29] , \G[28][28] ,
         \G[28][27] , \G[28][25] , \G[28][17] , \G[27][27] , \G[26][26] ,
         \G[26][25] , \G[25][25] , \G[24][24] , \G[24][23] , \G[24][21] ,
         \G[24][17] , \G[23][23] , \G[22][22] , \G[22][21] , \G[21][21] ,
         \G[20][20] , \G[20][19] , \G[20][17] , \G[19][19] , \G[18][18] ,
         \G[18][17] , \G[17][17] , \P[32][32] , \P[32][31] , \P[32][29] ,
         \P[32][25] , \P[32][17] , \P[31][31] , \P[30][30] , \P[30][29] ,
         \P[29][29] , \P[28][28] , \P[28][27] , \P[28][25] , \P[28][17] ,
         \P[27][27] , \P[26][26] , \P[26][25] , \P[25][25] , \P[24][24] ,
         \P[24][23] , \P[24][21] , \P[24][17] , \P[23][23] , \P[22][22] ,
         \P[22][21] , \P[21][21] , \P[20][20] , \P[20][19] , \P[20][17] ,
         \P[19][19] , \P[18][18] , \P[18][17] , \P[17][17] , n3, n1, n2;

  PG_net_0 PGnetblock_2 ( .a(A[2]), .b(B[2]), .p(\P[2][2] ), .g(\G[2][2] ) );
  PG_net_30 PGnetblock_3 ( .a(A[3]), .b(B[3]), .p(\P[3][3] ), .g(\G[3][3] ) );
  PG_net_29 PGnetblock_4 ( .a(A[4]), .b(B[4]), .p(\P[4][4] ), .g(\G[4][4] ) );
  PG_net_28 PGnetblock_5 ( .a(A[5]), .b(B[5]), .p(\P[5][5] ), .g(\G[5][5] ) );
  PG_net_27 PGnetblock_6 ( .a(A[6]), .b(B[6]), .p(\P[6][6] ), .g(\G[6][6] ) );
  PG_net_26 PGnetblock_7 ( .a(A[7]), .b(B[7]), .p(\P[7][7] ), .g(\G[7][7] ) );
  PG_net_25 PGnetblock_8 ( .a(A[8]), .b(B[8]), .p(\P[8][8] ), .g(\G[8][8] ) );
  PG_net_24 PGnetblock_9 ( .a(A[9]), .b(B[9]), .p(\P[9][9] ), .g(\G[9][9] ) );
  PG_net_23 PGnetblock_10 ( .a(A[10]), .b(B[10]), .p(\P[10][10] ), .g(
        \G[10][10] ) );
  PG_net_22 PGnetblock_11 ( .a(A[11]), .b(B[11]), .p(\P[11][11] ), .g(
        \G[11][11] ) );
  PG_net_21 PGnetblock_12 ( .a(A[12]), .b(B[12]), .p(\P[12][12] ), .g(
        \G[12][12] ) );
  PG_net_20 PGnetblock_13 ( .a(A[13]), .b(B[13]), .p(\P[13][13] ), .g(
        \G[13][13] ) );
  PG_net_19 PGnetblock_14 ( .a(A[14]), .b(B[14]), .p(\P[14][14] ), .g(
        \G[14][14] ) );
  PG_net_18 PGnetblock_15 ( .a(A[15]), .b(B[15]), .p(\P[15][15] ), .g(
        \G[15][15] ) );
  PG_net_17 PGnetblock_16 ( .a(A[16]), .b(B[16]), .p(\P[16][16] ), .g(
        \G[16][16] ) );
  PG_net_16 PGnetblock_17 ( .a(A[17]), .b(B[17]), .p(\P[17][17] ), .g(
        \G[17][17] ) );
  PG_net_15 PGnetblock_18 ( .a(A[18]), .b(B[18]), .p(\P[18][18] ), .g(
        \G[18][18] ) );
  PG_net_14 PGnetblock_19 ( .a(A[19]), .b(B[19]), .p(\P[19][19] ), .g(
        \G[19][19] ) );
  PG_net_13 PGnetblock_20 ( .a(A[20]), .b(B[20]), .p(\P[20][20] ), .g(
        \G[20][20] ) );
  PG_net_12 PGnetblock_21 ( .a(A[21]), .b(B[21]), .p(\P[21][21] ), .g(
        \G[21][21] ) );
  PG_net_11 PGnetblock_22 ( .a(A[22]), .b(B[22]), .p(\P[22][22] ), .g(
        \G[22][22] ) );
  PG_net_10 PGnetblock_23 ( .a(A[23]), .b(B[23]), .p(\P[23][23] ), .g(
        \G[23][23] ) );
  PG_net_9 PGnetblock_24 ( .a(A[24]), .b(B[24]), .p(\P[24][24] ), .g(
        \G[24][24] ) );
  PG_net_8 PGnetblock_25 ( .a(A[25]), .b(B[25]), .p(\P[25][25] ), .g(
        \G[25][25] ) );
  PG_net_7 PGnetblock_26 ( .a(A[26]), .b(B[26]), .p(\P[26][26] ), .g(
        \G[26][26] ) );
  PG_net_6 PGnetblock_27 ( .a(A[27]), .b(B[27]), .p(\P[27][27] ), .g(
        \G[27][27] ) );
  PG_net_5 PGnetblock_28 ( .a(A[28]), .b(B[28]), .p(\P[28][28] ), .g(
        \G[28][28] ) );
  PG_net_4 PGnetblock_29 ( .a(A[29]), .b(B[29]), .p(\P[29][29] ), .g(
        \G[29][29] ) );
  PG_net_3 PGnetblock_30 ( .a(A[30]), .b(B[30]), .p(\P[30][30] ), .g(
        \G[30][30] ) );
  PG_net_2 PGnetblock_31 ( .a(A[31]), .b(B[31]), .p(\P[31][31] ), .g(
        \G[31][31] ) );
  PG_net_1 PGnetblock_32 ( .a(A[32]), .b(B[32]), .p(\P[32][32] ), .g(
        \G[32][32] ) );
  Gblock_0 GB_low_1_2 ( .Pik(\P[2][2] ), .Gik(\G[2][2] ), .Gk_1j(\G[1][1] ), 
        .Gij(\G[2][1] ) );
  Gblock_8 GB_low_2_4 ( .Pik(\P[4][3] ), .Gik(\G[4][3] ), .Gk_1j(\G[2][1] ), 
        .Gij(Co[0]) );
  Gblock_7 GB_low_3_8 ( .Pik(\P[8][5] ), .Gik(\G[8][5] ), .Gk_1j(Co[0]), .Gij(
        Co[1]) );
  Gblock_6 GB_high_4_16_0 ( .Pik(\P[16][9] ), .Gik(\G[16][9] ), .Gk_1j(Co[1]), 
        .Gij(Co[3]) );
  Gblock_5 GB_high_4_16_1 ( .Pik(\P[12][9] ), .Gik(\G[12][9] ), .Gk_1j(Co[1]), 
        .Gij(Co[2]) );
  Gblock_4 GB_high_5_32_0 ( .Pik(\P[32][17] ), .Gik(\G[32][17] ), .Gk_1j(Co[3]), .Gij(Co[7]) );
  Gblock_3 GB_high_5_32_1 ( .Pik(\P[28][17] ), .Gik(\G[28][17] ), .Gk_1j(Co[3]), .Gij(Co[6]) );
  Gblock_2 GB_high_5_32_2 ( .Pik(\P[24][17] ), .Gik(\G[24][17] ), .Gk_1j(Co[3]), .Gij(Co[5]) );
  Gblock_1 GB_high_5_32_3 ( .Pik(\P[20][17] ), .Gik(\G[20][17] ), .Gk_1j(Co[3]), .Gij(Co[4]) );
  PGblock_0 PGB_low_1_4 ( .Pik(\P[4][4] ), .Gik(\G[4][4] ), .Pk_1j(\P[3][3] ), 
        .Gk_1j(\G[3][3] ), .Pij(\P[4][3] ), .Gij(\G[4][3] ) );
  PGblock_26 PGB_low_1_6 ( .Pik(\P[6][6] ), .Gik(\G[6][6] ), .Pk_1j(\P[5][5] ), 
        .Gk_1j(\G[5][5] ), .Pij(\P[6][5] ), .Gij(\G[6][5] ) );
  PGblock_25 PGB_low_1_8 ( .Pik(\P[8][8] ), .Gik(\G[8][8] ), .Pk_1j(\P[7][7] ), 
        .Gk_1j(\G[7][7] ), .Pij(\P[8][7] ), .Gij(\G[8][7] ) );
  PGblock_24 PGB_low_1_10 ( .Pik(\P[10][10] ), .Gik(\G[10][10] ), .Pk_1j(
        \P[9][9] ), .Gk_1j(\G[9][9] ), .Pij(\P[10][9] ), .Gij(\G[10][9] ) );
  PGblock_23 PGB_low_1_12 ( .Pik(\P[12][12] ), .Gik(\G[12][12] ), .Pk_1j(
        \P[11][11] ), .Gk_1j(\G[11][11] ), .Pij(\P[12][11] ), .Gij(\G[12][11] ) );
  PGblock_22 PGB_low_1_14 ( .Pik(\P[14][14] ), .Gik(\G[14][14] ), .Pk_1j(
        \P[13][13] ), .Gk_1j(\G[13][13] ), .Pij(\P[14][13] ), .Gij(\G[14][13] ) );
  PGblock_21 PGB_low_1_16 ( .Pik(\P[16][16] ), .Gik(\G[16][16] ), .Pk_1j(
        \P[15][15] ), .Gk_1j(\G[15][15] ), .Pij(\P[16][15] ), .Gij(\G[16][15] ) );
  PGblock_20 PGB_low_1_18 ( .Pik(\P[18][18] ), .Gik(\G[18][18] ), .Pk_1j(
        \P[17][17] ), .Gk_1j(\G[17][17] ), .Pij(\P[18][17] ), .Gij(\G[18][17] ) );
  PGblock_19 PGB_low_1_20 ( .Pik(\P[20][20] ), .Gik(\G[20][20] ), .Pk_1j(
        \P[19][19] ), .Gk_1j(\G[19][19] ), .Pij(\P[20][19] ), .Gij(\G[20][19] ) );
  PGblock_18 PGB_low_1_22 ( .Pik(\P[22][22] ), .Gik(\G[22][22] ), .Pk_1j(
        \P[21][21] ), .Gk_1j(\G[21][21] ), .Pij(\P[22][21] ), .Gij(\G[22][21] ) );
  PGblock_17 PGB_low_1_24 ( .Pik(\P[24][24] ), .Gik(\G[24][24] ), .Pk_1j(
        \P[23][23] ), .Gk_1j(\G[23][23] ), .Pij(\P[24][23] ), .Gij(\G[24][23] ) );
  PGblock_16 PGB_low_1_26 ( .Pik(\P[26][26] ), .Gik(\G[26][26] ), .Pk_1j(
        \P[25][25] ), .Gk_1j(\G[25][25] ), .Pij(\P[26][25] ), .Gij(\G[26][25] ) );
  PGblock_15 PGB_low_1_28 ( .Pik(\P[28][28] ), .Gik(\G[28][28] ), .Pk_1j(
        \P[27][27] ), .Gk_1j(\G[27][27] ), .Pij(\P[28][27] ), .Gij(\G[28][27] ) );
  PGblock_14 PGB_low_1_30 ( .Pik(\P[30][30] ), .Gik(\G[30][30] ), .Pk_1j(
        \P[29][29] ), .Gk_1j(\G[29][29] ), .Pij(\P[30][29] ), .Gij(\G[30][29] ) );
  PGblock_13 PGB_low_1_32 ( .Pik(\P[32][32] ), .Gik(\G[32][32] ), .Pk_1j(
        \P[31][31] ), .Gk_1j(\G[31][31] ), .Pij(\P[32][31] ), .Gij(\G[32][31] ) );
  PGblock_12 PGB_low_2_8 ( .Pik(\P[8][7] ), .Gik(\G[8][7] ), .Pk_1j(\P[6][5] ), 
        .Gk_1j(\G[6][5] ), .Pij(\P[8][5] ), .Gij(\G[8][5] ) );
  PGblock_11 PGB_low_2_12 ( .Pik(\P[12][11] ), .Gik(\G[12][11] ), .Pk_1j(
        \P[10][9] ), .Gk_1j(\G[10][9] ), .Pij(\P[12][9] ), .Gij(\G[12][9] ) );
  PGblock_10 PGB_low_2_16 ( .Pik(\P[16][15] ), .Gik(\G[16][15] ), .Pk_1j(
        \P[14][13] ), .Gk_1j(\G[14][13] ), .Pij(\P[16][13] ), .Gij(\G[16][13] ) );
  PGblock_9 PGB_low_2_20 ( .Pik(\P[20][19] ), .Gik(\G[20][19] ), .Pk_1j(
        \P[18][17] ), .Gk_1j(\G[18][17] ), .Pij(\P[20][17] ), .Gij(\G[20][17] ) );
  PGblock_8 PGB_low_2_24 ( .Pik(\P[24][23] ), .Gik(\G[24][23] ), .Pk_1j(
        \P[22][21] ), .Gk_1j(\G[22][21] ), .Pij(\P[24][21] ), .Gij(\G[24][21] ) );
  PGblock_7 PGB_low_2_28 ( .Pik(\P[28][27] ), .Gik(\G[28][27] ), .Pk_1j(
        \P[26][25] ), .Gk_1j(\G[26][25] ), .Pij(\P[28][25] ), .Gij(\G[28][25] ) );
  PGblock_6 PGB_low_2_32 ( .Pik(\P[32][31] ), .Gik(\G[32][31] ), .Pk_1j(
        \P[30][29] ), .Gk_1j(\G[30][29] ), .Pij(\P[32][29] ), .Gij(\G[32][29] ) );
  PGblock_5 PGB_low_3_16 ( .Pik(\P[16][13] ), .Gik(\G[16][13] ), .Pk_1j(
        \P[12][9] ), .Gk_1j(\G[12][9] ), .Pij(\P[16][9] ), .Gij(\G[16][9] ) );
  PGblock_4 PGB_low_3_24 ( .Pik(\P[24][21] ), .Gik(\G[24][21] ), .Pk_1j(
        \P[20][17] ), .Gk_1j(\G[20][17] ), .Pij(\P[24][17] ), .Gij(\G[24][17] ) );
  PGblock_3 PGB_low_3_32 ( .Pik(\P[32][29] ), .Gik(\G[32][29] ), .Pk_1j(
        \P[28][25] ), .Gk_1j(\G[28][25] ), .Pij(\P[32][25] ), .Gij(\G[32][25] ) );
  PGblock_2 PGB_high_4_32_0 ( .Pik(\P[32][25] ), .Gik(\G[32][25] ), .Pk_1j(
        \P[24][17] ), .Gk_1j(\G[24][17] ), .Pij(\P[32][17] ), .Gij(\G[32][17] ) );
  PGblock_1 PGB_high_4_32_1 ( .Pik(\P[28][25] ), .Gik(\G[28][25] ), .Pk_1j(
        \P[24][17] ), .Gk_1j(\G[24][17] ), .Pij(\P[28][17] ), .Gij(\G[28][17] ) );
  INV_X1 U1 ( .A(A[1]), .ZN(n1) );
  OAI21_X1 U2 ( .B1(n1), .B2(n2), .A(n3), .ZN(\G[1][1] ) );
  OAI21_X1 U3 ( .B1(A[1]), .B2(B[1]), .A(Cin), .ZN(n3) );
  INV_X1 U4 ( .A(B[1]), .ZN(n2) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_0 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n6, n7, n8, n9, n1;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_0 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_15 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(n7), .ZN(S[2]) );
  AOI22_X1 U4 ( .A1(Y1[2]), .A2(n1), .B1(Y2[2]), .B2(C_i), .ZN(n7) );
  INV_X1 U5 ( .A(n6), .ZN(S[3]) );
  AOI22_X1 U6 ( .A1(Y1[3]), .A2(n1), .B1(Y2[3]), .B2(C_i), .ZN(n6) );
  INV_X1 U7 ( .A(n9), .ZN(S[0]) );
  INV_X1 U8 ( .A(n8), .ZN(S[1]) );
  AOI22_X1 U9 ( .A1(Y1[1]), .A2(n1), .B1(Y2[1]), .B2(C_i), .ZN(n8) );
  AOI22_X1 U10 ( .A1(Y1[0]), .A2(n1), .B1(Y2[0]), .B2(C_i), .ZN(n9) );
  INV_X1 U11 ( .A(C_i), .ZN(n1) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_7 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_14 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_13 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U5 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U9 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_6 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_12 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_11 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U5 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U9 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_5 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_10 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_9 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U5 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U9 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_4 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_8 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_7 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U5 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U9 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_3 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_6 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_5 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U5 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U9 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_2 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_4 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_3 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U5 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U9 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_1 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_2 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_1 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U5 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U9 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_select_basic_N4_0 CSBI_1 ( .A(A[3:0]), .B(B[3:0]), .C_i(Ci[0]), .S(
        S[3:0]) );
  carry_select_basic_N4_7 CSBI_2 ( .A(A[7:4]), .B(B[7:4]), .C_i(Ci[1]), .S(
        S[7:4]) );
  carry_select_basic_N4_6 CSBI_3 ( .A(A[11:8]), .B(B[11:8]), .C_i(Ci[2]), .S(
        S[11:8]) );
  carry_select_basic_N4_5 CSBI_4 ( .A(A[15:12]), .B(B[15:12]), .C_i(Ci[3]), 
        .S(S[15:12]) );
  carry_select_basic_N4_4 CSBI_5 ( .A(A[19:16]), .B(B[19:16]), .C_i(Ci[4]), 
        .S(S[19:16]) );
  carry_select_basic_N4_3 CSBI_6 ( .A(A[23:20]), .B(B[23:20]), .C_i(Ci[5]), 
        .S(S[23:20]) );
  carry_select_basic_N4_2 CSBI_7 ( .A(A[27:24]), .B(B[27:24]), .C_i(Ci[6]), 
        .S(S[27:24]) );
  carry_select_basic_N4_1 CSBI_8 ( .A(A[31:28]), .B(B[31:28]), .C_i(Ci[7]), 
        .S(S[31:28]) );
endmodule


module P4Adder_NBIT32 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;

  wire   [7:1] Csum;

  carry_generator_NBIT32_NBIT_PER_BLOCK4 Carrygen0 ( .A(A), .B(B), .Cin(Cin), 
        .Co({Cout, Csum}) );
  SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 Sumgen0 ( .A(A), .B(B), .Ci({Csum, 
        Cin}), .S(S) );
endmodule


module mux41_NBIT32_1 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149;

  BUF_X1 U1 ( .A(n145), .Z(n72) );
  BUF_X1 U2 ( .A(n145), .Z(n73) );
  BUF_X1 U3 ( .A(n147), .Z(n78) );
  BUF_X1 U4 ( .A(n147), .Z(n79) );
  BUF_X1 U5 ( .A(n144), .Z(n1) );
  BUF_X1 U6 ( .A(n144), .Z(n70) );
  BUF_X1 U7 ( .A(n146), .Z(n75) );
  BUF_X1 U8 ( .A(n146), .Z(n76) );
  BUF_X1 U9 ( .A(n145), .Z(n74) );
  BUF_X1 U10 ( .A(n147), .Z(n80) );
  BUF_X1 U11 ( .A(n144), .Z(n71) );
  BUF_X1 U12 ( .A(n146), .Z(n77) );
  NOR2_X1 U13 ( .A1(S[0]), .A2(S[1]), .ZN(n144) );
  NOR2_X1 U14 ( .A1(n81), .A2(S[1]), .ZN(n145) );
  AND2_X1 U15 ( .A1(S[1]), .A2(S[0]), .ZN(n147) );
  AND2_X1 U16 ( .A1(S[1]), .A2(n81), .ZN(n146) );
  INV_X1 U17 ( .A(S[0]), .ZN(n81) );
  NAND2_X1 U18 ( .A1(n83), .A2(n82), .ZN(Z[0]) );
  AOI22_X1 U19 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n83) );
  AOI22_X1 U20 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n82) );
  NAND2_X1 U21 ( .A1(n131), .A2(n130), .ZN(Z[31]) );
  AOI22_X1 U22 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n130) );
  AOI22_X1 U23 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n131) );
  NAND2_X1 U24 ( .A1(n141), .A2(n140), .ZN(Z[7]) );
  AOI22_X1 U25 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n140) );
  AOI22_X1 U26 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n141) );
  NAND2_X1 U27 ( .A1(n143), .A2(n142), .ZN(Z[8]) );
  AOI22_X1 U28 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n142) );
  AOI22_X1 U29 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n143) );
  NAND2_X1 U30 ( .A1(n149), .A2(n148), .ZN(Z[9]) );
  AOI22_X1 U31 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n148) );
  AOI22_X1 U32 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n149) );
  NAND2_X1 U33 ( .A1(n89), .A2(n88), .ZN(Z[12]) );
  AOI22_X1 U34 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n88) );
  AOI22_X1 U35 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n89) );
  NAND2_X1 U36 ( .A1(n91), .A2(n90), .ZN(Z[13]) );
  AOI22_X1 U37 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n90) );
  AOI22_X1 U38 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n91) );
  NAND2_X1 U39 ( .A1(n93), .A2(n92), .ZN(Z[14]) );
  AOI22_X1 U40 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n92) );
  AOI22_X1 U41 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n93) );
  NAND2_X1 U42 ( .A1(n99), .A2(n98), .ZN(Z[17]) );
  AOI22_X1 U43 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n98) );
  AOI22_X1 U44 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n99) );
  NAND2_X1 U45 ( .A1(n95), .A2(n94), .ZN(Z[15]) );
  AOI22_X1 U46 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n94) );
  AOI22_X1 U47 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n95) );
  NAND2_X1 U48 ( .A1(n101), .A2(n100), .ZN(Z[18]) );
  AOI22_X1 U49 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n100) );
  AOI22_X1 U50 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n101) );
  NAND2_X1 U51 ( .A1(n97), .A2(n96), .ZN(Z[16]) );
  AOI22_X1 U52 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n96) );
  AOI22_X1 U53 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n97) );
  NAND2_X1 U54 ( .A1(n103), .A2(n102), .ZN(Z[19]) );
  AOI22_X1 U55 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n102) );
  AOI22_X1 U56 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n103) );
  NAND2_X1 U57 ( .A1(n107), .A2(n106), .ZN(Z[20]) );
  AOI22_X1 U58 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n106) );
  AOI22_X1 U59 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n107) );
  NAND2_X1 U60 ( .A1(n109), .A2(n108), .ZN(Z[21]) );
  AOI22_X1 U61 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n108) );
  AOI22_X1 U62 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n109) );
  NAND2_X1 U63 ( .A1(n111), .A2(n110), .ZN(Z[22]) );
  AOI22_X1 U64 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n110) );
  AOI22_X1 U65 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n111) );
  NAND2_X1 U66 ( .A1(n113), .A2(n112), .ZN(Z[23]) );
  AOI22_X1 U67 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n112) );
  AOI22_X1 U68 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n113) );
  NAND2_X1 U69 ( .A1(n115), .A2(n114), .ZN(Z[24]) );
  AOI22_X1 U70 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n114) );
  AOI22_X1 U71 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n115) );
  NAND2_X1 U72 ( .A1(n117), .A2(n116), .ZN(Z[25]) );
  AOI22_X1 U73 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n116) );
  AOI22_X1 U74 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n117) );
  NAND2_X1 U75 ( .A1(n139), .A2(n138), .ZN(Z[6]) );
  AOI22_X1 U76 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n138) );
  AOI22_X1 U77 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n139) );
  NAND2_X1 U78 ( .A1(n85), .A2(n84), .ZN(Z[10]) );
  AOI22_X1 U79 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n84) );
  AOI22_X1 U80 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n85) );
  NAND2_X1 U81 ( .A1(n87), .A2(n86), .ZN(Z[11]) );
  AOI22_X1 U82 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n86) );
  AOI22_X1 U83 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n87) );
  NAND2_X1 U84 ( .A1(n119), .A2(n118), .ZN(Z[26]) );
  AOI22_X1 U85 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n118) );
  AOI22_X1 U86 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n119) );
  NAND2_X1 U87 ( .A1(n121), .A2(n120), .ZN(Z[27]) );
  AOI22_X1 U88 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n120) );
  AOI22_X1 U89 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n121) );
  NAND2_X1 U90 ( .A1(n137), .A2(n136), .ZN(Z[5]) );
  AOI22_X1 U91 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n136) );
  AOI22_X1 U92 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n137) );
  NAND2_X1 U93 ( .A1(n123), .A2(n122), .ZN(Z[28]) );
  AOI22_X1 U94 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n122) );
  AOI22_X1 U95 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n123) );
  NAND2_X1 U96 ( .A1(n125), .A2(n124), .ZN(Z[29]) );
  AOI22_X1 U97 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n124) );
  AOI22_X1 U98 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n125) );
  NAND2_X1 U99 ( .A1(n129), .A2(n128), .ZN(Z[30]) );
  AOI22_X1 U100 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n128) );
  AOI22_X1 U101 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n129) );
  NAND2_X1 U102 ( .A1(n127), .A2(n126), .ZN(Z[2]) );
  AOI22_X1 U103 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n126) );
  AOI22_X1 U104 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n127) );
  NAND2_X1 U105 ( .A1(n105), .A2(n104), .ZN(Z[1]) );
  AOI22_X1 U106 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n104) );
  AOI22_X1 U107 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n105) );
  NAND2_X1 U108 ( .A1(n133), .A2(n132), .ZN(Z[3]) );
  AOI22_X1 U109 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n132) );
  AOI22_X1 U110 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n133) );
  NAND2_X1 U111 ( .A1(n135), .A2(n134), .ZN(Z[4]) );
  AOI22_X1 U112 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n134) );
  AOI22_X1 U113 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n135) );
endmodule


module mux21_NBIT32_1 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n11) );
  BUF_X1 U6 ( .A(n2), .Z(n9) );
  BUF_X1 U7 ( .A(n1), .Z(n8) );
  BUF_X1 U8 ( .A(n2), .Z(n10) );
  BUF_X1 U9 ( .A(n1), .Z(n7) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(S), .Z(n3) );
  BUF_X1 U13 ( .A(S), .Z(n2) );
  BUF_X1 U14 ( .A(S), .Z(n1) );
  INV_X1 U15 ( .A(n79), .ZN(Z[0]) );
  AOI22_X1 U16 ( .A1(A[0]), .A2(n4), .B1(B[0]), .B2(n13), .ZN(n79) );
  INV_X1 U17 ( .A(n90), .ZN(Z[1]) );
  AOI22_X1 U18 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(n10), .ZN(n90) );
  INV_X1 U19 ( .A(n101), .ZN(Z[2]) );
  AOI22_X1 U20 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n7), .ZN(n101) );
  INV_X1 U21 ( .A(n104), .ZN(Z[3]) );
  AOI22_X1 U22 ( .A1(A[3]), .A2(n4), .B1(B[3]), .B2(n7), .ZN(n104) );
  INV_X1 U23 ( .A(n105), .ZN(Z[4]) );
  AOI22_X1 U24 ( .A1(A[4]), .A2(n5), .B1(B[4]), .B2(n7), .ZN(n105) );
  INV_X1 U25 ( .A(n106), .ZN(Z[5]) );
  AOI22_X1 U26 ( .A1(A[5]), .A2(n4), .B1(B[5]), .B2(n6), .ZN(n106) );
  INV_X1 U27 ( .A(n107), .ZN(Z[6]) );
  AOI22_X1 U28 ( .A1(A[6]), .A2(n5), .B1(B[6]), .B2(n6), .ZN(n107) );
  INV_X1 U29 ( .A(n108), .ZN(Z[7]) );
  AOI22_X1 U30 ( .A1(A[7]), .A2(n4), .B1(B[7]), .B2(n6), .ZN(n108) );
  INV_X1 U31 ( .A(n109), .ZN(Z[8]) );
  AOI22_X1 U32 ( .A1(A[8]), .A2(n5), .B1(B[8]), .B2(n6), .ZN(n109) );
  INV_X1 U33 ( .A(n110), .ZN(Z[9]) );
  AOI22_X1 U34 ( .A1(A[9]), .A2(n4), .B1(n13), .B2(B[9]), .ZN(n110) );
  INV_X1 U35 ( .A(n80), .ZN(Z[10]) );
  AOI22_X1 U36 ( .A1(A[10]), .A2(n4), .B1(B[10]), .B2(n13), .ZN(n80) );
  INV_X1 U37 ( .A(n81), .ZN(Z[11]) );
  AOI22_X1 U38 ( .A1(A[11]), .A2(n4), .B1(B[11]), .B2(n13), .ZN(n81) );
  INV_X1 U39 ( .A(n82), .ZN(Z[12]) );
  AOI22_X1 U40 ( .A1(A[12]), .A2(n4), .B1(B[12]), .B2(n12), .ZN(n82) );
  INV_X1 U41 ( .A(n83), .ZN(Z[13]) );
  AOI22_X1 U42 ( .A1(A[13]), .A2(n4), .B1(B[13]), .B2(n12), .ZN(n83) );
  INV_X1 U43 ( .A(n84), .ZN(Z[14]) );
  AOI22_X1 U44 ( .A1(A[14]), .A2(n4), .B1(B[14]), .B2(n12), .ZN(n84) );
  INV_X1 U45 ( .A(n85), .ZN(Z[15]) );
  AOI22_X1 U46 ( .A1(A[15]), .A2(n4), .B1(B[15]), .B2(n12), .ZN(n85) );
  INV_X1 U47 ( .A(n86), .ZN(Z[16]) );
  AOI22_X1 U48 ( .A1(A[16]), .A2(n4), .B1(B[16]), .B2(n11), .ZN(n86) );
  INV_X1 U49 ( .A(n87), .ZN(Z[17]) );
  AOI22_X1 U50 ( .A1(A[17]), .A2(n4), .B1(B[17]), .B2(n11), .ZN(n87) );
  INV_X1 U51 ( .A(n88), .ZN(Z[18]) );
  AOI22_X1 U52 ( .A1(A[18]), .A2(n4), .B1(B[18]), .B2(n11), .ZN(n88) );
  INV_X1 U53 ( .A(n89), .ZN(Z[19]) );
  AOI22_X1 U54 ( .A1(A[19]), .A2(n4), .B1(B[19]), .B2(n11), .ZN(n89) );
  INV_X1 U55 ( .A(n91), .ZN(Z[20]) );
  AOI22_X1 U56 ( .A1(A[20]), .A2(n5), .B1(B[20]), .B2(n10), .ZN(n91) );
  INV_X1 U57 ( .A(n92), .ZN(Z[21]) );
  AOI22_X1 U58 ( .A1(A[21]), .A2(n5), .B1(B[21]), .B2(n10), .ZN(n92) );
  INV_X1 U59 ( .A(n93), .ZN(Z[22]) );
  AOI22_X1 U60 ( .A1(A[22]), .A2(n5), .B1(B[22]), .B2(n9), .ZN(n93) );
  INV_X1 U61 ( .A(n94), .ZN(Z[23]) );
  AOI22_X1 U62 ( .A1(A[23]), .A2(n5), .B1(B[23]), .B2(n9), .ZN(n94) );
  INV_X1 U63 ( .A(n95), .ZN(Z[24]) );
  AOI22_X1 U64 ( .A1(A[24]), .A2(n5), .B1(B[24]), .B2(n9), .ZN(n95) );
  INV_X1 U65 ( .A(n96), .ZN(Z[25]) );
  AOI22_X1 U66 ( .A1(A[25]), .A2(n5), .B1(B[25]), .B2(n9), .ZN(n96) );
  INV_X1 U67 ( .A(n97), .ZN(Z[26]) );
  AOI22_X1 U68 ( .A1(A[26]), .A2(n5), .B1(B[26]), .B2(n8), .ZN(n97) );
  INV_X1 U69 ( .A(n98), .ZN(Z[27]) );
  AOI22_X1 U70 ( .A1(A[27]), .A2(n5), .B1(B[27]), .B2(n8), .ZN(n98) );
  INV_X1 U71 ( .A(n99), .ZN(Z[28]) );
  AOI22_X1 U72 ( .A1(A[28]), .A2(n5), .B1(B[28]), .B2(n8), .ZN(n99) );
  INV_X1 U73 ( .A(n100), .ZN(Z[29]) );
  AOI22_X1 U74 ( .A1(A[29]), .A2(n5), .B1(B[29]), .B2(n8), .ZN(n100) );
  INV_X1 U75 ( .A(n102), .ZN(Z[30]) );
  AOI22_X1 U76 ( .A1(A[30]), .A2(n5), .B1(B[30]), .B2(n10), .ZN(n102) );
  INV_X1 U77 ( .A(n103), .ZN(Z[31]) );
  AOI22_X1 U78 ( .A1(A[31]), .A2(n5), .B1(B[31]), .B2(n7), .ZN(n103) );
endmodule


module ALU_NBIT32 ( OP1, OP2, .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , 
        \ALU_OPC[1] , \ALU_OPC[0] }), ALU_RES );
  input [31:0] OP1;
  input [31:0] OP2;
  output [31:0] ALU_RES;
  input \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] ;
  wire   select_zero_sig, LOGIC_ARITH, \OPSel[0] , n78, n79, n80, n81, n82,
         n83, n84, n85, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n86, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186;
  wire   [3:0] ALU_OPC;
  wire   [1:0] select_type_sig;
  wire   [31:0] A_SHF;
  wire   [31:0] B_SHF;
  wire   [31:0] A_ADD;
  wire   [31:0] B_ADD;
  wire   [31:0] LOGIC_RES;
  wire   [31:0] COMP_RES;
  wire   [31:0] SHIFT_RES;
  wire   [31:0] ADD_SUB_RES;
  wire   [31:0] sig_intraMux;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  NOR2_X2 U177 ( .A1(n13), .A2(n55), .ZN(A_SHF[31]) );
  NAND3_X1 U317 ( .A1(n185), .A2(n184), .A3(n186), .ZN(n79) );
  NAND3_X1 U318 ( .A1(n84), .A2(n83), .A3(n87), .ZN(\OPSel[0] ) );
  NAND3_X1 U319 ( .A1(ALU_OPC[3]), .A2(n186), .A3(n88), .ZN(n87) );
  NAND3_X1 U320 ( .A1(ALU_OPC[3]), .A2(n186), .A3(n89), .ZN(n83) );
  NAND3_X1 U321 ( .A1(ALU_OPC[3]), .A2(ALU_OPC[0]), .A3(n89), .ZN(n84) );
  NAND3_X1 U322 ( .A1(ALU_OPC[2]), .A2(ALU_OPC[1]), .A3(n155), .ZN(n157) );
  NAND3_X1 U323 ( .A1(ALU_OPC[2]), .A2(ALU_OPC[1]), .A3(n154), .ZN(n85) );
  NAND3_X1 U324 ( .A1(n185), .A2(n184), .A3(n155), .ZN(n156) );
  comparator_NBIT32 Comp ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .OPSel({n183, n182, 
        \OPSel[0] }), .RES({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, COMP_RES[0]}) );
  shifter_NBIT32 Shift ( .A(A_SHF), .B(B_SHF), .LOGIC_ARITH(LOGIC_ARITH), 
        .LEFT_RIGHT(n180), .RES(SHIFT_RES) );
  P4Adder_NBIT32 Add_Sub_unit ( .A(A_ADD), .B(B_ADD), .Cin(n1), .S(ADD_SUB_RES) );
  mux41_NBIT32_1 Res_mux ( .A(ADD_SUB_RES), .B(LOGIC_RES), .C(SHIFT_RES), .D({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, COMP_RES[0]}), .S(
        select_type_sig), .Z(sig_intraMux) );
  mux21_NBIT32_1 Zeros_mux ( .A(sig_intraMux), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .S(select_zero_sig), .Z(ALU_RES) );
  NOR2_X1 U2 ( .A1(n13), .A2(n58), .ZN(A_SHF[5]) );
  NOR2_X1 U3 ( .A1(n13), .A2(n59), .ZN(A_SHF[6]) );
  BUF_X1 U4 ( .A(n158), .Z(n23) );
  BUF_X1 U5 ( .A(n158), .Z(n24) );
  BUF_X1 U6 ( .A(n158), .Z(n25) );
  BUF_X1 U7 ( .A(n177), .Z(n5) );
  BUF_X1 U8 ( .A(n177), .Z(n6) );
  BUF_X1 U9 ( .A(n177), .Z(n7) );
  BUF_X1 U10 ( .A(n177), .Z(n9) );
  BUF_X1 U11 ( .A(n177), .Z(n8) );
  BUF_X1 U12 ( .A(n179), .Z(n17) );
  BUF_X1 U13 ( .A(n179), .Z(n18) );
  BUF_X1 U14 ( .A(n179), .Z(n21) );
  BUF_X1 U15 ( .A(n179), .Z(n20) );
  BUF_X1 U16 ( .A(n179), .Z(n19) );
  BUF_X1 U17 ( .A(n176), .Z(n2) );
  BUF_X1 U18 ( .A(n176), .Z(n3) );
  BUF_X1 U19 ( .A(n176), .Z(n4) );
  AND2_X1 U20 ( .A1(n28), .A2(n29), .ZN(n158) );
  NOR2_X1 U21 ( .A1(n15), .A2(n168), .ZN(B_SHF[3]) );
  NOR2_X1 U22 ( .A1(n12), .A2(n50), .ZN(A_SHF[27]) );
  NOR2_X1 U23 ( .A1(n12), .A2(n49), .ZN(A_SHF[26]) );
  NOR2_X1 U24 ( .A1(n13), .A2(n64), .ZN(B_SHF[10]) );
  NOR2_X1 U25 ( .A1(n16), .A2(n174), .ZN(B_SHF[9]) );
  NOR2_X1 U26 ( .A1(n16), .A2(n173), .ZN(B_SHF[8]) );
  NOR2_X1 U27 ( .A1(n11), .A2(n39), .ZN(A_SHF[17]) );
  NOR2_X1 U28 ( .A1(n13), .A2(n60), .ZN(A_SHF[7]) );
  NOR2_X1 U29 ( .A1(n15), .A2(n165), .ZN(B_SHF[2]) );
  NOR2_X1 U30 ( .A1(n11), .A2(n40), .ZN(A_SHF[18]) );
  NOR2_X1 U31 ( .A1(n12), .A2(n48), .ZN(A_SHF[25]) );
  NOR2_X1 U32 ( .A1(n13), .A2(n57), .ZN(A_SHF[4]) );
  NOR2_X1 U33 ( .A1(n12), .A2(n51), .ZN(A_SHF[28]) );
  NOR2_X1 U34 ( .A1(n15), .A2(n170), .ZN(B_SHF[5]) );
  NOR2_X1 U35 ( .A1(n16), .A2(n172), .ZN(B_SHF[7]) );
  NOR2_X1 U36 ( .A1(n16), .A2(n171), .ZN(B_SHF[6]) );
  NOR2_X1 U37 ( .A1(n23), .A2(n31), .ZN(A_ADD[0]) );
  NOR2_X1 U38 ( .A1(n13), .A2(n61), .ZN(A_SHF[8]) );
  NOR2_X1 U39 ( .A1(n12), .A2(n53), .ZN(A_SHF[2]) );
  NOR2_X1 U40 ( .A1(n25), .A2(n57), .ZN(A_ADD[4]) );
  NOR2_X1 U41 ( .A1(n25), .A2(n58), .ZN(A_ADD[5]) );
  NOR2_X1 U42 ( .A1(n25), .A2(n59), .ZN(A_ADD[6]) );
  NOR2_X1 U43 ( .A1(n25), .A2(n61), .ZN(A_ADD[8]) );
  NOR2_X1 U44 ( .A1(n25), .A2(n62), .ZN(A_ADD[9]) );
  NOR2_X1 U45 ( .A1(n25), .A2(n56), .ZN(A_ADD[3]) );
  NOR2_X1 U46 ( .A1(n25), .A2(n60), .ZN(A_ADD[7]) );
  NOR2_X1 U47 ( .A1(n25), .A2(n55), .ZN(A_ADD[31]) );
  NOR2_X1 U48 ( .A1(n23), .A2(n42), .ZN(A_ADD[1]) );
  NOR2_X1 U49 ( .A1(n24), .A2(n53), .ZN(A_ADD[2]) );
  NOR2_X1 U50 ( .A1(n23), .A2(n32), .ZN(A_ADD[10]) );
  NOR2_X1 U51 ( .A1(n23), .A2(n34), .ZN(A_ADD[12]) );
  NOR2_X1 U52 ( .A1(n23), .A2(n35), .ZN(A_ADD[13]) );
  NOR2_X1 U53 ( .A1(n23), .A2(n36), .ZN(A_ADD[14]) );
  NOR2_X1 U54 ( .A1(n23), .A2(n38), .ZN(A_ADD[16]) );
  NOR2_X1 U55 ( .A1(n23), .A2(n39), .ZN(A_ADD[17]) );
  NOR2_X1 U56 ( .A1(n23), .A2(n40), .ZN(A_ADD[18]) );
  NOR2_X1 U57 ( .A1(n24), .A2(n43), .ZN(A_ADD[20]) );
  NOR2_X1 U58 ( .A1(n24), .A2(n44), .ZN(A_ADD[21]) );
  NOR2_X1 U59 ( .A1(n24), .A2(n45), .ZN(A_ADD[22]) );
  NOR2_X1 U60 ( .A1(n24), .A2(n47), .ZN(A_ADD[24]) );
  NOR2_X1 U61 ( .A1(n24), .A2(n48), .ZN(A_ADD[25]) );
  NOR2_X1 U62 ( .A1(n24), .A2(n49), .ZN(A_ADD[26]) );
  NOR2_X1 U63 ( .A1(n24), .A2(n51), .ZN(A_ADD[28]) );
  NOR2_X1 U64 ( .A1(n24), .A2(n52), .ZN(A_ADD[29]) );
  NOR2_X1 U65 ( .A1(n24), .A2(n54), .ZN(A_ADD[30]) );
  NOR2_X1 U66 ( .A1(n23), .A2(n33), .ZN(A_ADD[11]) );
  NOR2_X1 U67 ( .A1(n23), .A2(n37), .ZN(A_ADD[15]) );
  NOR2_X1 U68 ( .A1(n23), .A2(n41), .ZN(A_ADD[19]) );
  NOR2_X1 U69 ( .A1(n24), .A2(n46), .ZN(A_ADD[23]) );
  NOR2_X1 U70 ( .A1(n24), .A2(n50), .ZN(A_ADD[27]) );
  NOR2_X1 U71 ( .A1(n14), .A2(n74), .ZN(B_SHF[1]) );
  NOR2_X1 U72 ( .A1(n12), .A2(n43), .ZN(A_SHF[20]) );
  NOR2_X1 U73 ( .A1(n11), .A2(n34), .ZN(A_SHF[12]) );
  NOR2_X1 U74 ( .A1(n12), .A2(n44), .ZN(A_SHF[21]) );
  NOR2_X1 U75 ( .A1(n11), .A2(n35), .ZN(A_SHF[13]) );
  NOR2_X1 U76 ( .A1(n11), .A2(n41), .ZN(A_SHF[19]) );
  NOR2_X1 U77 ( .A1(n12), .A2(n45), .ZN(A_SHF[22]) );
  NOR2_X1 U78 ( .A1(n11), .A2(n36), .ZN(A_SHF[14]) );
  NOR2_X1 U79 ( .A1(n12), .A2(n46), .ZN(A_SHF[23]) );
  NOR2_X1 U80 ( .A1(n12), .A2(n47), .ZN(A_SHF[24]) );
  NOR2_X1 U81 ( .A1(n15), .A2(n163), .ZN(B_SHF[28]) );
  NOR2_X1 U82 ( .A1(n15), .A2(n162), .ZN(B_SHF[27]) );
  NOR2_X1 U83 ( .A1(n15), .A2(n161), .ZN(B_SHF[26]) );
  NOR2_X1 U84 ( .A1(n11), .A2(n42), .ZN(A_SHF[1]) );
  NOR2_X1 U85 ( .A1(n13), .A2(n65), .ZN(B_SHF[11]) );
  NOR2_X1 U86 ( .A1(n13), .A2(n62), .ZN(A_SHF[9]) );
  NOR2_X1 U87 ( .A1(n11), .A2(n31), .ZN(A_SHF[0]) );
  NOR2_X1 U88 ( .A1(n11), .A2(n33), .ZN(A_SHF[11]) );
  NOR2_X1 U89 ( .A1(n11), .A2(n37), .ZN(A_SHF[15]) );
  NOR2_X1 U90 ( .A1(n12), .A2(n52), .ZN(A_SHF[29]) );
  NOR2_X1 U91 ( .A1(n11), .A2(n38), .ZN(A_SHF[16]) );
  NOR2_X1 U92 ( .A1(n13), .A2(n56), .ZN(A_SHF[3]) );
  NOR2_X1 U93 ( .A1(n14), .A2(n72), .ZN(B_SHF[18]) );
  BUF_X1 U94 ( .A(n178), .Z(n13) );
  BUF_X1 U95 ( .A(n178), .Z(n14) );
  BUF_X1 U96 ( .A(n178), .Z(n11) );
  BUF_X1 U97 ( .A(n178), .Z(n12) );
  BUF_X1 U98 ( .A(n178), .Z(n15) );
  NOR2_X1 U99 ( .A1(n15), .A2(n164), .ZN(B_SHF[29]) );
  NOR2_X1 U100 ( .A1(n15), .A2(n166), .ZN(B_SHF[30]) );
  NOR2_X1 U101 ( .A1(n15), .A2(n160), .ZN(B_SHF[25]) );
  NOR2_X1 U102 ( .A1(n13), .A2(n63), .ZN(B_SHF[0]) );
  NOR2_X1 U103 ( .A1(n14), .A2(n70), .ZN(B_SHF[16]) );
  NOR2_X1 U104 ( .A1(n11), .A2(n32), .ZN(A_SHF[10]) );
  NOR2_X1 U105 ( .A1(n14), .A2(n71), .ZN(B_SHF[17]) );
  NOR2_X1 U106 ( .A1(n14), .A2(n69), .ZN(B_SHF[15]) );
  BUF_X1 U107 ( .A(n156), .Z(n27) );
  BUF_X1 U108 ( .A(n156), .Z(n26) );
  NOR2_X1 U109 ( .A1(n15), .A2(n159), .ZN(B_SHF[24]) );
  NOR2_X1 U110 ( .A1(n14), .A2(n86), .ZN(B_SHF[23]) );
  NOR2_X1 U111 ( .A1(n14), .A2(n77), .ZN(B_SHF[22]) );
  NOR2_X1 U112 ( .A1(n15), .A2(n169), .ZN(B_SHF[4]) );
  NAND4_X1 U113 ( .A1(n80), .A2(n81), .A3(n82), .A4(n181), .ZN(
        select_type_sig[0]) );
  NOR2_X1 U114 ( .A1(n12), .A2(n54), .ZN(A_SHF[30]) );
  INV_X1 U115 ( .A(n81), .ZN(n179) );
  NOR2_X1 U116 ( .A1(n14), .A2(n73), .ZN(B_SHF[19]) );
  NOR2_X1 U117 ( .A1(n14), .A2(n67), .ZN(B_SHF[13]) );
  NOR2_X1 U118 ( .A1(n14), .A2(n76), .ZN(B_SHF[21]) );
  NOR2_X1 U119 ( .A1(n14), .A2(n68), .ZN(B_SHF[14]) );
  NOR2_X1 U120 ( .A1(n14), .A2(n75), .ZN(B_SHF[20]) );
  NOR2_X1 U121 ( .A1(n13), .A2(n66), .ZN(B_SHF[12]) );
  NAND2_X1 U122 ( .A1(n16), .A2(n181), .ZN(select_type_sig[1]) );
  BUF_X1 U123 ( .A(n156), .Z(n28) );
  INV_X1 U124 ( .A(n80), .ZN(n177) );
  INV_X1 U125 ( .A(n82), .ZN(n176) );
  NOR2_X1 U126 ( .A1(n15), .A2(n167), .ZN(B_SHF[31]) );
  OAI22_X1 U127 ( .A1(n63), .A2(n28), .B1(OP2[0]), .B2(n29), .ZN(B_ADD[0]) );
  OAI22_X1 U128 ( .A1(n74), .A2(n27), .B1(OP2[1]), .B2(n30), .ZN(B_ADD[1]) );
  OAI22_X1 U129 ( .A1(n165), .A2(n26), .B1(OP2[2]), .B2(n29), .ZN(B_ADD[2]) );
  OAI22_X1 U130 ( .A1(n169), .A2(n26), .B1(OP2[4]), .B2(n29), .ZN(B_ADD[4]) );
  OAI22_X1 U131 ( .A1(n170), .A2(n26), .B1(OP2[5]), .B2(n29), .ZN(B_ADD[5]) );
  OAI22_X1 U132 ( .A1(n171), .A2(n26), .B1(OP2[6]), .B2(n29), .ZN(B_ADD[6]) );
  OAI22_X1 U133 ( .A1(n173), .A2(n26), .B1(OP2[8]), .B2(n29), .ZN(B_ADD[8]) );
  OAI22_X1 U134 ( .A1(n174), .A2(n26), .B1(OP2[9]), .B2(n29), .ZN(B_ADD[9]) );
  OAI22_X1 U135 ( .A1(n71), .A2(n27), .B1(OP2[17]), .B2(n30), .ZN(B_ADD[17])
         );
  OAI22_X1 U136 ( .A1(n72), .A2(n27), .B1(OP2[18]), .B2(n30), .ZN(B_ADD[18])
         );
  OAI22_X1 U137 ( .A1(n75), .A2(n27), .B1(OP2[20]), .B2(n30), .ZN(B_ADD[20])
         );
  OAI22_X1 U138 ( .A1(n76), .A2(n27), .B1(OP2[21]), .B2(n30), .ZN(B_ADD[21])
         );
  OAI22_X1 U139 ( .A1(n77), .A2(n27), .B1(OP2[22]), .B2(n30), .ZN(B_ADD[22])
         );
  OAI22_X1 U140 ( .A1(n159), .A2(n27), .B1(OP2[24]), .B2(n30), .ZN(B_ADD[24])
         );
  OAI22_X1 U141 ( .A1(n160), .A2(n27), .B1(OP2[25]), .B2(n30), .ZN(B_ADD[25])
         );
  OAI22_X1 U142 ( .A1(n161), .A2(n27), .B1(OP2[26]), .B2(n30), .ZN(B_ADD[26])
         );
  OAI22_X1 U143 ( .A1(n163), .A2(n26), .B1(OP2[28]), .B2(n29), .ZN(B_ADD[28])
         );
  OAI22_X1 U144 ( .A1(n164), .A2(n26), .B1(OP2[29]), .B2(n29), .ZN(B_ADD[29])
         );
  OAI22_X1 U145 ( .A1(n166), .A2(n26), .B1(OP2[30]), .B2(n29), .ZN(B_ADD[30])
         );
  OAI22_X1 U146 ( .A1(n168), .A2(n26), .B1(OP2[3]), .B2(n29), .ZN(B_ADD[3]) );
  OAI22_X1 U147 ( .A1(n172), .A2(n26), .B1(OP2[7]), .B2(n29), .ZN(B_ADD[7]) );
  OAI22_X1 U148 ( .A1(n73), .A2(n27), .B1(OP2[19]), .B2(n30), .ZN(B_ADD[19])
         );
  OAI22_X1 U149 ( .A1(n86), .A2(n27), .B1(OP2[23]), .B2(n30), .ZN(B_ADD[23])
         );
  OAI22_X1 U150 ( .A1(n162), .A2(n27), .B1(OP2[27]), .B2(n30), .ZN(B_ADD[27])
         );
  OAI22_X1 U151 ( .A1(n167), .A2(n26), .B1(OP2[31]), .B2(n29), .ZN(B_ADD[31])
         );
  OAI22_X1 U152 ( .A1(n64), .A2(n28), .B1(OP2[10]), .B2(n30), .ZN(B_ADD[10])
         );
  OAI22_X1 U153 ( .A1(n66), .A2(n28), .B1(OP2[12]), .B2(n29), .ZN(B_ADD[12])
         );
  OAI22_X1 U154 ( .A1(n67), .A2(n28), .B1(OP2[13]), .B2(n30), .ZN(B_ADD[13])
         );
  OAI22_X1 U155 ( .A1(n68), .A2(n28), .B1(OP2[14]), .B2(n29), .ZN(B_ADD[14])
         );
  OAI22_X1 U156 ( .A1(n70), .A2(n28), .B1(OP2[16]), .B2(n30), .ZN(B_ADD[16])
         );
  OAI22_X1 U157 ( .A1(n65), .A2(n28), .B1(OP2[11]), .B2(n29), .ZN(B_ADD[11])
         );
  OAI22_X1 U158 ( .A1(n69), .A2(n28), .B1(OP2[15]), .B2(n30), .ZN(B_ADD[15])
         );
  OAI22_X1 U159 ( .A1(n152), .A2(n63), .B1(n153), .B2(n31), .ZN(LOGIC_RES[0])
         );
  AOI21_X1 U160 ( .B1(n7), .B2(n63), .A(n19), .ZN(n153) );
  AOI221_X1 U161 ( .B1(OP1[0]), .B2(n4), .C1(n5), .C2(n31), .A(n17), .ZN(n152)
         );
  OAI22_X1 U162 ( .A1(n130), .A2(n74), .B1(n131), .B2(n42), .ZN(LOGIC_RES[1])
         );
  AOI21_X1 U163 ( .B1(n9), .B2(n74), .A(n21), .ZN(n131) );
  AOI221_X1 U164 ( .B1(OP1[1]), .B2(n3), .C1(n6), .C2(n42), .A(n18), .ZN(n130)
         );
  OAI22_X1 U165 ( .A1(n108), .A2(n165), .B1(n109), .B2(n53), .ZN(LOGIC_RES[2])
         );
  AOI21_X1 U166 ( .B1(n8), .B2(n165), .A(n20), .ZN(n109) );
  AOI221_X1 U167 ( .B1(OP1[2]), .B2(n2), .C1(n7), .C2(n53), .A(n19), .ZN(n108)
         );
  OAI22_X1 U168 ( .A1(n102), .A2(n168), .B1(n103), .B2(n56), .ZN(LOGIC_RES[3])
         );
  AOI21_X1 U169 ( .B1(n8), .B2(n168), .A(n20), .ZN(n103) );
  AOI221_X1 U170 ( .B1(OP1[3]), .B2(n2), .C1(n6), .C2(n56), .A(n18), .ZN(n102)
         );
  OAI22_X1 U171 ( .A1(n100), .A2(n169), .B1(n101), .B2(n57), .ZN(LOGIC_RES[4])
         );
  AOI21_X1 U172 ( .B1(n8), .B2(n169), .A(n20), .ZN(n101) );
  AOI221_X1 U173 ( .B1(OP1[4]), .B2(n2), .C1(n6), .C2(n57), .A(n18), .ZN(n100)
         );
  OAI22_X1 U174 ( .A1(n98), .A2(n170), .B1(n99), .B2(n58), .ZN(LOGIC_RES[5])
         );
  AOI21_X1 U175 ( .B1(n7), .B2(n170), .A(n19), .ZN(n99) );
  AOI221_X1 U176 ( .B1(OP1[5]), .B2(n2), .C1(n6), .C2(n58), .A(n18), .ZN(n98)
         );
  OAI22_X1 U178 ( .A1(n96), .A2(n171), .B1(n97), .B2(n59), .ZN(LOGIC_RES[6])
         );
  AOI21_X1 U179 ( .B1(n7), .B2(n171), .A(n19), .ZN(n97) );
  AOI221_X1 U180 ( .B1(OP1[6]), .B2(n2), .C1(n5), .C2(n59), .A(n17), .ZN(n96)
         );
  OAI22_X1 U181 ( .A1(n94), .A2(n172), .B1(n95), .B2(n60), .ZN(LOGIC_RES[7])
         );
  AOI21_X1 U182 ( .B1(n8), .B2(n172), .A(n20), .ZN(n95) );
  AOI221_X1 U183 ( .B1(OP1[7]), .B2(n2), .C1(n5), .C2(n60), .A(n17), .ZN(n94)
         );
  OAI22_X1 U184 ( .A1(n92), .A2(n173), .B1(n93), .B2(n61), .ZN(LOGIC_RES[8])
         );
  AOI21_X1 U185 ( .B1(n7), .B2(n173), .A(n19), .ZN(n93) );
  AOI221_X1 U186 ( .B1(OP1[8]), .B2(n2), .C1(n5), .C2(n61), .A(n17), .ZN(n92)
         );
  OAI22_X1 U187 ( .A1(n90), .A2(n174), .B1(n91), .B2(n62), .ZN(LOGIC_RES[9])
         );
  AOI21_X1 U188 ( .B1(n8), .B2(n174), .A(n20), .ZN(n91) );
  AOI221_X1 U189 ( .B1(n2), .B2(OP1[9]), .C1(n5), .C2(n62), .A(n17), .ZN(n90)
         );
  OAI22_X1 U190 ( .A1(n150), .A2(n64), .B1(n151), .B2(n32), .ZN(LOGIC_RES[10])
         );
  AOI21_X1 U191 ( .B1(n10), .B2(n64), .A(n22), .ZN(n151) );
  AOI221_X1 U192 ( .B1(OP1[10]), .B2(n4), .C1(n5), .C2(n32), .A(n17), .ZN(n150) );
  OAI22_X1 U193 ( .A1(n148), .A2(n65), .B1(n149), .B2(n33), .ZN(LOGIC_RES[11])
         );
  AOI21_X1 U194 ( .B1(n10), .B2(n65), .A(n22), .ZN(n149) );
  AOI221_X1 U195 ( .B1(OP1[11]), .B2(n4), .C1(n5), .C2(n33), .A(n17), .ZN(n148) );
  OAI22_X1 U196 ( .A1(n146), .A2(n66), .B1(n147), .B2(n34), .ZN(LOGIC_RES[12])
         );
  AOI21_X1 U197 ( .B1(n10), .B2(n66), .A(n21), .ZN(n147) );
  AOI221_X1 U198 ( .B1(OP1[12]), .B2(n4), .C1(n5), .C2(n34), .A(n17), .ZN(n146) );
  OAI22_X1 U199 ( .A1(n144), .A2(n67), .B1(n145), .B2(n35), .ZN(LOGIC_RES[13])
         );
  AOI21_X1 U200 ( .B1(n10), .B2(n67), .A(n21), .ZN(n145) );
  AOI221_X1 U201 ( .B1(OP1[13]), .B2(n4), .C1(n5), .C2(n35), .A(n17), .ZN(n144) );
  OAI22_X1 U202 ( .A1(n142), .A2(n68), .B1(n143), .B2(n36), .ZN(LOGIC_RES[14])
         );
  AOI21_X1 U203 ( .B1(n9), .B2(n68), .A(n21), .ZN(n143) );
  AOI221_X1 U204 ( .B1(OP1[14]), .B2(n4), .C1(n5), .C2(n36), .A(n17), .ZN(n142) );
  OAI22_X1 U205 ( .A1(n140), .A2(n69), .B1(n141), .B2(n37), .ZN(LOGIC_RES[15])
         );
  AOI21_X1 U206 ( .B1(n9), .B2(n69), .A(n21), .ZN(n141) );
  AOI221_X1 U207 ( .B1(OP1[15]), .B2(n4), .C1(n5), .C2(n37), .A(n17), .ZN(n140) );
  OAI22_X1 U208 ( .A1(n138), .A2(n70), .B1(n139), .B2(n38), .ZN(LOGIC_RES[16])
         );
  AOI21_X1 U209 ( .B1(n9), .B2(n70), .A(n21), .ZN(n139) );
  AOI221_X1 U210 ( .B1(OP1[16]), .B2(n4), .C1(n5), .C2(n38), .A(n17), .ZN(n138) );
  OAI22_X1 U211 ( .A1(n136), .A2(n71), .B1(n137), .B2(n39), .ZN(LOGIC_RES[17])
         );
  AOI21_X1 U212 ( .B1(n9), .B2(n71), .A(n21), .ZN(n137) );
  AOI221_X1 U213 ( .B1(OP1[17]), .B2(n3), .C1(n6), .C2(n39), .A(n18), .ZN(n136) );
  OAI22_X1 U214 ( .A1(n134), .A2(n72), .B1(n135), .B2(n40), .ZN(LOGIC_RES[18])
         );
  AOI21_X1 U215 ( .B1(n9), .B2(n72), .A(n21), .ZN(n135) );
  AOI221_X1 U216 ( .B1(OP1[18]), .B2(n3), .C1(n6), .C2(n40), .A(n18), .ZN(n134) );
  OAI22_X1 U217 ( .A1(n132), .A2(n73), .B1(n133), .B2(n41), .ZN(LOGIC_RES[19])
         );
  AOI21_X1 U218 ( .B1(n9), .B2(n73), .A(n21), .ZN(n133) );
  AOI221_X1 U219 ( .B1(OP1[19]), .B2(n3), .C1(n6), .C2(n41), .A(n18), .ZN(n132) );
  OAI22_X1 U220 ( .A1(n128), .A2(n75), .B1(n129), .B2(n43), .ZN(LOGIC_RES[20])
         );
  AOI21_X1 U221 ( .B1(n9), .B2(n75), .A(n21), .ZN(n129) );
  AOI221_X1 U222 ( .B1(OP1[20]), .B2(n3), .C1(n6), .C2(n43), .A(n18), .ZN(n128) );
  OAI22_X1 U223 ( .A1(n126), .A2(n76), .B1(n127), .B2(n44), .ZN(LOGIC_RES[21])
         );
  AOI21_X1 U224 ( .B1(n9), .B2(n76), .A(n21), .ZN(n127) );
  AOI221_X1 U225 ( .B1(OP1[21]), .B2(n3), .C1(n6), .C2(n44), .A(n18), .ZN(n126) );
  OAI22_X1 U226 ( .A1(n124), .A2(n77), .B1(n125), .B2(n45), .ZN(LOGIC_RES[22])
         );
  AOI21_X1 U227 ( .B1(n9), .B2(n77), .A(n21), .ZN(n125) );
  AOI221_X1 U228 ( .B1(OP1[22]), .B2(n3), .C1(n6), .C2(n45), .A(n18), .ZN(n124) );
  OAI22_X1 U229 ( .A1(n122), .A2(n86), .B1(n123), .B2(n46), .ZN(LOGIC_RES[23])
         );
  AOI21_X1 U230 ( .B1(n9), .B2(n86), .A(n21), .ZN(n123) );
  AOI221_X1 U231 ( .B1(OP1[23]), .B2(n3), .C1(n6), .C2(n46), .A(n18), .ZN(n122) );
  OAI22_X1 U232 ( .A1(n120), .A2(n159), .B1(n121), .B2(n47), .ZN(LOGIC_RES[24]) );
  AOI21_X1 U233 ( .B1(n9), .B2(n159), .A(n20), .ZN(n121) );
  AOI221_X1 U234 ( .B1(OP1[24]), .B2(n3), .C1(n7), .C2(n47), .A(n19), .ZN(n120) );
  OAI22_X1 U235 ( .A1(n118), .A2(n160), .B1(n119), .B2(n48), .ZN(LOGIC_RES[25]) );
  AOI21_X1 U236 ( .B1(n8), .B2(n160), .A(n20), .ZN(n119) );
  AOI221_X1 U237 ( .B1(OP1[25]), .B2(n3), .C1(n7), .C2(n48), .A(n19), .ZN(n118) );
  OAI22_X1 U238 ( .A1(n116), .A2(n161), .B1(n117), .B2(n49), .ZN(LOGIC_RES[26]) );
  AOI21_X1 U239 ( .B1(n8), .B2(n161), .A(n20), .ZN(n117) );
  AOI221_X1 U240 ( .B1(OP1[26]), .B2(n3), .C1(n6), .C2(n49), .A(n18), .ZN(n116) );
  OAI22_X1 U241 ( .A1(n114), .A2(n162), .B1(n115), .B2(n50), .ZN(LOGIC_RES[27]) );
  AOI21_X1 U242 ( .B1(n8), .B2(n162), .A(n20), .ZN(n115) );
  AOI221_X1 U243 ( .B1(OP1[27]), .B2(n3), .C1(n7), .C2(n50), .A(n19), .ZN(n114) );
  OAI22_X1 U244 ( .A1(n112), .A2(n163), .B1(n113), .B2(n51), .ZN(LOGIC_RES[28]) );
  AOI21_X1 U245 ( .B1(n8), .B2(n163), .A(n20), .ZN(n113) );
  AOI221_X1 U246 ( .B1(OP1[28]), .B2(n2), .C1(n7), .C2(n51), .A(n19), .ZN(n112) );
  OAI22_X1 U247 ( .A1(n110), .A2(n164), .B1(n111), .B2(n52), .ZN(LOGIC_RES[29]) );
  AOI21_X1 U248 ( .B1(n8), .B2(n164), .A(n20), .ZN(n111) );
  AOI221_X1 U249 ( .B1(OP1[29]), .B2(n2), .C1(n7), .C2(n52), .A(n19), .ZN(n110) );
  OAI22_X1 U250 ( .A1(n106), .A2(n166), .B1(n107), .B2(n54), .ZN(LOGIC_RES[30]) );
  AOI21_X1 U251 ( .B1(n8), .B2(n166), .A(n20), .ZN(n107) );
  AOI221_X1 U252 ( .B1(OP1[30]), .B2(n2), .C1(n7), .C2(n54), .A(n19), .ZN(n106) );
  OAI22_X1 U253 ( .A1(n104), .A2(n167), .B1(n105), .B2(n55), .ZN(LOGIC_RES[31]) );
  AOI21_X1 U254 ( .B1(n8), .B2(n167), .A(n20), .ZN(n105) );
  AOI221_X1 U255 ( .B1(OP1[31]), .B2(n2), .C1(n7), .C2(n55), .A(n19), .ZN(n104) );
  INV_X1 U256 ( .A(n85), .ZN(n180) );
  INV_X1 U257 ( .A(\OPSel[0] ), .ZN(n181) );
  INV_X1 U258 ( .A(OP1[10]), .ZN(n32) );
  INV_X1 U259 ( .A(OP1[16]), .ZN(n38) );
  INV_X1 U260 ( .A(OP1[20]), .ZN(n43) );
  INV_X1 U261 ( .A(OP1[4]), .ZN(n57) );
  INV_X1 U262 ( .A(OP1[12]), .ZN(n34) );
  INV_X1 U263 ( .A(OP1[21]), .ZN(n44) );
  INV_X1 U264 ( .A(OP1[13]), .ZN(n35) );
  INV_X1 U265 ( .A(OP1[22]), .ZN(n45) );
  INV_X1 U266 ( .A(OP1[14]), .ZN(n36) );
  INV_X1 U267 ( .A(OP1[0]), .ZN(n31) );
  INV_X1 U268 ( .A(OP1[1]), .ZN(n42) );
  INV_X1 U269 ( .A(OP1[2]), .ZN(n53) );
  INV_X1 U270 ( .A(OP1[17]), .ZN(n39) );
  INV_X1 U271 ( .A(OP1[18]), .ZN(n40) );
  INV_X1 U272 ( .A(OP1[5]), .ZN(n58) );
  INV_X1 U273 ( .A(OP1[6]), .ZN(n59) );
  INV_X1 U274 ( .A(OP1[24]), .ZN(n47) );
  INV_X1 U275 ( .A(OP1[25]), .ZN(n48) );
  INV_X1 U276 ( .A(OP1[28]), .ZN(n51) );
  INV_X1 U277 ( .A(OP1[29]), .ZN(n52) );
  INV_X1 U278 ( .A(OP1[30]), .ZN(n54) );
  INV_X1 U279 ( .A(OP1[8]), .ZN(n61) );
  INV_X1 U280 ( .A(OP1[9]), .ZN(n62) );
  INV_X1 U281 ( .A(OP1[26]), .ZN(n49) );
  INV_X1 U282 ( .A(OP1[3]), .ZN(n56) );
  INV_X1 U283 ( .A(OP1[7]), .ZN(n60) );
  INV_X1 U284 ( .A(OP1[11]), .ZN(n33) );
  INV_X1 U285 ( .A(OP1[15]), .ZN(n37) );
  INV_X1 U286 ( .A(OP1[19]), .ZN(n41) );
  INV_X1 U287 ( .A(OP1[23]), .ZN(n46) );
  INV_X1 U288 ( .A(OP1[27]), .ZN(n50) );
  INV_X1 U289 ( .A(OP1[31]), .ZN(n55) );
  INV_X1 U290 ( .A(OP2[1]), .ZN(n74) );
  INV_X1 U291 ( .A(OP2[0]), .ZN(n63) );
  INV_X1 U292 ( .A(OP2[2]), .ZN(n165) );
  INV_X1 U293 ( .A(OP2[6]), .ZN(n171) );
  INV_X1 U294 ( .A(OP2[5]), .ZN(n170) );
  INV_X1 U295 ( .A(OP2[4]), .ZN(n169) );
  INV_X1 U296 ( .A(OP2[13]), .ZN(n67) );
  INV_X1 U297 ( .A(OP2[14]), .ZN(n68) );
  INV_X1 U298 ( .A(OP2[12]), .ZN(n66) );
  INV_X1 U299 ( .A(OP2[16]), .ZN(n70) );
  INV_X1 U300 ( .A(OP2[17]), .ZN(n71) );
  INV_X1 U301 ( .A(OP2[8]), .ZN(n173) );
  INV_X1 U302 ( .A(OP2[9]), .ZN(n174) );
  INV_X1 U303 ( .A(OP2[10]), .ZN(n64) );
  INV_X1 U304 ( .A(OP2[18]), .ZN(n72) );
  INV_X1 U305 ( .A(OP2[21]), .ZN(n76) );
  INV_X1 U306 ( .A(OP2[20]), .ZN(n75) );
  INV_X1 U307 ( .A(OP2[30]), .ZN(n166) );
  INV_X1 U308 ( .A(OP2[29]), .ZN(n164) );
  INV_X1 U309 ( .A(OP2[24]), .ZN(n159) );
  INV_X1 U310 ( .A(OP2[22]), .ZN(n77) );
  INV_X1 U311 ( .A(OP2[25]), .ZN(n160) );
  INV_X1 U312 ( .A(OP2[26]), .ZN(n161) );
  INV_X1 U313 ( .A(OP2[28]), .ZN(n163) );
  INV_X1 U314 ( .A(OP2[3]), .ZN(n168) );
  INV_X1 U315 ( .A(OP2[7]), .ZN(n172) );
  INV_X1 U316 ( .A(OP2[11]), .ZN(n65) );
  INV_X1 U325 ( .A(OP2[15]), .ZN(n69) );
  INV_X1 U326 ( .A(OP2[19]), .ZN(n73) );
  INV_X1 U327 ( .A(OP2[23]), .ZN(n86) );
  INV_X1 U328 ( .A(OP2[27]), .ZN(n162) );
  INV_X1 U329 ( .A(OP2[31]), .ZN(n167) );
  AND2_X1 U330 ( .A1(n154), .A2(n89), .ZN(n1) );
  INV_X1 U331 ( .A(n83), .ZN(n182) );
  INV_X1 U332 ( .A(LOGIC_ARITH), .ZN(n178) );
  NAND2_X1 U333 ( .A1(n155), .A2(n89), .ZN(n82) );
  NAND2_X1 U334 ( .A1(n155), .A2(n88), .ZN(n80) );
  NAND2_X1 U335 ( .A1(n154), .A2(n88), .ZN(n81) );
  INV_X1 U336 ( .A(n84), .ZN(n183) );
  NOR2_X1 U337 ( .A1(n185), .A2(ALU_OPC[2]), .ZN(n89) );
  NOR2_X1 U338 ( .A1(n186), .A2(ALU_OPC[3]), .ZN(n155) );
  NOR2_X1 U339 ( .A1(n184), .A2(ALU_OPC[1]), .ZN(n88) );
  NOR2_X1 U340 ( .A1(ALU_OPC[3]), .A2(ALU_OPC[0]), .ZN(n154) );
  NAND2_X1 U341 ( .A1(n85), .A2(n157), .ZN(LOGIC_ARITH) );
  OAI21_X1 U342 ( .B1(n78), .B2(n175), .A(n79), .ZN(select_zero_sig) );
  INV_X1 U343 ( .A(ALU_OPC[3]), .ZN(n175) );
  AOI22_X1 U344 ( .A1(ALU_OPC[0]), .A2(n185), .B1(ALU_OPC[2]), .B2(ALU_OPC[1]), 
        .ZN(n78) );
  INV_X1 U345 ( .A(ALU_OPC[1]), .ZN(n185) );
  INV_X1 U346 ( .A(ALU_OPC[0]), .ZN(n186) );
  INV_X1 U347 ( .A(ALU_OPC[2]), .ZN(n184) );
  CLKBUF_X1 U348 ( .A(n177), .Z(n10) );
  CLKBUF_X1 U349 ( .A(n178), .Z(n16) );
  CLKBUF_X1 U350 ( .A(n179), .Z(n22) );
  INV_X1 U351 ( .A(n1), .ZN(n29) );
  INV_X1 U352 ( .A(n1), .ZN(n30) );
endmodule


module regn_N32_6 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
endmodule


module regn_N32_5 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
endmodule


module regn_N5_2 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 \DOUT_reg[4]  ( .D(n16), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n21)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n17), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n22)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n18), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n23)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n19), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n24)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n20), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n25)
         );
  OAI21_X1 U2 ( .B1(n25), .B2(EN), .A(n30), .ZN(n20) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n30) );
  OAI21_X1 U4 ( .B1(n24), .B2(EN), .A(n29), .ZN(n19) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n29) );
  OAI21_X1 U6 ( .B1(n23), .B2(EN), .A(n28), .ZN(n18) );
  NAND2_X1 U7 ( .A1(DIN[2]), .A2(EN), .ZN(n28) );
  OAI21_X1 U8 ( .B1(n22), .B2(EN), .A(n27), .ZN(n17) );
  NAND2_X1 U9 ( .A1(DIN[3]), .A2(EN), .ZN(n27) );
  OAI21_X1 U10 ( .B1(n21), .B2(EN), .A(n26), .ZN(n16) );
  NAND2_X1 U11 ( .A1(DIN[4]), .A2(EN), .ZN(n26) );
endmodule


module regn_N32_4 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
endmodule


module regn_N32_3 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
endmodule


module Execute_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \B[0] , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57;
  assign SUM[1] = B[1];
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR2_X1 U1 ( .A(B[31]), .B(n57), .ZN(SUM[31]) );
  NAND2_X1 U2 ( .A1(B[30]), .A2(n56), .ZN(n57) );
  INV_X1 U3 ( .A(B[2]), .ZN(SUM[2]) );
  XOR2_X1 U4 ( .A(B[3]), .B(B[2]), .Z(SUM[3]) );
  XOR2_X1 U5 ( .A(B[4]), .B(n30), .Z(SUM[4]) );
  XOR2_X1 U6 ( .A(B[5]), .B(n31), .Z(SUM[5]) );
  XOR2_X1 U7 ( .A(B[6]), .B(n32), .Z(SUM[6]) );
  XOR2_X1 U8 ( .A(B[7]), .B(n33), .Z(SUM[7]) );
  XOR2_X1 U9 ( .A(B[8]), .B(n34), .Z(SUM[8]) );
  XOR2_X1 U10 ( .A(B[9]), .B(n35), .Z(SUM[9]) );
  XOR2_X1 U11 ( .A(B[10]), .B(n36), .Z(SUM[10]) );
  XOR2_X1 U12 ( .A(B[11]), .B(n37), .Z(SUM[11]) );
  XOR2_X1 U13 ( .A(B[12]), .B(n38), .Z(SUM[12]) );
  XOR2_X1 U14 ( .A(B[13]), .B(n39), .Z(SUM[13]) );
  XOR2_X1 U15 ( .A(B[14]), .B(n40), .Z(SUM[14]) );
  XOR2_X1 U16 ( .A(B[15]), .B(n41), .Z(SUM[15]) );
  XOR2_X1 U17 ( .A(B[16]), .B(n42), .Z(SUM[16]) );
  XOR2_X1 U18 ( .A(B[17]), .B(n43), .Z(SUM[17]) );
  XOR2_X1 U19 ( .A(B[18]), .B(n44), .Z(SUM[18]) );
  XOR2_X1 U20 ( .A(B[19]), .B(n45), .Z(SUM[19]) );
  XOR2_X1 U21 ( .A(B[20]), .B(n46), .Z(SUM[20]) );
  XOR2_X1 U22 ( .A(B[21]), .B(n47), .Z(SUM[21]) );
  XOR2_X1 U23 ( .A(B[22]), .B(n48), .Z(SUM[22]) );
  XOR2_X1 U24 ( .A(B[23]), .B(n49), .Z(SUM[23]) );
  XOR2_X1 U25 ( .A(B[24]), .B(n50), .Z(SUM[24]) );
  XOR2_X1 U26 ( .A(B[25]), .B(n51), .Z(SUM[25]) );
  XOR2_X1 U27 ( .A(B[26]), .B(n52), .Z(SUM[26]) );
  XOR2_X1 U28 ( .A(B[27]), .B(n53), .Z(SUM[27]) );
  XOR2_X1 U29 ( .A(B[28]), .B(n54), .Z(SUM[28]) );
  XOR2_X1 U30 ( .A(B[29]), .B(n55), .Z(SUM[29]) );
  XOR2_X1 U31 ( .A(B[30]), .B(n56), .Z(SUM[30]) );
  AND2_X1 U32 ( .A1(B[3]), .A2(B[2]), .ZN(n30) );
  AND2_X1 U33 ( .A1(B[4]), .A2(n30), .ZN(n31) );
  AND2_X1 U34 ( .A1(B[5]), .A2(n31), .ZN(n32) );
  AND2_X1 U35 ( .A1(B[6]), .A2(n32), .ZN(n33) );
  AND2_X1 U36 ( .A1(B[7]), .A2(n33), .ZN(n34) );
  AND2_X1 U37 ( .A1(B[8]), .A2(n34), .ZN(n35) );
  AND2_X1 U38 ( .A1(B[9]), .A2(n35), .ZN(n36) );
  AND2_X1 U39 ( .A1(B[10]), .A2(n36), .ZN(n37) );
  AND2_X1 U40 ( .A1(B[11]), .A2(n37), .ZN(n38) );
  AND2_X1 U41 ( .A1(B[12]), .A2(n38), .ZN(n39) );
  AND2_X1 U42 ( .A1(B[13]), .A2(n39), .ZN(n40) );
  AND2_X1 U43 ( .A1(B[14]), .A2(n40), .ZN(n41) );
  AND2_X1 U44 ( .A1(B[15]), .A2(n41), .ZN(n42) );
  AND2_X1 U45 ( .A1(B[16]), .A2(n42), .ZN(n43) );
  AND2_X1 U46 ( .A1(B[17]), .A2(n43), .ZN(n44) );
  AND2_X1 U47 ( .A1(B[18]), .A2(n44), .ZN(n45) );
  AND2_X1 U48 ( .A1(B[19]), .A2(n45), .ZN(n46) );
  AND2_X1 U49 ( .A1(B[20]), .A2(n46), .ZN(n47) );
  AND2_X1 U50 ( .A1(B[21]), .A2(n47), .ZN(n48) );
  AND2_X1 U51 ( .A1(B[22]), .A2(n48), .ZN(n49) );
  AND2_X1 U52 ( .A1(B[23]), .A2(n49), .ZN(n50) );
  AND2_X1 U53 ( .A1(B[24]), .A2(n50), .ZN(n51) );
  AND2_X1 U54 ( .A1(B[25]), .A2(n51), .ZN(n52) );
  AND2_X1 U55 ( .A1(B[26]), .A2(n52), .ZN(n53) );
  AND2_X1 U56 ( .A1(B[27]), .A2(n53), .ZN(n54) );
  AND2_X1 U57 ( .A1(B[28]), .A2(n54), .ZN(n55) );
  AND2_X1 U58 ( .A1(B[29]), .A2(n55), .ZN(n56) );
endmodule


module Execute_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module Execute ( CLK, RST, MUX_A_SEL, MUX_B_SEL, .ALU_OPC({\ALU_OPC[3] , 
        \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), ALU_OUTREG_EN, JUMP_TYPE, 
        PC_IN, A_IN, B_IN, IMM_IN, ADD_WR_IN, ADD_RS1_IN, ADD_RS2_IN, 
        ADD_WR_MEM, ADD_WR_WB, RF_WE_MEM, RF_WE_WB, OP_MEM, OP_WB, PC_SEL, 
        ZERO_FLAG, NPC_ABS, NPC_REL, ALU_RES, B_OUT, ADD_WR_OUT );
  input [1:0] MUX_B_SEL;
  input [1:0] JUMP_TYPE;
  input [31:0] PC_IN;
  input [31:0] A_IN;
  input [31:0] B_IN;
  input [31:0] IMM_IN;
  input [4:0] ADD_WR_IN;
  input [4:0] ADD_RS1_IN;
  input [4:0] ADD_RS2_IN;
  input [4:0] ADD_WR_MEM;
  input [4:0] ADD_WR_WB;
  input [31:0] OP_MEM;
  input [31:0] OP_WB;
  output [1:0] PC_SEL;
  output [31:0] NPC_ABS;
  output [31:0] NPC_REL;
  output [31:0] ALU_RES;
  output [31:0] B_OUT;
  output [4:0] ADD_WR_OUT;
  input CLK, RST, MUX_A_SEL, \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] ,
         \ALU_OPC[0] , ALU_OUTREG_EN, RF_WE_MEM, RF_WE_WB;
  output ZERO_FLAG;
  wire   sig_RST, sig_ZERO_FLAG, N9, N8, N7, N6, N5, N4, N31, N30, N3, N29,
         N28, N27, N26, N25, N24, N23, N22, N21, N20, N2, N19, N18, N17, N16,
         N15, N14, N13, N12, N11, N10, N1, N0, n1;
  wire   [3:0] ALU_OPC;
  wire   [31:0] sig_NPC_ABS;
  wire   [31:0] sig_NPC_REL;
  wire   [1:0] sig_PC_SEL;
  wire   [1:0] FWDA;
  wire   [1:0] FWDB;
  wire   [31:0] OP2_FW;
  wire   [31:0] sig_OP1;
  wire   [31:0] sig_OP2;
  wire   [31:0] sig_ALU_RES;

  Branch_Cond_Unit_NBIT32 Branch_Cond ( .RST(sig_RST), .A(sig_NPC_ABS), 
        .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), 
        .JUMP_TYPE(JUMP_TYPE), .PC_SEL(sig_PC_SEL), .ZERO(sig_ZERO_FLAG) );
  ff_1 ff0 ( .D(sig_ZERO_FLAG), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(ZERO_FLAG)
         );
  regn_N2 reg0 ( .DIN(sig_PC_SEL), .CLK(CLK), .EN(1'b1), .RST(RST), .DOUT(
        PC_SEL) );
  FWD_Unit FWD ( .RST(sig_RST), .ADD_RS1(ADD_RS1_IN), .ADD_RS2(ADD_RS2_IN), 
        .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_WB(ADD_WR_WB), .RF_WE_MEM(RF_WE_MEM), 
        .RF_WE_WB(RF_WE_WB), .FWDA(FWDA), .FWDB(FWDB) );
  mux41_NBIT32_0 FW1 ( .A(A_IN), .B(OP_WB), .C(OP_MEM), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(FWDA), .Z(sig_NPC_ABS) );
  mux41_NBIT32_4 FW2 ( .A(B_IN), .B(OP_WB), .C(OP_MEM), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(FWDB), .Z(OP2_FW) );
  mux21_NBIT32_3 muxA ( .A(sig_NPC_ABS), .B(PC_IN), .S(MUX_A_SEL), .Z(sig_OP1)
         );
  mux41_NBIT32_3 muxB ( .A(OP2_FW), .B(IMM_IN), .C({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(MUX_B_SEL), .Z(sig_OP2) );
  ALU_NBIT32 alu0 ( .OP1(sig_OP1), .OP2(sig_OP2), .ALU_OPC({\ALU_OPC[3] , 
        \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), .ALU_RES(sig_ALU_RES) );
  regn_N32_6 alureg ( .DIN(sig_ALU_RES), .CLK(CLK), .EN(ALU_OUTREG_EN), .RST(
        RST), .DOUT(ALU_RES) );
  regn_N32_5 B_reg ( .DIN(OP2_FW), .CLK(CLK), .EN(ALU_OUTREG_EN), .RST(RST), 
        .DOUT(B_OUT) );
  regn_N5_2 ADD_WR_reg ( .DIN(ADD_WR_IN), .CLK(CLK), .EN(ALU_OUTREG_EN), .RST(
        RST), .DOUT(ADD_WR_OUT) );
  regn_N32_4 NPC_ABS_reg ( .DIN(sig_NPC_ABS), .CLK(CLK), .EN(ALU_OUTREG_EN), 
        .RST(RST), .DOUT(NPC_ABS) );
  regn_N32_3 NPC_REL_reg ( .DIN(sig_NPC_REL), .CLK(CLK), .EN(ALU_OUTREG_EN), 
        .RST(RST), .DOUT(NPC_REL) );
  Execute_DW01_add_1 add_1_root_add_0_root_add_118_2 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .B(IMM_IN), .CI(1'b0), .SUM({N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0})
         );
  Execute_DW01_add_0 add_0_root_add_0_root_add_118_2 ( .A(PC_IN), .B({N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}), 
        .CI(1'b0), .SUM(sig_NPC_REL) );
  NOR2_X1 U3 ( .A1(ZERO_FLAG), .A2(n1), .ZN(sig_RST) );
  INV_X1 U4 ( .A(RST), .ZN(n1) );
endmodule


module ff_0 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n2, n3;

  DFFR_X1 Q_reg ( .D(n3), .CK(CLK), .RN(RST), .Q(Q), .QN(n2) );
  OAI21_X1 U2 ( .B1(n2), .B2(EN), .A(n1), .ZN(n3) );
  NAND2_X1 U3 ( .A1(EN), .A2(D), .ZN(n1) );
endmodule


module regn_N32_2 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  OAI21_X1 U2 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U4 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U6 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U7 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U8 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U9 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U10 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U11 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U12 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U13 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U14 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U15 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U16 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U17 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U18 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U19 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U20 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U21 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U22 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U23 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U24 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U25 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U26 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U27 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U28 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U29 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U30 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U31 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U32 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U33 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U34 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U35 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U36 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U37 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U38 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U39 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U40 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U41 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U42 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U43 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U44 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U45 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U46 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U47 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U48 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U49 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U50 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U51 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U52 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U53 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U54 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U55 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U56 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U57 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U58 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U59 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U60 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U61 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U62 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U63 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U64 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U65 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
  BUF_X1 U66 ( .A(RST), .Z(n97) );
  BUF_X1 U67 ( .A(RST), .Z(n98) );
  BUF_X1 U68 ( .A(RST), .Z(n99) );
endmodule


module regn_N5_1 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 \DOUT_reg[4]  ( .D(n16), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n21)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n17), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n22)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n18), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n23)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n19), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n24)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n20), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n25)
         );
  OAI21_X1 U2 ( .B1(n25), .B2(EN), .A(n30), .ZN(n20) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n30) );
  OAI21_X1 U4 ( .B1(n24), .B2(EN), .A(n29), .ZN(n19) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n29) );
  OAI21_X1 U6 ( .B1(n23), .B2(EN), .A(n28), .ZN(n18) );
  NAND2_X1 U7 ( .A1(DIN[2]), .A2(EN), .ZN(n28) );
  OAI21_X1 U8 ( .B1(n22), .B2(EN), .A(n27), .ZN(n17) );
  NAND2_X1 U9 ( .A1(DIN[3]), .A2(EN), .ZN(n27) );
  OAI21_X1 U10 ( .B1(n21), .B2(EN), .A(n26), .ZN(n16) );
  NAND2_X1 U11 ( .A1(DIN[4]), .A2(EN), .ZN(n26) );
endmodule


module regn_N32_1 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  OAI21_X1 U2 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U4 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U6 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U7 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U8 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U9 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U10 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U11 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U12 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U13 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U14 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U15 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U16 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U17 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U18 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U19 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U20 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U21 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U22 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U23 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U24 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U25 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U26 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U27 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U28 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U29 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U30 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U31 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U32 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U33 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U34 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U35 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U36 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U37 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U38 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U39 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U40 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U41 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U42 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U43 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U44 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U45 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U46 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U47 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U48 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U49 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U50 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U51 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U52 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U53 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U54 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U55 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U56 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U57 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U58 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U59 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U60 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U61 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U62 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U63 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U64 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U65 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
  BUF_X1 U66 ( .A(RST), .Z(n97) );
  BUF_X1 U67 ( .A(RST), .Z(n98) );
  BUF_X1 U68 ( .A(RST), .Z(n99) );
endmodule


module mux41_NBIT32_2 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n20, n21, n22, n23, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105;

  OAI221_X1 U1 ( .B1(n1), .B2(n9), .C1(n2), .C2(n3), .A(n105), .ZN(Z[7]) );
  INV_X1 U2 ( .A(B[7]), .ZN(n1) );
  INV_X1 U3 ( .A(A[7]), .ZN(n2) );
  INV_X1 U4 ( .A(n32), .ZN(n3) );
  OAI221_X1 U5 ( .B1(n4), .B2(n5), .C1(n6), .C2(n7), .A(n50), .ZN(Z[9]) );
  INV_X1 U6 ( .A(B[9]), .ZN(n4) );
  INV_X1 U7 ( .A(n34), .ZN(n5) );
  INV_X1 U8 ( .A(A[9]), .ZN(n6) );
  INV_X1 U9 ( .A(n32), .ZN(n7) );
  AOI22_X1 U10 ( .A1(B[27]), .A2(n34), .B1(A[27]), .B2(n32), .ZN(n82) );
  OAI221_X1 U11 ( .B1(n8), .B2(n9), .C1(n10), .C2(n7), .A(n78), .ZN(Z[25]) );
  INV_X1 U12 ( .A(B[25]), .ZN(n8) );
  INV_X1 U13 ( .A(n34), .ZN(n9) );
  INV_X1 U14 ( .A(A[25]), .ZN(n10) );
  OAI221_X1 U15 ( .B1(n20), .B2(n5), .C1(n21), .C2(n3), .A(n63), .ZN(Z[17]) );
  INV_X1 U16 ( .A(B[17]), .ZN(n20) );
  INV_X1 U17 ( .A(A[17]), .ZN(n21) );
  OAI221_X1 U18 ( .B1(n22), .B2(n5), .C1(n23), .C2(n7), .A(n51), .ZN(Z[10]) );
  INV_X1 U19 ( .A(B[10]), .ZN(n22) );
  INV_X1 U20 ( .A(A[10]), .ZN(n23) );
  OAI221_X1 U21 ( .B1(n26), .B2(n9), .C1(n27), .C2(n7), .A(n52), .ZN(Z[11]) );
  INV_X1 U22 ( .A(B[11]), .ZN(n26) );
  INV_X1 U23 ( .A(A[11]), .ZN(n27) );
  AOI221_X1 U24 ( .B1(B[19]), .B2(n34), .C1(A[19]), .C2(n32), .A(n28), .ZN(n29) );
  INV_X1 U25 ( .A(n66), .ZN(n28) );
  INV_X1 U26 ( .A(n29), .ZN(Z[19]) );
  OAI221_X1 U27 ( .B1(n30), .B2(n5), .C1(n31), .C2(n3), .A(n67), .ZN(Z[20]) );
  INV_X1 U28 ( .A(B[20]), .ZN(n30) );
  INV_X1 U29 ( .A(A[20]), .ZN(n31) );
  AOI22_X1 U30 ( .A1(B[28]), .A2(n34), .B1(A[28]), .B2(n32), .ZN(n84) );
  AOI22_X1 U31 ( .A1(B[31]), .A2(n34), .B1(A[31]), .B2(n32), .ZN(n90) );
  AOI22_X1 U32 ( .A1(B[15]), .A2(n34), .B1(A[15]), .B2(n32), .ZN(n60) );
  BUF_X1 U33 ( .A(n32), .Z(n41) );
  BUF_X1 U34 ( .A(n32), .Z(n40) );
  BUF_X1 U35 ( .A(n34), .Z(n43) );
  BUF_X1 U36 ( .A(n33), .Z(n37) );
  BUF_X1 U37 ( .A(n33), .Z(n36) );
  BUF_X1 U38 ( .A(n34), .Z(n42) );
  AND2_X1 U39 ( .A1(n44), .A2(n45), .ZN(n32) );
  BUF_X1 U40 ( .A(n35), .Z(n39) );
  BUF_X1 U41 ( .A(n35), .Z(n38) );
  NAND2_X1 U42 ( .A1(n92), .A2(n91), .ZN(Z[0]) );
  AOI22_X1 U43 ( .A1(D[0]), .A2(n38), .B1(C[0]), .B2(n36), .ZN(n91) );
  AOI22_X1 U44 ( .A1(B[0]), .A2(n42), .B1(A[0]), .B2(n40), .ZN(n92) );
  AND2_X1 U45 ( .A1(S[1]), .A2(n45), .ZN(n33) );
  AND2_X1 U46 ( .A1(S[0]), .A2(n44), .ZN(n34) );
  AOI22_X1 U47 ( .A1(D[7]), .A2(n38), .B1(C[7]), .B2(n36), .ZN(n105) );
  NAND2_X1 U48 ( .A1(n96), .A2(n95), .ZN(Z[2]) );
  AOI22_X1 U49 ( .A1(D[2]), .A2(n38), .B1(C[2]), .B2(n36), .ZN(n95) );
  AOI22_X1 U50 ( .A1(B[2]), .A2(n42), .B1(A[2]), .B2(n40), .ZN(n96) );
  NAND2_X1 U51 ( .A1(n104), .A2(n103), .ZN(Z[6]) );
  AOI22_X1 U52 ( .A1(D[6]), .A2(n38), .B1(C[6]), .B2(n36), .ZN(n103) );
  AOI22_X1 U53 ( .A1(B[6]), .A2(n42), .B1(A[6]), .B2(n40), .ZN(n104) );
  NAND2_X1 U54 ( .A1(n102), .A2(n101), .ZN(Z[5]) );
  AOI22_X1 U55 ( .A1(D[5]), .A2(n38), .B1(C[5]), .B2(n36), .ZN(n101) );
  AOI22_X1 U56 ( .A1(B[5]), .A2(n42), .B1(A[5]), .B2(n40), .ZN(n102) );
  NAND2_X1 U57 ( .A1(n94), .A2(n93), .ZN(Z[1]) );
  AOI22_X1 U58 ( .A1(D[1]), .A2(n38), .B1(C[1]), .B2(n36), .ZN(n93) );
  AOI22_X1 U59 ( .A1(B[1]), .A2(n42), .B1(A[1]), .B2(n40), .ZN(n94) );
  NAND2_X1 U60 ( .A1(n98), .A2(n97), .ZN(Z[3]) );
  AOI22_X1 U61 ( .A1(D[3]), .A2(n38), .B1(C[3]), .B2(n36), .ZN(n97) );
  AOI22_X1 U62 ( .A1(B[3]), .A2(n42), .B1(A[3]), .B2(n40), .ZN(n98) );
  NAND2_X1 U63 ( .A1(n100), .A2(n99), .ZN(Z[4]) );
  AOI22_X1 U64 ( .A1(D[4]), .A2(n38), .B1(C[4]), .B2(n36), .ZN(n99) );
  AOI22_X1 U65 ( .A1(B[4]), .A2(n42), .B1(A[4]), .B2(n40), .ZN(n100) );
  AND2_X1 U66 ( .A1(S[0]), .A2(S[1]), .ZN(n35) );
  INV_X1 U67 ( .A(S[1]), .ZN(n44) );
  INV_X1 U68 ( .A(S[0]), .ZN(n45) );
  AOI22_X1 U69 ( .A1(B[8]), .A2(n43), .B1(A[8]), .B2(n41), .ZN(n49) );
  AOI22_X1 U70 ( .A1(D[8]), .A2(n39), .B1(C[8]), .B2(n37), .ZN(n48) );
  NAND2_X1 U71 ( .A1(n49), .A2(n48), .ZN(Z[8]) );
  AOI22_X1 U72 ( .A1(D[9]), .A2(n39), .B1(C[9]), .B2(n37), .ZN(n50) );
  AOI22_X1 U73 ( .A1(D[10]), .A2(n39), .B1(C[10]), .B2(n37), .ZN(n51) );
  AOI22_X1 U74 ( .A1(D[11]), .A2(n39), .B1(C[11]), .B2(n37), .ZN(n52) );
  AOI22_X1 U75 ( .A1(B[12]), .A2(n43), .B1(A[12]), .B2(n41), .ZN(n54) );
  AOI22_X1 U76 ( .A1(D[12]), .A2(n39), .B1(C[12]), .B2(n37), .ZN(n53) );
  NAND2_X1 U77 ( .A1(n54), .A2(n53), .ZN(Z[12]) );
  AOI22_X1 U78 ( .A1(B[13]), .A2(n43), .B1(A[13]), .B2(n41), .ZN(n56) );
  AOI22_X1 U79 ( .A1(D[13]), .A2(n39), .B1(C[13]), .B2(n37), .ZN(n55) );
  NAND2_X1 U80 ( .A1(n56), .A2(n55), .ZN(Z[13]) );
  AOI22_X1 U81 ( .A1(B[14]), .A2(n43), .B1(A[14]), .B2(n41), .ZN(n58) );
  AOI22_X1 U82 ( .A1(D[14]), .A2(n39), .B1(C[14]), .B2(n37), .ZN(n57) );
  NAND2_X1 U83 ( .A1(n58), .A2(n57), .ZN(Z[14]) );
  AOI22_X1 U84 ( .A1(D[15]), .A2(n39), .B1(C[15]), .B2(n37), .ZN(n59) );
  NAND2_X1 U85 ( .A1(n60), .A2(n59), .ZN(Z[15]) );
  AOI22_X1 U86 ( .A1(B[16]), .A2(n43), .B1(A[16]), .B2(n41), .ZN(n62) );
  AOI22_X1 U87 ( .A1(D[16]), .A2(n39), .B1(C[16]), .B2(n37), .ZN(n61) );
  NAND2_X1 U88 ( .A1(n62), .A2(n61), .ZN(Z[16]) );
  AOI22_X1 U89 ( .A1(D[17]), .A2(n39), .B1(C[17]), .B2(n37), .ZN(n63) );
  AOI22_X1 U90 ( .A1(B[18]), .A2(n43), .B1(A[18]), .B2(n41), .ZN(n65) );
  AOI22_X1 U91 ( .A1(D[18]), .A2(n39), .B1(C[18]), .B2(n37), .ZN(n64) );
  NAND2_X1 U92 ( .A1(n65), .A2(n64), .ZN(Z[18]) );
  AOI22_X1 U93 ( .A1(D[19]), .A2(n39), .B1(C[19]), .B2(n37), .ZN(n66) );
  AOI22_X1 U94 ( .A1(D[20]), .A2(n39), .B1(C[20]), .B2(n37), .ZN(n67) );
  AOI22_X1 U95 ( .A1(B[21]), .A2(n43), .B1(A[21]), .B2(n41), .ZN(n71) );
  AOI22_X1 U96 ( .A1(D[21]), .A2(n39), .B1(C[21]), .B2(n37), .ZN(n70) );
  NAND2_X1 U97 ( .A1(n71), .A2(n70), .ZN(Z[21]) );
  AOI22_X1 U98 ( .A1(B[22]), .A2(n43), .B1(A[22]), .B2(n41), .ZN(n73) );
  AOI22_X1 U99 ( .A1(D[22]), .A2(n39), .B1(C[22]), .B2(n37), .ZN(n72) );
  NAND2_X1 U100 ( .A1(n73), .A2(n72), .ZN(Z[22]) );
  AOI22_X1 U101 ( .A1(B[23]), .A2(n43), .B1(A[23]), .B2(n41), .ZN(n75) );
  AOI22_X1 U102 ( .A1(D[23]), .A2(n39), .B1(C[23]), .B2(n37), .ZN(n74) );
  NAND2_X1 U103 ( .A1(n75), .A2(n74), .ZN(Z[23]) );
  AOI22_X1 U104 ( .A1(B[24]), .A2(n43), .B1(A[24]), .B2(n41), .ZN(n77) );
  AOI22_X1 U105 ( .A1(D[24]), .A2(n39), .B1(C[24]), .B2(n37), .ZN(n76) );
  NAND2_X1 U106 ( .A1(n77), .A2(n76), .ZN(Z[24]) );
  AOI22_X1 U107 ( .A1(D[25]), .A2(n38), .B1(C[25]), .B2(n36), .ZN(n78) );
  AOI22_X1 U108 ( .A1(B[26]), .A2(n42), .B1(A[26]), .B2(n40), .ZN(n80) );
  AOI22_X1 U109 ( .A1(D[26]), .A2(n38), .B1(C[26]), .B2(n36), .ZN(n79) );
  NAND2_X1 U110 ( .A1(n80), .A2(n79), .ZN(Z[26]) );
  AOI22_X1 U111 ( .A1(D[27]), .A2(n38), .B1(C[27]), .B2(n36), .ZN(n81) );
  NAND2_X1 U112 ( .A1(n82), .A2(n81), .ZN(Z[27]) );
  AOI22_X1 U113 ( .A1(D[28]), .A2(n38), .B1(C[28]), .B2(n36), .ZN(n83) );
  NAND2_X1 U114 ( .A1(n84), .A2(n83), .ZN(Z[28]) );
  AOI22_X1 U115 ( .A1(B[29]), .A2(n42), .B1(A[29]), .B2(n40), .ZN(n86) );
  AOI22_X1 U116 ( .A1(D[29]), .A2(n38), .B1(C[29]), .B2(n36), .ZN(n85) );
  NAND2_X1 U117 ( .A1(n86), .A2(n85), .ZN(Z[29]) );
  AOI22_X1 U118 ( .A1(B[30]), .A2(n42), .B1(A[30]), .B2(n40), .ZN(n88) );
  AOI22_X1 U119 ( .A1(D[30]), .A2(n38), .B1(C[30]), .B2(n36), .ZN(n87) );
  NAND2_X1 U120 ( .A1(n88), .A2(n87), .ZN(Z[30]) );
  AOI22_X1 U121 ( .A1(D[31]), .A2(n38), .B1(C[31]), .B2(n36), .ZN(n89) );
  NAND2_X1 U122 ( .A1(n90), .A2(n89), .ZN(Z[31]) );
endmodule


module Memory ( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, DRAM_EN_IN, PC_SEL, 
        NPC_IN, NPC_ABS, NPC_REL, ALU_RES_IN, B_IN, ADD_WR_IN, DRAM_DATA_IN, 
        PC_OUT, DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, DRAM_ADDR_OUT, 
        DRAM_DATA_OUT, DATA_OUT, ALU_RES_OUT, OP_MEM, ADD_WR_MEM, ADD_WR_OUT
 );
  input [1:0] PC_SEL;
  input [31:0] NPC_IN;
  input [31:0] NPC_ABS;
  input [31:0] NPC_REL;
  input [31:0] ALU_RES_IN;
  input [31:0] B_IN;
  input [4:0] ADD_WR_IN;
  input [31:0] DRAM_DATA_IN;
  output [31:0] PC_OUT;
  output [31:0] DRAM_ADDR_OUT;
  output [31:0] DRAM_DATA_OUT;
  output [31:0] DATA_OUT;
  output [31:0] ALU_RES_OUT;
  output [31:0] OP_MEM;
  output [4:0] ADD_WR_MEM;
  output [4:0] ADD_WR_OUT;
  input CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, DRAM_EN_IN;
  output DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT;
  wire   DRAM_EN_IN, DRAM_R_IN, DRAM_W_IN;
  assign DRAM_EN_OUT = DRAM_EN_IN;
  assign DRAM_R_OUT = DRAM_R_IN;
  assign DRAM_W_OUT = DRAM_W_IN;
  assign OP_MEM[31] = ALU_RES_IN[31];
  assign DRAM_ADDR_OUT[31] = ALU_RES_IN[31];
  assign OP_MEM[30] = ALU_RES_IN[30];
  assign DRAM_ADDR_OUT[30] = ALU_RES_IN[30];
  assign OP_MEM[29] = ALU_RES_IN[29];
  assign DRAM_ADDR_OUT[29] = ALU_RES_IN[29];
  assign OP_MEM[28] = ALU_RES_IN[28];
  assign DRAM_ADDR_OUT[28] = ALU_RES_IN[28];
  assign OP_MEM[27] = ALU_RES_IN[27];
  assign DRAM_ADDR_OUT[27] = ALU_RES_IN[27];
  assign OP_MEM[26] = ALU_RES_IN[26];
  assign DRAM_ADDR_OUT[26] = ALU_RES_IN[26];
  assign OP_MEM[25] = ALU_RES_IN[25];
  assign DRAM_ADDR_OUT[25] = ALU_RES_IN[25];
  assign OP_MEM[24] = ALU_RES_IN[24];
  assign DRAM_ADDR_OUT[24] = ALU_RES_IN[24];
  assign OP_MEM[23] = ALU_RES_IN[23];
  assign DRAM_ADDR_OUT[23] = ALU_RES_IN[23];
  assign OP_MEM[22] = ALU_RES_IN[22];
  assign DRAM_ADDR_OUT[22] = ALU_RES_IN[22];
  assign OP_MEM[21] = ALU_RES_IN[21];
  assign DRAM_ADDR_OUT[21] = ALU_RES_IN[21];
  assign OP_MEM[20] = ALU_RES_IN[20];
  assign DRAM_ADDR_OUT[20] = ALU_RES_IN[20];
  assign OP_MEM[19] = ALU_RES_IN[19];
  assign DRAM_ADDR_OUT[19] = ALU_RES_IN[19];
  assign OP_MEM[18] = ALU_RES_IN[18];
  assign DRAM_ADDR_OUT[18] = ALU_RES_IN[18];
  assign OP_MEM[17] = ALU_RES_IN[17];
  assign DRAM_ADDR_OUT[17] = ALU_RES_IN[17];
  assign OP_MEM[16] = ALU_RES_IN[16];
  assign DRAM_ADDR_OUT[16] = ALU_RES_IN[16];
  assign OP_MEM[15] = ALU_RES_IN[15];
  assign DRAM_ADDR_OUT[15] = ALU_RES_IN[15];
  assign OP_MEM[14] = ALU_RES_IN[14];
  assign DRAM_ADDR_OUT[14] = ALU_RES_IN[14];
  assign OP_MEM[13] = ALU_RES_IN[13];
  assign DRAM_ADDR_OUT[13] = ALU_RES_IN[13];
  assign OP_MEM[12] = ALU_RES_IN[12];
  assign DRAM_ADDR_OUT[12] = ALU_RES_IN[12];
  assign OP_MEM[11] = ALU_RES_IN[11];
  assign DRAM_ADDR_OUT[11] = ALU_RES_IN[11];
  assign OP_MEM[10] = ALU_RES_IN[10];
  assign DRAM_ADDR_OUT[10] = ALU_RES_IN[10];
  assign OP_MEM[9] = ALU_RES_IN[9];
  assign DRAM_ADDR_OUT[9] = ALU_RES_IN[9];
  assign OP_MEM[8] = ALU_RES_IN[8];
  assign DRAM_ADDR_OUT[8] = ALU_RES_IN[8];
  assign OP_MEM[7] = ALU_RES_IN[7];
  assign DRAM_ADDR_OUT[7] = ALU_RES_IN[7];
  assign OP_MEM[6] = ALU_RES_IN[6];
  assign DRAM_ADDR_OUT[6] = ALU_RES_IN[6];
  assign OP_MEM[5] = ALU_RES_IN[5];
  assign DRAM_ADDR_OUT[5] = ALU_RES_IN[5];
  assign OP_MEM[4] = ALU_RES_IN[4];
  assign DRAM_ADDR_OUT[4] = ALU_RES_IN[4];
  assign OP_MEM[3] = ALU_RES_IN[3];
  assign DRAM_ADDR_OUT[3] = ALU_RES_IN[3];
  assign OP_MEM[2] = ALU_RES_IN[2];
  assign DRAM_ADDR_OUT[2] = ALU_RES_IN[2];
  assign OP_MEM[1] = ALU_RES_IN[1];
  assign DRAM_ADDR_OUT[1] = ALU_RES_IN[1];
  assign OP_MEM[0] = ALU_RES_IN[0];
  assign DRAM_ADDR_OUT[0] = ALU_RES_IN[0];
  assign DRAM_DATA_OUT[31] = B_IN[31];
  assign DRAM_DATA_OUT[30] = B_IN[30];
  assign DRAM_DATA_OUT[29] = B_IN[29];
  assign DRAM_DATA_OUT[28] = B_IN[28];
  assign DRAM_DATA_OUT[27] = B_IN[27];
  assign DRAM_DATA_OUT[26] = B_IN[26];
  assign DRAM_DATA_OUT[25] = B_IN[25];
  assign DRAM_DATA_OUT[24] = B_IN[24];
  assign DRAM_DATA_OUT[23] = B_IN[23];
  assign DRAM_DATA_OUT[22] = B_IN[22];
  assign DRAM_DATA_OUT[21] = B_IN[21];
  assign DRAM_DATA_OUT[20] = B_IN[20];
  assign DRAM_DATA_OUT[19] = B_IN[19];
  assign DRAM_DATA_OUT[18] = B_IN[18];
  assign DRAM_DATA_OUT[17] = B_IN[17];
  assign DRAM_DATA_OUT[16] = B_IN[16];
  assign DRAM_DATA_OUT[15] = B_IN[15];
  assign DRAM_DATA_OUT[14] = B_IN[14];
  assign DRAM_DATA_OUT[13] = B_IN[13];
  assign DRAM_DATA_OUT[12] = B_IN[12];
  assign DRAM_DATA_OUT[11] = B_IN[11];
  assign DRAM_DATA_OUT[10] = B_IN[10];
  assign DRAM_DATA_OUT[9] = B_IN[9];
  assign DRAM_DATA_OUT[8] = B_IN[8];
  assign DRAM_DATA_OUT[7] = B_IN[7];
  assign DRAM_DATA_OUT[6] = B_IN[6];
  assign DRAM_DATA_OUT[5] = B_IN[5];
  assign DRAM_DATA_OUT[4] = B_IN[4];
  assign DRAM_DATA_OUT[3] = B_IN[3];
  assign DRAM_DATA_OUT[2] = B_IN[2];
  assign DRAM_DATA_OUT[1] = B_IN[1];
  assign DRAM_DATA_OUT[0] = B_IN[0];
  assign ADD_WR_MEM[4] = ADD_WR_IN[4];
  assign ADD_WR_MEM[3] = ADD_WR_IN[3];
  assign ADD_WR_MEM[2] = ADD_WR_IN[2];
  assign ADD_WR_MEM[1] = ADD_WR_IN[1];
  assign ADD_WR_MEM[0] = ADD_WR_IN[0];

  regn_N32_2 LMD ( .DIN(DRAM_DATA_IN), .CLK(CLK), .EN(MEM_EN_IN), .RST(RST), 
        .DOUT(DATA_OUT) );
  regn_N5_1 reg0 ( .DIN(ADD_WR_IN), .CLK(CLK), .EN(MEM_EN_IN), .RST(RST), 
        .DOUT(ADD_WR_OUT) );
  regn_N32_1 reg1 ( .DIN(ALU_RES_IN), .CLK(CLK), .EN(MEM_EN_IN), .RST(RST), 
        .DOUT(ALU_RES_OUT) );
  mux41_NBIT32_2 PCsel ( .A(NPC_IN), .B(NPC_REL), .C(NPC_ABS), .D({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(PC_SEL), .Z(PC_OUT) );
endmodule


module ff_2 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n4, n5, n6;

  DFFR_X1 Q_reg ( .D(n4), .CK(CLK), .RN(RST), .Q(Q), .QN(n5) );
  OAI21_X1 U2 ( .B1(n5), .B2(EN), .A(n6), .ZN(n4) );
  NAND2_X1 U3 ( .A1(EN), .A2(D), .ZN(n6) );
endmodule


module mux21_NBIT32_2 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100;

  BUF_X1 U1 ( .A(n68), .Z(n1) );
  BUF_X1 U2 ( .A(n68), .Z(n2) );
  BUF_X1 U3 ( .A(n68), .Z(n3) );
  INV_X1 U4 ( .A(n81), .ZN(Z[20]) );
  AOI22_X1 U5 ( .A1(A[20]), .A2(n2), .B1(B[20]), .B2(S), .ZN(n81) );
  INV_X1 U6 ( .A(n82), .ZN(Z[21]) );
  AOI22_X1 U7 ( .A1(A[21]), .A2(n2), .B1(B[21]), .B2(S), .ZN(n82) );
  INV_X1 U8 ( .A(n83), .ZN(Z[22]) );
  AOI22_X1 U9 ( .A1(A[22]), .A2(n2), .B1(B[22]), .B2(S), .ZN(n83) );
  INV_X1 U10 ( .A(n84), .ZN(Z[23]) );
  AOI22_X1 U11 ( .A1(A[23]), .A2(n2), .B1(B[23]), .B2(S), .ZN(n84) );
  INV_X1 U12 ( .A(n77), .ZN(Z[17]) );
  AOI22_X1 U13 ( .A1(A[17]), .A2(n1), .B1(B[17]), .B2(S), .ZN(n77) );
  INV_X1 U14 ( .A(n78), .ZN(Z[18]) );
  AOI22_X1 U15 ( .A1(A[18]), .A2(n1), .B1(B[18]), .B2(S), .ZN(n78) );
  INV_X1 U16 ( .A(n79), .ZN(Z[19]) );
  AOI22_X1 U17 ( .A1(A[19]), .A2(n1), .B1(B[19]), .B2(S), .ZN(n79) );
  INV_X1 U18 ( .A(n80), .ZN(Z[1]) );
  AOI22_X1 U19 ( .A1(A[1]), .A2(n1), .B1(B[1]), .B2(S), .ZN(n80) );
  INV_X1 U20 ( .A(n73), .ZN(Z[13]) );
  AOI22_X1 U21 ( .A1(A[13]), .A2(n1), .B1(B[13]), .B2(S), .ZN(n73) );
  INV_X1 U22 ( .A(n74), .ZN(Z[14]) );
  AOI22_X1 U23 ( .A1(A[14]), .A2(n1), .B1(B[14]), .B2(S), .ZN(n74) );
  INV_X1 U24 ( .A(n75), .ZN(Z[15]) );
  AOI22_X1 U25 ( .A1(A[15]), .A2(n1), .B1(B[15]), .B2(S), .ZN(n75) );
  INV_X1 U26 ( .A(n76), .ZN(Z[16]) );
  AOI22_X1 U27 ( .A1(A[16]), .A2(n1), .B1(B[16]), .B2(S), .ZN(n76) );
  INV_X1 U28 ( .A(n69), .ZN(Z[0]) );
  AOI22_X1 U29 ( .A1(A[0]), .A2(n1), .B1(B[0]), .B2(S), .ZN(n69) );
  INV_X1 U30 ( .A(n70), .ZN(Z[10]) );
  AOI22_X1 U31 ( .A1(A[10]), .A2(n1), .B1(B[10]), .B2(S), .ZN(n70) );
  INV_X1 U32 ( .A(n71), .ZN(Z[11]) );
  AOI22_X1 U33 ( .A1(A[11]), .A2(n1), .B1(B[11]), .B2(S), .ZN(n71) );
  INV_X1 U34 ( .A(n72), .ZN(Z[12]) );
  AOI22_X1 U35 ( .A1(A[12]), .A2(n1), .B1(B[12]), .B2(S), .ZN(n72) );
  INV_X1 U36 ( .A(n97), .ZN(Z[6]) );
  AOI22_X1 U37 ( .A1(A[6]), .A2(n3), .B1(B[6]), .B2(S), .ZN(n97) );
  INV_X1 U38 ( .A(n98), .ZN(Z[7]) );
  AOI22_X1 U39 ( .A1(A[7]), .A2(n3), .B1(B[7]), .B2(S), .ZN(n98) );
  INV_X1 U40 ( .A(n99), .ZN(Z[8]) );
  AOI22_X1 U41 ( .A1(A[8]), .A2(n3), .B1(B[8]), .B2(S), .ZN(n99) );
  INV_X1 U42 ( .A(n94), .ZN(Z[3]) );
  AOI22_X1 U43 ( .A1(A[3]), .A2(n3), .B1(B[3]), .B2(S), .ZN(n94) );
  INV_X1 U44 ( .A(n95), .ZN(Z[4]) );
  AOI22_X1 U45 ( .A1(A[4]), .A2(n3), .B1(B[4]), .B2(S), .ZN(n95) );
  INV_X1 U46 ( .A(n96), .ZN(Z[5]) );
  AOI22_X1 U47 ( .A1(A[5]), .A2(n3), .B1(B[5]), .B2(S), .ZN(n96) );
  INV_X1 U48 ( .A(n89), .ZN(Z[28]) );
  AOI22_X1 U49 ( .A1(A[28]), .A2(n2), .B1(B[28]), .B2(S), .ZN(n89) );
  INV_X1 U50 ( .A(n90), .ZN(Z[29]) );
  AOI22_X1 U51 ( .A1(A[29]), .A2(n2), .B1(B[29]), .B2(S), .ZN(n90) );
  INV_X1 U52 ( .A(n91), .ZN(Z[2]) );
  AOI22_X1 U53 ( .A1(A[2]), .A2(n2), .B1(B[2]), .B2(S), .ZN(n91) );
  INV_X1 U54 ( .A(n92), .ZN(Z[30]) );
  AOI22_X1 U55 ( .A1(A[30]), .A2(n2), .B1(B[30]), .B2(S), .ZN(n92) );
  INV_X1 U56 ( .A(n85), .ZN(Z[24]) );
  AOI22_X1 U57 ( .A1(A[24]), .A2(n2), .B1(B[24]), .B2(S), .ZN(n85) );
  INV_X1 U58 ( .A(n86), .ZN(Z[25]) );
  AOI22_X1 U59 ( .A1(A[25]), .A2(n2), .B1(B[25]), .B2(S), .ZN(n86) );
  INV_X1 U60 ( .A(n87), .ZN(Z[26]) );
  AOI22_X1 U61 ( .A1(A[26]), .A2(n2), .B1(B[26]), .B2(S), .ZN(n87) );
  INV_X1 U62 ( .A(n88), .ZN(Z[27]) );
  AOI22_X1 U63 ( .A1(A[27]), .A2(n2), .B1(B[27]), .B2(S), .ZN(n88) );
  INV_X1 U64 ( .A(n93), .ZN(Z[31]) );
  AOI22_X1 U65 ( .A1(A[31]), .A2(n3), .B1(B[31]), .B2(S), .ZN(n93) );
  INV_X1 U66 ( .A(n100), .ZN(Z[9]) );
  AOI22_X1 U67 ( .A1(A[9]), .A2(n3), .B1(S), .B2(B[9]), .ZN(n100) );
  INV_X1 U68 ( .A(S), .ZN(n68) );
endmodule


module Writeback ( WB_MUX_SEL, DATA_IN, ALU_RES_IN, ADD_WR_IN, DATA_OUT, 
        ADD_WR_OUT );
  input [31:0] DATA_IN;
  input [31:0] ALU_RES_IN;
  input [4:0] ADD_WR_IN;
  output [31:0] DATA_OUT;
  output [4:0] ADD_WR_OUT;
  input WB_MUX_SEL;

  assign ADD_WR_OUT[4] = ADD_WR_IN[4];
  assign ADD_WR_OUT[3] = ADD_WR_IN[3];
  assign ADD_WR_OUT[2] = ADD_WR_IN[2];
  assign ADD_WR_OUT[1] = ADD_WR_IN[1];
  assign ADD_WR_OUT[0] = ADD_WR_IN[0];

  mux21_NBIT32_2 WBmux ( .A(DATA_IN), .B(ALU_RES_IN), .S(WB_MUX_SEL), .Z(
        DATA_OUT) );
endmodule


module HazardDetection_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \A[0] , n1, n2;
  wire   [32:0] carry;
  assign DIFF[1] = A[1];
  assign DIFF[0] = \A[0] ;
  assign \A[0]  = A[0];

  XNOR2_X1 U1 ( .A(A[4]), .B(carry[4]), .ZN(DIFF[4]) );
  XNOR2_X1 U2 ( .A(A[21]), .B(carry[21]), .ZN(DIFF[21]) );
  XNOR2_X1 U3 ( .A(A[22]), .B(carry[22]), .ZN(DIFF[22]) );
  XNOR2_X1 U4 ( .A(A[23]), .B(carry[23]), .ZN(DIFF[23]) );
  XNOR2_X1 U5 ( .A(A[28]), .B(carry[28]), .ZN(DIFF[28]) );
  XNOR2_X1 U6 ( .A(A[29]), .B(carry[29]), .ZN(DIFF[29]) );
  XNOR2_X1 U7 ( .A(A[30]), .B(carry[30]), .ZN(DIFF[30]) );
  XNOR2_X1 U8 ( .A(A[31]), .B(carry[31]), .ZN(DIFF[31]) );
  NAND2_X1 U9 ( .A1(n1), .A2(n2), .ZN(carry[31]) );
  INV_X1 U10 ( .A(carry[30]), .ZN(n2) );
  INV_X1 U11 ( .A(A[30]), .ZN(n1) );
  XNOR2_X1 U12 ( .A(A[3]), .B(A[2]), .ZN(DIFF[3]) );
  XNOR2_X1 U13 ( .A(A[5]), .B(carry[5]), .ZN(DIFF[5]) );
  XNOR2_X1 U14 ( .A(A[6]), .B(carry[6]), .ZN(DIFF[6]) );
  XNOR2_X1 U15 ( .A(A[7]), .B(carry[7]), .ZN(DIFF[7]) );
  OR2_X1 U16 ( .A1(A[3]), .A2(A[2]), .ZN(carry[4]) );
  XNOR2_X1 U17 ( .A(A[25]), .B(carry[25]), .ZN(DIFF[25]) );
  XNOR2_X1 U18 ( .A(A[9]), .B(carry[9]), .ZN(DIFF[9]) );
  OR2_X1 U19 ( .A1(A[4]), .A2(carry[4]), .ZN(carry[5]) );
  OR2_X1 U20 ( .A1(A[5]), .A2(carry[5]), .ZN(carry[6]) );
  OR2_X1 U21 ( .A1(A[6]), .A2(carry[6]), .ZN(carry[7]) );
  OR2_X1 U22 ( .A1(A[7]), .A2(carry[7]), .ZN(carry[8]) );
  OR2_X1 U23 ( .A1(A[8]), .A2(carry[8]), .ZN(carry[9]) );
  OR2_X1 U24 ( .A1(A[9]), .A2(carry[9]), .ZN(carry[10]) );
  OR2_X1 U25 ( .A1(A[10]), .A2(carry[10]), .ZN(carry[11]) );
  OR2_X1 U26 ( .A1(A[11]), .A2(carry[11]), .ZN(carry[12]) );
  OR2_X1 U27 ( .A1(A[12]), .A2(carry[12]), .ZN(carry[13]) );
  OR2_X1 U28 ( .A1(A[13]), .A2(carry[13]), .ZN(carry[14]) );
  OR2_X1 U29 ( .A1(A[14]), .A2(carry[14]), .ZN(carry[15]) );
  OR2_X1 U30 ( .A1(A[15]), .A2(carry[15]), .ZN(carry[16]) );
  OR2_X1 U31 ( .A1(A[16]), .A2(carry[16]), .ZN(carry[17]) );
  OR2_X1 U32 ( .A1(A[17]), .A2(carry[17]), .ZN(carry[18]) );
  OR2_X1 U33 ( .A1(A[18]), .A2(carry[18]), .ZN(carry[19]) );
  OR2_X1 U34 ( .A1(A[19]), .A2(carry[19]), .ZN(carry[20]) );
  OR2_X1 U35 ( .A1(A[20]), .A2(carry[20]), .ZN(carry[21]) );
  OR2_X1 U36 ( .A1(A[21]), .A2(carry[21]), .ZN(carry[22]) );
  OR2_X1 U37 ( .A1(A[22]), .A2(carry[22]), .ZN(carry[23]) );
  OR2_X1 U38 ( .A1(A[23]), .A2(carry[23]), .ZN(carry[24]) );
  OR2_X1 U39 ( .A1(A[24]), .A2(carry[24]), .ZN(carry[25]) );
  OR2_X1 U40 ( .A1(A[25]), .A2(carry[25]), .ZN(carry[26]) );
  OR2_X1 U41 ( .A1(A[26]), .A2(carry[26]), .ZN(carry[27]) );
  OR2_X1 U42 ( .A1(A[27]), .A2(carry[27]), .ZN(carry[28]) );
  OR2_X1 U43 ( .A1(A[28]), .A2(carry[28]), .ZN(carry[29]) );
  OR2_X1 U44 ( .A1(A[29]), .A2(carry[29]), .ZN(carry[30]) );
  XNOR2_X1 U45 ( .A(A[8]), .B(carry[8]), .ZN(DIFF[8]) );
  XNOR2_X1 U46 ( .A(A[10]), .B(carry[10]), .ZN(DIFF[10]) );
  XNOR2_X1 U47 ( .A(A[11]), .B(carry[11]), .ZN(DIFF[11]) );
  XNOR2_X1 U48 ( .A(A[12]), .B(carry[12]), .ZN(DIFF[12]) );
  XNOR2_X1 U49 ( .A(A[13]), .B(carry[13]), .ZN(DIFF[13]) );
  XNOR2_X1 U50 ( .A(A[14]), .B(carry[14]), .ZN(DIFF[14]) );
  XNOR2_X1 U51 ( .A(A[15]), .B(carry[15]), .ZN(DIFF[15]) );
  XNOR2_X1 U52 ( .A(A[16]), .B(carry[16]), .ZN(DIFF[16]) );
  XNOR2_X1 U53 ( .A(A[17]), .B(carry[17]), .ZN(DIFF[17]) );
  XNOR2_X1 U54 ( .A(A[18]), .B(carry[18]), .ZN(DIFF[18]) );
  XNOR2_X1 U55 ( .A(A[19]), .B(carry[19]), .ZN(DIFF[19]) );
  XNOR2_X1 U56 ( .A(A[20]), .B(carry[20]), .ZN(DIFF[20]) );
  XNOR2_X1 U57 ( .A(A[24]), .B(carry[24]), .ZN(DIFF[24]) );
  XNOR2_X1 U58 ( .A(A[26]), .B(carry[26]), .ZN(DIFF[26]) );
  XNOR2_X1 U59 ( .A(A[27]), .B(carry[27]), .ZN(DIFF[27]) );
  INV_X1 U60 ( .A(A[2]), .ZN(DIFF[2]) );
endmodule


module HazardDetection ( RST, ADD_RS1, ADD_RS2, ADD_WR, DRAM_R, INS_IN, PC_IN, 
        Bubble, HDU_INS_OUT, HDU_PC_OUT, HDU_NPC_OUT );
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [4:0] ADD_WR;
  input [31:0] INS_IN;
  input [31:0] PC_IN;
  output [31:0] HDU_INS_OUT;
  output [31:0] HDU_PC_OUT;
  output [31:0] HDU_NPC_OUT;
  input RST, DRAM_R;
  output Bubble;
  wire   n1, n2, n3, n4, n5, n6, n9, n10, n12, n13, n14, n15, n16;
  assign HDU_INS_OUT[31] = INS_IN[31];
  assign HDU_INS_OUT[30] = INS_IN[30];
  assign HDU_INS_OUT[29] = INS_IN[29];
  assign HDU_INS_OUT[28] = INS_IN[28];
  assign HDU_INS_OUT[27] = INS_IN[27];
  assign HDU_INS_OUT[26] = INS_IN[26];
  assign HDU_INS_OUT[25] = INS_IN[25];
  assign HDU_INS_OUT[24] = INS_IN[24];
  assign HDU_INS_OUT[23] = INS_IN[23];
  assign HDU_INS_OUT[22] = INS_IN[22];
  assign HDU_INS_OUT[21] = INS_IN[21];
  assign HDU_INS_OUT[20] = INS_IN[20];
  assign HDU_INS_OUT[19] = INS_IN[19];
  assign HDU_INS_OUT[18] = INS_IN[18];
  assign HDU_INS_OUT[17] = INS_IN[17];
  assign HDU_INS_OUT[16] = INS_IN[16];
  assign HDU_INS_OUT[15] = INS_IN[15];
  assign HDU_INS_OUT[14] = INS_IN[14];
  assign HDU_INS_OUT[13] = INS_IN[13];
  assign HDU_INS_OUT[12] = INS_IN[12];
  assign HDU_INS_OUT[11] = INS_IN[11];
  assign HDU_INS_OUT[10] = INS_IN[10];
  assign HDU_INS_OUT[9] = INS_IN[9];
  assign HDU_INS_OUT[8] = INS_IN[8];
  assign HDU_INS_OUT[7] = INS_IN[7];
  assign HDU_INS_OUT[6] = INS_IN[6];
  assign HDU_INS_OUT[5] = INS_IN[5];
  assign HDU_INS_OUT[4] = INS_IN[4];
  assign HDU_INS_OUT[3] = INS_IN[3];
  assign HDU_INS_OUT[2] = INS_IN[2];
  assign HDU_INS_OUT[1] = INS_IN[1];
  assign HDU_INS_OUT[0] = INS_IN[0];
  assign HDU_NPC_OUT[31] = PC_IN[31];
  assign HDU_NPC_OUT[30] = PC_IN[30];
  assign HDU_NPC_OUT[29] = PC_IN[29];
  assign HDU_NPC_OUT[28] = PC_IN[28];
  assign HDU_NPC_OUT[27] = PC_IN[27];
  assign HDU_NPC_OUT[26] = PC_IN[26];
  assign HDU_NPC_OUT[25] = PC_IN[25];
  assign HDU_NPC_OUT[24] = PC_IN[24];
  assign HDU_NPC_OUT[23] = PC_IN[23];
  assign HDU_NPC_OUT[22] = PC_IN[22];
  assign HDU_NPC_OUT[21] = PC_IN[21];
  assign HDU_NPC_OUT[20] = PC_IN[20];
  assign HDU_NPC_OUT[19] = PC_IN[19];
  assign HDU_NPC_OUT[18] = PC_IN[18];
  assign HDU_NPC_OUT[17] = PC_IN[17];
  assign HDU_NPC_OUT[16] = PC_IN[16];
  assign HDU_NPC_OUT[15] = PC_IN[15];
  assign HDU_NPC_OUT[14] = PC_IN[14];
  assign HDU_NPC_OUT[13] = PC_IN[13];
  assign HDU_NPC_OUT[12] = PC_IN[12];
  assign HDU_NPC_OUT[11] = PC_IN[11];
  assign HDU_NPC_OUT[10] = PC_IN[10];
  assign HDU_NPC_OUT[9] = PC_IN[9];
  assign HDU_NPC_OUT[8] = PC_IN[8];
  assign HDU_NPC_OUT[7] = PC_IN[7];
  assign HDU_NPC_OUT[6] = PC_IN[6];
  assign HDU_NPC_OUT[5] = PC_IN[5];
  assign HDU_NPC_OUT[4] = PC_IN[4];
  assign HDU_NPC_OUT[3] = PC_IN[3];
  assign HDU_NPC_OUT[2] = PC_IN[2];
  assign HDU_NPC_OUT[1] = PC_IN[1];
  assign HDU_NPC_OUT[0] = PC_IN[0];

  HazardDetection_DW01_sub_0 sub_25 ( .A(PC_IN), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .DIFF(HDU_PC_OUT) );
  AND3_X1 U4 ( .A1(DRAM_R), .A2(n1), .A3(RST), .ZN(Bubble) );
  OAI33_X1 U5 ( .A1(n2), .A2(n3), .A3(n4), .B1(n5), .B2(n6), .B3(n9), .ZN(n1)
         );
  XOR2_X1 U6 ( .A(ADD_WR[4]), .B(ADD_RS2[4]), .Z(n9) );
  XOR2_X1 U8 ( .A(ADD_WR[2]), .B(ADD_RS2[2]), .Z(n6) );
  NAND3_X1 U9 ( .A1(n10), .A2(n12), .A3(n13), .ZN(n5) );
  XNOR2_X1 U11 ( .A(ADD_WR[0]), .B(ADD_RS2[0]), .ZN(n13) );
  XNOR2_X1 U12 ( .A(ADD_WR[1]), .B(ADD_RS2[1]), .ZN(n12) );
  XNOR2_X1 U13 ( .A(ADD_WR[3]), .B(ADD_RS2[3]), .ZN(n10) );
  XOR2_X1 U14 ( .A(ADD_WR[4]), .B(ADD_RS1[4]), .Z(n4) );
  XOR2_X1 U15 ( .A(ADD_WR[2]), .B(ADD_RS1[2]), .Z(n3) );
  NAND3_X1 U16 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n2) );
  XNOR2_X1 U17 ( .A(ADD_WR[0]), .B(ADD_RS1[0]), .ZN(n16) );
  XNOR2_X1 U18 ( .A(ADD_WR[1]), .B(ADD_RS1[1]), .ZN(n15) );
  XNOR2_X1 U19 ( .A(ADD_WR[3]), .B(ADD_RS1[3]), .ZN(n14) );
endmodule


module Datapath ( CLK, RST, INS_IN, DATA_IN, REG_LATCH_EN, RD1, RD2, MUX_A_SEL, 
        MUX_B_SEL, .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , 
        \ALU_OPC[0] }), ALU_OUTREG_EN, JUMP_TYPE, DRAM_R_IN, MEM_EN_IN, 
        DRAM_W_IN, RF_WE, DRAM_EN_IN, WB_MUX_SEL, INS_OUT, IRAM_ADDR_OUT, 
        DRAM_ADDR_OUT, DATA_OUT, DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, 
        Bubble_out );
  input [31:0] INS_IN;
  input [31:0] DATA_IN;
  input [1:0] MUX_B_SEL;
  input [1:0] JUMP_TYPE;
  output [31:0] INS_OUT;
  output [31:0] IRAM_ADDR_OUT;
  output [31:0] DRAM_ADDR_OUT;
  output [31:0] DATA_OUT;
  input CLK, RST, REG_LATCH_EN, RD1, RD2, MUX_A_SEL, \ALU_OPC[3] ,
         \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] , ALU_OUTREG_EN, DRAM_R_IN,
         MEM_EN_IN, DRAM_W_IN, RF_WE, DRAM_EN_IN, WB_MUX_SEL;
  output DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble_out;
  wire   n2, ZERO_FLAG_EX, RF_WE_WB, DRAM_R_MEM;
  wire   [3:0] ALU_OPC;
  wire   [31:0] PC_MEM_OUT;
  wire   [31:0] sig_HDU_INS_OUT;
  wire   [31:0] sig_HDU_PC_OUT;
  wire   [31:0] sig_HDU_NPC_OUT;
  wire   [31:0] PC_FETCH_OUT;
  wire   [31:0] NPC_FETCH_OUT;
  wire   [4:0] ADD_WR_WB;
  wire   [31:0] OP_WB;
  wire   [31:0] PC_DECODE_OUT;
  wire   [31:0] A_DECODE_OUT;
  wire   [31:0] B_DECODE_OUT;
  wire   [31:0] IMM_DECODE_OUT;
  wire   [4:0] ADD_RS1_HDU;
  wire   [4:0] ADD_RS2_HDU;
  wire   [4:0] ADD_WR_DECODE_OUT;
  wire   [4:0] ADD_RS1_DECODE_OUT;
  wire   [4:0] ADD_RS2_DECODE_OUT;
  wire   [4:0] ADD_WR_MEM;
  wire   [31:0] OP_MEM;
  wire   [1:0] PC_SEL_EX;
  wire   [31:0] NPC_ABS_EX;
  wire   [31:0] NPC_REL_EX;
  wire   [31:0] ALU_RES_EX;
  wire   [31:0] B_EX_OUT;
  wire   [4:0] ADD_WR_EX_OUT;
  wire   [31:0] DATA_MEM_OUT;
  wire   [31:0] ALU_RES_MEM;
  wire   [4:0] ADD_WR_MEM_OUT;

  Fetch FetchStage ( .CLK(CLK), .RST(RST), .ZERO_FLAG(ZERO_FLAG_EX), .PC_EXT(
        PC_MEM_OUT), .INS_IN(INS_IN), .Bubble_in(Bubble_out), .HDU_INS_IN(
        sig_HDU_INS_OUT), .HDU_PC_IN(sig_HDU_PC_OUT), .HDU_NPC_IN(
        sig_HDU_NPC_OUT), .PC_OUT(PC_FETCH_OUT), .ADDR_OUT(IRAM_ADDR_OUT), 
        .NPC_OUT(NPC_FETCH_OUT), .INS_OUT(INS_OUT) );
  Decode DecodeStage ( .CLK(CLK), .RST(RST), .REG_LATCH_EN(REG_LATCH_EN), 
        .RD1(RD1), .RD2(RD2), .RF_WE(RF_WE_WB), .ZERO_FLAG(ZERO_FLAG_EX), 
        .PC_IN(PC_FETCH_OUT), .INS_IN(INS_OUT), .ADD_WR(ADD_WR_WB), 
        .DATA_WR_IN(OP_WB), .PC_OUT(PC_DECODE_OUT), .A_OUT(A_DECODE_OUT), 
        .B_OUT(B_DECODE_OUT), .IMM_OUT(IMM_DECODE_OUT), .ADD_RS1_HDU(
        ADD_RS1_HDU), .ADD_RS2_HDU(ADD_RS2_HDU), .ADD_WR_OUT(ADD_WR_DECODE_OUT), .ADD_RS1_OUT(ADD_RS1_DECODE_OUT), .ADD_RS2_OUT(ADD_RS2_DECODE_OUT) );
  Execute ExecuteStage ( .CLK(CLK), .RST(RST), .MUX_A_SEL(MUX_A_SEL), 
        .MUX_B_SEL(MUX_B_SEL), .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , 
        \ALU_OPC[1] , \ALU_OPC[0] }), .ALU_OUTREG_EN(ALU_OUTREG_EN), 
        .JUMP_TYPE(JUMP_TYPE), .PC_IN(PC_DECODE_OUT), .A_IN(A_DECODE_OUT), 
        .B_IN(B_DECODE_OUT), .IMM_IN(IMM_DECODE_OUT), .ADD_WR_IN(
        ADD_WR_DECODE_OUT), .ADD_RS1_IN(ADD_RS1_DECODE_OUT), .ADD_RS2_IN(
        ADD_RS2_DECODE_OUT), .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_WB(ADD_WR_WB), 
        .RF_WE_MEM(RF_WE), .RF_WE_WB(RF_WE_WB), .OP_MEM(OP_MEM), .OP_WB(OP_WB), 
        .PC_SEL(PC_SEL_EX), .ZERO_FLAG(ZERO_FLAG_EX), .NPC_ABS(NPC_ABS_EX), 
        .NPC_REL(NPC_REL_EX), .ALU_RES(ALU_RES_EX), .B_OUT(B_EX_OUT), 
        .ADD_WR_OUT(ADD_WR_EX_OUT) );
  ff_0 DRAM_R_ff ( .D(DRAM_R_IN), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(
        DRAM_R_MEM) );
  Memory MemoryStage ( .CLK(CLK), .RST(RST), .MEM_EN_IN(MEM_EN_IN), 
        .DRAM_R_IN(DRAM_R_MEM), .DRAM_W_IN(DRAM_W_IN), .DRAM_EN_IN(DRAM_EN_IN), 
        .PC_SEL(PC_SEL_EX), .NPC_IN(NPC_FETCH_OUT), .NPC_ABS(NPC_ABS_EX), 
        .NPC_REL(NPC_REL_EX), .ALU_RES_IN(ALU_RES_EX), .B_IN(B_EX_OUT), 
        .ADD_WR_IN(ADD_WR_EX_OUT), .DRAM_DATA_IN(DATA_IN), .PC_OUT(PC_MEM_OUT), 
        .DRAM_EN_OUT(DRAM_EN_OUT), .DRAM_R_OUT(DRAM_R_OUT), .DRAM_W_OUT(
        DRAM_W_OUT), .DRAM_ADDR_OUT(DRAM_ADDR_OUT), .DRAM_DATA_OUT(DATA_OUT), 
        .DATA_OUT(DATA_MEM_OUT), .ALU_RES_OUT(ALU_RES_MEM), .OP_MEM(OP_MEM), 
        .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_OUT(ADD_WR_MEM_OUT) );
  ff_2 RF_WE_ff ( .D(RF_WE), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(RF_WE_WB) );
  Writeback WritebackStage ( .WB_MUX_SEL(WB_MUX_SEL), .DATA_IN(DATA_MEM_OUT), 
        .ALU_RES_IN(ALU_RES_MEM), .ADD_WR_IN(ADD_WR_MEM_OUT), .DATA_OUT(OP_WB), 
        .ADD_WR_OUT(ADD_WR_WB) );
  HazardDetection HDU ( .RST(RST), .ADD_RS1(ADD_RS1_HDU), .ADD_RS2(ADD_RS2_HDU), .ADD_WR(ADD_WR_DECODE_OUT), .DRAM_R(DRAM_R_IN), .INS_IN(INS_OUT), .PC_IN(
        PC_FETCH_OUT), .Bubble(n2), .HDU_INS_OUT(sig_HDU_INS_OUT), 
        .HDU_PC_OUT(sig_HDU_PC_OUT), .HDU_NPC_OUT(sig_HDU_NPC_OUT) );
  BUF_X1 U2 ( .A(n2), .Z(Bubble_out) );
endmodule


module hardwired_cu_NBIT32 ( REG_LATCH_EN, RD1, RD2, MUX_A_SEL, MUX_B_SEL, 
    .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), 
        ALU_OUTREG_EN, DRAM_R_IN, JUMP_TYPE, MEM_EN_IN, DRAM_W_IN, RF_WE, 
        DRAM_EN_IN, WB_MUX_SEL, INS_IN, Bubble, Clk, Rst );
  output [1:0] MUX_B_SEL;
  output [1:0] JUMP_TYPE;
  input [31:0] INS_IN;
  input Bubble, Clk, Rst;
  output REG_LATCH_EN, RD1, RD2, MUX_A_SEL, \ALU_OPC[3] , \ALU_OPC[2] ,
         \ALU_OPC[1] , \ALU_OPC[0] , ALU_OUTREG_EN, DRAM_R_IN, MEM_EN_IN,
         DRAM_W_IN, RF_WE, DRAM_EN_IN, WB_MUX_SEL;
  wire   INS_IN_31, INS_IN_30, INS_IN_29, INS_IN_28, INS_IN_27, INS_IN_26, N24,
         N25, N26, N27, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n58,
         n59, n60, n61, n62, n63, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18;
  wire   [3:0] ALU_OPC;
  wire   [3:0] AluOP_E;
  assign REG_LATCH_EN = 1'b0;
  assign RD1 = 1'b0;
  assign RD2 = 1'b0;
  assign MUX_A_SEL = 1'b0;
  assign MUX_B_SEL[1] = 1'b0;
  assign MUX_B_SEL[0] = 1'b0;
  assign ALU_OUTREG_EN = 1'b0;
  assign DRAM_R_IN = 1'b0;
  assign JUMP_TYPE[1] = 1'b0;
  assign JUMP_TYPE[0] = 1'b0;
  assign MEM_EN_IN = 1'b0;
  assign DRAM_W_IN = 1'b0;
  assign RF_WE = 1'b0;
  assign DRAM_EN_IN = 1'b0;
  assign WB_MUX_SEL = 1'b0;
  assign INS_IN_31 = INS_IN[31];
  assign INS_IN_30 = INS_IN[30];
  assign INS_IN_29 = INS_IN[29];
  assign INS_IN_28 = INS_IN[28];
  assign INS_IN_27 = INS_IN[27];
  assign INS_IN_26 = INS_IN[26];

  DFFR_X1 \AluOP_E_reg[3]  ( .D(N27), .CK(Clk), .RN(Rst), .Q(AluOP_E[3]) );
  DFFR_X1 \AluOP_E_reg[2]  ( .D(N26), .CK(Clk), .RN(Rst), .Q(AluOP_E[2]) );
  DFFR_X1 \AluOP_E_reg[1]  ( .D(N25), .CK(Clk), .RN(Rst), .Q(AluOP_E[1]) );
  DFFR_X1 \AluOP_E_reg[0]  ( .D(N24), .CK(Clk), .RN(Rst), .Q(AluOP_E[0]) );
  XOR2_X1 U74 ( .A(n2), .B(INS_IN[1]), .Z(n33) );
  NAND3_X1 U75 ( .A1(n16), .A2(n13), .A3(INS_IN_30), .ZN(n37) );
  OAI33_X1 U76 ( .A1(n26), .A2(n13), .A3(n17), .B1(n46), .B2(INS_IN_30), .B3(
        INS_IN_28), .ZN(n43) );
  OAI33_X1 U77 ( .A1(n24), .A2(n25), .A3(n17), .B1(n3), .B2(n8), .B3(n34), 
        .ZN(n50) );
  OAI33_X1 U78 ( .A1(n12), .A2(n56), .A3(n11), .B1(n27), .B2(INS_IN_30), .B3(
        n25), .ZN(n55) );
  NAND3_X1 U79 ( .A1(n51), .A2(n7), .A3(INS_IN[5]), .ZN(n35) );
  OAI33_X1 U80 ( .A1(n58), .A2(n13), .A3(n17), .B1(n59), .B2(n39), .B3(n6), 
        .ZN(n48) );
  NAND3_X1 U81 ( .A1(INS_IN[3]), .A2(n51), .A3(INS_IN[5]), .ZN(n39) );
  NAND3_X1 U82 ( .A1(n15), .A2(n18), .A3(INS_IN_28), .ZN(n24) );
  NAND3_X1 U83 ( .A1(n10), .A2(n13), .A3(n63), .ZN(n34) );
  NAND3_X1 U84 ( .A1(n16), .A2(n17), .A3(INS_IN_28), .ZN(n36) );
  DFFR_X1 \ALU_OPC_reg[3]  ( .D(AluOP_E[3]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[3]) );
  DFFR_X1 \ALU_OPC_reg[2]  ( .D(AluOP_E[2]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[2]) );
  DFFR_X1 \ALU_OPC_reg[1]  ( .D(AluOP_E[1]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[1]) );
  DFFR_X1 \ALU_OPC_reg[0]  ( .D(AluOP_E[0]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[0]) );
  INV_X1 U18 ( .A(n25), .ZN(n10) );
  NAND2_X1 U19 ( .A1(n12), .A2(n11), .ZN(n25) );
  AOI21_X1 U20 ( .B1(n40), .B2(n41), .A(Bubble), .ZN(N25) );
  AOI211_X1 U21 ( .C1(n14), .C2(n10), .A(n38), .B(n48), .ZN(n40) );
  AOI221_X1 U22 ( .B1(n42), .B2(n5), .C1(n16), .C2(n43), .A(n44), .ZN(n41) );
  INV_X1 U23 ( .A(n47), .ZN(n5) );
  AOI21_X1 U24 ( .B1(n28), .B2(n29), .A(Bubble), .ZN(N26) );
  AOI21_X1 U25 ( .B1(n20), .B2(n6), .A(n38), .ZN(n28) );
  NOR3_X1 U26 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n29) );
  AOI21_X1 U27 ( .B1(n36), .B2(n37), .A(n26), .ZN(n30) );
  INV_X1 U28 ( .A(n36), .ZN(n14) );
  INV_X1 U29 ( .A(n27), .ZN(n16) );
  OR2_X1 U30 ( .A1(n49), .A2(n50), .ZN(n38) );
  INV_X1 U31 ( .A(n52), .ZN(n3) );
  INV_X1 U32 ( .A(n51), .ZN(n8) );
  NAND2_X1 U33 ( .A1(n16), .A2(n10), .ZN(n58) );
  OR3_X1 U34 ( .A1(INS_IN[0]), .A2(INS_IN[1]), .A3(n34), .ZN(n59) );
  NOR4_X1 U35 ( .A1(INS_IN[6]), .A2(INS_IN[4]), .A3(INS_IN[10]), .A4(n62), 
        .ZN(n51) );
  OR3_X1 U36 ( .A1(INS_IN[9]), .A2(INS_IN[8]), .A3(INS_IN[7]), .ZN(n62) );
  NAND2_X1 U37 ( .A1(INS_IN_27), .A2(n11), .ZN(n46) );
  NOR3_X1 U38 ( .A1(INS_IN_29), .A2(INS_IN_31), .A3(INS_IN_30), .ZN(n63) );
  NOR4_X1 U39 ( .A1(n2), .A2(n39), .A3(n34), .A4(INS_IN[1]), .ZN(n20) );
  NOR4_X1 U40 ( .A1(n6), .A2(INS_IN[0]), .A3(INS_IN[3]), .A4(INS_IN[5]), .ZN(
        n52) );
  NOR4_X1 U41 ( .A1(n33), .A2(n34), .A3(n6), .A4(n35), .ZN(n32) );
  NOR4_X1 U42 ( .A1(INS_IN[1]), .A2(n4), .A3(n34), .A4(n6), .ZN(n44) );
  INV_X1 U43 ( .A(n45), .ZN(n4) );
  OAI21_X1 U44 ( .B1(n35), .B2(INS_IN[0]), .A(n39), .ZN(n45) );
  NOR3_X1 U45 ( .A1(n34), .A2(INS_IN[0]), .A3(n35), .ZN(n42) );
  INV_X1 U46 ( .A(INS_IN[3]), .ZN(n7) );
  NOR3_X1 U47 ( .A1(n36), .A2(INS_IN_26), .A3(n12), .ZN(n31) );
  INV_X1 U48 ( .A(INS_IN[2]), .ZN(n6) );
  INV_X1 U49 ( .A(INS_IN_30), .ZN(n17) );
  AOI22_X1 U50 ( .A1(n15), .A2(n18), .B1(INS_IN_31), .B2(n17), .ZN(n56) );
  NAND2_X1 U51 ( .A1(INS_IN_26), .A2(n12), .ZN(n26) );
  INV_X1 U52 ( .A(INS_IN_27), .ZN(n12) );
  AOI21_X1 U53 ( .B1(n53), .B2(n54), .A(Bubble), .ZN(N24) );
  AOI211_X1 U54 ( .C1(n14), .C2(n10), .A(n49), .B(n23), .ZN(n53) );
  AOI221_X1 U55 ( .B1(n42), .B2(n47), .C1(n55), .C2(n13), .A(n31), .ZN(n54) );
  INV_X1 U56 ( .A(INS_IN_28), .ZN(n13) );
  NAND2_X1 U57 ( .A1(INS_IN_29), .A2(n18), .ZN(n27) );
  OR2_X1 U58 ( .A1(n48), .A2(n1), .ZN(n23) );
  NOR3_X1 U59 ( .A1(n26), .A2(INS_IN_30), .A3(n24), .ZN(n1) );
  NAND2_X1 U60 ( .A1(INS_IN[1]), .A2(n6), .ZN(n47) );
  INV_X1 U61 ( .A(INS_IN_31), .ZN(n18) );
  INV_X1 U62 ( .A(INS_IN_26), .ZN(n11) );
  NAND2_X1 U63 ( .A1(n60), .A2(n61), .ZN(n49) );
  OR4_X1 U64 ( .A1(n12), .A2(n24), .A3(n17), .A4(INS_IN_26), .ZN(n61) );
  NAND4_X1 U65 ( .A1(INS_IN[1]), .A2(n52), .A3(n9), .A4(n51), .ZN(n60) );
  INV_X1 U66 ( .A(n34), .ZN(n9) );
  NOR2_X1 U67 ( .A1(Bubble), .A2(n19), .ZN(N27) );
  NOR4_X1 U68 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n19) );
  NOR3_X1 U69 ( .A1(n26), .A2(n27), .A3(n17), .ZN(n21) );
  NOR3_X1 U70 ( .A1(n24), .A2(INS_IN_30), .A3(n25), .ZN(n22) );
  INV_X1 U71 ( .A(INS_IN[0]), .ZN(n2) );
  INV_X1 U72 ( .A(INS_IN_29), .ZN(n15) );
endmodule


module DLX ( Clk, Rst );
  input Clk, Rst;
  wire   DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble;
  wire   [31:0] INS_IN;
  wire   [31:0] DATA_IN;
  wire   [1:0] MUX_B_SEL;
  wire   [3:0] ALU_OPC;
  wire   [1:0] JUMP_TYPE;
  wire   [31:0] IRAM_ADDR_OUT;
  wire   [31:0] DRAM_ADDR_OUT;
  wire   [31:0] DATA_OUT;

  Datapath DP ( .CLK(Clk), .RST(Rst), .INS_IN(INS_IN), .DATA_IN(DATA_IN), 
        .REG_LATCH_EN(1'b0), .RD1(1'b0), .RD2(1'b0), .MUX_A_SEL(1'b0), 
        .MUX_B_SEL({1'b0, 1'b0}), .ALU_OPC(ALU_OPC), .ALU_OUTREG_EN(1'b0), 
        .JUMP_TYPE({1'b0, 1'b0}), .DRAM_R_IN(1'b0), .MEM_EN_IN(1'b0), 
        .DRAM_W_IN(1'b0), .RF_WE(1'b0), .DRAM_EN_IN(1'b0), .WB_MUX_SEL(1'b0), 
        .IRAM_ADDR_OUT(IRAM_ADDR_OUT), .DRAM_ADDR_OUT(DRAM_ADDR_OUT), 
        .DATA_OUT(DATA_OUT), .DRAM_EN_OUT(DRAM_EN_OUT), .DRAM_R_OUT(DRAM_R_OUT), .DRAM_W_OUT(DRAM_W_OUT), .Bubble_out(Bubble) );
  hardwired_cu_NBIT32 CU ( .ALU_OPC(ALU_OPC), .INS_IN(INS_IN), .Bubble(Bubble), 
        .Clk(Clk), .Rst(Rst) );
  IRAM IRAM_I ( .Rst(Rst), .Addr(IRAM_ADDR_OUT), .Iout(INS_IN) );
  DRAM DRAM_I ( .En(DRAM_EN_OUT), .Rst(Rst), .ADDR_IN(DRAM_ADDR_OUT), 
        .DATA_IN(DATA_OUT), .DRAM_W(DRAM_W_OUT), .DRAM_R(DRAM_R_OUT), 
        .DATA_OUT(DATA_IN) );
endmodule

