
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type VHDLOUT_TYPE is range 0 to 5;
type aluOp is (NOP, ADDS, SUBS, ANDS, ORS, XORS, SLLS, SRLS, BEQZS, BNEZS, 
   SGES, SLES, NEQS);
attribute ENUM_ENCODING of aluOp : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010 1011 1100";
   
   -- Declarations for conversion functions.
   function integer_to_unsigned(arg, size : in INTEGER) return std_logic_vector
               ;
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 4 )) 
               return aluOp;
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX;

package body CONV_PACK_DLX is
   
   -- integer type to std_logic_vector function
   function integer_to_unsigned(arg, size : in INTEGER) return std_logic_vector
   is 
      variable result: std_logic_vector(size-1 downto 0);
      variable temp: INTEGER;
      -- synopsys built_in SYN_INTEGER_TO_UNSIGNED
   begin
      temp := arg;
      for i in 0 to size-1 loop
         if (temp mod 2) = 1 then
            result(i) := '1';
         else
            result(i) := '0';
         end if;
         temp := temp / 2;
      end loop;
      return result;
   end;
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 4 )) 
   return aluOp is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "0000" => return NOP;
         when "0001" => return ADDS;
         when "0010" => return SUBS;
         when "0011" => return ANDS;
         when "0100" => return ORS;
         when "0101" => return XORS;
         when "0110" => return SLLS;
         when "0111" => return SRLS;
         when "1000" => return BEQZS;
         when "1001" => return BNEZS;
         when "1010" => return SGES;
         when "1011" => return SLES;
         when "1100" => return NEQS;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "0000";
         when ADDS => return "0001";
         when SUBS => return "0010";
         when ANDS => return "0011";
         when ORS => return "0100";
         when XORS => return "0101";
         when SLLS => return "0110";
         when SRLS => return "0111";
         when BEQZS => return "1000";
         when BNEZS => return "1001";
         when SGES => return "1010";
         when SLES => return "1011";
         when NEQS => return "1100";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Fetch_DW01_add_3 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Fetch_DW01_add_3;

architecture SYN_cla of Fetch_DW01_add_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, n1, n2, n3, n4, n5, n6, 
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116 : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U2 : XNOR2_X1 port map( A => n116, B => n69, ZN => SUM_5_port);
   U3 : XOR2_X1 port map( A => n1, B => n3, Z => SUM_14_port);
   U4 : AND2_X1 port map( A1 => n109, A2 => n59, ZN => n1);
   U5 : AND2_X1 port map( A1 => n2, A2 => n109, ZN => n107);
   U6 : AND2_X1 port map( A1 => n59, A2 => n3, ZN => n2);
   U7 : INV_X1 port map( A => n108, ZN => n3);
   U8 : BUF_X1 port map( A => n58, Z => n26);
   U9 : AND2_X1 port map( A1 => A(24), A2 => A(25), ZN => n4);
   U10 : AND2_X1 port map( A1 => n70, A2 => n31, ZN => n5);
   U11 : BUF_X1 port map( A => A(4), Z => n20);
   U12 : INV_X1 port map( A => n10, ZN => n6);
   U13 : XOR2_X1 port map( A => n7, B => n35, Z => SUM_9_port);
   U14 : NOR2_X1 port map( A1 => n76, A2 => n22, ZN => n7);
   U15 : CLKBUF_X1 port map( A => A(16), Z => n8);
   U16 : AND2_X1 port map( A1 => n57, A2 => n41, ZN => n9);
   U17 : INV_X1 port map( A => n53, ZN => n10);
   U18 : AND2_X1 port map( A1 => n69, A2 => n11, ZN => n13);
   U19 : NOR2_X1 port map( A1 => n116, A2 => n10, ZN => n11);
   U20 : XOR2_X1 port map( A => n12, B => n72, Z => SUM_8_port);
   U21 : NOR2_X1 port map( A1 => n76, A2 => n75, ZN => n12);
   U22 : NOR2_X1 port map( A1 => n78, A2 => n116, ZN => n77);
   U23 : XOR2_X1 port map( A => n13, B => n36, Z => SUM_7_port);
   U24 : XOR2_X1 port map( A => A(12), B => n14, Z => SUM_12_port);
   U25 : NOR2_X1 port map( A1 => n62, A2 => n19, ZN => n14);
   U26 : XNOR2_X1 port map( A => n15, B => n111, ZN => SUM_13_port);
   U27 : AND2_X1 port map( A1 => n23, A2 => n12, ZN => n15);
   U28 : BUF_X1 port map( A => n113, Z => n16);
   U29 : NOR2_X1 port map( A1 => n76, A2 => n17, ZN => n59);
   U30 : NAND2_X1 port map( A1 => n18, A2 => n60, ZN => n17);
   U31 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n18);
   U32 : AND2_X1 port map( A1 => A(2), A2 => A(3), ZN => n79);
   U33 : NAND4_X1 port map( A1 => n112, A2 => n46, A3 => n31, A4 => n35, ZN => 
                           n19);
   U34 : XOR2_X1 port map( A => n21, B => n43, Z => SUM_21_port);
   U35 : AND2_X1 port map( A1 => n26, A2 => n9, ZN => n21);
   U36 : NAND2_X1 port map( A1 => n18, A2 => A(8), ZN => n22);
   U37 : NOR2_X1 port map( A1 => n19, A2 => n105, ZN => n23);
   U38 : NAND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n24);
   U39 : CLKBUF_X1 port map( A => A(2), Z => n25);
   U40 : XOR2_X1 port map( A => n54, B => A(31), Z => SUM_31_port);
   U41 : CLKBUF_X1 port map( A => n57, Z => n27);
   U42 : XNOR2_X1 port map( A => n28, B => n88, ZN => SUM_29_port);
   U43 : NOR2_X1 port map( A1 => n71, A2 => n86, ZN => n28);
   U44 : XOR2_X1 port map( A => n48, B => n29, Z => SUM_17_port);
   U45 : AND2_X1 port map( A1 => n26, A2 => n8, ZN => n29);
   U46 : NAND2_X1 port map( A1 => n114, A2 => n115, ZN => n30);
   U47 : BUF_X1 port map( A => A(10), Z => n31);
   U48 : AND2_X1 port map( A1 => n45, A2 => n85, ZN => n89);
   U49 : AND2_X1 port map( A1 => n61, A2 => n4, ZN => n92);
   U50 : NOR3_X1 port map( A1 => n83, A2 => n82, A3 => n81, ZN => n54);
   U51 : CLKBUF_X1 port map( A => A(3), Z => n32);
   U52 : CLKBUF_X1 port map( A => A(15), Z => n33);
   U53 : CLKBUF_X1 port map( A => A(23), Z => n34);
   U54 : BUF_X1 port map( A => A(9), Z => n35);
   U55 : CLKBUF_X1 port map( A => A(7), Z => n36);
   U56 : CLKBUF_X1 port map( A => A(22), Z => n37);
   U57 : XNOR2_X1 port map( A => n38, B => n90, ZN => SUM_28_port);
   U58 : NOR2_X1 port map( A1 => n71, A2 => n44, ZN => n38);
   U59 : AND2_X1 port map( A1 => n4, A2 => A(26), ZN => n39);
   U60 : AND2_X1 port map( A1 => n61, A2 => n39, ZN => n66);
   U61 : XOR2_X1 port map( A => n40, B => n41, Z => SUM_20_port);
   U62 : AND2_X1 port map( A1 => n27, A2 => n58, ZN => n40);
   U63 : AND2_X1 port map( A1 => n101, A2 => n102, ZN => n45);
   U64 : BUF_X1 port map( A => A(20), Z => n41);
   U65 : NOR2_X1 port map( A1 => n87, A2 => n90, ZN => n42);
   U66 : CLKBUF_X1 port map( A => A(21), Z => n43);
   U67 : CLKBUF_X1 port map( A => n87, Z => n44);
   U68 : INV_X1 port map( A => n113, ZN => n46);
   U69 : AND3_X1 port map( A1 => A(22), A2 => A(21), A3 => A(23), ZN => n47);
   U70 : AND2_X1 port map( A1 => n47, A2 => n41, ZN => n63);
   U71 : CLKBUF_X1 port map( A => A(17), Z => n48);
   U72 : NAND2_X1 port map( A1 => A(19), A2 => A(18), ZN => n96);
   U73 : AND2_X1 port map( A1 => A(5), A2 => A(4), ZN => n114);
   U74 : CLKBUF_X1 port map( A => A(6), Z => n53);
   U75 : AND2_X1 port map( A1 => n63, A2 => n94, ZN => n49);
   U76 : OR2_X1 port map( A1 => n87, A2 => n90, ZN => n86);
   U77 : AND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n50);
   U78 : AND2_X1 port map( A1 => n45, A2 => n50, ZN => n64);
   U79 : XNOR2_X1 port map( A => n92, B => n93, ZN => SUM_26_port);
   U80 : AND3_X1 port map( A1 => n45, A2 => n9, A3 => n43, ZN => n51);
   U81 : AND3_X1 port map( A1 => n9, A2 => n45, A3 => n43, ZN => n65);
   U82 : XOR2_X1 port map( A => n52, B => A(25), Z => SUM_25_port);
   U83 : AND2_X1 port map( A1 => A(24), A2 => n89, ZN => n52);
   U84 : NOR2_X1 port map( A1 => n55, A2 => n56, ZN => n102);
   U85 : NAND4_X1 port map( A1 => A(3), A2 => A(5), A3 => A(6), A4 => A(7), ZN 
                           => n55);
   U86 : NAND3_X1 port map( A1 => A(4), A2 => A(2), A3 => A(9), ZN => n56);
   U87 : NOR2_X1 port map( A1 => n96, A2 => n97, ZN => n57);
   U88 : AND2_X1 port map( A1 => A(7), A2 => A(6), ZN => n115);
   U89 : AND2_X1 port map( A1 => n101, A2 => n102, ZN => n58);
   U90 : INV_X1 port map( A => n111, ZN => n60);
   U91 : AND2_X1 port map( A1 => n45, A2 => n85, ZN => n61);
   U92 : OR2_X1 port map( A1 => n30, A2 => n75, ZN => n62);
   U93 : NOR2_X1 port map( A1 => n110, A2 => n105, ZN => n109);
   U94 : AND2_X1 port map( A1 => n63, A2 => n94, ZN => n85);
   U95 : XNOR2_X1 port map( A => n95, B => n34, ZN => SUM_23_port);
   U96 : NOR2_X1 port map( A1 => n30, A2 => n75, ZN => n73);
   U97 : NOR2_X1 port map( A1 => n24, A2 => n96, ZN => n94);
   U98 : INV_X1 port map( A => n74, ZN => n72);
   U99 : AND2_X1 port map( A1 => n64, A2 => n98, ZN => n67);
   U100 : INV_X1 port map( A => A(27), ZN => n91);
   U101 : INV_X1 port map( A => n33, ZN => n106);
   U102 : INV_X1 port map( A => n74, ZN => n112);
   U103 : XNOR2_X1 port map( A => n68, B => n80, ZN => SUM_30_port);
   U104 : OR2_X1 port map( A1 => n83, A2 => n82, ZN => n68);
   U105 : XOR2_X1 port map( A => n64, B => n98, Z => SUM_18_port);
   U106 : XOR2_X1 port map( A => n26, B => n8, Z => SUM_16_port);
   U107 : XOR2_X1 port map( A => n77, B => n6, Z => SUM_6_port);
   U108 : XOR2_X1 port map( A => n25, B => n32, Z => SUM_3_port);
   U109 : XOR2_X1 port map( A => n18, B => n20, Z => SUM_4_port);
   U110 : XOR2_X1 port map( A => n70, B => n31, Z => SUM_10_port);
   U111 : XOR2_X1 port map( A => n89, B => A(24), Z => SUM_24_port);
   U112 : XOR2_X1 port map( A => n51, B => n37, Z => SUM_22_port);
   U113 : INV_X1 port map( A => n100, ZN => n98);
   U114 : AND2_X1 port map( A1 => n79, A2 => n20, ZN => n69);
   U115 : INV_X1 port map( A => A(26), ZN => n93);
   U116 : INV_X1 port map( A => A(28), ZN => n90);
   U117 : INV_X1 port map( A => n81, ZN => n80);
   U118 : INV_X1 port map( A => A(30), ZN => n81);
   U119 : AND3_X1 port map( A1 => n73, A2 => n35, A3 => A(8), ZN => n70);
   U120 : INV_X1 port map( A => n88, ZN => n84);
   U121 : INV_X1 port map( A => A(29), ZN => n88);
   U122 : INV_X1 port map( A => A(11), ZN => n113);
   U123 : INV_X1 port map( A => A(8), ZN => n74);
   U124 : INV_X1 port map( A => n25, ZN => SUM_2_port);
   U125 : NAND4_X1 port map( A1 => A(24), A2 => A(25), A3 => A(26), A4 => A(27)
                           , ZN => n87);
   U126 : INV_X1 port map( A => A(19), ZN => n99);
   U127 : INV_X1 port map( A => A(18), ZN => n100);
   U128 : NAND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n97);
   U129 : XNOR2_X1 port map( A => n66, B => n91, ZN => SUM_27_port);
   U130 : INV_X1 port map( A => A(13), ZN => n111);
   U131 : NAND2_X1 port map( A1 => n65, A2 => n37, ZN => n95);
   U132 : INV_X1 port map( A => A(5), ZN => n116);
   U133 : XNOR2_X1 port map( A => n67, B => n99, ZN => SUM_19_port);
   U134 : NAND2_X1 port map( A1 => n114, A2 => n115, ZN => n76);
   U135 : NAND2_X1 port map( A1 => n58, A2 => n85, ZN => n71);
   U136 : NOR2_X1 port map( A1 => n103, A2 => n104, ZN => n101);
   U137 : INV_X1 port map( A => A(12), ZN => n105);
   U138 : NAND4_X1 port map( A1 => n112, A2 => n46, A3 => n31, A4 => n35, ZN =>
                           n110);
   U139 : NAND4_X1 port map( A1 => A(14), A2 => A(15), A3 => A(13), A4 => A(10)
                           , ZN => n103);
   U140 : XNOR2_X1 port map( A => n5, B => n16, ZN => SUM_11_port);
   U141 : INV_X1 port map( A => n69, ZN => n78);
   U142 : INV_X1 port map( A => n58, ZN => n83);
   U143 : NAND3_X1 port map( A1 => n49, A2 => n42, A3 => n84, ZN => n82);
   U144 : NAND3_X1 port map( A1 => A(8), A2 => A(11), A3 => A(12), ZN => n104);
   U145 : XNOR2_X1 port map( A => n107, B => n106, ZN => SUM_15_port);
   U146 : INV_X1 port map( A => A(14), ZN => n108);
   U147 : INV_X1 port map( A => n79, ZN => n75);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute_DW01_add_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Execute_DW01_add_1;

architecture SYN_rpl of Execute_DW01_add_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_3_port, SUM_4_port, SUM_5_port, SUM_6_port, 
      SUM_7_port, SUM_8_port, SUM_9_port, SUM_10_port, SUM_11_port, SUM_12_port
      , SUM_13_port, SUM_14_port, SUM_15_port, SUM_16_port, SUM_17_port, 
      SUM_18_port, SUM_19_port, SUM_20_port, SUM_21_port, SUM_22_port, 
      SUM_23_port, SUM_24_port, SUM_25_port, SUM_26_port, SUM_27_port, 
      SUM_28_port, SUM_29_port, SUM_30_port, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n54, n55, n56, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, B(1), B(0) );
   
   U1 : XNOR2_X1 port map( A => B(31), B => n57, ZN => SUM_31_port);
   U2 : NAND2_X1 port map( A1 => B(30), A2 => n56, ZN => n57);
   U3 : INV_X1 port map( A => B(2), ZN => SUM_2_port);
   U4 : XOR2_X1 port map( A => B(3), B => B(2), Z => SUM_3_port);
   U5 : XOR2_X1 port map( A => B(4), B => n30, Z => SUM_4_port);
   U6 : XOR2_X1 port map( A => B(5), B => n31, Z => SUM_5_port);
   U7 : XOR2_X1 port map( A => B(6), B => n32, Z => SUM_6_port);
   U8 : XOR2_X1 port map( A => B(7), B => n33, Z => SUM_7_port);
   U9 : XOR2_X1 port map( A => B(8), B => n34, Z => SUM_8_port);
   U10 : XOR2_X1 port map( A => B(9), B => n35, Z => SUM_9_port);
   U11 : XOR2_X1 port map( A => B(10), B => n36, Z => SUM_10_port);
   U12 : XOR2_X1 port map( A => B(11), B => n37, Z => SUM_11_port);
   U13 : XOR2_X1 port map( A => B(12), B => n38, Z => SUM_12_port);
   U14 : XOR2_X1 port map( A => B(13), B => n39, Z => SUM_13_port);
   U15 : XOR2_X1 port map( A => B(14), B => n40, Z => SUM_14_port);
   U16 : XOR2_X1 port map( A => B(15), B => n41, Z => SUM_15_port);
   U17 : XOR2_X1 port map( A => B(16), B => n42, Z => SUM_16_port);
   U18 : XOR2_X1 port map( A => B(17), B => n43, Z => SUM_17_port);
   U19 : XOR2_X1 port map( A => B(18), B => n44, Z => SUM_18_port);
   U20 : XOR2_X1 port map( A => B(19), B => n45, Z => SUM_19_port);
   U21 : XOR2_X1 port map( A => B(20), B => n46, Z => SUM_20_port);
   U22 : XOR2_X1 port map( A => B(21), B => n47, Z => SUM_21_port);
   U23 : XOR2_X1 port map( A => B(22), B => n48, Z => SUM_22_port);
   U24 : XOR2_X1 port map( A => B(23), B => n49, Z => SUM_23_port);
   U25 : XOR2_X1 port map( A => B(24), B => n50, Z => SUM_24_port);
   U26 : XOR2_X1 port map( A => B(25), B => n51, Z => SUM_25_port);
   U27 : XOR2_X1 port map( A => B(26), B => n52, Z => SUM_26_port);
   U28 : XOR2_X1 port map( A => B(27), B => n53, Z => SUM_27_port);
   U29 : XOR2_X1 port map( A => B(28), B => n54, Z => SUM_28_port);
   U30 : XOR2_X1 port map( A => B(29), B => n55, Z => SUM_29_port);
   U31 : XOR2_X1 port map( A => B(30), B => n56, Z => SUM_30_port);
   U32 : AND2_X1 port map( A1 => B(3), A2 => B(2), ZN => n30);
   U33 : AND2_X1 port map( A1 => B(4), A2 => n30, ZN => n31);
   U34 : AND2_X1 port map( A1 => B(5), A2 => n31, ZN => n32);
   U35 : AND2_X1 port map( A1 => B(6), A2 => n32, ZN => n33);
   U36 : AND2_X1 port map( A1 => B(7), A2 => n33, ZN => n34);
   U37 : AND2_X1 port map( A1 => B(8), A2 => n34, ZN => n35);
   U38 : AND2_X1 port map( A1 => B(9), A2 => n35, ZN => n36);
   U39 : AND2_X1 port map( A1 => B(10), A2 => n36, ZN => n37);
   U40 : AND2_X1 port map( A1 => B(11), A2 => n37, ZN => n38);
   U41 : AND2_X1 port map( A1 => B(12), A2 => n38, ZN => n39);
   U42 : AND2_X1 port map( A1 => B(13), A2 => n39, ZN => n40);
   U43 : AND2_X1 port map( A1 => B(14), A2 => n40, ZN => n41);
   U44 : AND2_X1 port map( A1 => B(15), A2 => n41, ZN => n42);
   U45 : AND2_X1 port map( A1 => B(16), A2 => n42, ZN => n43);
   U46 : AND2_X1 port map( A1 => B(17), A2 => n43, ZN => n44);
   U47 : AND2_X1 port map( A1 => B(18), A2 => n44, ZN => n45);
   U48 : AND2_X1 port map( A1 => B(19), A2 => n45, ZN => n46);
   U49 : AND2_X1 port map( A1 => B(20), A2 => n46, ZN => n47);
   U50 : AND2_X1 port map( A1 => B(21), A2 => n47, ZN => n48);
   U51 : AND2_X1 port map( A1 => B(22), A2 => n48, ZN => n49);
   U52 : AND2_X1 port map( A1 => B(23), A2 => n49, ZN => n50);
   U53 : AND2_X1 port map( A1 => B(24), A2 => n50, ZN => n51);
   U54 : AND2_X1 port map( A1 => B(25), A2 => n51, ZN => n52);
   U55 : AND2_X1 port map( A1 => B(26), A2 => n52, ZN => n53);
   U56 : AND2_X1 port map( A1 => B(27), A2 => n53, ZN => n54);
   U57 : AND2_X1 port map( A1 => B(28), A2 => n54, ZN => n55);
   U58 : AND2_X1 port map( A1 => B(29), A2 => n55, ZN => n56);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Execute_DW01_add_0;

architecture SYN_rpl of Execute_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n2, n_1070 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1070, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n2, CO => carry_2_port, S
                           => SUM(1));
   U1 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U2 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n2);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity comparator_NBIT32_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end comparator_NBIT32_DW01_cmp6_0;

architecture SYN_rpl of comparator_NBIT32_DW01_cmp6_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal GT_port, GE_port, NE_port, n3, LE_port, n5, n6, n7, n8, n9, n10, n11,
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55
      , n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, 
      n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84
      , n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, 
      n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202 : std_logic;

begin
   GT <= GT_port;
   LE <= LE_port;
   GE <= GE_port;
   NE <= NE_port;
   
   U1 : INV_X1 port map( A => n142, ZN => n10);
   U2 : INV_X1 port map( A => n130, ZN => n14);
   U3 : INV_X1 port map( A => n118, ZN => n18);
   U4 : INV_X1 port map( A => n106, ZN => n22);
   U5 : INV_X1 port map( A => n94, ZN => n26);
   U6 : INV_X1 port map( A => n82, ZN => n30);
   U7 : INV_X1 port map( A => GE_port, ZN => LT);
   U8 : INV_X1 port map( A => NE_port, ZN => EQ);
   U9 : INV_X1 port map( A => n139, ZN => n12);
   U10 : INV_X1 port map( A => n127, ZN => n16);
   U11 : INV_X1 port map( A => n115, ZN => n20);
   U12 : INV_X1 port map( A => n103, ZN => n24);
   U13 : INV_X1 port map( A => n91, ZN => n28);
   U14 : INV_X1 port map( A => n79, ZN => n32);
   U15 : INV_X1 port map( A => GT_port, ZN => LE_port);
   U16 : INV_X1 port map( A => n144, ZN => n9);
   U17 : INV_X1 port map( A => n132, ZN => n13);
   U18 : INV_X1 port map( A => n120, ZN => n17);
   U19 : INV_X1 port map( A => n108, ZN => n21);
   U20 : INV_X1 port map( A => n96, ZN => n25);
   U21 : INV_X1 port map( A => n84, ZN => n29);
   U22 : INV_X1 port map( A => n154, ZN => n7);
   U23 : INV_X1 port map( A => n141, ZN => n11);
   U24 : INV_X1 port map( A => n129, ZN => n15);
   U25 : INV_X1 port map( A => n117, ZN => n19);
   U26 : INV_X1 port map( A => n105, ZN => n23);
   U27 : INV_X1 port map( A => n93, ZN => n27);
   U28 : INV_X1 port map( A => n81, ZN => n31);
   U29 : INV_X1 port map( A => n68, ZN => n3);
   U30 : INV_X1 port map( A => A(30), ZN => n65);
   U31 : INV_X1 port map( A => n72, ZN => n33);
   U32 : INV_X1 port map( A => n151, ZN => n8);
   U33 : INV_X1 port map( A => n202, ZN => n5);
   U34 : INV_X1 port map( A => B(30), ZN => n34);
   U35 : INV_X1 port map( A => A(0), ZN => n36);
   U36 : INV_X1 port map( A => A(3), ZN => n38);
   U37 : INV_X1 port map( A => A(5), ZN => n40);
   U38 : INV_X1 port map( A => A(7), ZN => n42);
   U39 : INV_X1 port map( A => A(9), ZN => n44);
   U40 : INV_X1 port map( A => A(11), ZN => n46);
   U41 : INV_X1 port map( A => A(13), ZN => n48);
   U42 : INV_X1 port map( A => A(15), ZN => n50);
   U43 : INV_X1 port map( A => A(17), ZN => n52);
   U44 : INV_X1 port map( A => A(19), ZN => n54);
   U45 : INV_X1 port map( A => A(21), ZN => n56);
   U46 : INV_X1 port map( A => A(23), ZN => n58);
   U47 : INV_X1 port map( A => A(25), ZN => n60);
   U48 : INV_X1 port map( A => A(27), ZN => n62);
   U49 : INV_X1 port map( A => A(29), ZN => n64);
   U50 : INV_X1 port map( A => B(31), ZN => n35);
   U51 : INV_X1 port map( A => B(1), ZN => n6);
   U52 : INV_X1 port map( A => A(4), ZN => n39);
   U53 : INV_X1 port map( A => A(8), ZN => n43);
   U54 : INV_X1 port map( A => A(12), ZN => n47);
   U55 : INV_X1 port map( A => A(16), ZN => n51);
   U56 : INV_X1 port map( A => A(20), ZN => n55);
   U57 : INV_X1 port map( A => A(24), ZN => n59);
   U58 : INV_X1 port map( A => A(28), ZN => n63);
   U59 : INV_X1 port map( A => A(2), ZN => n37);
   U60 : INV_X1 port map( A => A(6), ZN => n41);
   U61 : INV_X1 port map( A => A(10), ZN => n45);
   U62 : INV_X1 port map( A => A(14), ZN => n49);
   U63 : INV_X1 port map( A => A(18), ZN => n53);
   U64 : INV_X1 port map( A => A(22), ZN => n57);
   U65 : INV_X1 port map( A => A(26), ZN => n61);
   U66 : NAND2_X1 port map( A1 => LE_port, A2 => GE_port, ZN => NE_port);
   U67 : AOI21_X1 port map( B1 => n66, B2 => n3, A => n67, ZN => GE_port);
   U68 : AOI22_X1 port map( A1 => B(30), A2 => n65, B1 => n69, B2 => n70, ZN =>
                           n68);
   U69 : AOI21_X1 port map( B1 => n71, B2 => n72, A => n73, ZN => n69);
   U70 : AOI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => n71);
   U71 : AOI21_X1 port map( B1 => n77, B2 => n78, A => n79, ZN => n74);
   U72 : AOI21_X1 port map( B1 => n80, B2 => n30, A => n31, ZN => n77);
   U73 : AOI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n80);
   U74 : AOI21_X1 port map( B1 => n86, B2 => n87, A => n88, ZN => n83);
   U75 : AOI21_X1 port map( B1 => n89, B2 => n90, A => n91, ZN => n86);
   U76 : AOI21_X1 port map( B1 => n92, B2 => n26, A => n27, ZN => n89);
   U77 : AOI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n92);
   U78 : AOI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => n95);
   U79 : AOI21_X1 port map( B1 => n101, B2 => n102, A => n103, ZN => n98);
   U80 : AOI21_X1 port map( B1 => n104, B2 => n22, A => n23, ZN => n101);
   U81 : AOI21_X1 port map( B1 => n107, B2 => n108, A => n109, ZN => n104);
   U82 : AOI21_X1 port map( B1 => n110, B2 => n111, A => n112, ZN => n107);
   U83 : AOI21_X1 port map( B1 => n113, B2 => n114, A => n115, ZN => n110);
   U84 : AOI21_X1 port map( B1 => n116, B2 => n18, A => n19, ZN => n113);
   U85 : AOI21_X1 port map( B1 => n119, B2 => n120, A => n121, ZN => n116);
   U86 : AOI21_X1 port map( B1 => n122, B2 => n123, A => n124, ZN => n119);
   U87 : AOI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n122);
   U88 : AOI21_X1 port map( B1 => n128, B2 => n14, A => n15, ZN => n125);
   U89 : AOI21_X1 port map( B1 => n131, B2 => n132, A => n133, ZN => n128);
   U90 : AOI21_X1 port map( B1 => n134, B2 => n135, A => n136, ZN => n131);
   U91 : AOI21_X1 port map( B1 => n137, B2 => n138, A => n139, ZN => n134);
   U92 : AOI21_X1 port map( B1 => n140, B2 => n10, A => n11, ZN => n137);
   U93 : AOI21_X1 port map( B1 => n143, B2 => n144, A => n145, ZN => n140);
   U94 : AOI21_X1 port map( B1 => n146, B2 => n147, A => n148, ZN => n143);
   U95 : AOI21_X1 port map( B1 => n149, B2 => n150, A => n151, ZN => n146);
   U96 : AOI21_X1 port map( B1 => n152, B2 => n153, A => n7, ZN => n149);
   U97 : AOI22_X1 port map( A1 => n155, A2 => n6, B1 => A(1), B2 => n156, ZN =>
                           n152);
   U98 : OR2_X1 port map( A1 => n156, A2 => A(1), ZN => n155);
   U99 : NAND2_X1 port map( A1 => B(0), A2 => n36, ZN => n156);
   U100 : OAI21_X1 port map( B1 => n67, B2 => n157, A => n66, ZN => GT_port);
   U101 : NAND2_X1 port map( A1 => A(31), A2 => n35, ZN => n66);
   U102 : AOI22_X1 port map( A1 => A(30), A2 => n34, B1 => n158, B2 => n70, ZN 
                           => n157);
   U103 : XOR2_X1 port map( A => A(30), B => n34, Z => n70);
   U104 : AOI21_X1 port map( B1 => n159, B2 => n160, A => n33, ZN => n158);
   U105 : NAND2_X1 port map( A1 => B(29), A2 => n64, ZN => n72);
   U106 : OAI211_X1 port map( C1 => n161, C2 => n162, A => n78, B => n75, ZN =>
                           n160);
   U107 : NOR2_X1 port map( A1 => n163, A2 => n76, ZN => n75);
   U108 : AND2_X1 port map( A1 => B(28), A2 => n63, ZN => n76);
   U109 : NAND2_X1 port map( A1 => B(27), A2 => n62, ZN => n78);
   U110 : NAND2_X1 port map( A1 => n32, A2 => n164, ZN => n162);
   U111 : NOR2_X1 port map( A1 => n62, A2 => B(27), ZN => n79);
   U112 : AOI211_X1 port map( C1 => n165, C2 => n166, A => n82, B => n29, ZN =>
                           n161);
   U113 : NAND2_X1 port map( A1 => B(25), A2 => n60, ZN => n84);
   U114 : NAND2_X1 port map( A1 => n164, A2 => n81, ZN => n82);
   U115 : NAND2_X1 port map( A1 => B(26), A2 => n61, ZN => n81);
   U116 : OR2_X1 port map( A1 => n61, A2 => B(26), ZN => n164);
   U117 : OAI211_X1 port map( C1 => n167, C2 => n168, A => n90, B => n87, ZN =>
                           n166);
   U118 : NOR2_X1 port map( A1 => n169, A2 => n88, ZN => n87);
   U119 : AND2_X1 port map( A1 => B(24), A2 => n59, ZN => n88);
   U120 : NAND2_X1 port map( A1 => B(23), A2 => n58, ZN => n90);
   U121 : NAND2_X1 port map( A1 => n28, A2 => n170, ZN => n168);
   U122 : NOR2_X1 port map( A1 => n58, A2 => B(23), ZN => n91);
   U123 : AOI211_X1 port map( C1 => n171, C2 => n172, A => n94, B => n25, ZN =>
                           n167);
   U124 : NAND2_X1 port map( A1 => B(21), A2 => n56, ZN => n96);
   U125 : NAND2_X1 port map( A1 => n170, A2 => n93, ZN => n94);
   U126 : NAND2_X1 port map( A1 => B(22), A2 => n57, ZN => n93);
   U127 : OR2_X1 port map( A1 => n57, A2 => B(22), ZN => n170);
   U128 : OAI211_X1 port map( C1 => n173, C2 => n174, A => n102, B => n99, ZN 
                           => n172);
   U129 : NOR2_X1 port map( A1 => n175, A2 => n100, ZN => n99);
   U130 : AND2_X1 port map( A1 => B(20), A2 => n55, ZN => n100);
   U131 : NAND2_X1 port map( A1 => B(19), A2 => n54, ZN => n102);
   U132 : NAND2_X1 port map( A1 => n24, A2 => n176, ZN => n174);
   U133 : NOR2_X1 port map( A1 => n54, A2 => B(19), ZN => n103);
   U134 : AOI211_X1 port map( C1 => n177, C2 => n178, A => n106, B => n21, ZN 
                           => n173);
   U135 : NAND2_X1 port map( A1 => B(17), A2 => n52, ZN => n108);
   U136 : NAND2_X1 port map( A1 => n176, A2 => n105, ZN => n106);
   U137 : NAND2_X1 port map( A1 => B(18), A2 => n53, ZN => n105);
   U138 : OR2_X1 port map( A1 => n53, A2 => B(18), ZN => n176);
   U139 : OAI211_X1 port map( C1 => n179, C2 => n180, A => n114, B => n111, ZN 
                           => n178);
   U140 : NOR2_X1 port map( A1 => n181, A2 => n112, ZN => n111);
   U141 : AND2_X1 port map( A1 => B(16), A2 => n51, ZN => n112);
   U142 : NAND2_X1 port map( A1 => B(15), A2 => n50, ZN => n114);
   U143 : NAND2_X1 port map( A1 => n20, A2 => n182, ZN => n180);
   U144 : NOR2_X1 port map( A1 => n50, A2 => B(15), ZN => n115);
   U145 : AOI211_X1 port map( C1 => n183, C2 => n184, A => n118, B => n17, ZN 
                           => n179);
   U146 : NAND2_X1 port map( A1 => B(13), A2 => n48, ZN => n120);
   U147 : NAND2_X1 port map( A1 => n182, A2 => n117, ZN => n118);
   U148 : NAND2_X1 port map( A1 => B(14), A2 => n49, ZN => n117);
   U149 : OR2_X1 port map( A1 => n49, A2 => B(14), ZN => n182);
   U150 : OAI211_X1 port map( C1 => n185, C2 => n186, A => n126, B => n123, ZN 
                           => n184);
   U151 : NOR2_X1 port map( A1 => n187, A2 => n124, ZN => n123);
   U152 : AND2_X1 port map( A1 => B(12), A2 => n47, ZN => n124);
   U153 : NAND2_X1 port map( A1 => B(11), A2 => n46, ZN => n126);
   U154 : NAND2_X1 port map( A1 => n16, A2 => n188, ZN => n186);
   U155 : NOR2_X1 port map( A1 => n46, A2 => B(11), ZN => n127);
   U156 : AOI211_X1 port map( C1 => n189, C2 => n190, A => n130, B => n13, ZN 
                           => n185);
   U157 : NAND2_X1 port map( A1 => B(9), A2 => n44, ZN => n132);
   U158 : NAND2_X1 port map( A1 => n188, A2 => n129, ZN => n130);
   U159 : NAND2_X1 port map( A1 => B(10), A2 => n45, ZN => n129);
   U160 : OR2_X1 port map( A1 => n45, A2 => B(10), ZN => n188);
   U161 : OAI211_X1 port map( C1 => n191, C2 => n192, A => n138, B => n135, ZN 
                           => n190);
   U162 : NOR2_X1 port map( A1 => n193, A2 => n136, ZN => n135);
   U163 : AND2_X1 port map( A1 => B(8), A2 => n43, ZN => n136);
   U164 : NAND2_X1 port map( A1 => B(7), A2 => n42, ZN => n138);
   U165 : NAND2_X1 port map( A1 => n12, A2 => n194, ZN => n192);
   U166 : NOR2_X1 port map( A1 => n42, A2 => B(7), ZN => n139);
   U167 : AOI211_X1 port map( C1 => n195, C2 => n196, A => n142, B => n9, ZN =>
                           n191);
   U168 : NAND2_X1 port map( A1 => B(5), A2 => n40, ZN => n144);
   U169 : NAND2_X1 port map( A1 => n194, A2 => n141, ZN => n142);
   U170 : NAND2_X1 port map( A1 => B(6), A2 => n41, ZN => n141);
   U171 : OR2_X1 port map( A1 => n41, A2 => B(6), ZN => n194);
   U172 : NAND3_X1 port map( A1 => n197, A2 => n150, A3 => n147, ZN => n196);
   U173 : NOR2_X1 port map( A1 => n198, A2 => n148, ZN => n147);
   U174 : AND2_X1 port map( A1 => B(4), A2 => n39, ZN => n148);
   U175 : NAND2_X1 port map( A1 => B(3), A2 => n38, ZN => n150);
   U176 : NAND3_X1 port map( A1 => n8, A2 => n199, A3 => n200, ZN => n197);
   U177 : OAI211_X1 port map( C1 => A(1), C2 => n201, A => n5, B => n153, ZN =>
                           n200);
   U178 : AND2_X1 port map( A1 => n199, A2 => n154, ZN => n153);
   U179 : NAND2_X1 port map( A1 => B(2), A2 => n37, ZN => n154);
   U180 : AOI21_X1 port map( B1 => A(1), B2 => n201, A => n6, ZN => n202);
   U181 : NOR2_X1 port map( A1 => n36, A2 => B(0), ZN => n201);
   U182 : OR2_X1 port map( A1 => n37, A2 => B(2), ZN => n199);
   U183 : NOR2_X1 port map( A1 => n38, A2 => B(3), ZN => n151);
   U184 : NOR2_X1 port map( A1 => n198, A2 => n145, ZN => n195);
   U185 : NOR2_X1 port map( A1 => n40, A2 => B(5), ZN => n145);
   U186 : NOR2_X1 port map( A1 => n39, A2 => B(4), ZN => n198);
   U187 : NOR2_X1 port map( A1 => n193, A2 => n133, ZN => n189);
   U188 : NOR2_X1 port map( A1 => n44, A2 => B(9), ZN => n133);
   U189 : NOR2_X1 port map( A1 => n43, A2 => B(8), ZN => n193);
   U190 : NOR2_X1 port map( A1 => n187, A2 => n121, ZN => n183);
   U191 : NOR2_X1 port map( A1 => n48, A2 => B(13), ZN => n121);
   U192 : NOR2_X1 port map( A1 => n47, A2 => B(12), ZN => n187);
   U193 : NOR2_X1 port map( A1 => n181, A2 => n109, ZN => n177);
   U194 : NOR2_X1 port map( A1 => n52, A2 => B(17), ZN => n109);
   U195 : NOR2_X1 port map( A1 => n51, A2 => B(16), ZN => n181);
   U196 : NOR2_X1 port map( A1 => n175, A2 => n97, ZN => n171);
   U197 : NOR2_X1 port map( A1 => n56, A2 => B(21), ZN => n97);
   U198 : NOR2_X1 port map( A1 => n55, A2 => B(20), ZN => n175);
   U199 : NOR2_X1 port map( A1 => n169, A2 => n85, ZN => n165);
   U200 : NOR2_X1 port map( A1 => n60, A2 => B(25), ZN => n85);
   U201 : NOR2_X1 port map( A1 => n59, A2 => B(24), ZN => n169);
   U202 : NOR2_X1 port map( A1 => n163, A2 => n73, ZN => n159);
   U203 : NOR2_X1 port map( A1 => n64, A2 => B(29), ZN => n73);
   U204 : NOR2_X1 port map( A1 => n63, A2 => B(28), ZN => n163);
   U205 : NOR2_X1 port map( A1 => n35, A2 => A(31), ZN => n67);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HazardDetection_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end HazardDetection_DW01_sub_0;

architecture SYN_rpl of HazardDetection_DW01_sub_0 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port,
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, carry_31_port, 
      carry_30_port, carry_29_port, carry_28_port, carry_27_port, carry_26_port
      , carry_25_port, carry_24_port, carry_23_port, carry_22_port, 
      carry_21_port, carry_20_port, carry_19_port, carry_18_port, carry_17_port
      , carry_16_port, carry_15_port, carry_14_port, carry_13_port, 
      carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, DIFF_2_port : 
      std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, A(1), A(0) );
   
   U1 : XNOR2_X1 port map( A => A(5), B => carry_5_port, ZN => DIFF_5_port);
   U2 : XNOR2_X1 port map( A => A(6), B => carry_6_port, ZN => DIFF_6_port);
   U3 : XNOR2_X1 port map( A => A(10), B => carry_10_port, ZN => DIFF_10_port);
   U4 : XNOR2_X1 port map( A => A(13), B => carry_13_port, ZN => DIFF_13_port);
   U5 : XNOR2_X1 port map( A => A(11), B => carry_11_port, ZN => DIFF_11_port);
   U6 : XNOR2_X1 port map( A => A(14), B => carry_14_port, ZN => DIFF_14_port);
   U7 : XNOR2_X1 port map( A => A(15), B => carry_15_port, ZN => DIFF_15_port);
   U8 : XNOR2_X1 port map( A => A(17), B => carry_17_port, ZN => DIFF_17_port);
   U9 : XNOR2_X1 port map( A => A(4), B => carry_4_port, ZN => DIFF_4_port);
   U10 : XNOR2_X1 port map( A => A(8), B => carry_8_port, ZN => DIFF_8_port);
   U11 : XNOR2_X1 port map( A => A(9), B => carry_9_port, ZN => DIFF_9_port);
   U12 : INV_X1 port map( A => A(2), ZN => DIFF_2_port);
   U13 : XNOR2_X1 port map( A => A(20), B => carry_20_port, ZN => DIFF_20_port)
                           ;
   U14 : XNOR2_X1 port map( A => A(21), B => carry_21_port, ZN => DIFF_21_port)
                           ;
   U15 : XNOR2_X1 port map( A => A(22), B => carry_22_port, ZN => DIFF_22_port)
                           ;
   U16 : XNOR2_X1 port map( A => A(23), B => carry_23_port, ZN => DIFF_23_port)
                           ;
   U17 : XNOR2_X1 port map( A => A(24), B => carry_24_port, ZN => DIFF_24_port)
                           ;
   U18 : XNOR2_X1 port map( A => A(25), B => carry_25_port, ZN => DIFF_25_port)
                           ;
   U19 : XNOR2_X1 port map( A => A(26), B => carry_26_port, ZN => DIFF_26_port)
                           ;
   U20 : XNOR2_X1 port map( A => A(28), B => carry_28_port, ZN => DIFF_28_port)
                           ;
   U21 : XNOR2_X1 port map( A => A(29), B => carry_29_port, ZN => DIFF_29_port)
                           ;
   U22 : XNOR2_X1 port map( A => A(30), B => carry_30_port, ZN => DIFF_30_port)
                           ;
   U23 : XNOR2_X1 port map( A => A(31), B => carry_31_port, ZN => DIFF_31_port)
                           ;
   U24 : XNOR2_X1 port map( A => A(7), B => carry_7_port, ZN => DIFF_7_port);
   U25 : XNOR2_X1 port map( A => A(12), B => carry_12_port, ZN => DIFF_12_port)
                           ;
   U26 : XNOR2_X1 port map( A => A(16), B => carry_16_port, ZN => DIFF_16_port)
                           ;
   U27 : XNOR2_X1 port map( A => A(3), B => A(2), ZN => DIFF_3_port);
   U28 : XNOR2_X1 port map( A => A(18), B => carry_18_port, ZN => DIFF_18_port)
                           ;
   U29 : XNOR2_X1 port map( A => A(19), B => carry_19_port, ZN => DIFF_19_port)
                           ;
   U30 : XNOR2_X1 port map( A => A(27), B => carry_27_port, ZN => DIFF_27_port)
                           ;
   U31 : OR2_X1 port map( A1 => A(3), A2 => A(2), ZN => carry_4_port);
   U32 : OR2_X1 port map( A1 => A(4), A2 => carry_4_port, ZN => carry_5_port);
   U33 : OR2_X1 port map( A1 => A(5), A2 => carry_5_port, ZN => carry_6_port);
   U34 : OR2_X1 port map( A1 => A(6), A2 => carry_6_port, ZN => carry_7_port);
   U35 : OR2_X1 port map( A1 => A(7), A2 => carry_7_port, ZN => carry_8_port);
   U36 : OR2_X1 port map( A1 => A(8), A2 => carry_8_port, ZN => carry_9_port);
   U37 : OR2_X1 port map( A1 => A(9), A2 => carry_9_port, ZN => carry_10_port);
   U38 : OR2_X1 port map( A1 => A(10), A2 => carry_10_port, ZN => carry_11_port
                           );
   U39 : OR2_X1 port map( A1 => A(11), A2 => carry_11_port, ZN => carry_12_port
                           );
   U40 : OR2_X1 port map( A1 => A(12), A2 => carry_12_port, ZN => carry_13_port
                           );
   U41 : OR2_X1 port map( A1 => A(13), A2 => carry_13_port, ZN => carry_14_port
                           );
   U42 : OR2_X1 port map( A1 => A(14), A2 => carry_14_port, ZN => carry_15_port
                           );
   U43 : OR2_X1 port map( A1 => A(15), A2 => carry_15_port, ZN => carry_16_port
                           );
   U44 : OR2_X1 port map( A1 => A(16), A2 => carry_16_port, ZN => carry_17_port
                           );
   U45 : OR2_X1 port map( A1 => A(17), A2 => carry_17_port, ZN => carry_18_port
                           );
   U46 : OR2_X1 port map( A1 => A(18), A2 => carry_18_port, ZN => carry_19_port
                           );
   U47 : OR2_X1 port map( A1 => A(19), A2 => carry_19_port, ZN => carry_20_port
                           );
   U48 : OR2_X1 port map( A1 => A(20), A2 => carry_20_port, ZN => carry_21_port
                           );
   U49 : OR2_X1 port map( A1 => A(21), A2 => carry_21_port, ZN => carry_22_port
                           );
   U50 : OR2_X1 port map( A1 => A(22), A2 => carry_22_port, ZN => carry_23_port
                           );
   U51 : OR2_X1 port map( A1 => A(23), A2 => carry_23_port, ZN => carry_24_port
                           );
   U52 : OR2_X1 port map( A1 => A(24), A2 => carry_24_port, ZN => carry_25_port
                           );
   U53 : OR2_X1 port map( A1 => A(25), A2 => carry_25_port, ZN => carry_26_port
                           );
   U54 : OR2_X1 port map( A1 => A(26), A2 => carry_26_port, ZN => carry_27_port
                           );
   U55 : OR2_X1 port map( A1 => A(27), A2 => carry_27_port, ZN => carry_28_port
                           );
   U56 : OR2_X1 port map( A1 => A(28), A2 => carry_28_port, ZN => carry_29_port
                           );
   U57 : OR2_X1 port map( A1 => A(29), A2 => carry_29_port, ZN => carry_30_port
                           );
   U58 : OR2_X1 port map( A1 => A(30), A2 => carry_30_port, ZN => carry_31_port
                           );

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_15;

architecture SYN_STRUCTURAL of RCA_N4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_14;

architecture SYN_STRUCTURAL of RCA_N4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_13;

architecture SYN_STRUCTURAL of RCA_N4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_12;

architecture SYN_STRUCTURAL of RCA_N4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_11;

architecture SYN_STRUCTURAL of RCA_N4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_10;

architecture SYN_STRUCTURAL of RCA_N4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_9;

architecture SYN_STRUCTURAL of RCA_N4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_8;

architecture SYN_STRUCTURAL of RCA_N4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_7;

architecture SYN_STRUCTURAL of RCA_N4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_6;

architecture SYN_STRUCTURAL of RCA_N4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_5;

architecture SYN_STRUCTURAL of RCA_N4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_4;

architecture SYN_STRUCTURAL of RCA_N4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_3;

architecture SYN_STRUCTURAL of RCA_N4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_2;

architecture SYN_STRUCTURAL of RCA_N4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_1;

architecture SYN_STRUCTURAL of RCA_N4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_7;

architecture SYN_struct of carry_select_basic_N4_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1106, n_1107 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1106);
   RCA1 : RCA_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1107);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n11, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_6;

architecture SYN_struct of carry_select_basic_N4_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1108, n_1109 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1108);
   RCA1 : RCA_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1109);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n11, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_5;

architecture SYN_struct of carry_select_basic_N4_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1110, n_1111 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1110);
   RCA1 : RCA_N4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1111);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n11, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_4;

architecture SYN_struct of carry_select_basic_N4_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1112, n_1113 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1112);
   RCA1 : RCA_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1113);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n11, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_3;

architecture SYN_struct of carry_select_basic_N4_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1114, n_1115 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1114);
   RCA1 : RCA_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1115);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n11, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_2;

architecture SYN_struct of carry_select_basic_N4_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1116, n_1117 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1116);
   RCA1 : RCA_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1117);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n11, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_1;

architecture SYN_struct of carry_select_basic_N4_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1118, n_1119 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1118);
   RCA1 : RCA_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1119);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n11, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_26 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_26;

architecture SYN_bhv of PGblock_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_25 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_25;

architecture SYN_bhv of PGblock_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_24 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_24;

architecture SYN_bhv of PGblock_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_23 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_23;

architecture SYN_bhv of PGblock_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_22 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_22;

architecture SYN_bhv of PGblock_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_21 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_21;

architecture SYN_bhv of PGblock_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_20 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_20;

architecture SYN_bhv of PGblock_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_19 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_19;

architecture SYN_bhv of PGblock_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_18 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_18;

architecture SYN_bhv of PGblock_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_17 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_17;

architecture SYN_bhv of PGblock_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_16 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_16;

architecture SYN_bhv of PGblock_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_15 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_15;

architecture SYN_bhv of PGblock_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_14 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_14;

architecture SYN_bhv of PGblock_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_13 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_13;

architecture SYN_bhv of PGblock_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_12 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_12;

architecture SYN_bhv of PGblock_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_11 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_11;

architecture SYN_bhv of PGblock_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_10 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_10;

architecture SYN_bhv of PGblock_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_9 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_9;

architecture SYN_bhv of PGblock_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_8 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_8;

architecture SYN_bhv of PGblock_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_7 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_7;

architecture SYN_bhv of PGblock_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_6 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_6;

architecture SYN_bhv of PGblock_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_5 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_5;

architecture SYN_bhv of PGblock_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_4 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_4;

architecture SYN_bhv of PGblock_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_3 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_3;

architecture SYN_bhv of PGblock_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_2 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_2;

architecture SYN_bhv of PGblock_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_1 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_1;

architecture SYN_bhv of PGblock_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_8 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_8;

architecture SYN_bhv of Gblock_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_7 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_7;

architecture SYN_bhv of Gblock_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_6 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_6;

architecture SYN_bhv of Gblock_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_5 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_5;

architecture SYN_bhv of Gblock_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_4 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_4;

architecture SYN_bhv of Gblock_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_3 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_3;

architecture SYN_bhv of Gblock_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_2 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_2;

architecture SYN_bhv of Gblock_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_1 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_1;

architecture SYN_bhv of Gblock_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_30 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_30;

architecture SYN_bhv of PG_net_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_29 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_29;

architecture SYN_bhv of PG_net_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_28 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_28;

architecture SYN_bhv of PG_net_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_27 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_27;

architecture SYN_bhv of PG_net_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_26 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_26;

architecture SYN_bhv of PG_net_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_25 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_25;

architecture SYN_bhv of PG_net_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_24 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_24;

architecture SYN_bhv of PG_net_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_23 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_23;

architecture SYN_bhv of PG_net_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_22 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_22;

architecture SYN_bhv of PG_net_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_21 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_21;

architecture SYN_bhv of PG_net_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_20 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_20;

architecture SYN_bhv of PG_net_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_19 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_19;

architecture SYN_bhv of PG_net_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_18 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_18;

architecture SYN_bhv of PG_net_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_17 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_17;

architecture SYN_bhv of PG_net_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_16 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_16;

architecture SYN_bhv of PG_net_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_15 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_15;

architecture SYN_bhv of PG_net_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_14 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_14;

architecture SYN_bhv of PG_net_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_13 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_13;

architecture SYN_bhv of PG_net_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_12 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_12;

architecture SYN_bhv of PG_net_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_11 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_11;

architecture SYN_bhv of PG_net_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_10 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_10;

architecture SYN_bhv of PG_net_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_9 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_9;

architecture SYN_bhv of PG_net_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_8 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_8;

architecture SYN_bhv of PG_net_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_7 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_7;

architecture SYN_bhv of PG_net_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_6 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_6;

architecture SYN_bhv of PG_net_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_5 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_5;

architecture SYN_bhv of PG_net_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_4 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_4;

architecture SYN_bhv of PG_net_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_3 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_3;

architecture SYN_bhv of PG_net_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_2 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_2;

architecture SYN_bhv of PG_net_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_1 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_1;

architecture SYN_bhv of PG_net_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_4 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_4;

architecture SYN_bhv of mux41_NBIT32_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n145, Z => n72);
   U2 : BUF_X1 port map( A => n145, Z => n73);
   U3 : BUF_X1 port map( A => n147, Z => n78);
   U4 : BUF_X1 port map( A => n147, Z => n79);
   U5 : BUF_X1 port map( A => n144, Z => n1);
   U6 : BUF_X1 port map( A => n144, Z => n70);
   U7 : BUF_X1 port map( A => n146, Z => n75);
   U8 : BUF_X1 port map( A => n146, Z => n76);
   U9 : BUF_X1 port map( A => n145, Z => n74);
   U10 : BUF_X1 port map( A => n147, Z => n80);
   U11 : BUF_X1 port map( A => n144, Z => n71);
   U12 : BUF_X1 port map( A => n146, Z => n77);
   U13 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n145);
   U14 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n144);
   U15 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n147);
   U16 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n146);
   U17 : INV_X1 port map( A => S(0), ZN => n81);
   U18 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(1));
   U19 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN =>
                           n104);
   U20 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN => 
                           n105);
   U21 : NAND2_X1 port map( A1 => n83, A2 => n82, ZN => Z(0));
   U22 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n82);
   U23 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n83);
   U24 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(2));
   U25 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN =>
                           n126);
   U26 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN =>
                           n127);
   U27 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(6));
   U28 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n138);
   U29 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n139);
   U30 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(5));
   U31 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN =>
                           n136);
   U32 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN =>
                           n137);
   U33 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(4));
   U34 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN =>
                           n134);
   U35 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN =>
                           n135);
   U36 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => Z(13));
   U37 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN 
                           => n90);
   U38 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n91);
   U39 : NAND2_X1 port map( A1 => n93, A2 => n92, ZN => Z(14));
   U40 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN 
                           => n92);
   U41 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n93);
   U42 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => Z(12));
   U43 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN 
                           => n88);
   U44 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n89);
   U45 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(16));
   U46 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n96);
   U47 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n97);
   U48 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(17));
   U49 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n98);
   U50 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n99);
   U51 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(8));
   U52 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n142);
   U53 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n143);
   U54 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(9));
   U55 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN =>
                           n148);
   U56 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN =>
                           n149);
   U57 : NAND2_X1 port map( A1 => n85, A2 => n84, ZN => Z(10));
   U58 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN 
                           => n84);
   U59 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n85);
   U60 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(18));
   U61 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n100);
   U62 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n101);
   U63 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(21));
   U64 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n108);
   U65 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n109);
   U66 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(20));
   U67 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN 
                           => n106);
   U68 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN 
                           => n107);
   U69 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(30));
   U70 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN 
                           => n128);
   U71 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN 
                           => n129);
   U72 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(29));
   U73 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n124);
   U74 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n125);
   U75 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(24));
   U76 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN 
                           => n114);
   U77 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN 
                           => n115);
   U78 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(22));
   U79 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n110);
   U80 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n111);
   U81 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(25));
   U82 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n116);
   U83 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n117);
   U84 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(26));
   U85 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n118);
   U86 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n119);
   U87 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(28));
   U88 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n122);
   U89 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n123);
   U90 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(3));
   U91 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN =>
                           n132);
   U92 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN =>
                           n133);
   U93 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(7));
   U94 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n140);
   U95 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n141);
   U96 : NAND2_X1 port map( A1 => n87, A2 => n86, ZN => Z(11));
   U97 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN 
                           => n86);
   U98 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n87);
   U99 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => Z(15));
   U100 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN
                           => n94);
   U101 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n95);
   U102 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(19));
   U103 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN
                           => n102);
   U104 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n103);
   U105 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(23));
   U106 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN
                           => n112);
   U107 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN
                           => n113);
   U108 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(27));
   U109 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN
                           => n120);
   U110 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN
                           => n121);
   U111 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(31));
   U112 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN
                           => n130);
   U113 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN
                           => n131);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_3 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_3;

architecture SYN_bhv of mux41_NBIT32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n145, Z => n72);
   U2 : BUF_X1 port map( A => n147, Z => n78);
   U3 : BUF_X1 port map( A => n145, Z => n73);
   U4 : BUF_X1 port map( A => n147, Z => n79);
   U5 : BUF_X1 port map( A => n144, Z => n1);
   U6 : BUF_X1 port map( A => n146, Z => n75);
   U7 : BUF_X1 port map( A => n144, Z => n70);
   U8 : BUF_X1 port map( A => n146, Z => n76);
   U9 : BUF_X1 port map( A => n145, Z => n74);
   U10 : BUF_X1 port map( A => n147, Z => n80);
   U11 : BUF_X1 port map( A => n144, Z => n71);
   U12 : BUF_X1 port map( A => n146, Z => n77);
   U13 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(1));
   U14 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN =>
                           n104);
   U15 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN => 
                           n105);
   U16 : NAND2_X1 port map( A1 => n83, A2 => n82, ZN => Z(0));
   U17 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n82);
   U18 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n83);
   U19 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(2));
   U20 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN =>
                           n126);
   U21 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN =>
                           n127);
   U22 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(6));
   U23 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n138);
   U24 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n139);
   U25 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(5));
   U26 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN =>
                           n136);
   U27 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN =>
                           n137);
   U28 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(4));
   U29 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN =>
                           n134);
   U30 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN =>
                           n135);
   U31 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => Z(13));
   U32 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN 
                           => n90);
   U33 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n91);
   U34 : NAND2_X1 port map( A1 => n93, A2 => n92, ZN => Z(14));
   U35 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN 
                           => n92);
   U36 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n93);
   U37 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => Z(12));
   U38 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN 
                           => n88);
   U39 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n89);
   U40 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(16));
   U41 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n96);
   U42 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n97);
   U43 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(17));
   U44 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n98);
   U45 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n99);
   U46 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(8));
   U47 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n142);
   U48 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n143);
   U49 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(9));
   U50 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN =>
                           n148);
   U51 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN =>
                           n149);
   U52 : NAND2_X1 port map( A1 => n85, A2 => n84, ZN => Z(10));
   U53 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN 
                           => n84);
   U54 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n85);
   U55 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(18));
   U56 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n100);
   U57 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n101);
   U58 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(21));
   U59 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n108);
   U60 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n109);
   U61 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(20));
   U62 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN 
                           => n106);
   U63 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN 
                           => n107);
   U64 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(30));
   U65 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN 
                           => n128);
   U66 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN 
                           => n129);
   U67 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(29));
   U68 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n124);
   U69 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n125);
   U70 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(24));
   U71 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN 
                           => n114);
   U72 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN 
                           => n115);
   U73 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(22));
   U74 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n110);
   U75 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n111);
   U76 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(25));
   U77 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n116);
   U78 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n117);
   U79 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(26));
   U80 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n118);
   U81 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n119);
   U82 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(28));
   U83 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n122);
   U84 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n123);
   U85 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(3));
   U86 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN =>
                           n132);
   U87 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN =>
                           n133);
   U88 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(7));
   U89 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n140);
   U90 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n141);
   U91 : NAND2_X1 port map( A1 => n87, A2 => n86, ZN => Z(11));
   U92 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN 
                           => n86);
   U93 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n87);
   U94 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => Z(15));
   U95 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN 
                           => n94);
   U96 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n95);
   U97 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(19));
   U98 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN 
                           => n102);
   U99 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n103);
   U100 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(23));
   U101 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN
                           => n112);
   U102 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN
                           => n113);
   U103 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(27));
   U104 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN
                           => n120);
   U105 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN
                           => n121);
   U106 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(31));
   U107 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN
                           => n130);
   U108 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN
                           => n131);
   U109 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n145);
   U110 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n144);
   U111 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n147);
   U112 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n146);
   U113 : INV_X1 port map( A => S(0), ZN => n81);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_2 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_2;

architecture SYN_bhv of mux41_NBIT32_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => S(1), Z => n1);
   U2 : BUF_X1 port map( A => n30, Z => n2);
   U3 : BUF_X1 port map( A => n30, Z => n3);
   U4 : BUF_X2 port map( A => n28, Z => n4);
   U5 : BUF_X2 port map( A => n28, Z => n5);
   U6 : BUF_X1 port map( A => n30, Z => n38);
   U7 : BUF_X1 port map( A => n30, Z => n6);
   U8 : BUF_X1 port map( A => n30, Z => n40);
   U9 : BUF_X1 port map( A => n30, Z => n7);
   U10 : AND2_X2 port map( A1 => n44, A2 => n45, ZN => n28);
   U11 : AND2_X2 port map( A1 => S(0), A2 => n45, ZN => n30);
   U12 : AND2_X1 port map( A1 => n99, A2 => n26, ZN => n8);
   U13 : OAI221_X1 port map( B1 => n9, B2 => n10, C1 => n11, C2 => n12, A => 
                           n72, ZN => Z(14));
   U14 : INV_X1 port map( A => A(14), ZN => n9);
   U15 : INV_X1 port map( A => n28, ZN => n10);
   U16 : INV_X1 port map( A => B(14), ZN => n11);
   U17 : INV_X1 port map( A => n30, ZN => n12);
   U18 : OAI211_X1 port map( C1 => n13, C2 => n15, A => n27, B => n101, ZN => 
                           Z(30));
   U19 : INV_X1 port map( A => A(30), ZN => n13);
   U20 : AOI22_X1 port map( A1 => A(15), A2 => n28, B1 => B(15), B2 => n40, ZN 
                           => n73);
   U21 : OAI221_X1 port map( B1 => n14, B2 => n15, C1 => n16, C2 => n17, A => 
                           n100, ZN => Z(29));
   U22 : INV_X1 port map( A => A(29), ZN => n14);
   U23 : INV_X1 port map( A => n28, ZN => n15);
   U24 : INV_X1 port map( A => B(29), ZN => n16);
   U25 : INV_X1 port map( A => n30, ZN => n17);
   U26 : OAI221_X1 port map( B1 => n18, B2 => n19, C1 => n20, C2 => n21, A => 
                           n64, ZN => Z(9));
   U27 : INV_X1 port map( A => A(9), ZN => n18);
   U28 : INV_X1 port map( A => n28, ZN => n19);
   U29 : INV_X1 port map( A => B(9), ZN => n20);
   U30 : INV_X1 port map( A => n30, ZN => n21);
   U31 : OAI221_X1 port map( B1 => n22, B2 => n23, C1 => n24, C2 => n17, A => 
                           n71, ZN => Z(13));
   U32 : INV_X1 port map( A => A(13), ZN => n22);
   U33 : INV_X1 port map( A => n28, ZN => n23);
   U34 : INV_X1 port map( A => B(13), ZN => n24);
   U35 : NAND2_X1 port map( A1 => A(28), A2 => n36, ZN => n25);
   U36 : NAND2_X1 port map( A1 => B(28), A2 => n38, ZN => n26);
   U37 : BUF_X2 port map( A => n28, Z => n35);
   U38 : NAND2_X1 port map( A1 => B(30), A2 => n40, ZN => n27);
   U39 : BUF_X2 port map( A => n29, Z => n33);
   U40 : BUF_X2 port map( A => n29, Z => n34);
   U41 : BUF_X1 port map( A => n28, Z => n36);
   U42 : BUF_X1 port map( A => n28, Z => n37);
   U43 : BUF_X1 port map( A => n29, Z => n32);
   U44 : BUF_X1 port map( A => n30, Z => n39);
   U45 : BUF_X1 port map( A => n31, Z => n41);
   U46 : BUF_X1 port map( A => n31, Z => n42);
   U47 : BUF_X1 port map( A => n31, Z => n43);
   U48 : AND2_X1 port map( A1 => n44, A2 => n1, ZN => n29);
   U49 : AND2_X1 port map( A1 => S(0), A2 => n1, ZN => n31);
   U50 : INV_X1 port map( A => S(0), ZN => n44);
   U51 : AOI22_X1 port map( A1 => C(0), A2 => n33, B1 => D(0), B2 => n42, ZN =>
                           n47);
   U52 : INV_X1 port map( A => S(1), ZN => n45);
   U53 : AOI22_X1 port map( A1 => A(0), A2 => n36, B1 => B(0), B2 => n39, ZN =>
                           n46);
   U54 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => Z(0));
   U55 : AOI22_X1 port map( A1 => C(1), A2 => n34, B1 => D(1), B2 => n41, ZN =>
                           n49);
   U56 : AOI22_X1 port map( A1 => A(1), A2 => n35, B1 => B(1), B2 => n2, ZN => 
                           n48);
   U57 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => Z(1));
   U58 : AOI22_X1 port map( A1 => C(2), A2 => n34, B1 => D(2), B2 => n43, ZN =>
                           n51);
   U59 : AOI22_X1 port map( A1 => A(2), A2 => n35, B1 => n6, B2 => B(2), ZN => 
                           n50);
   U60 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => Z(2));
   U61 : AOI22_X1 port map( A1 => C(3), A2 => n34, B1 => D(3), B2 => n43, ZN =>
                           n53);
   U62 : AOI22_X1 port map( A1 => A(3), A2 => n35, B1 => n7, B2 => B(3), ZN => 
                           n52);
   U63 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => Z(3));
   U64 : AOI22_X1 port map( A1 => C(4), A2 => n34, B1 => D(4), B2 => n43, ZN =>
                           n55);
   U65 : AOI22_X1 port map( A1 => A(4), A2 => n35, B1 => n30, B2 => B(4), ZN =>
                           n54);
   U66 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => Z(4));
   U67 : AOI22_X1 port map( A1 => C(5), A2 => n33, B1 => D(5), B2 => n43, ZN =>
                           n57);
   U68 : AOI22_X1 port map( A1 => A(5), A2 => n35, B1 => B(5), B2 => n6, ZN => 
                           n56);
   U69 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => Z(5));
   U70 : AOI22_X1 port map( A1 => C(6), A2 => n33, B1 => D(6), B2 => n43, ZN =>
                           n59);
   U71 : AOI22_X1 port map( A1 => A(6), A2 => n4, B1 => B(6), B2 => n3, ZN => 
                           n58);
   U72 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => Z(6));
   U73 : AOI22_X1 port map( A1 => C(7), A2 => n33, B1 => D(7), B2 => n43, ZN =>
                           n61);
   U74 : AOI22_X1 port map( A1 => A(7), A2 => n36, B1 => B(7), B2 => n3, ZN => 
                           n60);
   U75 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => Z(7));
   U76 : AOI22_X1 port map( A1 => C(8), A2 => n33, B1 => D(8), B2 => n42, ZN =>
                           n63);
   U77 : AOI22_X1 port map( A1 => A(8), A2 => n37, B1 => B(8), B2 => n40, ZN =>
                           n62);
   U78 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => Z(8));
   U79 : AOI22_X1 port map( A1 => C(9), A2 => n33, B1 => D(9), B2 => n43, ZN =>
                           n64);
   U80 : AOI22_X1 port map( A1 => C(10), A2 => n33, B1 => D(10), B2 => n42, ZN 
                           => n66);
   U81 : AOI22_X1 port map( A1 => A(10), A2 => n5, B1 => B(10), B2 => n7, ZN =>
                           n65);
   U82 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => Z(10));
   U83 : AOI22_X1 port map( A1 => C(11), A2 => n33, B1 => D(11), B2 => n42, ZN 
                           => n68);
   U84 : AOI22_X1 port map( A1 => A(11), A2 => n5, B1 => B(11), B2 => n2, ZN =>
                           n67);
   U85 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => Z(11));
   U86 : AOI22_X1 port map( A1 => C(12), A2 => n33, B1 => D(12), B2 => n42, ZN 
                           => n70);
   U87 : AOI22_X1 port map( A1 => A(12), A2 => n5, B1 => B(12), B2 => n38, ZN 
                           => n69);
   U88 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => Z(12));
   U89 : AOI22_X1 port map( A1 => C(13), A2 => n33, B1 => D(13), B2 => n42, ZN 
                           => n71);
   U90 : AOI22_X1 port map( A1 => C(14), A2 => n33, B1 => D(14), B2 => n42, ZN 
                           => n72);
   U91 : AOI22_X1 port map( A1 => C(15), A2 => n33, B1 => D(15), B2 => n42, ZN 
                           => n74);
   U92 : NAND2_X1 port map( A1 => n73, A2 => n74, ZN => Z(15));
   U93 : AOI22_X1 port map( A1 => C(16), A2 => n32, B1 => D(16), B2 => n42, ZN 
                           => n76);
   U94 : AOI22_X1 port map( A1 => A(16), A2 => n37, B1 => B(16), B2 => n38, ZN 
                           => n75);
   U95 : NAND2_X1 port map( A1 => n75, A2 => n76, ZN => Z(16));
   U96 : AOI22_X1 port map( A1 => C(17), A2 => n32, B1 => D(17), B2 => n42, ZN 
                           => n78);
   U97 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n7, ZN =>
                           n77);
   U98 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => Z(17));
   U99 : AOI22_X1 port map( A1 => C(18), A2 => n32, B1 => D(18), B2 => n42, ZN 
                           => n80);
   U100 : AOI22_X1 port map( A1 => A(18), A2 => n5, B1 => B(18), B2 => n3, ZN 
                           => n79);
   U101 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => Z(18));
   U102 : AOI22_X1 port map( A1 => A(19), A2 => n37, B1 => C(19), B2 => n34, ZN
                           => n82);
   U103 : AOI22_X1 port map( A1 => D(19), A2 => n41, B1 => B(19), B2 => n40, ZN
                           => n81);
   U104 : NAND2_X1 port map( A1 => n82, A2 => n81, ZN => Z(19));
   U105 : AOI22_X1 port map( A1 => C(20), A2 => n32, B1 => D(20), B2 => n42, ZN
                           => n84);
   U106 : AOI22_X1 port map( A1 => A(20), A2 => n36, B1 => B(20), B2 => n2, ZN 
                           => n83);
   U107 : NAND2_X1 port map( A1 => n83, A2 => n84, ZN => Z(20));
   U108 : AOI22_X1 port map( A1 => C(21), A2 => n32, B1 => D(21), B2 => n41, ZN
                           => n86);
   U109 : AOI22_X1 port map( A1 => A(21), A2 => n4, B1 => B(21), B2 => n6, ZN 
                           => n85);
   U110 : NAND2_X1 port map( A1 => n85, A2 => n86, ZN => Z(21));
   U111 : AOI22_X1 port map( A1 => C(22), A2 => n32, B1 => D(22), B2 => n41, ZN
                           => n88);
   U112 : AOI22_X1 port map( A1 => A(22), A2 => n4, B1 => B(22), B2 => n38, ZN 
                           => n87);
   U113 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => Z(22));
   U114 : NAND2_X1 port map( A1 => A(23), A2 => n5, ZN => n90);
   U115 : AOI222_X1 port map( A1 => B(23), A2 => n3, B1 => C(23), B2 => n34, C1
                           => D(23), C2 => n43, ZN => n89);
   U116 : NAND2_X1 port map( A1 => n90, A2 => n89, ZN => Z(23));
   U117 : AOI22_X1 port map( A1 => C(24), A2 => n32, B1 => D(24), B2 => n41, ZN
                           => n92);
   U118 : AOI22_X1 port map( A1 => A(24), A2 => n36, B1 => B(24), B2 => n39, ZN
                           => n91);
   U119 : NAND2_X1 port map( A1 => n91, A2 => n92, ZN => Z(24));
   U120 : AOI22_X1 port map( A1 => C(25), A2 => n32, B1 => D(25), B2 => n41, ZN
                           => n94);
   U121 : AOI22_X1 port map( A1 => A(25), A2 => n37, B1 => B(25), B2 => n6, ZN 
                           => n93);
   U122 : NAND2_X1 port map( A1 => n93, A2 => n94, ZN => Z(25));
   U123 : AOI22_X1 port map( A1 => C(26), A2 => n32, B1 => D(26), B2 => n41, ZN
                           => n96);
   U124 : AOI22_X1 port map( A1 => A(26), A2 => n37, B1 => B(26), B2 => n39, ZN
                           => n95);
   U125 : NAND2_X1 port map( A1 => n95, A2 => n96, ZN => Z(26));
   U126 : AOI22_X1 port map( A1 => A(27), A2 => n5, B1 => C(27), B2 => n34, ZN 
                           => n98);
   U127 : AOI22_X1 port map( A1 => D(27), A2 => n41, B1 => B(27), B2 => n39, ZN
                           => n97);
   U128 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => Z(27));
   U129 : AOI22_X1 port map( A1 => C(28), A2 => n32, B1 => D(28), B2 => n41, ZN
                           => n99);
   U130 : NAND2_X1 port map( A1 => n25, A2 => n8, ZN => Z(28));
   U131 : AOI22_X1 port map( A1 => C(29), A2 => n32, B1 => D(29), B2 => n41, ZN
                           => n100);
   U132 : AOI22_X1 port map( A1 => C(30), A2 => n32, B1 => D(30), B2 => n41, ZN
                           => n101);
   U133 : AOI22_X1 port map( A1 => A(31), A2 => n4, B1 => C(31), B2 => n34, ZN 
                           => n103);
   U134 : AOI22_X1 port map( A1 => D(31), A2 => n41, B1 => B(31), B2 => n7, ZN 
                           => n102);
   U135 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(31));

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_1 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_1;

architecture SYN_bhv of mux41_NBIT32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n145, Z => n72);
   U2 : BUF_X1 port map( A => n145, Z => n73);
   U3 : BUF_X1 port map( A => n147, Z => n78);
   U4 : BUF_X1 port map( A => n147, Z => n79);
   U5 : BUF_X1 port map( A => n144, Z => n1);
   U6 : BUF_X1 port map( A => n144, Z => n70);
   U7 : BUF_X1 port map( A => n146, Z => n75);
   U8 : BUF_X1 port map( A => n146, Z => n76);
   U9 : BUF_X1 port map( A => n145, Z => n74);
   U10 : BUF_X1 port map( A => n147, Z => n80);
   U11 : BUF_X1 port map( A => n144, Z => n71);
   U12 : BUF_X1 port map( A => n146, Z => n77);
   U13 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n144);
   U14 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n145);
   U15 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n147);
   U16 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n146);
   U17 : INV_X1 port map( A => S(0), ZN => n81);
   U18 : NAND2_X1 port map( A1 => n83, A2 => n82, ZN => Z(0));
   U19 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n83);
   U20 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n82);
   U21 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(31));
   U22 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN 
                           => n130);
   U23 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN 
                           => n131);
   U24 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(7));
   U25 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n140);
   U26 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n141);
   U27 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(8));
   U28 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n142);
   U29 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n143);
   U30 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(9));
   U31 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN =>
                           n148);
   U32 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN =>
                           n149);
   U33 : NAND2_X1 port map( A1 => n87, A2 => n86, ZN => Z(11));
   U34 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN 
                           => n86);
   U35 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n87);
   U36 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => Z(12));
   U37 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN 
                           => n88);
   U38 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n89);
   U39 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => Z(13));
   U40 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN 
                           => n90);
   U41 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n91);
   U42 : NAND2_X1 port map( A1 => n93, A2 => n92, ZN => Z(14));
   U43 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN 
                           => n92);
   U44 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n93);
   U45 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(17));
   U46 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n98);
   U47 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n99);
   U48 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => Z(15));
   U49 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN 
                           => n94);
   U50 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n95);
   U51 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(18));
   U52 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n100);
   U53 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n101);
   U54 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(19));
   U55 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN 
                           => n102);
   U56 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n103);
   U57 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(20));
   U58 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN 
                           => n106);
   U59 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN 
                           => n107);
   U60 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(21));
   U61 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n108);
   U62 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n109);
   U63 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(22));
   U64 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n110);
   U65 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n111);
   U66 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(23));
   U67 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN 
                           => n112);
   U68 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN 
                           => n113);
   U69 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(24));
   U70 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN 
                           => n114);
   U71 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN 
                           => n115);
   U72 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(25));
   U73 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n116);
   U74 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n117);
   U75 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(5));
   U76 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN =>
                           n136);
   U77 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN =>
                           n137);
   U78 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(6));
   U79 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n138);
   U80 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n139);
   U81 : NAND2_X1 port map( A1 => n85, A2 => n84, ZN => Z(10));
   U82 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN 
                           => n84);
   U83 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n85);
   U84 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(16));
   U85 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n96);
   U86 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n97);
   U87 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(26));
   U88 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n118);
   U89 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n119);
   U90 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(27));
   U91 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN 
                           => n120);
   U92 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN 
                           => n121);
   U93 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(28));
   U94 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n122);
   U95 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n123);
   U96 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(29));
   U97 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n124);
   U98 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n125);
   U99 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(30));
   U100 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN
                           => n128);
   U101 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN
                           => n129);
   U102 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(2));
   U103 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN 
                           => n126);
   U104 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN 
                           => n127);
   U105 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(1));
   U106 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN 
                           => n104);
   U107 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN =>
                           n105);
   U108 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(3));
   U109 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN 
                           => n132);
   U110 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN 
                           => n133);
   U111 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(4));
   U112 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN 
                           => n134);
   U113 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN 
                           => n135);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_4 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_4;

architecture SYN_bhv of regn_N5_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DOUT_0_port, DOUT_1_port, DOUT_2_port, DOUT_3_port, DOUT_4_port, n6, 
      n7, n8, n9, n10, n_1120, n_1121, n_1122, n_1123, n_1124 : std_logic;

begin
   DOUT <= ( DOUT_4_port, DOUT_3_port, DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n6, CK => CLK, RN => RST, Q => 
                           DOUT_4_port, QN => n_1120);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n7, CK => CLK, RN => RST, Q => 
                           DOUT_3_port, QN => n_1121);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n8, CK => CLK, RN => RST, Q => 
                           DOUT_2_port, QN => n_1122);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n9, CK => CLK, RN => RST, Q => 
                           DOUT_1_port, QN => n_1123);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n10, CK => CLK, RN => RST, Q => 
                           DOUT_0_port, QN => n_1124);
   U2 : MUX2_X1 port map( A => DOUT_0_port, B => DIN(0), S => EN, Z => n10);
   U3 : MUX2_X1 port map( A => DOUT_1_port, B => DIN(1), S => EN, Z => n9);
   U4 : MUX2_X1 port map( A => DOUT_2_port, B => DIN(2), S => EN, Z => n8);
   U5 : MUX2_X1 port map( A => DOUT_3_port, B => DIN(3), S => EN, Z => n7);
   U6 : MUX2_X1 port map( A => DOUT_4_port, B => DIN(4), S => EN, Z => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_3 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_3;

architecture SYN_bhv of regn_N5_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DOUT_0_port, DOUT_1_port, DOUT_2_port, DOUT_3_port, DOUT_4_port, n6, 
      n7, n8, n9, n10, n_1125, n_1126, n_1127, n_1128, n_1129 : std_logic;

begin
   DOUT <= ( DOUT_4_port, DOUT_3_port, DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n6, CK => CLK, RN => RST, Q => 
                           DOUT_4_port, QN => n_1125);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n7, CK => CLK, RN => RST, Q => 
                           DOUT_3_port, QN => n_1126);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n8, CK => CLK, RN => RST, Q => 
                           DOUT_2_port, QN => n_1127);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n9, CK => CLK, RN => RST, Q => 
                           DOUT_1_port, QN => n_1128);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n10, CK => CLK, RN => RST, Q => 
                           DOUT_0_port, QN => n_1129);
   U2 : MUX2_X1 port map( A => DOUT_0_port, B => DIN(0), S => EN, Z => n10);
   U3 : MUX2_X1 port map( A => DOUT_1_port, B => DIN(1), S => EN, Z => n9);
   U4 : MUX2_X1 port map( A => DOUT_2_port, B => DIN(2), S => EN, Z => n8);
   U5 : MUX2_X1 port map( A => DOUT_3_port, B => DIN(3), S => EN, Z => n7);
   U6 : MUX2_X1 port map( A => DOUT_4_port, B => DIN(4), S => EN, Z => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_2 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_2;

architecture SYN_bhv of regn_N5_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DOUT_0_port, DOUT_1_port, DOUT_2_port, DOUT_3_port, DOUT_4_port, n6, 
      n7, n8, n9, n10, n_1130, n_1131, n_1132, n_1133, n_1134 : std_logic;

begin
   DOUT <= ( DOUT_4_port, DOUT_3_port, DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n6, CK => CLK, RN => RST, Q => 
                           DOUT_4_port, QN => n_1130);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n7, CK => CLK, RN => RST, Q => 
                           DOUT_3_port, QN => n_1131);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n8, CK => CLK, RN => RST, Q => 
                           DOUT_2_port, QN => n_1132);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n9, CK => CLK, RN => RST, Q => 
                           DOUT_1_port, QN => n_1133);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n10, CK => CLK, RN => RST, Q => 
                           DOUT_0_port, QN => n_1134);
   U2 : MUX2_X1 port map( A => DOUT_0_port, B => DIN(0), S => EN, Z => n10);
   U3 : MUX2_X1 port map( A => DOUT_1_port, B => DIN(1), S => EN, Z => n9);
   U4 : MUX2_X1 port map( A => DOUT_2_port, B => DIN(2), S => EN, Z => n8);
   U5 : MUX2_X1 port map( A => DOUT_3_port, B => DIN(3), S => EN, Z => n7);
   U6 : MUX2_X1 port map( A => DOUT_4_port, B => DIN(4), S => EN, Z => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_1 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_1;

architecture SYN_bhv of regn_N5_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DOUT_0_port, DOUT_1_port, DOUT_2_port, DOUT_3_port, DOUT_4_port, n6, 
      n7, n8, n9, n10, n_1135, n_1136, n_1137, n_1138, n_1139 : std_logic;

begin
   DOUT <= ( DOUT_4_port, DOUT_3_port, DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n6, CK => CLK, RN => RST, Q => 
                           DOUT_4_port, QN => n_1135);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n7, CK => CLK, RN => RST, Q => 
                           DOUT_3_port, QN => n_1136);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n8, CK => CLK, RN => RST, Q => 
                           DOUT_2_port, QN => n_1137);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n9, CK => CLK, RN => RST, Q => 
                           DOUT_1_port, QN => n_1138);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n10, CK => CLK, RN => RST, Q => 
                           DOUT_0_port, QN => n_1139);
   U2 : MUX2_X1 port map( A => DOUT_0_port, B => DIN(0), S => EN, Z => n10);
   U3 : MUX2_X1 port map( A => DOUT_1_port, B => DIN(1), S => EN, Z => n9);
   U4 : MUX2_X1 port map( A => DOUT_2_port, B => DIN(2), S => EN, Z => n8);
   U5 : MUX2_X1 port map( A => DOUT_3_port, B => DIN(3), S => EN, Z => n7);
   U6 : MUX2_X1 port map( A => DOUT_4_port, B => DIN(4), S => EN, Z => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_10 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_10;

architecture SYN_bhv of regn_N32_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, DOUT_0_port, DOUT_1_port, DOUT_2_port, DOUT_3_port, 
      DOUT_4_port, DOUT_5_port, DOUT_6_port, DOUT_7_port, DOUT_8_port, 
      DOUT_9_port, DOUT_10_port, DOUT_11_port, DOUT_12_port, DOUT_13_port, 
      DOUT_14_port, DOUT_15_port, DOUT_16_port, DOUT_17_port, DOUT_18_port, 
      DOUT_19_port, DOUT_20_port, DOUT_21_port, DOUT_22_port, DOUT_23_port, 
      DOUT_24_port, DOUT_25_port, DOUT_26_port, DOUT_27_port, DOUT_28_port, 
      DOUT_29_port, DOUT_30_port, DOUT_31_port, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n68, n69, n70, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, 
      n_1169, n_1170, n_1171 : std_logic;

begin
   DOUT <= ( DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, 
      DOUT_27_port, DOUT_26_port, DOUT_25_port, DOUT_24_port, DOUT_23_port, 
      DOUT_22_port, DOUT_21_port, DOUT_20_port, DOUT_19_port, DOUT_18_port, 
      DOUT_17_port, DOUT_16_port, DOUT_15_port, DOUT_14_port, DOUT_13_port, 
      DOUT_12_port, DOUT_11_port, DOUT_10_port, DOUT_9_port, DOUT_8_port, 
      DOUT_7_port, DOUT_6_port, DOUT_5_port, DOUT_4_port, DOUT_3_port, 
      DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n36, CK => CLK, RN => n3, Q => 
                           DOUT_31_port, QN => n_1140);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n37, CK => CLK, RN => n3, Q => 
                           DOUT_30_port, QN => n_1141);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n38, CK => CLK, RN => n3, Q => 
                           DOUT_29_port, QN => n_1142);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n39, CK => CLK, RN => n3, Q => 
                           DOUT_28_port, QN => n_1143);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n40, CK => CLK, RN => n3, Q => 
                           DOUT_27_port, QN => n_1144);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n41, CK => CLK, RN => n3, Q => 
                           DOUT_26_port, QN => n_1145);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n42, CK => CLK, RN => n3, Q => 
                           DOUT_25_port, QN => n_1146);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n43, CK => CLK, RN => n3, Q => 
                           DOUT_24_port, QN => n_1147);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n44, CK => CLK, RN => n2, Q => 
                           DOUT_23_port, QN => n_1148);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n45, CK => CLK, RN => n2, Q => 
                           DOUT_22_port, QN => n_1149);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n46, CK => CLK, RN => n2, Q => 
                           DOUT_21_port, QN => n_1150);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n47, CK => CLK, RN => n2, Q => 
                           DOUT_20_port, QN => n_1151);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n48, CK => CLK, RN => n2, Q => 
                           DOUT_19_port, QN => n_1152);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n49, CK => CLK, RN => n2, Q => 
                           DOUT_18_port, QN => n_1153);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n50, CK => CLK, RN => n2, Q => 
                           DOUT_17_port, QN => n_1154);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n51, CK => CLK, RN => n2, Q => 
                           DOUT_16_port, QN => n_1155);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n52, CK => CLK, RN => n2, Q => 
                           DOUT_15_port, QN => n_1156);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n53, CK => CLK, RN => n2, Q => 
                           DOUT_14_port, QN => n_1157);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n54, CK => CLK, RN => n2, Q => 
                           DOUT_13_port, QN => n_1158);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n55, CK => CLK, RN => n2, Q => 
                           DOUT_12_port, QN => n_1159);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n56, CK => CLK, RN => n1, Q => 
                           DOUT_11_port, QN => n_1160);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n57, CK => CLK, RN => n1, Q => 
                           DOUT_10_port, QN => n_1161);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n58, CK => CLK, RN => n1, Q => 
                           DOUT_9_port, QN => n_1162);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n59, CK => CLK, RN => n1, Q => 
                           DOUT_8_port, QN => n_1163);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n60, CK => CLK, RN => n1, Q => 
                           DOUT_7_port, QN => n_1164);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n61, CK => CLK, RN => n1, Q => 
                           DOUT_6_port, QN => n_1165);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n62, CK => CLK, RN => n1, Q => 
                           DOUT_5_port, QN => n_1166);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n63, CK => CLK, RN => n1, Q => 
                           DOUT_4_port, QN => n_1167);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n64, CK => CLK, RN => n1, Q => 
                           DOUT_3_port, QN => n_1168);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n68, CK => CLK, RN => n1, Q => 
                           DOUT_2_port, QN => n_1169);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n69, CK => CLK, RN => n1, Q => 
                           DOUT_1_port, QN => n_1170);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n70, CK => CLK, RN => n1, Q => 
                           DOUT_0_port, QN => n_1171);
   U2 : BUF_X1 port map( A => RST, Z => n1);
   U3 : BUF_X1 port map( A => RST, Z => n2);
   U4 : BUF_X1 port map( A => RST, Z => n3);
   U5 : MUX2_X1 port map( A => DOUT_0_port, B => DIN(0), S => EN, Z => n70);
   U6 : MUX2_X1 port map( A => DOUT_1_port, B => DIN(1), S => EN, Z => n69);
   U7 : MUX2_X1 port map( A => DOUT_2_port, B => DIN(2), S => EN, Z => n68);
   U8 : MUX2_X1 port map( A => DOUT_3_port, B => DIN(3), S => EN, Z => n64);
   U9 : MUX2_X1 port map( A => DOUT_4_port, B => DIN(4), S => EN, Z => n63);
   U10 : MUX2_X1 port map( A => DOUT_5_port, B => DIN(5), S => EN, Z => n62);
   U11 : MUX2_X1 port map( A => DOUT_6_port, B => DIN(6), S => EN, Z => n61);
   U12 : MUX2_X1 port map( A => DOUT_7_port, B => DIN(7), S => EN, Z => n60);
   U13 : MUX2_X1 port map( A => DOUT_8_port, B => DIN(8), S => EN, Z => n59);
   U14 : MUX2_X1 port map( A => DOUT_9_port, B => DIN(9), S => EN, Z => n58);
   U15 : MUX2_X1 port map( A => DOUT_10_port, B => DIN(10), S => EN, Z => n57);
   U16 : MUX2_X1 port map( A => DOUT_11_port, B => DIN(11), S => EN, Z => n56);
   U17 : MUX2_X1 port map( A => DOUT_12_port, B => DIN(12), S => EN, Z => n55);
   U18 : MUX2_X1 port map( A => DOUT_13_port, B => DIN(13), S => EN, Z => n54);
   U19 : MUX2_X1 port map( A => DOUT_14_port, B => DIN(14), S => EN, Z => n53);
   U20 : MUX2_X1 port map( A => DOUT_15_port, B => DIN(15), S => EN, Z => n52);
   U21 : MUX2_X1 port map( A => DOUT_16_port, B => DIN(16), S => EN, Z => n51);
   U22 : MUX2_X1 port map( A => DOUT_17_port, B => DIN(17), S => EN, Z => n50);
   U23 : MUX2_X1 port map( A => DOUT_18_port, B => DIN(18), S => EN, Z => n49);
   U24 : MUX2_X1 port map( A => DOUT_19_port, B => DIN(19), S => EN, Z => n48);
   U25 : MUX2_X1 port map( A => DOUT_20_port, B => DIN(20), S => EN, Z => n47);
   U26 : MUX2_X1 port map( A => DOUT_21_port, B => DIN(21), S => EN, Z => n46);
   U27 : MUX2_X1 port map( A => DOUT_22_port, B => DIN(22), S => EN, Z => n45);
   U28 : MUX2_X1 port map( A => DOUT_23_port, B => DIN(23), S => EN, Z => n44);
   U29 : MUX2_X1 port map( A => DOUT_24_port, B => DIN(24), S => EN, Z => n43);
   U30 : MUX2_X1 port map( A => DOUT_25_port, B => DIN(25), S => EN, Z => n42);
   U31 : MUX2_X1 port map( A => DOUT_26_port, B => DIN(26), S => EN, Z => n41);
   U32 : MUX2_X1 port map( A => DOUT_27_port, B => DIN(27), S => EN, Z => n40);
   U33 : MUX2_X1 port map( A => DOUT_28_port, B => DIN(28), S => EN, Z => n39);
   U34 : MUX2_X1 port map( A => DOUT_29_port, B => DIN(29), S => EN, Z => n38);
   U35 : MUX2_X1 port map( A => DOUT_30_port, B => DIN(30), S => EN, Z => n37);
   U36 : MUX2_X1 port map( A => DOUT_31_port, B => DIN(31), S => EN, Z => n36);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_9 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_9;

architecture SYN_bhv of regn_N32_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U6 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U7 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U8 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U9 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U10 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U11 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U12 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U13 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U14 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U15 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U16 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U17 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U18 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U19 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U20 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U21 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U22 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U23 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U24 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U25 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U26 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U27 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U28 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U29 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U30 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U31 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U32 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U33 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U34 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U35 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U36 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U37 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U38 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U39 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U40 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U41 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U42 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U43 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U44 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U45 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U46 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U47 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U48 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U49 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U50 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U51 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U52 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U53 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U54 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U55 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U56 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U57 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U58 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U59 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U60 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U61 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U62 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U63 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U64 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);
   U65 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U66 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U67 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U68 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_8 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_8;

architecture SYN_bhv of regn_N32_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, DOUT_0_port, DOUT_1_port, DOUT_2_port, DOUT_3_port, 
      DOUT_4_port, DOUT_5_port, DOUT_6_port, DOUT_7_port, DOUT_8_port, 
      DOUT_9_port, DOUT_10_port, DOUT_11_port, DOUT_12_port, DOUT_13_port, 
      DOUT_14_port, DOUT_15_port, DOUT_16_port, DOUT_17_port, DOUT_18_port, 
      DOUT_19_port, DOUT_20_port, DOUT_21_port, DOUT_22_port, DOUT_23_port, 
      DOUT_24_port, DOUT_25_port, DOUT_26_port, DOUT_27_port, DOUT_28_port, 
      DOUT_29_port, DOUT_30_port, DOUT_31_port, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n68, n69, n70, n_1172, n_1173, 
      n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, 
      n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, 
      n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, 
      n_1201, n_1202, n_1203 : std_logic;

begin
   DOUT <= ( DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, 
      DOUT_27_port, DOUT_26_port, DOUT_25_port, DOUT_24_port, DOUT_23_port, 
      DOUT_22_port, DOUT_21_port, DOUT_20_port, DOUT_19_port, DOUT_18_port, 
      DOUT_17_port, DOUT_16_port, DOUT_15_port, DOUT_14_port, DOUT_13_port, 
      DOUT_12_port, DOUT_11_port, DOUT_10_port, DOUT_9_port, DOUT_8_port, 
      DOUT_7_port, DOUT_6_port, DOUT_5_port, DOUT_4_port, DOUT_3_port, 
      DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n36, CK => CLK, RN => n3, Q => 
                           DOUT_31_port, QN => n_1172);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n37, CK => CLK, RN => n3, Q => 
                           DOUT_30_port, QN => n_1173);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n38, CK => CLK, RN => n3, Q => 
                           DOUT_29_port, QN => n_1174);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n39, CK => CLK, RN => n3, Q => 
                           DOUT_28_port, QN => n_1175);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n40, CK => CLK, RN => n3, Q => 
                           DOUT_27_port, QN => n_1176);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n41, CK => CLK, RN => n3, Q => 
                           DOUT_26_port, QN => n_1177);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n42, CK => CLK, RN => n3, Q => 
                           DOUT_25_port, QN => n_1178);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n43, CK => CLK, RN => n3, Q => 
                           DOUT_24_port, QN => n_1179);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n44, CK => CLK, RN => n2, Q => 
                           DOUT_23_port, QN => n_1180);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n45, CK => CLK, RN => n2, Q => 
                           DOUT_22_port, QN => n_1181);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n46, CK => CLK, RN => n2, Q => 
                           DOUT_21_port, QN => n_1182);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n47, CK => CLK, RN => n2, Q => 
                           DOUT_20_port, QN => n_1183);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n48, CK => CLK, RN => n2, Q => 
                           DOUT_19_port, QN => n_1184);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n49, CK => CLK, RN => n2, Q => 
                           DOUT_18_port, QN => n_1185);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n50, CK => CLK, RN => n2, Q => 
                           DOUT_17_port, QN => n_1186);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n51, CK => CLK, RN => n2, Q => 
                           DOUT_16_port, QN => n_1187);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n52, CK => CLK, RN => n2, Q => 
                           DOUT_15_port, QN => n_1188);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n53, CK => CLK, RN => n2, Q => 
                           DOUT_14_port, QN => n_1189);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n54, CK => CLK, RN => n2, Q => 
                           DOUT_13_port, QN => n_1190);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n55, CK => CLK, RN => n2, Q => 
                           DOUT_12_port, QN => n_1191);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n56, CK => CLK, RN => n1, Q => 
                           DOUT_11_port, QN => n_1192);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n57, CK => CLK, RN => n1, Q => 
                           DOUT_10_port, QN => n_1193);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n58, CK => CLK, RN => n1, Q => 
                           DOUT_9_port, QN => n_1194);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n59, CK => CLK, RN => n1, Q => 
                           DOUT_8_port, QN => n_1195);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n60, CK => CLK, RN => n1, Q => 
                           DOUT_7_port, QN => n_1196);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n61, CK => CLK, RN => n1, Q => 
                           DOUT_6_port, QN => n_1197);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n62, CK => CLK, RN => n1, Q => 
                           DOUT_5_port, QN => n_1198);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n63, CK => CLK, RN => n1, Q => 
                           DOUT_4_port, QN => n_1199);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n64, CK => CLK, RN => n1, Q => 
                           DOUT_3_port, QN => n_1200);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n68, CK => CLK, RN => n1, Q => 
                           DOUT_2_port, QN => n_1201);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n69, CK => CLK, RN => n1, Q => 
                           DOUT_1_port, QN => n_1202);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n70, CK => CLK, RN => n1, Q => 
                           DOUT_0_port, QN => n_1203);
   U2 : BUF_X1 port map( A => RST, Z => n1);
   U3 : BUF_X1 port map( A => RST, Z => n2);
   U4 : BUF_X1 port map( A => RST, Z => n3);
   U5 : MUX2_X1 port map( A => DOUT_0_port, B => DIN(0), S => EN, Z => n70);
   U6 : MUX2_X1 port map( A => DOUT_1_port, B => DIN(1), S => EN, Z => n69);
   U7 : MUX2_X1 port map( A => DOUT_2_port, B => DIN(2), S => EN, Z => n68);
   U8 : MUX2_X1 port map( A => DOUT_3_port, B => DIN(3), S => EN, Z => n64);
   U9 : MUX2_X1 port map( A => DOUT_4_port, B => DIN(4), S => EN, Z => n63);
   U10 : MUX2_X1 port map( A => DOUT_5_port, B => DIN(5), S => EN, Z => n62);
   U11 : MUX2_X1 port map( A => DOUT_6_port, B => DIN(6), S => EN, Z => n61);
   U12 : MUX2_X1 port map( A => DOUT_7_port, B => DIN(7), S => EN, Z => n60);
   U13 : MUX2_X1 port map( A => DOUT_8_port, B => DIN(8), S => EN, Z => n59);
   U14 : MUX2_X1 port map( A => DOUT_9_port, B => DIN(9), S => EN, Z => n58);
   U15 : MUX2_X1 port map( A => DOUT_10_port, B => DIN(10), S => EN, Z => n57);
   U16 : MUX2_X1 port map( A => DOUT_11_port, B => DIN(11), S => EN, Z => n56);
   U17 : MUX2_X1 port map( A => DOUT_12_port, B => DIN(12), S => EN, Z => n55);
   U18 : MUX2_X1 port map( A => DOUT_13_port, B => DIN(13), S => EN, Z => n54);
   U19 : MUX2_X1 port map( A => DOUT_14_port, B => DIN(14), S => EN, Z => n53);
   U20 : MUX2_X1 port map( A => DOUT_15_port, B => DIN(15), S => EN, Z => n52);
   U21 : MUX2_X1 port map( A => DOUT_16_port, B => DIN(16), S => EN, Z => n51);
   U22 : MUX2_X1 port map( A => DOUT_17_port, B => DIN(17), S => EN, Z => n50);
   U23 : MUX2_X1 port map( A => DOUT_18_port, B => DIN(18), S => EN, Z => n49);
   U24 : MUX2_X1 port map( A => DOUT_19_port, B => DIN(19), S => EN, Z => n48);
   U25 : MUX2_X1 port map( A => DOUT_20_port, B => DIN(20), S => EN, Z => n47);
   U26 : MUX2_X1 port map( A => DOUT_21_port, B => DIN(21), S => EN, Z => n46);
   U27 : MUX2_X1 port map( A => DOUT_22_port, B => DIN(22), S => EN, Z => n45);
   U28 : MUX2_X1 port map( A => DOUT_23_port, B => DIN(23), S => EN, Z => n44);
   U29 : MUX2_X1 port map( A => DOUT_24_port, B => DIN(24), S => EN, Z => n43);
   U30 : MUX2_X1 port map( A => DOUT_25_port, B => DIN(25), S => EN, Z => n42);
   U31 : MUX2_X1 port map( A => DOUT_26_port, B => DIN(26), S => EN, Z => n41);
   U32 : MUX2_X1 port map( A => DOUT_27_port, B => DIN(27), S => EN, Z => n40);
   U33 : MUX2_X1 port map( A => DOUT_28_port, B => DIN(28), S => EN, Z => n39);
   U34 : MUX2_X1 port map( A => DOUT_29_port, B => DIN(29), S => EN, Z => n38);
   U35 : MUX2_X1 port map( A => DOUT_30_port, B => DIN(30), S => EN, Z => n37);
   U36 : MUX2_X1 port map( A => DOUT_31_port, B => DIN(31), S => EN, Z => n36);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_7 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_7;

architecture SYN_bhv of regn_N32_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, DOUT_0_port, DOUT_1_port, DOUT_2_port, DOUT_3_port, 
      DOUT_4_port, DOUT_5_port, DOUT_6_port, DOUT_7_port, DOUT_8_port, 
      DOUT_9_port, DOUT_10_port, DOUT_11_port, DOUT_12_port, DOUT_13_port, 
      DOUT_14_port, DOUT_15_port, DOUT_16_port, DOUT_17_port, DOUT_18_port, 
      DOUT_19_port, DOUT_20_port, DOUT_21_port, DOUT_22_port, DOUT_23_port, 
      DOUT_24_port, DOUT_25_port, DOUT_26_port, DOUT_27_port, DOUT_28_port, 
      DOUT_29_port, DOUT_30_port, DOUT_31_port, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n68, n69, n70, n_1204, n_1205, 
      n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, 
      n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, 
      n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, 
      n_1233, n_1234, n_1235 : std_logic;

begin
   DOUT <= ( DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, 
      DOUT_27_port, DOUT_26_port, DOUT_25_port, DOUT_24_port, DOUT_23_port, 
      DOUT_22_port, DOUT_21_port, DOUT_20_port, DOUT_19_port, DOUT_18_port, 
      DOUT_17_port, DOUT_16_port, DOUT_15_port, DOUT_14_port, DOUT_13_port, 
      DOUT_12_port, DOUT_11_port, DOUT_10_port, DOUT_9_port, DOUT_8_port, 
      DOUT_7_port, DOUT_6_port, DOUT_5_port, DOUT_4_port, DOUT_3_port, 
      DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n36, CK => CLK, RN => n3, Q => 
                           DOUT_31_port, QN => n_1204);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n37, CK => CLK, RN => n3, Q => 
                           DOUT_30_port, QN => n_1205);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n38, CK => CLK, RN => n3, Q => 
                           DOUT_29_port, QN => n_1206);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n39, CK => CLK, RN => n3, Q => 
                           DOUT_28_port, QN => n_1207);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n40, CK => CLK, RN => n3, Q => 
                           DOUT_27_port, QN => n_1208);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n41, CK => CLK, RN => n3, Q => 
                           DOUT_26_port, QN => n_1209);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n42, CK => CLK, RN => n3, Q => 
                           DOUT_25_port, QN => n_1210);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n43, CK => CLK, RN => n3, Q => 
                           DOUT_24_port, QN => n_1211);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n44, CK => CLK, RN => n2, Q => 
                           DOUT_23_port, QN => n_1212);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n45, CK => CLK, RN => n2, Q => 
                           DOUT_22_port, QN => n_1213);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n46, CK => CLK, RN => n2, Q => 
                           DOUT_21_port, QN => n_1214);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n47, CK => CLK, RN => n2, Q => 
                           DOUT_20_port, QN => n_1215);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n48, CK => CLK, RN => n2, Q => 
                           DOUT_19_port, QN => n_1216);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n49, CK => CLK, RN => n2, Q => 
                           DOUT_18_port, QN => n_1217);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n50, CK => CLK, RN => n2, Q => 
                           DOUT_17_port, QN => n_1218);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n51, CK => CLK, RN => n2, Q => 
                           DOUT_16_port, QN => n_1219);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n52, CK => CLK, RN => n2, Q => 
                           DOUT_15_port, QN => n_1220);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n53, CK => CLK, RN => n2, Q => 
                           DOUT_14_port, QN => n_1221);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n54, CK => CLK, RN => n2, Q => 
                           DOUT_13_port, QN => n_1222);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n55, CK => CLK, RN => n2, Q => 
                           DOUT_12_port, QN => n_1223);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n56, CK => CLK, RN => n1, Q => 
                           DOUT_11_port, QN => n_1224);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n57, CK => CLK, RN => n1, Q => 
                           DOUT_10_port, QN => n_1225);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n58, CK => CLK, RN => n1, Q => 
                           DOUT_9_port, QN => n_1226);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n59, CK => CLK, RN => n1, Q => 
                           DOUT_8_port, QN => n_1227);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n60, CK => CLK, RN => n1, Q => 
                           DOUT_7_port, QN => n_1228);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n61, CK => CLK, RN => n1, Q => 
                           DOUT_6_port, QN => n_1229);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n62, CK => CLK, RN => n1, Q => 
                           DOUT_5_port, QN => n_1230);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n63, CK => CLK, RN => n1, Q => 
                           DOUT_4_port, QN => n_1231);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n64, CK => CLK, RN => n1, Q => 
                           DOUT_3_port, QN => n_1232);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n68, CK => CLK, RN => n1, Q => 
                           DOUT_2_port, QN => n_1233);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n69, CK => CLK, RN => n1, Q => 
                           DOUT_1_port, QN => n_1234);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n70, CK => CLK, RN => n1, Q => 
                           DOUT_0_port, QN => n_1235);
   U2 : BUF_X1 port map( A => RST, Z => n1);
   U3 : BUF_X1 port map( A => RST, Z => n2);
   U4 : BUF_X1 port map( A => RST, Z => n3);
   U5 : MUX2_X1 port map( A => DOUT_0_port, B => DIN(0), S => EN, Z => n70);
   U6 : MUX2_X1 port map( A => DOUT_1_port, B => DIN(1), S => EN, Z => n69);
   U7 : MUX2_X1 port map( A => DOUT_2_port, B => DIN(2), S => EN, Z => n68);
   U8 : MUX2_X1 port map( A => DOUT_3_port, B => DIN(3), S => EN, Z => n64);
   U9 : MUX2_X1 port map( A => DOUT_4_port, B => DIN(4), S => EN, Z => n63);
   U10 : MUX2_X1 port map( A => DOUT_5_port, B => DIN(5), S => EN, Z => n62);
   U11 : MUX2_X1 port map( A => DOUT_6_port, B => DIN(6), S => EN, Z => n61);
   U12 : MUX2_X1 port map( A => DOUT_7_port, B => DIN(7), S => EN, Z => n60);
   U13 : MUX2_X1 port map( A => DOUT_8_port, B => DIN(8), S => EN, Z => n59);
   U14 : MUX2_X1 port map( A => DOUT_9_port, B => DIN(9), S => EN, Z => n58);
   U15 : MUX2_X1 port map( A => DOUT_10_port, B => DIN(10), S => EN, Z => n57);
   U16 : MUX2_X1 port map( A => DOUT_11_port, B => DIN(11), S => EN, Z => n56);
   U17 : MUX2_X1 port map( A => DOUT_12_port, B => DIN(12), S => EN, Z => n55);
   U18 : MUX2_X1 port map( A => DOUT_13_port, B => DIN(13), S => EN, Z => n54);
   U19 : MUX2_X1 port map( A => DOUT_14_port, B => DIN(14), S => EN, Z => n53);
   U20 : MUX2_X1 port map( A => DOUT_15_port, B => DIN(15), S => EN, Z => n52);
   U21 : MUX2_X1 port map( A => DOUT_16_port, B => DIN(16), S => EN, Z => n51);
   U22 : MUX2_X1 port map( A => DOUT_17_port, B => DIN(17), S => EN, Z => n50);
   U23 : MUX2_X1 port map( A => DOUT_18_port, B => DIN(18), S => EN, Z => n49);
   U24 : MUX2_X1 port map( A => DOUT_19_port, B => DIN(19), S => EN, Z => n48);
   U25 : MUX2_X1 port map( A => DOUT_20_port, B => DIN(20), S => EN, Z => n47);
   U26 : MUX2_X1 port map( A => DOUT_21_port, B => DIN(21), S => EN, Z => n46);
   U27 : MUX2_X1 port map( A => DOUT_22_port, B => DIN(22), S => EN, Z => n45);
   U28 : MUX2_X1 port map( A => DOUT_23_port, B => DIN(23), S => EN, Z => n44);
   U29 : MUX2_X1 port map( A => DOUT_24_port, B => DIN(24), S => EN, Z => n43);
   U30 : MUX2_X1 port map( A => DOUT_25_port, B => DIN(25), S => EN, Z => n42);
   U31 : MUX2_X1 port map( A => DOUT_26_port, B => DIN(26), S => EN, Z => n41);
   U32 : MUX2_X1 port map( A => DOUT_27_port, B => DIN(27), S => EN, Z => n40);
   U33 : MUX2_X1 port map( A => DOUT_28_port, B => DIN(28), S => EN, Z => n39);
   U34 : MUX2_X1 port map( A => DOUT_29_port, B => DIN(29), S => EN, Z => n38);
   U35 : MUX2_X1 port map( A => DOUT_30_port, B => DIN(30), S => EN, Z => n37);
   U36 : MUX2_X1 port map( A => DOUT_31_port, B => DIN(31), S => EN, Z => n36);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_6 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_6;

architecture SYN_bhv of regn_N32_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, DOUT_0_port, DOUT_1_port, DOUT_2_port, DOUT_3_port, 
      DOUT_4_port, DOUT_5_port, DOUT_6_port, DOUT_7_port, DOUT_8_port, 
      DOUT_9_port, DOUT_10_port, DOUT_11_port, DOUT_12_port, DOUT_13_port, 
      DOUT_14_port, DOUT_15_port, DOUT_16_port, DOUT_17_port, DOUT_18_port, 
      DOUT_19_port, DOUT_20_port, DOUT_21_port, DOUT_22_port, DOUT_23_port, 
      DOUT_24_port, DOUT_25_port, DOUT_26_port, DOUT_27_port, DOUT_28_port, 
      DOUT_29_port, DOUT_30_port, DOUT_31_port, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n68, n69, n70, n_1236, n_1237, 
      n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, 
      n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, 
      n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, 
      n_1265, n_1266, n_1267 : std_logic;

begin
   DOUT <= ( DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, 
      DOUT_27_port, DOUT_26_port, DOUT_25_port, DOUT_24_port, DOUT_23_port, 
      DOUT_22_port, DOUT_21_port, DOUT_20_port, DOUT_19_port, DOUT_18_port, 
      DOUT_17_port, DOUT_16_port, DOUT_15_port, DOUT_14_port, DOUT_13_port, 
      DOUT_12_port, DOUT_11_port, DOUT_10_port, DOUT_9_port, DOUT_8_port, 
      DOUT_7_port, DOUT_6_port, DOUT_5_port, DOUT_4_port, DOUT_3_port, 
      DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n36, CK => CLK, RN => n3, Q => 
                           DOUT_31_port, QN => n_1236);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n37, CK => CLK, RN => n3, Q => 
                           DOUT_30_port, QN => n_1237);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n38, CK => CLK, RN => n3, Q => 
                           DOUT_29_port, QN => n_1238);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n39, CK => CLK, RN => n3, Q => 
                           DOUT_28_port, QN => n_1239);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n40, CK => CLK, RN => n3, Q => 
                           DOUT_27_port, QN => n_1240);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n41, CK => CLK, RN => n3, Q => 
                           DOUT_26_port, QN => n_1241);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n42, CK => CLK, RN => n3, Q => 
                           DOUT_25_port, QN => n_1242);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n43, CK => CLK, RN => n3, Q => 
                           DOUT_24_port, QN => n_1243);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n44, CK => CLK, RN => n2, Q => 
                           DOUT_23_port, QN => n_1244);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n45, CK => CLK, RN => n2, Q => 
                           DOUT_22_port, QN => n_1245);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n46, CK => CLK, RN => n2, Q => 
                           DOUT_21_port, QN => n_1246);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n47, CK => CLK, RN => n2, Q => 
                           DOUT_20_port, QN => n_1247);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n48, CK => CLK, RN => n2, Q => 
                           DOUT_19_port, QN => n_1248);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n49, CK => CLK, RN => n2, Q => 
                           DOUT_18_port, QN => n_1249);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n50, CK => CLK, RN => n2, Q => 
                           DOUT_17_port, QN => n_1250);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n51, CK => CLK, RN => n2, Q => 
                           DOUT_16_port, QN => n_1251);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n52, CK => CLK, RN => n2, Q => 
                           DOUT_15_port, QN => n_1252);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n53, CK => CLK, RN => n2, Q => 
                           DOUT_14_port, QN => n_1253);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n54, CK => CLK, RN => n2, Q => 
                           DOUT_13_port, QN => n_1254);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n55, CK => CLK, RN => n2, Q => 
                           DOUT_12_port, QN => n_1255);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n56, CK => CLK, RN => n1, Q => 
                           DOUT_11_port, QN => n_1256);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n57, CK => CLK, RN => n1, Q => 
                           DOUT_10_port, QN => n_1257);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n58, CK => CLK, RN => n1, Q => 
                           DOUT_9_port, QN => n_1258);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n59, CK => CLK, RN => n1, Q => 
                           DOUT_8_port, QN => n_1259);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n60, CK => CLK, RN => n1, Q => 
                           DOUT_7_port, QN => n_1260);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n61, CK => CLK, RN => n1, Q => 
                           DOUT_6_port, QN => n_1261);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n62, CK => CLK, RN => n1, Q => 
                           DOUT_5_port, QN => n_1262);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n63, CK => CLK, RN => n1, Q => 
                           DOUT_4_port, QN => n_1263);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n64, CK => CLK, RN => n1, Q => 
                           DOUT_3_port, QN => n_1264);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n68, CK => CLK, RN => n1, Q => 
                           DOUT_2_port, QN => n_1265);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n69, CK => CLK, RN => n1, Q => 
                           DOUT_1_port, QN => n_1266);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n70, CK => CLK, RN => n1, Q => 
                           DOUT_0_port, QN => n_1267);
   U2 : BUF_X1 port map( A => RST, Z => n1);
   U3 : BUF_X1 port map( A => RST, Z => n2);
   U4 : BUF_X1 port map( A => RST, Z => n3);
   U5 : MUX2_X1 port map( A => DOUT_0_port, B => DIN(0), S => EN, Z => n70);
   U6 : MUX2_X1 port map( A => DOUT_1_port, B => DIN(1), S => EN, Z => n69);
   U7 : MUX2_X1 port map( A => DOUT_2_port, B => DIN(2), S => EN, Z => n68);
   U8 : MUX2_X1 port map( A => DOUT_3_port, B => DIN(3), S => EN, Z => n64);
   U9 : MUX2_X1 port map( A => DOUT_4_port, B => DIN(4), S => EN, Z => n63);
   U10 : MUX2_X1 port map( A => DOUT_5_port, B => DIN(5), S => EN, Z => n62);
   U11 : MUX2_X1 port map( A => DOUT_6_port, B => DIN(6), S => EN, Z => n61);
   U12 : MUX2_X1 port map( A => DOUT_7_port, B => DIN(7), S => EN, Z => n60);
   U13 : MUX2_X1 port map( A => DOUT_8_port, B => DIN(8), S => EN, Z => n59);
   U14 : MUX2_X1 port map( A => DOUT_9_port, B => DIN(9), S => EN, Z => n58);
   U15 : MUX2_X1 port map( A => DOUT_10_port, B => DIN(10), S => EN, Z => n57);
   U16 : MUX2_X1 port map( A => DOUT_11_port, B => DIN(11), S => EN, Z => n56);
   U17 : MUX2_X1 port map( A => DOUT_12_port, B => DIN(12), S => EN, Z => n55);
   U18 : MUX2_X1 port map( A => DOUT_13_port, B => DIN(13), S => EN, Z => n54);
   U19 : MUX2_X1 port map( A => DOUT_14_port, B => DIN(14), S => EN, Z => n53);
   U20 : MUX2_X1 port map( A => DOUT_15_port, B => DIN(15), S => EN, Z => n52);
   U21 : MUX2_X1 port map( A => DOUT_16_port, B => DIN(16), S => EN, Z => n51);
   U22 : MUX2_X1 port map( A => DOUT_17_port, B => DIN(17), S => EN, Z => n50);
   U23 : MUX2_X1 port map( A => DOUT_18_port, B => DIN(18), S => EN, Z => n49);
   U24 : MUX2_X1 port map( A => DOUT_19_port, B => DIN(19), S => EN, Z => n48);
   U25 : MUX2_X1 port map( A => DOUT_20_port, B => DIN(20), S => EN, Z => n47);
   U26 : MUX2_X1 port map( A => DOUT_21_port, B => DIN(21), S => EN, Z => n46);
   U27 : MUX2_X1 port map( A => DOUT_22_port, B => DIN(22), S => EN, Z => n45);
   U28 : MUX2_X1 port map( A => DOUT_23_port, B => DIN(23), S => EN, Z => n44);
   U29 : MUX2_X1 port map( A => DOUT_24_port, B => DIN(24), S => EN, Z => n43);
   U30 : MUX2_X1 port map( A => DOUT_25_port, B => DIN(25), S => EN, Z => n42);
   U31 : MUX2_X1 port map( A => DOUT_26_port, B => DIN(26), S => EN, Z => n41);
   U32 : MUX2_X1 port map( A => DOUT_27_port, B => DIN(27), S => EN, Z => n40);
   U33 : MUX2_X1 port map( A => DOUT_28_port, B => DIN(28), S => EN, Z => n39);
   U34 : MUX2_X1 port map( A => DOUT_29_port, B => DIN(29), S => EN, Z => n38);
   U35 : MUX2_X1 port map( A => DOUT_30_port, B => DIN(30), S => EN, Z => n37);
   U36 : MUX2_X1 port map( A => DOUT_31_port, B => DIN(31), S => EN, Z => n36);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_5 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_5;

architecture SYN_bhv of regn_N32_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, DOUT_0_port, DOUT_1_port, DOUT_2_port, DOUT_3_port, 
      DOUT_4_port, DOUT_5_port, DOUT_6_port, DOUT_7_port, DOUT_8_port, 
      DOUT_9_port, DOUT_10_port, DOUT_11_port, DOUT_12_port, DOUT_13_port, 
      DOUT_14_port, DOUT_15_port, DOUT_16_port, DOUT_17_port, DOUT_18_port, 
      DOUT_19_port, DOUT_20_port, DOUT_21_port, DOUT_22_port, DOUT_23_port, 
      DOUT_24_port, DOUT_25_port, DOUT_26_port, DOUT_27_port, DOUT_28_port, 
      DOUT_29_port, DOUT_30_port, DOUT_31_port, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n68, n69, n70, n_1268, n_1269, 
      n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, 
      n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, 
      n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, 
      n_1297, n_1298, n_1299 : std_logic;

begin
   DOUT <= ( DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, 
      DOUT_27_port, DOUT_26_port, DOUT_25_port, DOUT_24_port, DOUT_23_port, 
      DOUT_22_port, DOUT_21_port, DOUT_20_port, DOUT_19_port, DOUT_18_port, 
      DOUT_17_port, DOUT_16_port, DOUT_15_port, DOUT_14_port, DOUT_13_port, 
      DOUT_12_port, DOUT_11_port, DOUT_10_port, DOUT_9_port, DOUT_8_port, 
      DOUT_7_port, DOUT_6_port, DOUT_5_port, DOUT_4_port, DOUT_3_port, 
      DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n36, CK => CLK, RN => n3, Q => 
                           DOUT_31_port, QN => n_1268);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n37, CK => CLK, RN => n3, Q => 
                           DOUT_30_port, QN => n_1269);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n38, CK => CLK, RN => n3, Q => 
                           DOUT_29_port, QN => n_1270);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n39, CK => CLK, RN => n3, Q => 
                           DOUT_28_port, QN => n_1271);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n40, CK => CLK, RN => n3, Q => 
                           DOUT_27_port, QN => n_1272);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n41, CK => CLK, RN => n3, Q => 
                           DOUT_26_port, QN => n_1273);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n42, CK => CLK, RN => n3, Q => 
                           DOUT_25_port, QN => n_1274);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n43, CK => CLK, RN => n3, Q => 
                           DOUT_24_port, QN => n_1275);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n44, CK => CLK, RN => n2, Q => 
                           DOUT_23_port, QN => n_1276);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n45, CK => CLK, RN => n2, Q => 
                           DOUT_22_port, QN => n_1277);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n46, CK => CLK, RN => n2, Q => 
                           DOUT_21_port, QN => n_1278);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n47, CK => CLK, RN => n2, Q => 
                           DOUT_20_port, QN => n_1279);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n48, CK => CLK, RN => n2, Q => 
                           DOUT_19_port, QN => n_1280);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n49, CK => CLK, RN => n2, Q => 
                           DOUT_18_port, QN => n_1281);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n50, CK => CLK, RN => n2, Q => 
                           DOUT_17_port, QN => n_1282);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n51, CK => CLK, RN => n2, Q => 
                           DOUT_16_port, QN => n_1283);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n52, CK => CLK, RN => n2, Q => 
                           DOUT_15_port, QN => n_1284);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n53, CK => CLK, RN => n2, Q => 
                           DOUT_14_port, QN => n_1285);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n54, CK => CLK, RN => n2, Q => 
                           DOUT_13_port, QN => n_1286);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n55, CK => CLK, RN => n2, Q => 
                           DOUT_12_port, QN => n_1287);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n56, CK => CLK, RN => n1, Q => 
                           DOUT_11_port, QN => n_1288);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n57, CK => CLK, RN => n1, Q => 
                           DOUT_10_port, QN => n_1289);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n58, CK => CLK, RN => n1, Q => 
                           DOUT_9_port, QN => n_1290);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n59, CK => CLK, RN => n1, Q => 
                           DOUT_8_port, QN => n_1291);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n60, CK => CLK, RN => n1, Q => 
                           DOUT_7_port, QN => n_1292);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n61, CK => CLK, RN => n1, Q => 
                           DOUT_6_port, QN => n_1293);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n62, CK => CLK, RN => n1, Q => 
                           DOUT_5_port, QN => n_1294);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n63, CK => CLK, RN => n1, Q => 
                           DOUT_4_port, QN => n_1295);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n64, CK => CLK, RN => n1, Q => 
                           DOUT_3_port, QN => n_1296);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n68, CK => CLK, RN => n1, Q => 
                           DOUT_2_port, QN => n_1297);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n69, CK => CLK, RN => n1, Q => 
                           DOUT_1_port, QN => n_1298);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n70, CK => CLK, RN => n1, Q => 
                           DOUT_0_port, QN => n_1299);
   U2 : BUF_X1 port map( A => RST, Z => n1);
   U3 : BUF_X1 port map( A => RST, Z => n2);
   U4 : BUF_X1 port map( A => RST, Z => n3);
   U5 : MUX2_X1 port map( A => DOUT_0_port, B => DIN(0), S => EN, Z => n70);
   U6 : MUX2_X1 port map( A => DOUT_1_port, B => DIN(1), S => EN, Z => n69);
   U7 : MUX2_X1 port map( A => DOUT_2_port, B => DIN(2), S => EN, Z => n68);
   U8 : MUX2_X1 port map( A => DOUT_3_port, B => DIN(3), S => EN, Z => n64);
   U9 : MUX2_X1 port map( A => DOUT_4_port, B => DIN(4), S => EN, Z => n63);
   U10 : MUX2_X1 port map( A => DOUT_5_port, B => DIN(5), S => EN, Z => n62);
   U11 : MUX2_X1 port map( A => DOUT_6_port, B => DIN(6), S => EN, Z => n61);
   U12 : MUX2_X1 port map( A => DOUT_7_port, B => DIN(7), S => EN, Z => n60);
   U13 : MUX2_X1 port map( A => DOUT_8_port, B => DIN(8), S => EN, Z => n59);
   U14 : MUX2_X1 port map( A => DOUT_9_port, B => DIN(9), S => EN, Z => n58);
   U15 : MUX2_X1 port map( A => DOUT_10_port, B => DIN(10), S => EN, Z => n57);
   U16 : MUX2_X1 port map( A => DOUT_11_port, B => DIN(11), S => EN, Z => n56);
   U17 : MUX2_X1 port map( A => DOUT_12_port, B => DIN(12), S => EN, Z => n55);
   U18 : MUX2_X1 port map( A => DOUT_13_port, B => DIN(13), S => EN, Z => n54);
   U19 : MUX2_X1 port map( A => DOUT_14_port, B => DIN(14), S => EN, Z => n53);
   U20 : MUX2_X1 port map( A => DOUT_15_port, B => DIN(15), S => EN, Z => n52);
   U21 : MUX2_X1 port map( A => DOUT_16_port, B => DIN(16), S => EN, Z => n51);
   U22 : MUX2_X1 port map( A => DOUT_17_port, B => DIN(17), S => EN, Z => n50);
   U23 : MUX2_X1 port map( A => DOUT_18_port, B => DIN(18), S => EN, Z => n49);
   U24 : MUX2_X1 port map( A => DOUT_19_port, B => DIN(19), S => EN, Z => n48);
   U25 : MUX2_X1 port map( A => DOUT_20_port, B => DIN(20), S => EN, Z => n47);
   U26 : MUX2_X1 port map( A => DOUT_21_port, B => DIN(21), S => EN, Z => n46);
   U27 : MUX2_X1 port map( A => DOUT_22_port, B => DIN(22), S => EN, Z => n45);
   U28 : MUX2_X1 port map( A => DOUT_23_port, B => DIN(23), S => EN, Z => n44);
   U29 : MUX2_X1 port map( A => DOUT_24_port, B => DIN(24), S => EN, Z => n43);
   U30 : MUX2_X1 port map( A => DOUT_25_port, B => DIN(25), S => EN, Z => n42);
   U31 : MUX2_X1 port map( A => DOUT_26_port, B => DIN(26), S => EN, Z => n41);
   U32 : MUX2_X1 port map( A => DOUT_27_port, B => DIN(27), S => EN, Z => n40);
   U33 : MUX2_X1 port map( A => DOUT_28_port, B => DIN(28), S => EN, Z => n39);
   U34 : MUX2_X1 port map( A => DOUT_29_port, B => DIN(29), S => EN, Z => n38);
   U35 : MUX2_X1 port map( A => DOUT_30_port, B => DIN(30), S => EN, Z => n37);
   U36 : MUX2_X1 port map( A => DOUT_31_port, B => DIN(31), S => EN, Z => n36);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_4 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_4;

architecture SYN_bhv of regn_N32_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, DOUT_27_port,
      DOUT_26_port, DOUT_25_port, DOUT_24_port, DOUT_22_port, DOUT_21_port, 
      DOUT_20_port, DOUT_19_port, DOUT_18_port, DOUT_16_port, DOUT_15_port, 
      DOUT_14_port, DOUT_13_port, DOUT_12_port, DOUT_11_port, DOUT_10_port, 
      DOUT_8_port, DOUT_7_port, DOUT_6_port, DOUT_5_port, DOUT_4_port, 
      DOUT_3_port, DOUT_2_port, n1, n2, n3, DOUT_0_port, DOUT_1_port, n6, n7, 
      n8, n9, n10, n11, n12, DOUT_9_port, n14, n15, n16, n17, n18, n19, n20, 
      DOUT_17_port, n22, n23, n24, n25, n26, DOUT_23_port, n28, n29, n30, n31, 
      n32, n33, n34, n42, n50, n56, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n_1300, n_1301, n_1302, n_1303, n_1304 : std_logic;

begin
   DOUT <= ( DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, 
      DOUT_27_port, DOUT_26_port, DOUT_25_port, DOUT_24_port, DOUT_23_port, 
      DOUT_22_port, DOUT_21_port, DOUT_20_port, DOUT_19_port, DOUT_18_port, 
      DOUT_17_port, DOUT_16_port, DOUT_15_port, DOUT_14_port, DOUT_13_port, 
      DOUT_12_port, DOUT_11_port, DOUT_10_port, DOUT_9_port, DOUT_8_port, 
      DOUT_7_port, DOUT_6_port, DOUT_5_port, DOUT_4_port, DOUT_3_port, 
      DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n50, CK => CLK, RN => n3, Q => 
                           DOUT_31_port, QN => n125);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n56, CK => CLK, RN => n3, Q => 
                           DOUT_30_port, QN => n126);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n95, CK => CLK, RN => n3, Q => 
                           DOUT_29_port, QN => n127);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n96, CK => CLK, RN => n3, Q => 
                           DOUT_28_port, QN => n128);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n97, CK => CLK, RN => n3, Q => 
                           DOUT_27_port, QN => n129);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n98, CK => CLK, RN => n3, Q => 
                           DOUT_26_port, QN => n130);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n99, CK => CLK, RN => n3, Q => 
                           DOUT_25_port, QN => n131);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n3, Q => 
                           DOUT_24_port, QN => n132);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n2, Q => 
                           DOUT_23_port, QN => n_1300);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n2, Q => 
                           DOUT_22_port, QN => n133);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n2, Q => 
                           DOUT_21_port, QN => n134);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n2, Q => 
                           DOUT_20_port, QN => n135);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n2, Q => 
                           DOUT_19_port, QN => n136);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n2, Q => 
                           DOUT_18_port, QN => n137);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n2, Q => 
                           DOUT_17_port, QN => n_1301);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n2, Q => 
                           DOUT_16_port, QN => n138);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n2, Q => 
                           DOUT_15_port, QN => n139);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n2, Q => 
                           DOUT_14_port, QN => n140);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n2, Q => 
                           DOUT_13_port, QN => n141);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n2, Q => 
                           DOUT_12_port, QN => n142);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n1, Q => 
                           DOUT_11_port, QN => n143);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n1, Q => 
                           DOUT_10_port, QN => n144);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n1, Q => 
                           DOUT_9_port, QN => n_1302);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n1, Q => 
                           DOUT_8_port, QN => n145);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n1, Q => 
                           DOUT_7_port, QN => n146);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n1, Q => 
                           DOUT_6_port, QN => n147);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n1, Q => 
                           DOUT_5_port, QN => n148);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n1, Q => 
                           DOUT_4_port, QN => n149);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n1, Q => 
                           DOUT_3_port, QN => n150);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n1, Q => 
                           DOUT_2_port, QN => n151);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n1, Q => 
                           DOUT_1_port, QN => n_1303);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n1, Q => 
                           DOUT_0_port, QN => n_1304);
   U2 : BUF_X1 port map( A => RST, Z => n1);
   U3 : BUF_X1 port map( A => RST, Z => n2);
   U4 : BUF_X1 port map( A => RST, Z => n3);
   U5 : MUX2_X1 port map( A => DOUT_0_port, B => DIN(0), S => EN, Z => n124);
   U6 : MUX2_X1 port map( A => DOUT_1_port, B => DIN(1), S => EN, Z => n123);
   U7 : INV_X1 port map( A => n151, ZN => n6);
   U8 : MUX2_X1 port map( A => n6, B => DIN(2), S => EN, Z => n122);
   U9 : INV_X1 port map( A => n150, ZN => n7);
   U10 : MUX2_X1 port map( A => n7, B => DIN(3), S => EN, Z => n121);
   U11 : INV_X1 port map( A => n149, ZN => n8);
   U12 : MUX2_X1 port map( A => n8, B => DIN(4), S => EN, Z => n120);
   U13 : INV_X1 port map( A => n148, ZN => n9);
   U14 : MUX2_X1 port map( A => n9, B => DIN(5), S => EN, Z => n119);
   U15 : INV_X1 port map( A => n147, ZN => n10);
   U16 : MUX2_X1 port map( A => n10, B => DIN(6), S => EN, Z => n118);
   U17 : INV_X1 port map( A => n146, ZN => n11);
   U18 : MUX2_X1 port map( A => n11, B => DIN(7), S => EN, Z => n117);
   U19 : INV_X1 port map( A => n145, ZN => n12);
   U20 : MUX2_X1 port map( A => n12, B => DIN(8), S => EN, Z => n116);
   U21 : MUX2_X1 port map( A => DOUT_9_port, B => DIN(9), S => EN, Z => n115);
   U22 : INV_X1 port map( A => n144, ZN => n14);
   U23 : MUX2_X1 port map( A => n14, B => DIN(10), S => EN, Z => n114);
   U24 : INV_X1 port map( A => n143, ZN => n15);
   U25 : MUX2_X1 port map( A => n15, B => DIN(11), S => EN, Z => n113);
   U26 : INV_X1 port map( A => n142, ZN => n16);
   U27 : MUX2_X1 port map( A => n16, B => DIN(12), S => EN, Z => n112);
   U28 : INV_X1 port map( A => n141, ZN => n17);
   U29 : MUX2_X1 port map( A => n17, B => DIN(13), S => EN, Z => n111);
   U30 : INV_X1 port map( A => n140, ZN => n18);
   U31 : MUX2_X1 port map( A => n18, B => DIN(14), S => EN, Z => n110);
   U32 : INV_X1 port map( A => n139, ZN => n19);
   U33 : MUX2_X1 port map( A => n19, B => DIN(15), S => EN, Z => n109);
   U34 : INV_X1 port map( A => n138, ZN => n20);
   U35 : MUX2_X1 port map( A => n20, B => DIN(16), S => EN, Z => n108);
   U36 : MUX2_X1 port map( A => DOUT_17_port, B => DIN(17), S => EN, Z => n107)
                           ;
   U37 : INV_X1 port map( A => n137, ZN => n22);
   U38 : MUX2_X1 port map( A => n22, B => DIN(18), S => EN, Z => n106);
   U39 : INV_X1 port map( A => n136, ZN => n23);
   U40 : MUX2_X1 port map( A => n23, B => DIN(19), S => EN, Z => n105);
   U41 : INV_X1 port map( A => n135, ZN => n24);
   U42 : MUX2_X1 port map( A => n24, B => DIN(20), S => EN, Z => n104);
   U43 : INV_X1 port map( A => n134, ZN => n25);
   U44 : MUX2_X1 port map( A => n25, B => DIN(21), S => EN, Z => n103);
   U45 : INV_X1 port map( A => n133, ZN => n26);
   U46 : MUX2_X1 port map( A => n26, B => DIN(22), S => EN, Z => n102);
   U47 : MUX2_X1 port map( A => DOUT_23_port, B => DIN(23), S => EN, Z => n101)
                           ;
   U48 : INV_X1 port map( A => n132, ZN => n28);
   U49 : MUX2_X1 port map( A => n28, B => DIN(24), S => EN, Z => n100);
   U50 : INV_X1 port map( A => n131, ZN => n29);
   U51 : MUX2_X1 port map( A => n29, B => DIN(25), S => EN, Z => n99);
   U52 : INV_X1 port map( A => n130, ZN => n30);
   U53 : MUX2_X1 port map( A => n30, B => DIN(26), S => EN, Z => n98);
   U54 : INV_X1 port map( A => n129, ZN => n31);
   U55 : MUX2_X1 port map( A => n31, B => DIN(27), S => EN, Z => n97);
   U56 : INV_X1 port map( A => n128, ZN => n32);
   U57 : MUX2_X1 port map( A => n32, B => DIN(28), S => EN, Z => n96);
   U58 : INV_X1 port map( A => n127, ZN => n33);
   U59 : MUX2_X1 port map( A => n33, B => DIN(29), S => EN, Z => n95);
   U60 : INV_X1 port map( A => n126, ZN => n34);
   U61 : MUX2_X1 port map( A => n34, B => DIN(30), S => EN, Z => n56);
   U62 : INV_X1 port map( A => n125, ZN => n42);
   U63 : MUX2_X1 port map( A => n42, B => DIN(31), S => EN, Z => n50);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_3 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_3;

architecture SYN_bhv of regn_N32_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n3, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n3, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n3, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n3, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n3, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n3, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n3, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n3, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n2, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n2, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n2, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n2, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n2, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n2, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n2, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n2, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n2, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n2, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n2, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n2, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n1, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n1, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n1, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n1, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n1, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n1, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n1, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n1, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n1, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n1, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n1, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n1, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n1);
   U3 : BUF_X1 port map( A => RST, Z => n2);
   U4 : BUF_X1 port map( A => RST, Z => n3);
   U5 : INV_X1 port map( A => n163, ZN => n4);
   U6 : MUX2_X1 port map( A => n4, B => DIN(0), S => EN, Z => n131);
   U7 : INV_X1 port map( A => n162, ZN => n5);
   U8 : MUX2_X1 port map( A => n5, B => DIN(1), S => EN, Z => n130);
   U9 : INV_X1 port map( A => n161, ZN => n6);
   U10 : MUX2_X1 port map( A => n6, B => DIN(2), S => EN, Z => n129);
   U11 : INV_X1 port map( A => n160, ZN => n7);
   U12 : MUX2_X1 port map( A => n7, B => DIN(3), S => EN, Z => n128);
   U13 : INV_X1 port map( A => n159, ZN => n8);
   U14 : MUX2_X1 port map( A => n8, B => DIN(4), S => EN, Z => n127);
   U15 : INV_X1 port map( A => n158, ZN => n9);
   U16 : MUX2_X1 port map( A => n9, B => DIN(5), S => EN, Z => n126);
   U17 : INV_X1 port map( A => n157, ZN => n10);
   U18 : MUX2_X1 port map( A => n10, B => DIN(6), S => EN, Z => n125);
   U19 : INV_X1 port map( A => n156, ZN => n11);
   U20 : MUX2_X1 port map( A => n11, B => DIN(7), S => EN, Z => n124);
   U21 : INV_X1 port map( A => n155, ZN => n12);
   U22 : MUX2_X1 port map( A => n12, B => DIN(8), S => EN, Z => n123);
   U23 : INV_X1 port map( A => n154, ZN => n13);
   U24 : MUX2_X1 port map( A => n13, B => DIN(9), S => EN, Z => n122);
   U25 : INV_X1 port map( A => n153, ZN => n14);
   U26 : MUX2_X1 port map( A => n14, B => DIN(10), S => EN, Z => n121);
   U27 : INV_X1 port map( A => n152, ZN => n15);
   U28 : MUX2_X1 port map( A => n15, B => DIN(11), S => EN, Z => n120);
   U29 : INV_X1 port map( A => n151, ZN => n16);
   U30 : MUX2_X1 port map( A => n16, B => DIN(12), S => EN, Z => n119);
   U31 : INV_X1 port map( A => n150, ZN => n17);
   U32 : MUX2_X1 port map( A => n17, B => DIN(13), S => EN, Z => n118);
   U33 : INV_X1 port map( A => n149, ZN => n18);
   U34 : MUX2_X1 port map( A => n18, B => DIN(14), S => EN, Z => n117);
   U35 : INV_X1 port map( A => n148, ZN => n19);
   U36 : MUX2_X1 port map( A => n19, B => DIN(15), S => EN, Z => n116);
   U37 : INV_X1 port map( A => n147, ZN => n20);
   U38 : MUX2_X1 port map( A => n20, B => DIN(16), S => EN, Z => n115);
   U39 : INV_X1 port map( A => n146, ZN => n21);
   U40 : MUX2_X1 port map( A => n21, B => DIN(17), S => EN, Z => n114);
   U41 : INV_X1 port map( A => n145, ZN => n22);
   U42 : MUX2_X1 port map( A => n22, B => DIN(18), S => EN, Z => n113);
   U43 : INV_X1 port map( A => n144, ZN => n23);
   U44 : MUX2_X1 port map( A => n23, B => DIN(19), S => EN, Z => n112);
   U45 : INV_X1 port map( A => n143, ZN => n24);
   U46 : MUX2_X1 port map( A => n24, B => DIN(20), S => EN, Z => n111);
   U47 : INV_X1 port map( A => n142, ZN => n25);
   U48 : MUX2_X1 port map( A => n25, B => DIN(21), S => EN, Z => n110);
   U49 : INV_X1 port map( A => n141, ZN => n26);
   U50 : MUX2_X1 port map( A => n26, B => DIN(22), S => EN, Z => n109);
   U51 : INV_X1 port map( A => n140, ZN => n27);
   U52 : MUX2_X1 port map( A => n27, B => DIN(23), S => EN, Z => n108);
   U53 : INV_X1 port map( A => n139, ZN => n28);
   U54 : MUX2_X1 port map( A => n28, B => DIN(24), S => EN, Z => n107);
   U55 : INV_X1 port map( A => n138, ZN => n29);
   U56 : MUX2_X1 port map( A => n29, B => DIN(25), S => EN, Z => n106);
   U57 : INV_X1 port map( A => n137, ZN => n30);
   U58 : MUX2_X1 port map( A => n30, B => DIN(26), S => EN, Z => n105);
   U59 : INV_X1 port map( A => n136, ZN => n31);
   U60 : MUX2_X1 port map( A => n31, B => DIN(27), S => EN, Z => n104);
   U61 : INV_X1 port map( A => n135, ZN => n32);
   U62 : MUX2_X1 port map( A => n32, B => DIN(28), S => EN, Z => n103);
   U63 : INV_X1 port map( A => n134, ZN => n97);
   U64 : MUX2_X1 port map( A => n97, B => DIN(29), S => EN, Z => n102);
   U65 : INV_X1 port map( A => n133, ZN => n98);
   U66 : MUX2_X1 port map( A => n98, B => DIN(30), S => EN, Z => n101);
   U67 : INV_X1 port map( A => n132, ZN => n99);
   U68 : MUX2_X1 port map( A => n99, B => DIN(31), S => EN, Z => n100);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_2 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_2;

architecture SYN_bhv of regn_N32_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, DOUT_0_port, DOUT_1_port, DOUT_2_port, DOUT_3_port, 
      DOUT_4_port, DOUT_5_port, DOUT_6_port, DOUT_7_port, DOUT_8_port, 
      DOUT_9_port, DOUT_10_port, DOUT_11_port, DOUT_12_port, DOUT_13_port, 
      DOUT_14_port, DOUT_15_port, DOUT_16_port, DOUT_17_port, DOUT_18_port, 
      DOUT_19_port, DOUT_20_port, DOUT_21_port, DOUT_22_port, DOUT_23_port, 
      DOUT_24_port, DOUT_25_port, DOUT_26_port, DOUT_27_port, DOUT_28_port, 
      DOUT_29_port, DOUT_30_port, DOUT_31_port, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n68, n69, n70, n_1305, n_1306, 
      n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, 
      n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, 
      n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, 
      n_1334, n_1335, n_1336 : std_logic;

begin
   DOUT <= ( DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, 
      DOUT_27_port, DOUT_26_port, DOUT_25_port, DOUT_24_port, DOUT_23_port, 
      DOUT_22_port, DOUT_21_port, DOUT_20_port, DOUT_19_port, DOUT_18_port, 
      DOUT_17_port, DOUT_16_port, DOUT_15_port, DOUT_14_port, DOUT_13_port, 
      DOUT_12_port, DOUT_11_port, DOUT_10_port, DOUT_9_port, DOUT_8_port, 
      DOUT_7_port, DOUT_6_port, DOUT_5_port, DOUT_4_port, DOUT_3_port, 
      DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n36, CK => CLK, RN => n3, Q => 
                           DOUT_31_port, QN => n_1305);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n37, CK => CLK, RN => n3, Q => 
                           DOUT_30_port, QN => n_1306);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n38, CK => CLK, RN => n3, Q => 
                           DOUT_29_port, QN => n_1307);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n39, CK => CLK, RN => n3, Q => 
                           DOUT_28_port, QN => n_1308);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n40, CK => CLK, RN => n3, Q => 
                           DOUT_27_port, QN => n_1309);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n41, CK => CLK, RN => n3, Q => 
                           DOUT_26_port, QN => n_1310);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n42, CK => CLK, RN => n3, Q => 
                           DOUT_25_port, QN => n_1311);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n43, CK => CLK, RN => n3, Q => 
                           DOUT_24_port, QN => n_1312);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n44, CK => CLK, RN => n2, Q => 
                           DOUT_23_port, QN => n_1313);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n45, CK => CLK, RN => n2, Q => 
                           DOUT_22_port, QN => n_1314);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n46, CK => CLK, RN => n2, Q => 
                           DOUT_21_port, QN => n_1315);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n47, CK => CLK, RN => n2, Q => 
                           DOUT_20_port, QN => n_1316);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n48, CK => CLK, RN => n2, Q => 
                           DOUT_19_port, QN => n_1317);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n49, CK => CLK, RN => n2, Q => 
                           DOUT_18_port, QN => n_1318);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n50, CK => CLK, RN => n2, Q => 
                           DOUT_17_port, QN => n_1319);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n51, CK => CLK, RN => n2, Q => 
                           DOUT_16_port, QN => n_1320);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n52, CK => CLK, RN => n2, Q => 
                           DOUT_15_port, QN => n_1321);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n53, CK => CLK, RN => n2, Q => 
                           DOUT_14_port, QN => n_1322);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n54, CK => CLK, RN => n2, Q => 
                           DOUT_13_port, QN => n_1323);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n55, CK => CLK, RN => n2, Q => 
                           DOUT_12_port, QN => n_1324);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n56, CK => CLK, RN => n1, Q => 
                           DOUT_11_port, QN => n_1325);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n57, CK => CLK, RN => n1, Q => 
                           DOUT_10_port, QN => n_1326);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n58, CK => CLK, RN => n1, Q => 
                           DOUT_9_port, QN => n_1327);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n59, CK => CLK, RN => n1, Q => 
                           DOUT_8_port, QN => n_1328);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n60, CK => CLK, RN => n1, Q => 
                           DOUT_7_port, QN => n_1329);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n61, CK => CLK, RN => n1, Q => 
                           DOUT_6_port, QN => n_1330);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n62, CK => CLK, RN => n1, Q => 
                           DOUT_5_port, QN => n_1331);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n63, CK => CLK, RN => n1, Q => 
                           DOUT_4_port, QN => n_1332);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n64, CK => CLK, RN => n1, Q => 
                           DOUT_3_port, QN => n_1333);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n68, CK => CLK, RN => n1, Q => 
                           DOUT_2_port, QN => n_1334);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n69, CK => CLK, RN => n1, Q => 
                           DOUT_1_port, QN => n_1335);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n70, CK => CLK, RN => n1, Q => 
                           DOUT_0_port, QN => n_1336);
   U2 : BUF_X1 port map( A => RST, Z => n1);
   U3 : BUF_X1 port map( A => RST, Z => n2);
   U4 : BUF_X1 port map( A => RST, Z => n3);
   U5 : MUX2_X1 port map( A => DOUT_0_port, B => DIN(0), S => EN, Z => n70);
   U6 : MUX2_X1 port map( A => DOUT_1_port, B => DIN(1), S => EN, Z => n69);
   U7 : MUX2_X1 port map( A => DOUT_2_port, B => DIN(2), S => EN, Z => n68);
   U8 : MUX2_X1 port map( A => DOUT_3_port, B => DIN(3), S => EN, Z => n64);
   U9 : MUX2_X1 port map( A => DOUT_4_port, B => DIN(4), S => EN, Z => n63);
   U10 : MUX2_X1 port map( A => DOUT_5_port, B => DIN(5), S => EN, Z => n62);
   U11 : MUX2_X1 port map( A => DOUT_6_port, B => DIN(6), S => EN, Z => n61);
   U12 : MUX2_X1 port map( A => DOUT_7_port, B => DIN(7), S => EN, Z => n60);
   U13 : MUX2_X1 port map( A => DOUT_8_port, B => DIN(8), S => EN, Z => n59);
   U14 : MUX2_X1 port map( A => DOUT_9_port, B => DIN(9), S => EN, Z => n58);
   U15 : MUX2_X1 port map( A => DOUT_10_port, B => DIN(10), S => EN, Z => n57);
   U16 : MUX2_X1 port map( A => DOUT_11_port, B => DIN(11), S => EN, Z => n56);
   U17 : MUX2_X1 port map( A => DOUT_12_port, B => DIN(12), S => EN, Z => n55);
   U18 : MUX2_X1 port map( A => DOUT_13_port, B => DIN(13), S => EN, Z => n54);
   U19 : MUX2_X1 port map( A => DOUT_14_port, B => DIN(14), S => EN, Z => n53);
   U20 : MUX2_X1 port map( A => DOUT_15_port, B => DIN(15), S => EN, Z => n52);
   U21 : MUX2_X1 port map( A => DOUT_16_port, B => DIN(16), S => EN, Z => n51);
   U22 : MUX2_X1 port map( A => DOUT_17_port, B => DIN(17), S => EN, Z => n50);
   U23 : MUX2_X1 port map( A => DOUT_18_port, B => DIN(18), S => EN, Z => n49);
   U24 : MUX2_X1 port map( A => DOUT_19_port, B => DIN(19), S => EN, Z => n48);
   U25 : MUX2_X1 port map( A => DOUT_20_port, B => DIN(20), S => EN, Z => n47);
   U26 : MUX2_X1 port map( A => DOUT_21_port, B => DIN(21), S => EN, Z => n46);
   U27 : MUX2_X1 port map( A => DOUT_22_port, B => DIN(22), S => EN, Z => n45);
   U28 : MUX2_X1 port map( A => DOUT_23_port, B => DIN(23), S => EN, Z => n44);
   U29 : MUX2_X1 port map( A => DOUT_24_port, B => DIN(24), S => EN, Z => n43);
   U30 : MUX2_X1 port map( A => DOUT_25_port, B => DIN(25), S => EN, Z => n42);
   U31 : MUX2_X1 port map( A => DOUT_26_port, B => DIN(26), S => EN, Z => n41);
   U32 : MUX2_X1 port map( A => DOUT_27_port, B => DIN(27), S => EN, Z => n40);
   U33 : MUX2_X1 port map( A => DOUT_28_port, B => DIN(28), S => EN, Z => n39);
   U34 : MUX2_X1 port map( A => DOUT_29_port, B => DIN(29), S => EN, Z => n38);
   U35 : MUX2_X1 port map( A => DOUT_30_port, B => DIN(30), S => EN, Z => n37);
   U36 : MUX2_X1 port map( A => DOUT_31_port, B => DIN(31), S => EN, Z => n36);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_1 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_1;

architecture SYN_bhv of regn_N32_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, DOUT_0_port, DOUT_1_port, DOUT_2_port, DOUT_3_port, 
      DOUT_4_port, DOUT_5_port, DOUT_6_port, DOUT_7_port, DOUT_8_port, 
      DOUT_9_port, DOUT_10_port, DOUT_11_port, DOUT_12_port, DOUT_13_port, 
      DOUT_14_port, DOUT_15_port, DOUT_16_port, DOUT_17_port, DOUT_18_port, 
      DOUT_19_port, DOUT_20_port, DOUT_21_port, DOUT_22_port, DOUT_23_port, 
      DOUT_24_port, DOUT_25_port, DOUT_26_port, DOUT_27_port, DOUT_28_port, 
      DOUT_29_port, DOUT_30_port, DOUT_31_port, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n68, n69, n70, n_1337, n_1338, 
      n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, 
      n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, 
      n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, 
      n_1366, n_1367, n_1368 : std_logic;

begin
   DOUT <= ( DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, 
      DOUT_27_port, DOUT_26_port, DOUT_25_port, DOUT_24_port, DOUT_23_port, 
      DOUT_22_port, DOUT_21_port, DOUT_20_port, DOUT_19_port, DOUT_18_port, 
      DOUT_17_port, DOUT_16_port, DOUT_15_port, DOUT_14_port, DOUT_13_port, 
      DOUT_12_port, DOUT_11_port, DOUT_10_port, DOUT_9_port, DOUT_8_port, 
      DOUT_7_port, DOUT_6_port, DOUT_5_port, DOUT_4_port, DOUT_3_port, 
      DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n36, CK => CLK, RN => n3, Q => 
                           DOUT_31_port, QN => n_1337);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n37, CK => CLK, RN => n3, Q => 
                           DOUT_30_port, QN => n_1338);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n38, CK => CLK, RN => n3, Q => 
                           DOUT_29_port, QN => n_1339);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n39, CK => CLK, RN => n3, Q => 
                           DOUT_28_port, QN => n_1340);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n40, CK => CLK, RN => n3, Q => 
                           DOUT_27_port, QN => n_1341);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n41, CK => CLK, RN => n3, Q => 
                           DOUT_26_port, QN => n_1342);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n42, CK => CLK, RN => n3, Q => 
                           DOUT_25_port, QN => n_1343);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n43, CK => CLK, RN => n3, Q => 
                           DOUT_24_port, QN => n_1344);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n44, CK => CLK, RN => n2, Q => 
                           DOUT_23_port, QN => n_1345);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n45, CK => CLK, RN => n2, Q => 
                           DOUT_22_port, QN => n_1346);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n46, CK => CLK, RN => n2, Q => 
                           DOUT_21_port, QN => n_1347);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n47, CK => CLK, RN => n2, Q => 
                           DOUT_20_port, QN => n_1348);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n48, CK => CLK, RN => n2, Q => 
                           DOUT_19_port, QN => n_1349);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n49, CK => CLK, RN => n2, Q => 
                           DOUT_18_port, QN => n_1350);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n50, CK => CLK, RN => n2, Q => 
                           DOUT_17_port, QN => n_1351);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n51, CK => CLK, RN => n2, Q => 
                           DOUT_16_port, QN => n_1352);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n52, CK => CLK, RN => n2, Q => 
                           DOUT_15_port, QN => n_1353);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n53, CK => CLK, RN => n2, Q => 
                           DOUT_14_port, QN => n_1354);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n54, CK => CLK, RN => n2, Q => 
                           DOUT_13_port, QN => n_1355);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n55, CK => CLK, RN => n2, Q => 
                           DOUT_12_port, QN => n_1356);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n56, CK => CLK, RN => n1, Q => 
                           DOUT_11_port, QN => n_1357);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n57, CK => CLK, RN => n1, Q => 
                           DOUT_10_port, QN => n_1358);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n58, CK => CLK, RN => n1, Q => 
                           DOUT_9_port, QN => n_1359);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n59, CK => CLK, RN => n1, Q => 
                           DOUT_8_port, QN => n_1360);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n60, CK => CLK, RN => n1, Q => 
                           DOUT_7_port, QN => n_1361);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n61, CK => CLK, RN => n1, Q => 
                           DOUT_6_port, QN => n_1362);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n62, CK => CLK, RN => n1, Q => 
                           DOUT_5_port, QN => n_1363);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n63, CK => CLK, RN => n1, Q => 
                           DOUT_4_port, QN => n_1364);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n64, CK => CLK, RN => n1, Q => 
                           DOUT_3_port, QN => n_1365);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n68, CK => CLK, RN => n1, Q => 
                           DOUT_2_port, QN => n_1366);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n69, CK => CLK, RN => n1, Q => 
                           DOUT_1_port, QN => n_1367);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n70, CK => CLK, RN => n1, Q => 
                           DOUT_0_port, QN => n_1368);
   U2 : BUF_X1 port map( A => RST, Z => n1);
   U3 : BUF_X1 port map( A => RST, Z => n2);
   U4 : BUF_X1 port map( A => RST, Z => n3);
   U5 : MUX2_X1 port map( A => DOUT_0_port, B => DIN(0), S => EN, Z => n70);
   U6 : MUX2_X1 port map( A => DOUT_1_port, B => DIN(1), S => EN, Z => n69);
   U7 : MUX2_X1 port map( A => DOUT_2_port, B => DIN(2), S => EN, Z => n68);
   U8 : MUX2_X1 port map( A => DOUT_3_port, B => DIN(3), S => EN, Z => n64);
   U9 : MUX2_X1 port map( A => DOUT_4_port, B => DIN(4), S => EN, Z => n63);
   U10 : MUX2_X1 port map( A => DOUT_5_port, B => DIN(5), S => EN, Z => n62);
   U11 : MUX2_X1 port map( A => DOUT_6_port, B => DIN(6), S => EN, Z => n61);
   U12 : MUX2_X1 port map( A => DOUT_7_port, B => DIN(7), S => EN, Z => n60);
   U13 : MUX2_X1 port map( A => DOUT_8_port, B => DIN(8), S => EN, Z => n59);
   U14 : MUX2_X1 port map( A => DOUT_9_port, B => DIN(9), S => EN, Z => n58);
   U15 : MUX2_X1 port map( A => DOUT_10_port, B => DIN(10), S => EN, Z => n57);
   U16 : MUX2_X1 port map( A => DOUT_11_port, B => DIN(11), S => EN, Z => n56);
   U17 : MUX2_X1 port map( A => DOUT_12_port, B => DIN(12), S => EN, Z => n55);
   U18 : MUX2_X1 port map( A => DOUT_13_port, B => DIN(13), S => EN, Z => n54);
   U19 : MUX2_X1 port map( A => DOUT_14_port, B => DIN(14), S => EN, Z => n53);
   U20 : MUX2_X1 port map( A => DOUT_15_port, B => DIN(15), S => EN, Z => n52);
   U21 : MUX2_X1 port map( A => DOUT_16_port, B => DIN(16), S => EN, Z => n51);
   U22 : MUX2_X1 port map( A => DOUT_17_port, B => DIN(17), S => EN, Z => n50);
   U23 : MUX2_X1 port map( A => DOUT_18_port, B => DIN(18), S => EN, Z => n49);
   U24 : MUX2_X1 port map( A => DOUT_19_port, B => DIN(19), S => EN, Z => n48);
   U25 : MUX2_X1 port map( A => DOUT_20_port, B => DIN(20), S => EN, Z => n47);
   U26 : MUX2_X1 port map( A => DOUT_21_port, B => DIN(21), S => EN, Z => n46);
   U27 : MUX2_X1 port map( A => DOUT_22_port, B => DIN(22), S => EN, Z => n45);
   U28 : MUX2_X1 port map( A => DOUT_23_port, B => DIN(23), S => EN, Z => n44);
   U29 : MUX2_X1 port map( A => DOUT_24_port, B => DIN(24), S => EN, Z => n43);
   U30 : MUX2_X1 port map( A => DOUT_25_port, B => DIN(25), S => EN, Z => n42);
   U31 : MUX2_X1 port map( A => DOUT_26_port, B => DIN(26), S => EN, Z => n41);
   U32 : MUX2_X1 port map( A => DOUT_27_port, B => DIN(27), S => EN, Z => n40);
   U33 : MUX2_X1 port map( A => DOUT_28_port, B => DIN(28), S => EN, Z => n39);
   U34 : MUX2_X1 port map( A => DOUT_29_port, B => DIN(29), S => EN, Z => n38);
   U35 : MUX2_X1 port map( A => DOUT_30_port, B => DIN(30), S => EN, Z => n37);
   U36 : MUX2_X1 port map( A => DOUT_31_port, B => DIN(31), S => EN, Z => n36);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_5;

architecture SYN_bhv of mux21_NBIT32_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => S, Z => n1);
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n3);
   U4 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Z(0));
   U5 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Z(1));
   U6 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Z(2));
   U7 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Z(3));
   U8 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Z(4));
   U9 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Z(5));
   U10 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Z(6));
   U11 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Z(7));
   U12 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Z(8));
   U13 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Z(9));
   U14 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Z(10));
   U15 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Z(11));
   U16 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Z(12));
   U17 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Z(13));
   U18 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Z(14));
   U19 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Z(15));
   U20 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Z(16));
   U21 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Z(17));
   U22 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Z(18));
   U23 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Z(19));
   U24 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Z(20));
   U25 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Z(21));
   U26 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Z(22));
   U27 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Z(23));
   U28 : MUX2_X1 port map( A => A(24), B => B(24), S => n3, Z => Z(24));
   U29 : MUX2_X1 port map( A => A(25), B => B(25), S => n3, Z => Z(25));
   U30 : MUX2_X1 port map( A => A(26), B => B(26), S => n3, Z => Z(26));
   U31 : MUX2_X1 port map( A => A(27), B => B(27), S => n3, Z => Z(27));
   U32 : MUX2_X1 port map( A => A(28), B => B(28), S => n3, Z => Z(28));
   U33 : MUX2_X1 port map( A => A(29), B => B(29), S => n3, Z => Z(29));
   U34 : MUX2_X1 port map( A => A(30), B => B(30), S => n3, Z => Z(30));
   U35 : MUX2_X1 port map( A => A(31), B => B(31), S => n3, Z => Z(31));

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_4;

architecture SYN_bhv of mux21_NBIT32_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n15, ZN => n4);
   U2 : INV_X1 port map( A => n15, ZN => n5);
   U3 : BUF_X1 port map( A => n1, Z => n7);
   U4 : BUF_X1 port map( A => n3, Z => n13);
   U5 : BUF_X1 port map( A => n2, Z => n12);
   U6 : BUF_X1 port map( A => n2, Z => n10);
   U7 : BUF_X1 port map( A => n1, Z => n9);
   U8 : BUF_X1 port map( A => n2, Z => n11);
   U9 : BUF_X1 port map( A => n1, Z => n8);
   U10 : BUF_X1 port map( A => n3, Z => n15);
   U11 : BUF_X1 port map( A => n3, Z => n14);
   U12 : BUF_X1 port map( A => S, Z => n3);
   U13 : BUF_X1 port map( A => S, Z => n2);
   U14 : BUF_X1 port map( A => S, Z => n1);
   U15 : INV_X1 port map( A => n91, ZN => Z(1));
   U16 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n11, ZN => 
                           n91);
   U17 : INV_X1 port map( A => n102, ZN => Z(2));
   U18 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => n8, ZN => 
                           n102);
   U19 : INV_X1 port map( A => n105, ZN => Z(3));
   U20 : AOI22_X1 port map( A1 => A(3), A2 => n6, B1 => B(3), B2 => n8, ZN => 
                           n105);
   U21 : INV_X1 port map( A => n106, ZN => Z(4));
   U22 : AOI22_X1 port map( A1 => A(4), A2 => n6, B1 => B(4), B2 => n8, ZN => 
                           n106);
   U23 : INV_X1 port map( A => n107, ZN => Z(5));
   U24 : AOI22_X1 port map( A1 => A(5), A2 => n6, B1 => B(5), B2 => n7, ZN => 
                           n107);
   U25 : INV_X1 port map( A => n108, ZN => Z(6));
   U26 : AOI22_X1 port map( A1 => A(6), A2 => n6, B1 => B(6), B2 => n7, ZN => 
                           n108);
   U27 : INV_X1 port map( A => n109, ZN => Z(7));
   U28 : AOI22_X1 port map( A1 => A(7), A2 => n6, B1 => B(7), B2 => n7, ZN => 
                           n109);
   U29 : INV_X1 port map( A => n110, ZN => Z(8));
   U30 : AOI22_X1 port map( A1 => A(8), A2 => n6, B1 => B(8), B2 => n7, ZN => 
                           n110);
   U31 : INV_X1 port map( A => n81, ZN => Z(10));
   U32 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => B(10), B2 => n14, ZN 
                           => n81);
   U33 : INV_X1 port map( A => n82, ZN => Z(11));
   U34 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => B(11), B2 => n14, ZN 
                           => n82);
   U35 : INV_X1 port map( A => n83, ZN => Z(12));
   U36 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => B(12), B2 => n13, ZN 
                           => n83);
   U37 : INV_X1 port map( A => n84, ZN => Z(13));
   U38 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n13, ZN 
                           => n84);
   U39 : INV_X1 port map( A => n85, ZN => Z(14));
   U40 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n13, ZN 
                           => n85);
   U41 : INV_X1 port map( A => n86, ZN => Z(15));
   U42 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n13, ZN 
                           => n86);
   U43 : INV_X1 port map( A => n87, ZN => Z(16));
   U44 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => B(16), B2 => n12, ZN 
                           => n87);
   U45 : INV_X1 port map( A => n88, ZN => Z(17));
   U46 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n12, ZN 
                           => n88);
   U47 : INV_X1 port map( A => n89, ZN => Z(18));
   U48 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => B(18), B2 => n12, ZN 
                           => n89);
   U49 : INV_X1 port map( A => n90, ZN => Z(19));
   U50 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => B(19), B2 => n12, ZN 
                           => n90);
   U51 : INV_X1 port map( A => n92, ZN => Z(20));
   U52 : AOI22_X1 port map( A1 => A(20), A2 => n5, B1 => B(20), B2 => n11, ZN 
                           => n92);
   U53 : INV_X1 port map( A => n93, ZN => Z(21));
   U54 : AOI22_X1 port map( A1 => A(21), A2 => n5, B1 => B(21), B2 => n11, ZN 
                           => n93);
   U55 : INV_X1 port map( A => n94, ZN => Z(22));
   U56 : AOI22_X1 port map( A1 => A(22), A2 => n5, B1 => B(22), B2 => n10, ZN 
                           => n94);
   U57 : INV_X1 port map( A => n95, ZN => Z(23));
   U58 : AOI22_X1 port map( A1 => A(23), A2 => n5, B1 => B(23), B2 => n10, ZN 
                           => n95);
   U59 : INV_X1 port map( A => n96, ZN => Z(24));
   U60 : AOI22_X1 port map( A1 => A(24), A2 => n5, B1 => B(24), B2 => n10, ZN 
                           => n96);
   U61 : INV_X1 port map( A => n97, ZN => Z(25));
   U62 : AOI22_X1 port map( A1 => A(25), A2 => n5, B1 => B(25), B2 => n10, ZN 
                           => n97);
   U63 : INV_X1 port map( A => n98, ZN => Z(26));
   U64 : AOI22_X1 port map( A1 => A(26), A2 => n5, B1 => B(26), B2 => n9, ZN =>
                           n98);
   U65 : INV_X1 port map( A => n99, ZN => Z(27));
   U66 : AOI22_X1 port map( A1 => A(27), A2 => n5, B1 => B(27), B2 => n9, ZN =>
                           n99);
   U67 : INV_X1 port map( A => n100, ZN => Z(28));
   U68 : AOI22_X1 port map( A1 => A(28), A2 => n5, B1 => B(28), B2 => n9, ZN =>
                           n100);
   U69 : INV_X1 port map( A => n101, ZN => Z(29));
   U70 : AOI22_X1 port map( A1 => A(29), A2 => n5, B1 => B(29), B2 => n9, ZN =>
                           n101);
   U71 : INV_X1 port map( A => n103, ZN => Z(30));
   U72 : AOI22_X1 port map( A1 => A(30), A2 => n5, B1 => B(30), B2 => n11, ZN 
                           => n103);
   U73 : INV_X1 port map( A => n104, ZN => Z(31));
   U74 : AOI22_X1 port map( A1 => A(31), A2 => n6, B1 => B(31), B2 => n8, ZN =>
                           n104);
   U75 : INV_X1 port map( A => n111, ZN => Z(9));
   U76 : AOI22_X1 port map( A1 => A(9), A2 => n6, B1 => n14, B2 => B(9), ZN => 
                           n111);
   U77 : INV_X1 port map( A => n80, ZN => Z(0));
   U78 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => n14, ZN => 
                           n80);
   U79 : INV_X1 port map( A => n15, ZN => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_3;

architecture SYN_bhv of mux21_NBIT32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n68, Z => n1);
   U2 : BUF_X1 port map( A => n68, Z => n2);
   U3 : BUF_X1 port map( A => n68, Z => n3);
   U4 : INV_X1 port map( A => n81, ZN => Z(20));
   U5 : AOI22_X1 port map( A1 => A(20), A2 => n2, B1 => B(20), B2 => S, ZN => 
                           n81);
   U6 : INV_X1 port map( A => n73, ZN => Z(13));
   U7 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => S, ZN => 
                           n73);
   U8 : INV_X1 port map( A => n69, ZN => Z(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => S, ZN => n69
                           );
   U10 : INV_X1 port map( A => n77, ZN => Z(17));
   U11 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => S, ZN => 
                           n77);
   U12 : INV_X1 port map( A => n97, ZN => Z(6));
   U13 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => S, ZN => 
                           n97);
   U14 : INV_X1 port map( A => n85, ZN => Z(24));
   U15 : AOI22_X1 port map( A1 => A(24), A2 => n2, B1 => B(24), B2 => S, ZN => 
                           n85);
   U16 : INV_X1 port map( A => n89, ZN => Z(28));
   U17 : AOI22_X1 port map( A1 => A(28), A2 => n2, B1 => B(28), B2 => S, ZN => 
                           n89);
   U18 : INV_X1 port map( A => n93, ZN => Z(31));
   U19 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => S, ZN => 
                           n93);
   U20 : INV_X1 port map( A => n70, ZN => Z(10));
   U21 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => S, ZN => 
                           n70);
   U22 : INV_X1 port map( A => n82, ZN => Z(21));
   U23 : AOI22_X1 port map( A1 => A(21), A2 => n2, B1 => B(21), B2 => S, ZN => 
                           n82);
   U24 : INV_X1 port map( A => n74, ZN => Z(14));
   U25 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => S, ZN => 
                           n74);
   U26 : INV_X1 port map( A => n78, ZN => Z(18));
   U27 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => S, ZN => 
                           n78);
   U28 : INV_X1 port map( A => n86, ZN => Z(25));
   U29 : AOI22_X1 port map( A1 => A(25), A2 => n2, B1 => B(25), B2 => S, ZN => 
                           n86);
   U30 : INV_X1 port map( A => n90, ZN => Z(29));
   U31 : AOI22_X1 port map( A1 => A(29), A2 => n2, B1 => B(29), B2 => S, ZN => 
                           n90);
   U32 : INV_X1 port map( A => n94, ZN => Z(3));
   U33 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => S, ZN => 
                           n94);
   U34 : INV_X1 port map( A => n98, ZN => Z(7));
   U35 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => S, ZN => 
                           n98);
   U36 : INV_X1 port map( A => n95, ZN => Z(4));
   U37 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => S, ZN => 
                           n95);
   U38 : INV_X1 port map( A => n83, ZN => Z(22));
   U39 : AOI22_X1 port map( A1 => A(22), A2 => n2, B1 => B(22), B2 => S, ZN => 
                           n83);
   U40 : INV_X1 port map( A => n91, ZN => Z(2));
   U41 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => S, ZN => 
                           n91);
   U42 : INV_X1 port map( A => n99, ZN => Z(8));
   U43 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => S, ZN => 
                           n99);
   U44 : INV_X1 port map( A => n87, ZN => Z(26));
   U45 : AOI22_X1 port map( A1 => A(26), A2 => n2, B1 => B(26), B2 => S, ZN => 
                           n87);
   U46 : INV_X1 port map( A => n71, ZN => Z(11));
   U47 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => S, ZN => 
                           n71);
   U48 : INV_X1 port map( A => n75, ZN => Z(15));
   U49 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => S, ZN => 
                           n75);
   U50 : INV_X1 port map( A => n79, ZN => Z(19));
   U51 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => S, ZN => 
                           n79);
   U52 : INV_X1 port map( A => n76, ZN => Z(16));
   U53 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => S, ZN => 
                           n76);
   U54 : INV_X1 port map( A => n72, ZN => Z(12));
   U55 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => S, ZN => 
                           n72);
   U56 : INV_X1 port map( A => n80, ZN => Z(1));
   U57 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => S, ZN => 
                           n80);
   U58 : INV_X1 port map( A => n96, ZN => Z(5));
   U59 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => S, ZN => 
                           n96);
   U60 : INV_X1 port map( A => n92, ZN => Z(30));
   U61 : AOI22_X1 port map( A1 => A(30), A2 => n2, B1 => B(30), B2 => S, ZN => 
                           n92);
   U62 : INV_X1 port map( A => n84, ZN => Z(23));
   U63 : AOI22_X1 port map( A1 => A(23), A2 => n2, B1 => B(23), B2 => S, ZN => 
                           n84);
   U64 : INV_X1 port map( A => n88, ZN => Z(27));
   U65 : AOI22_X1 port map( A1 => A(27), A2 => n2, B1 => B(27), B2 => S, ZN => 
                           n88);
   U66 : INV_X1 port map( A => n100, ZN => Z(9));
   U67 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => S, B2 => B(9), ZN => 
                           n100);
   U68 : INV_X1 port map( A => S, ZN => n68);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_2;

architecture SYN_bhv of mux21_NBIT32_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n68, Z => n1);
   U2 : BUF_X1 port map( A => n68, Z => n2);
   U3 : BUF_X1 port map( A => n68, Z => n3);
   U4 : INV_X1 port map( A => n81, ZN => Z(20));
   U5 : AOI22_X1 port map( A1 => A(20), A2 => n2, B1 => B(20), B2 => S, ZN => 
                           n81);
   U6 : INV_X1 port map( A => n82, ZN => Z(21));
   U7 : AOI22_X1 port map( A1 => A(21), A2 => n2, B1 => B(21), B2 => S, ZN => 
                           n82);
   U8 : INV_X1 port map( A => n83, ZN => Z(22));
   U9 : AOI22_X1 port map( A1 => A(22), A2 => n2, B1 => B(22), B2 => S, ZN => 
                           n83);
   U10 : INV_X1 port map( A => n84, ZN => Z(23));
   U11 : AOI22_X1 port map( A1 => A(23), A2 => n2, B1 => B(23), B2 => S, ZN => 
                           n84);
   U12 : INV_X1 port map( A => n77, ZN => Z(17));
   U13 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => S, ZN => 
                           n77);
   U14 : INV_X1 port map( A => n78, ZN => Z(18));
   U15 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => S, ZN => 
                           n78);
   U16 : INV_X1 port map( A => n79, ZN => Z(19));
   U17 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => S, ZN => 
                           n79);
   U18 : INV_X1 port map( A => n80, ZN => Z(1));
   U19 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => S, ZN => 
                           n80);
   U20 : INV_X1 port map( A => n73, ZN => Z(13));
   U21 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => S, ZN => 
                           n73);
   U22 : INV_X1 port map( A => n74, ZN => Z(14));
   U23 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => S, ZN => 
                           n74);
   U24 : INV_X1 port map( A => n75, ZN => Z(15));
   U25 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => S, ZN => 
                           n75);
   U26 : INV_X1 port map( A => n76, ZN => Z(16));
   U27 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => S, ZN => 
                           n76);
   U28 : INV_X1 port map( A => n69, ZN => Z(0));
   U29 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => S, ZN => 
                           n69);
   U30 : INV_X1 port map( A => n70, ZN => Z(10));
   U31 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => S, ZN => 
                           n70);
   U32 : INV_X1 port map( A => n71, ZN => Z(11));
   U33 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => S, ZN => 
                           n71);
   U34 : INV_X1 port map( A => n72, ZN => Z(12));
   U35 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => S, ZN => 
                           n72);
   U36 : INV_X1 port map( A => n97, ZN => Z(6));
   U37 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => S, ZN => 
                           n97);
   U38 : INV_X1 port map( A => n98, ZN => Z(7));
   U39 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => S, ZN => 
                           n98);
   U40 : INV_X1 port map( A => n99, ZN => Z(8));
   U41 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => S, ZN => 
                           n99);
   U42 : INV_X1 port map( A => n94, ZN => Z(3));
   U43 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => S, ZN => 
                           n94);
   U44 : INV_X1 port map( A => n95, ZN => Z(4));
   U45 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => S, ZN => 
                           n95);
   U46 : INV_X1 port map( A => n96, ZN => Z(5));
   U47 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => S, ZN => 
                           n96);
   U48 : INV_X1 port map( A => n89, ZN => Z(28));
   U49 : AOI22_X1 port map( A1 => A(28), A2 => n2, B1 => B(28), B2 => S, ZN => 
                           n89);
   U50 : INV_X1 port map( A => n90, ZN => Z(29));
   U51 : AOI22_X1 port map( A1 => A(29), A2 => n2, B1 => B(29), B2 => S, ZN => 
                           n90);
   U52 : INV_X1 port map( A => n91, ZN => Z(2));
   U53 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => S, ZN => 
                           n91);
   U54 : INV_X1 port map( A => n92, ZN => Z(30));
   U55 : AOI22_X1 port map( A1 => A(30), A2 => n2, B1 => B(30), B2 => S, ZN => 
                           n92);
   U56 : INV_X1 port map( A => n85, ZN => Z(24));
   U57 : AOI22_X1 port map( A1 => A(24), A2 => n2, B1 => B(24), B2 => S, ZN => 
                           n85);
   U58 : INV_X1 port map( A => n86, ZN => Z(25));
   U59 : AOI22_X1 port map( A1 => A(25), A2 => n2, B1 => B(25), B2 => S, ZN => 
                           n86);
   U60 : INV_X1 port map( A => n87, ZN => Z(26));
   U61 : AOI22_X1 port map( A1 => A(26), A2 => n2, B1 => B(26), B2 => S, ZN => 
                           n87);
   U62 : INV_X1 port map( A => n88, ZN => Z(27));
   U63 : AOI22_X1 port map( A1 => A(27), A2 => n2, B1 => B(27), B2 => S, ZN => 
                           n88);
   U64 : INV_X1 port map( A => n93, ZN => Z(31));
   U65 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => S, ZN => 
                           n93);
   U66 : INV_X1 port map( A => n100, ZN => Z(9));
   U67 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => S, B2 => B(9), ZN => 
                           n100);
   U68 : INV_X1 port map( A => S, ZN => n68);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_1;

architecture SYN_bhv of mux21_NBIT32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => n4);
   U2 : INV_X1 port map( A => n14, ZN => n5);
   U3 : BUF_X1 port map( A => n1, Z => n6);
   U4 : BUF_X1 port map( A => n3, Z => n12);
   U5 : BUF_X1 port map( A => n2, Z => n11);
   U6 : BUF_X1 port map( A => n2, Z => n9);
   U7 : BUF_X1 port map( A => n1, Z => n8);
   U8 : BUF_X1 port map( A => n2, Z => n10);
   U9 : BUF_X1 port map( A => n1, Z => n7);
   U10 : BUF_X1 port map( A => n3, Z => n14);
   U11 : BUF_X1 port map( A => n3, Z => n13);
   U12 : BUF_X1 port map( A => S, Z => n3);
   U13 : BUF_X1 port map( A => S, Z => n2);
   U14 : BUF_X1 port map( A => S, Z => n1);
   U15 : INV_X1 port map( A => n79, ZN => Z(0));
   U16 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => n13, ZN => 
                           n79);
   U17 : INV_X1 port map( A => n90, ZN => Z(1));
   U18 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n10, ZN => 
                           n90);
   U19 : INV_X1 port map( A => n101, ZN => Z(2));
   U20 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           n101);
   U21 : INV_X1 port map( A => n104, ZN => Z(3));
   U22 : AOI22_X1 port map( A1 => A(3), A2 => n4, B1 => B(3), B2 => n7, ZN => 
                           n104);
   U23 : INV_X1 port map( A => n105, ZN => Z(4));
   U24 : AOI22_X1 port map( A1 => A(4), A2 => n5, B1 => B(4), B2 => n7, ZN => 
                           n105);
   U25 : INV_X1 port map( A => n106, ZN => Z(5));
   U26 : AOI22_X1 port map( A1 => A(5), A2 => n4, B1 => B(5), B2 => n6, ZN => 
                           n106);
   U27 : INV_X1 port map( A => n107, ZN => Z(6));
   U28 : AOI22_X1 port map( A1 => A(6), A2 => n5, B1 => B(6), B2 => n6, ZN => 
                           n107);
   U29 : INV_X1 port map( A => n108, ZN => Z(7));
   U30 : AOI22_X1 port map( A1 => A(7), A2 => n4, B1 => B(7), B2 => n6, ZN => 
                           n108);
   U31 : INV_X1 port map( A => n109, ZN => Z(8));
   U32 : AOI22_X1 port map( A1 => A(8), A2 => n5, B1 => B(8), B2 => n6, ZN => 
                           n109);
   U33 : INV_X1 port map( A => n110, ZN => Z(9));
   U34 : AOI22_X1 port map( A1 => A(9), A2 => n4, B1 => n13, B2 => B(9), ZN => 
                           n110);
   U35 : INV_X1 port map( A => n80, ZN => Z(10));
   U36 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => B(10), B2 => n13, ZN 
                           => n80);
   U37 : INV_X1 port map( A => n81, ZN => Z(11));
   U38 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => B(11), B2 => n13, ZN 
                           => n81);
   U39 : INV_X1 port map( A => n82, ZN => Z(12));
   U40 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => B(12), B2 => n12, ZN 
                           => n82);
   U41 : INV_X1 port map( A => n83, ZN => Z(13));
   U42 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n12, ZN 
                           => n83);
   U43 : INV_X1 port map( A => n84, ZN => Z(14));
   U44 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n12, ZN 
                           => n84);
   U45 : INV_X1 port map( A => n85, ZN => Z(15));
   U46 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n12, ZN 
                           => n85);
   U47 : INV_X1 port map( A => n86, ZN => Z(16));
   U48 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => B(16), B2 => n11, ZN 
                           => n86);
   U49 : INV_X1 port map( A => n87, ZN => Z(17));
   U50 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n11, ZN 
                           => n87);
   U51 : INV_X1 port map( A => n88, ZN => Z(18));
   U52 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => B(18), B2 => n11, ZN 
                           => n88);
   U53 : INV_X1 port map( A => n89, ZN => Z(19));
   U54 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => B(19), B2 => n11, ZN 
                           => n89);
   U55 : INV_X1 port map( A => n91, ZN => Z(20));
   U56 : AOI22_X1 port map( A1 => A(20), A2 => n5, B1 => B(20), B2 => n10, ZN 
                           => n91);
   U57 : INV_X1 port map( A => n92, ZN => Z(21));
   U58 : AOI22_X1 port map( A1 => A(21), A2 => n5, B1 => B(21), B2 => n10, ZN 
                           => n92);
   U59 : INV_X1 port map( A => n93, ZN => Z(22));
   U60 : AOI22_X1 port map( A1 => A(22), A2 => n5, B1 => B(22), B2 => n9, ZN =>
                           n93);
   U61 : INV_X1 port map( A => n94, ZN => Z(23));
   U62 : AOI22_X1 port map( A1 => A(23), A2 => n5, B1 => B(23), B2 => n9, ZN =>
                           n94);
   U63 : INV_X1 port map( A => n95, ZN => Z(24));
   U64 : AOI22_X1 port map( A1 => A(24), A2 => n5, B1 => B(24), B2 => n9, ZN =>
                           n95);
   U65 : INV_X1 port map( A => n96, ZN => Z(25));
   U66 : AOI22_X1 port map( A1 => A(25), A2 => n5, B1 => B(25), B2 => n9, ZN =>
                           n96);
   U67 : INV_X1 port map( A => n97, ZN => Z(26));
   U68 : AOI22_X1 port map( A1 => A(26), A2 => n5, B1 => B(26), B2 => n8, ZN =>
                           n97);
   U69 : INV_X1 port map( A => n98, ZN => Z(27));
   U70 : AOI22_X1 port map( A1 => A(27), A2 => n5, B1 => B(27), B2 => n8, ZN =>
                           n98);
   U71 : INV_X1 port map( A => n99, ZN => Z(28));
   U72 : AOI22_X1 port map( A1 => A(28), A2 => n5, B1 => B(28), B2 => n8, ZN =>
                           n99);
   U73 : INV_X1 port map( A => n100, ZN => Z(29));
   U74 : AOI22_X1 port map( A1 => A(29), A2 => n5, B1 => B(29), B2 => n8, ZN =>
                           n100);
   U75 : INV_X1 port map( A => n102, ZN => Z(30));
   U76 : AOI22_X1 port map( A1 => A(30), A2 => n5, B1 => B(30), B2 => n10, ZN 
                           => n102);
   U77 : INV_X1 port map( A => n103, ZN => Z(31));
   U78 : AOI22_X1 port map( A1 => A(31), A2 => n5, B1 => B(31), B2 => n7, ZN =>
                           n103);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ff_2 is

   port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);

end ff_2;

architecture SYN_bhv of ff_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CLK, RN => RST, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => EN, A => n6, ZN => n4);
   U3 : NAND2_X1 port map( A1 => EN, A2 => D, ZN => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ff_1 is

   port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);

end ff_1;

architecture SYN_bhv of ff_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CLK, RN => RST, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => EN, A => n6, ZN => n4);
   U3 : NAND2_X1 port map( A1 => EN, A2 => D, ZN => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_0;

architecture SYN_STRUCTURAL of RCA_N4_0 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_0;

architecture SYN_struct of carry_select_basic_N4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n6, n7, n8, n9, n1
      , n_1369, n_1370 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1369);
   RCA1 : RCA_N4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1370);
   U3 : INV_X1 port map( A => n7, ZN => S(2));
   U4 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n1, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n7);
   U5 : INV_X1 port map( A => n6, ZN => S(3));
   U6 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n1, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n6);
   U7 : INV_X1 port map( A => n9, ZN => S(0));
   U8 : INV_X1 port map( A => n8, ZN => S(1));
   U9 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n1, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n8);
   U10 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n1, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n9);
   U11 : INV_X1 port map( A => C_i, ZN => n1);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_0 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_0;

architecture SYN_bhv of PGblock_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n2);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_0 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_0;

architecture SYN_bhv of Gblock_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_0 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_0;

architecture SYN_bhv of PG_net_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8;

architecture SYN_structural of SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   component carry_select_basic_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CSBI_1 : carry_select_basic_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) 
                           => A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), 
                           B(1) => B(1), B(0) => B(0), C_i => Ci(0), S(3) => 
                           S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CSBI_2 : carry_select_basic_N4_7 port map( A(3) => A(7), A(2) => A(6), A(1) 
                           => A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), 
                           B(1) => B(5), B(0) => B(4), C_i => Ci(1), S(3) => 
                           S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   CSBI_3 : carry_select_basic_N4_6 port map( A(3) => A(11), A(2) => A(10), 
                           A(1) => A(9), A(0) => A(8), B(3) => B(11), B(2) => 
                           B(10), B(1) => B(9), B(0) => B(8), C_i => Ci(2), 
                           S(3) => S(11), S(2) => S(10), S(1) => S(9), S(0) => 
                           S(8));
   CSBI_4 : carry_select_basic_N4_5 port map( A(3) => A(15), A(2) => A(14), 
                           A(1) => A(13), A(0) => A(12), B(3) => B(15), B(2) =>
                           B(14), B(1) => B(13), B(0) => B(12), C_i => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   CSBI_5 : carry_select_basic_N4_4 port map( A(3) => A(19), A(2) => A(18), 
                           A(1) => A(17), A(0) => A(16), B(3) => B(19), B(2) =>
                           B(18), B(1) => B(17), B(0) => B(16), C_i => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   CSBI_6 : carry_select_basic_N4_3 port map( A(3) => A(23), A(2) => A(22), 
                           A(1) => A(21), A(0) => A(20), B(3) => B(23), B(2) =>
                           B(22), B(1) => B(21), B(0) => B(20), C_i => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   CSBI_7 : carry_select_basic_N4_2 port map( A(3) => A(27), A(2) => A(26), 
                           A(1) => A(25), A(0) => A(24), B(3) => B(27), B(2) =>
                           B(26), B(1) => B(25), B(0) => B(24), C_i => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   CSBI_8 : carry_select_basic_N4_1 port map( A(3) => A(31), A(2) => A(30), 
                           A(1) => A(29), A(0) => A(28), B(3) => B(31), B(2) =>
                           B(30), B(1) => B(29), B(0) => B(28), C_i => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_generator_NBIT32_NBIT_PER_BLOCK4 is

   port( A, B : in std_logic_vector (32 downto 1);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end carry_generator_NBIT32_NBIT_PER_BLOCK4;

architecture SYN_struct of carry_generator_NBIT32_NBIT_PER_BLOCK4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component PGblock_1
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_2
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_3
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_4
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_5
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_6
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_7
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_8
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_9
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_10
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_11
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_12
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_13
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_14
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_15
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_16
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_17
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_18
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_19
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_20
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_21
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_22
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_23
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_24
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_25
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_26
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_0
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component Gblock_1
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_2
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_3
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_4
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_5
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_6
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_7
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_8
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_0
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_net_1
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_2
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_3
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_4
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_5
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_6
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_7
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_8
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_9
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_10
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_11
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_12
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_13
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_14
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_15
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_16
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_17
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_18
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_19
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_20
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_21
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_22
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_23
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_24
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_25
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_26
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_27
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_28
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_29
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_30
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_0
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   signal Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port, G_16_16_port, G_16_15_port, G_16_13_port, 
      G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, G_13_13_port, 
      G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, G_10_10_port, 
      G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port, G_7_7_port, 
      G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port, G_3_3_port, 
      G_2_2_port, G_2_1_port, G_1_1_port, P_16_16_port, P_16_15_port, 
      P_16_13_port, P_16_9_port, P_15_15_port, P_14_14_port, P_14_13_port, 
      P_13_13_port, P_12_12_port, P_12_11_port, P_12_9_port, P_11_11_port, 
      P_10_10_port, P_10_9_port, P_9_9_port, P_8_8_port, P_8_7_port, P_8_5_port
      , P_7_7_port, P_6_6_port, P_6_5_port, P_5_5_port, P_4_4_port, P_4_3_port,
      P_3_3_port, P_2_2_port, G_32_32_port, G_32_31_port, G_32_29_port, 
      G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, G_30_29_port, 
      G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, G_28_17_port, 
      G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, G_24_24_port, 
      G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, G_22_22_port, 
      G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, G_20_17_port, 
      G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, P_32_32_port, 
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n3, n1, n2 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port );
   
   PGnetblock_2 : PG_net_0 port map( a => A(2), b => B(2), p => P_2_2_port, g 
                           => G_2_2_port);
   PGnetblock_3 : PG_net_30 port map( a => A(3), b => B(3), p => P_3_3_port, g 
                           => G_3_3_port);
   PGnetblock_4 : PG_net_29 port map( a => A(4), b => B(4), p => P_4_4_port, g 
                           => G_4_4_port);
   PGnetblock_5 : PG_net_28 port map( a => A(5), b => B(5), p => P_5_5_port, g 
                           => G_5_5_port);
   PGnetblock_6 : PG_net_27 port map( a => A(6), b => B(6), p => P_6_6_port, g 
                           => G_6_6_port);
   PGnetblock_7 : PG_net_26 port map( a => A(7), b => B(7), p => P_7_7_port, g 
                           => G_7_7_port);
   PGnetblock_8 : PG_net_25 port map( a => A(8), b => B(8), p => P_8_8_port, g 
                           => G_8_8_port);
   PGnetblock_9 : PG_net_24 port map( a => A(9), b => B(9), p => P_9_9_port, g 
                           => G_9_9_port);
   PGnetblock_10 : PG_net_23 port map( a => A(10), b => B(10), p => 
                           P_10_10_port, g => G_10_10_port);
   PGnetblock_11 : PG_net_22 port map( a => A(11), b => B(11), p => 
                           P_11_11_port, g => G_11_11_port);
   PGnetblock_12 : PG_net_21 port map( a => A(12), b => B(12), p => 
                           P_12_12_port, g => G_12_12_port);
   PGnetblock_13 : PG_net_20 port map( a => A(13), b => B(13), p => 
                           P_13_13_port, g => G_13_13_port);
   PGnetblock_14 : PG_net_19 port map( a => A(14), b => B(14), p => 
                           P_14_14_port, g => G_14_14_port);
   PGnetblock_15 : PG_net_18 port map( a => A(15), b => B(15), p => 
                           P_15_15_port, g => G_15_15_port);
   PGnetblock_16 : PG_net_17 port map( a => A(16), b => B(16), p => 
                           P_16_16_port, g => G_16_16_port);
   PGnetblock_17 : PG_net_16 port map( a => A(17), b => B(17), p => 
                           P_17_17_port, g => G_17_17_port);
   PGnetblock_18 : PG_net_15 port map( a => A(18), b => B(18), p => 
                           P_18_18_port, g => G_18_18_port);
   PGnetblock_19 : PG_net_14 port map( a => A(19), b => B(19), p => 
                           P_19_19_port, g => G_19_19_port);
   PGnetblock_20 : PG_net_13 port map( a => A(20), b => B(20), p => 
                           P_20_20_port, g => G_20_20_port);
   PGnetblock_21 : PG_net_12 port map( a => A(21), b => B(21), p => 
                           P_21_21_port, g => G_21_21_port);
   PGnetblock_22 : PG_net_11 port map( a => A(22), b => B(22), p => 
                           P_22_22_port, g => G_22_22_port);
   PGnetblock_23 : PG_net_10 port map( a => A(23), b => B(23), p => 
                           P_23_23_port, g => G_23_23_port);
   PGnetblock_24 : PG_net_9 port map( a => A(24), b => B(24), p => P_24_24_port
                           , g => G_24_24_port);
   PGnetblock_25 : PG_net_8 port map( a => A(25), b => B(25), p => P_25_25_port
                           , g => G_25_25_port);
   PGnetblock_26 : PG_net_7 port map( a => A(26), b => B(26), p => P_26_26_port
                           , g => G_26_26_port);
   PGnetblock_27 : PG_net_6 port map( a => A(27), b => B(27), p => P_27_27_port
                           , g => G_27_27_port);
   PGnetblock_28 : PG_net_5 port map( a => A(28), b => B(28), p => P_28_28_port
                           , g => G_28_28_port);
   PGnetblock_29 : PG_net_4 port map( a => A(29), b => B(29), p => P_29_29_port
                           , g => G_29_29_port);
   PGnetblock_30 : PG_net_3 port map( a => A(30), b => B(30), p => P_30_30_port
                           , g => G_30_30_port);
   PGnetblock_31 : PG_net_2 port map( a => A(31), b => B(31), p => P_31_31_port
                           , g => G_31_31_port);
   PGnetblock_32 : PG_net_1 port map( a => A(32), b => B(32), p => P_32_32_port
                           , g => G_32_32_port);
   GB_low_1_2 : Gblock_0 port map( Pik => P_2_2_port, Gik => G_2_2_port, Gk_1j 
                           => G_1_1_port, Gij => G_2_1_port);
   GB_low_2_4 : Gblock_8 port map( Pik => P_4_3_port, Gik => G_4_3_port, Gk_1j 
                           => G_2_1_port, Gij => Co_0_port);
   GB_low_3_8 : Gblock_7 port map( Pik => P_8_5_port, Gik => G_8_5_port, Gk_1j 
                           => Co_0_port, Gij => Co_1_port);
   GB_high_4_16_0 : Gblock_6 port map( Pik => P_16_9_port, Gik => G_16_9_port, 
                           Gk_1j => Co_1_port, Gij => Co_3_port);
   GB_high_4_16_1 : Gblock_5 port map( Pik => P_12_9_port, Gik => G_12_9_port, 
                           Gk_1j => Co_1_port, Gij => Co_2_port);
   GB_high_5_32_0 : Gblock_4 port map( Pik => P_32_17_port, Gik => G_32_17_port
                           , Gk_1j => Co_3_port, Gij => Co_7_port);
   GB_high_5_32_1 : Gblock_3 port map( Pik => P_28_17_port, Gik => G_28_17_port
                           , Gk_1j => Co_3_port, Gij => Co_6_port);
   GB_high_5_32_2 : Gblock_2 port map( Pik => P_24_17_port, Gik => G_24_17_port
                           , Gk_1j => Co_3_port, Gij => Co_5_port);
   GB_high_5_32_3 : Gblock_1 port map( Pik => P_20_17_port, Gik => G_20_17_port
                           , Gk_1j => Co_3_port, Gij => Co_4_port);
   PGB_low_1_4 : PGblock_0 port map( Pik => P_4_4_port, Gik => G_4_4_port, 
                           Pk_1j => P_3_3_port, Gk_1j => G_3_3_port, Pij => 
                           P_4_3_port, Gij => G_4_3_port);
   PGB_low_1_6 : PGblock_26 port map( Pik => P_6_6_port, Gik => G_6_6_port, 
                           Pk_1j => P_5_5_port, Gk_1j => G_5_5_port, Pij => 
                           P_6_5_port, Gij => G_6_5_port);
   PGB_low_1_8 : PGblock_25 port map( Pik => P_8_8_port, Gik => G_8_8_port, 
                           Pk_1j => P_7_7_port, Gk_1j => G_7_7_port, Pij => 
                           P_8_7_port, Gij => G_8_7_port);
   PGB_low_1_10 : PGblock_24 port map( Pik => P_10_10_port, Gik => G_10_10_port
                           , Pk_1j => P_9_9_port, Gk_1j => G_9_9_port, Pij => 
                           P_10_9_port, Gij => G_10_9_port);
   PGB_low_1_12 : PGblock_23 port map( Pik => P_12_12_port, Gik => G_12_12_port
                           , Pk_1j => P_11_11_port, Gk_1j => G_11_11_port, Pij 
                           => P_12_11_port, Gij => G_12_11_port);
   PGB_low_1_14 : PGblock_22 port map( Pik => P_14_14_port, Gik => G_14_14_port
                           , Pk_1j => P_13_13_port, Gk_1j => G_13_13_port, Pij 
                           => P_14_13_port, Gij => G_14_13_port);
   PGB_low_1_16 : PGblock_21 port map( Pik => P_16_16_port, Gik => G_16_16_port
                           , Pk_1j => P_15_15_port, Gk_1j => G_15_15_port, Pij 
                           => P_16_15_port, Gij => G_16_15_port);
   PGB_low_1_18 : PGblock_20 port map( Pik => P_18_18_port, Gik => G_18_18_port
                           , Pk_1j => P_17_17_port, Gk_1j => G_17_17_port, Pij 
                           => P_18_17_port, Gij => G_18_17_port);
   PGB_low_1_20 : PGblock_19 port map( Pik => P_20_20_port, Gik => G_20_20_port
                           , Pk_1j => P_19_19_port, Gk_1j => G_19_19_port, Pij 
                           => P_20_19_port, Gij => G_20_19_port);
   PGB_low_1_22 : PGblock_18 port map( Pik => P_22_22_port, Gik => G_22_22_port
                           , Pk_1j => P_21_21_port, Gk_1j => G_21_21_port, Pij 
                           => P_22_21_port, Gij => G_22_21_port);
   PGB_low_1_24 : PGblock_17 port map( Pik => P_24_24_port, Gik => G_24_24_port
                           , Pk_1j => P_23_23_port, Gk_1j => G_23_23_port, Pij 
                           => P_24_23_port, Gij => G_24_23_port);
   PGB_low_1_26 : PGblock_16 port map( Pik => P_26_26_port, Gik => G_26_26_port
                           , Pk_1j => P_25_25_port, Gk_1j => G_25_25_port, Pij 
                           => P_26_25_port, Gij => G_26_25_port);
   PGB_low_1_28 : PGblock_15 port map( Pik => P_28_28_port, Gik => G_28_28_port
                           , Pk_1j => P_27_27_port, Gk_1j => G_27_27_port, Pij 
                           => P_28_27_port, Gij => G_28_27_port);
   PGB_low_1_30 : PGblock_14 port map( Pik => P_30_30_port, Gik => G_30_30_port
                           , Pk_1j => P_29_29_port, Gk_1j => G_29_29_port, Pij 
                           => P_30_29_port, Gij => G_30_29_port);
   PGB_low_1_32 : PGblock_13 port map( Pik => P_32_32_port, Gik => G_32_32_port
                           , Pk_1j => P_31_31_port, Gk_1j => G_31_31_port, Pij 
                           => P_32_31_port, Gij => G_32_31_port);
   PGB_low_2_8 : PGblock_12 port map( Pik => P_8_7_port, Gik => G_8_7_port, 
                           Pk_1j => P_6_5_port, Gk_1j => G_6_5_port, Pij => 
                           P_8_5_port, Gij => G_8_5_port);
   PGB_low_2_12 : PGblock_11 port map( Pik => P_12_11_port, Gik => G_12_11_port
                           , Pk_1j => P_10_9_port, Gk_1j => G_10_9_port, Pij =>
                           P_12_9_port, Gij => G_12_9_port);
   PGB_low_2_16 : PGblock_10 port map( Pik => P_16_15_port, Gik => G_16_15_port
                           , Pk_1j => P_14_13_port, Gk_1j => G_14_13_port, Pij 
                           => P_16_13_port, Gij => G_16_13_port);
   PGB_low_2_20 : PGblock_9 port map( Pik => P_20_19_port, Gik => G_20_19_port,
                           Pk_1j => P_18_17_port, Gk_1j => G_18_17_port, Pij =>
                           P_20_17_port, Gij => G_20_17_port);
   PGB_low_2_24 : PGblock_8 port map( Pik => P_24_23_port, Gik => G_24_23_port,
                           Pk_1j => P_22_21_port, Gk_1j => G_22_21_port, Pij =>
                           P_24_21_port, Gij => G_24_21_port);
   PGB_low_2_28 : PGblock_7 port map( Pik => P_28_27_port, Gik => G_28_27_port,
                           Pk_1j => P_26_25_port, Gk_1j => G_26_25_port, Pij =>
                           P_28_25_port, Gij => G_28_25_port);
   PGB_low_2_32 : PGblock_6 port map( Pik => P_32_31_port, Gik => G_32_31_port,
                           Pk_1j => P_30_29_port, Gk_1j => G_30_29_port, Pij =>
                           P_32_29_port, Gij => G_32_29_port);
   PGB_low_3_16 : PGblock_5 port map( Pik => P_16_13_port, Gik => G_16_13_port,
                           Pk_1j => P_12_9_port, Gk_1j => G_12_9_port, Pij => 
                           P_16_9_port, Gij => G_16_9_port);
   PGB_low_3_24 : PGblock_4 port map( Pik => P_24_21_port, Gik => G_24_21_port,
                           Pk_1j => P_20_17_port, Gk_1j => G_20_17_port, Pij =>
                           P_24_17_port, Gij => G_24_17_port);
   PGB_low_3_32 : PGblock_3 port map( Pik => P_32_29_port, Gik => G_32_29_port,
                           Pk_1j => P_28_25_port, Gk_1j => G_28_25_port, Pij =>
                           P_32_25_port, Gij => G_32_25_port);
   PGB_high_4_32_0 : PGblock_2 port map( Pik => P_32_25_port, Gik => 
                           G_32_25_port, Pk_1j => P_24_17_port, Gk_1j => 
                           G_24_17_port, Pij => P_32_17_port, Gij => 
                           G_32_17_port);
   PGB_high_4_32_1 : PGblock_1 port map( Pik => P_28_25_port, Gik => 
                           G_28_25_port, Pk_1j => P_24_17_port, Gk_1j => 
                           G_24_17_port, Pij => P_28_17_port, Gij => 
                           G_28_17_port);
   U1 : INV_X1 port map( A => A(1), ZN => n1);
   U2 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => G_1_1_port);
   U3 : OAI21_X1 port map( B1 => A(1), B2 => B(1), A => Cin, ZN => n3);
   U4 : INV_X1 port map( A => B(1), ZN => n2);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity P4Adder_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (31 downto 0);  Cout : out std_logic);

end P4Adder_NBIT32;

architecture SYN_struct of P4Adder_NBIT32 is

   component SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component carry_generator_NBIT32_NBIT_PER_BLOCK4
      port( A, B : in std_logic_vector (32 downto 1);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal Csum_7_port, Csum_6_port, Csum_5_port, Csum_4_port, Csum_3_port, 
      Csum_2_port, Csum_1_port : std_logic;

begin
   
   Carrygen0 : carry_generator_NBIT32_NBIT_PER_BLOCK4 port map( A(32) => A(31),
                           A(31) => A(30), A(30) => A(29), A(29) => A(28), 
                           A(28) => A(27), A(27) => A(26), A(26) => A(25), 
                           A(25) => A(24), A(24) => A(23), A(23) => A(22), 
                           A(22) => A(21), A(21) => A(20), A(20) => A(19), 
                           A(19) => A(18), A(18) => A(17), A(17) => A(16), 
                           A(16) => A(15), A(15) => A(14), A(14) => A(13), 
                           A(13) => A(12), A(12) => A(11), A(11) => A(10), 
                           A(10) => A(9), A(9) => A(8), A(8) => A(7), A(7) => 
                           A(6), A(6) => A(5), A(5) => A(4), A(4) => A(3), A(3)
                           => A(2), A(2) => A(1), A(1) => A(0), B(32) => B(31),
                           B(31) => B(30), B(30) => B(29), B(29) => B(28), 
                           B(28) => B(27), B(27) => B(26), B(26) => B(25), 
                           B(25) => B(24), B(24) => B(23), B(23) => B(22), 
                           B(22) => B(21), B(21) => B(20), B(20) => B(19), 
                           B(19) => B(18), B(18) => B(17), B(17) => B(16), 
                           B(16) => B(15), B(15) => B(14), B(14) => B(13), 
                           B(13) => B(12), B(12) => B(11), B(11) => B(10), 
                           B(10) => B(9), B(9) => B(8), B(8) => B(7), B(7) => 
                           B(6), B(6) => B(5), B(5) => B(4), B(4) => B(3), B(3)
                           => B(2), B(2) => B(1), B(1) => B(0), Cin => Cin, 
                           Co(7) => Cout, Co(6) => Csum_7_port, Co(5) => 
                           Csum_6_port, Co(4) => Csum_5_port, Co(3) => 
                           Csum_4_port, Co(2) => Csum_3_port, Co(1) => 
                           Csum_2_port, Co(0) => Csum_1_port);
   Sumgen0 : SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), Ci(7) => 
                           Csum_7_port, Ci(6) => Csum_6_port, Ci(5) => 
                           Csum_5_port, Ci(4) => Csum_4_port, Ci(3) => 
                           Csum_3_port, Ci(2) => Csum_2_port, Ci(1) => 
                           Csum_1_port, Ci(0) => Cin, S(31) => S(31), S(30) => 
                           S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           S(21), S(20) => S(20), S(19) => S(19), S(18) => 
                           S(18), S(17) => S(17), S(16) => S(16), S(15) => 
                           S(15), S(14) => S(14), S(13) => S(13), S(12) => 
                           S(12), S(11) => S(11), S(10) => S(10), S(9) => S(9),
                           S(8) => S(8), S(7) => S(7), S(6) => S(6), S(5) => 
                           S(5), S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1)
                           => S(1), S(0) => S(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity shifter_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  LOGIC_ARITH, LEFT_RIGHT : 
         in std_logic;  RES : out std_logic_vector (31 downto 0));

end shifter_NBIT32;

architecture SYN_bhv of shifter_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X4
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X2
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, 
      n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
      n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, 
      n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, 
      n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n1, n2, n3, n4, n5, n6, 
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n266, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648 : std_logic;

begin
   
   U264 : AOI21_X2 port map( B1 => A(31), B2 => B(18), A => n483, ZN => n282);
   U267 : OAI21_X2 port map( B1 => n612, B2 => n628, A => n486, ZN => n285);
   U269 : AOI21_X2 port map( B1 => A(31), B2 => n38, A => n487, ZN => n288);
   U388 : AOI221_X2 port map( B1 => n30, B2 => A(18), C1 => n21, C2 => A(17), A
                           => n568, ZN => n196);
   U428 : NOR2_X2 port map( A1 => n638, A2 => n38, ZN => n165);
   U461 : NOR2_X2 port map( A1 => n642, A2 => n38, ZN => n199);
   U637 : NAND3_X1 port map( A1 => n227, A2 => n646, A3 => n228, ZN => n226);
   U638 : NAND3_X1 port map( A1 => n227, A2 => n646, A3 => B(4), ZN => n428);
   U639 : NAND3_X1 port map( A1 => n445, A2 => n199, A3 => LEFT_RIGHT, ZN => 
                           n240);
   U641 : NAND3_X1 port map( A1 => n489, A2 => n628, A3 => n579, ZN => n255);
   U642 : NAND3_X1 port map( A1 => n7, A2 => n199, A3 => n445, ZN => n138);
   U2 : NOR4_X1 port map( A1 => B(20), A2 => B(21), A3 => B(19), A4 => n594, ZN
                           => n484);
   U3 : NOR2_X2 port map( A1 => n639, A2 => B(3), ZN => n262);
   U4 : AOI221_X1 port map( B1 => n29, B2 => A(6), C1 => n19, C2 => A(7), A => 
                           n525, ZN => n363);
   U5 : AOI221_X1 port map( B1 => n30, B2 => A(7), C1 => n20, C2 => A(8), A => 
                           n570, ZN => n405);
   U6 : AOI221_X1 port map( B1 => n29, B2 => A(8), C1 => n21, C2 => A(9), A => 
                           n552, ZN => n387);
   U7 : AOI222_X1 port map( A1 => n11, A2 => A(1), B1 => A(0), B2 => n18, C1 =>
                           n7, C2 => A(2), ZN => n293);
   U8 : OAI21_X2 port map( B1 => n266, B2 => n632, A => n481, ZN => n279);
   U9 : INV_X1 port map( A => n167, ZN => n635);
   U10 : NOR2_X1 port map( A1 => n636, A2 => B(4), ZN => n167);
   U11 : INV_X1 port map( A => n169, ZN => n644);
   U12 : INV_X1 port map( A => n165, ZN => n637);
   U13 : INV_X1 port map( A => n199, ZN => n641);
   U14 : INV_X1 port map( A => n28, ZN => n26);
   U15 : INV_X1 port map( A => n31, ZN => n24);
   U16 : INV_X1 port map( A => n31, ZN => n25);
   U17 : INV_X1 port map( A => n21, ZN => n14);
   U18 : INV_X1 port map( A => n19, ZN => n16);
   U19 : INV_X1 port map( A => n19, ZN => n15);
   U20 : INV_X1 port map( A => n505, ZN => n643);
   U21 : INV_X1 port map( A => n29, ZN => n27);
   U22 : INV_X1 port map( A => n493, ZN => n640);
   U23 : NOR2_X1 port map( A1 => n645, A2 => n38, ZN => n169);
   U24 : NAND2_X1 port map( A1 => n488, A2 => n454, ZN => n161);
   U25 : INV_X1 port map( A => n41, ZN => n38);
   U26 : OAI222_X1 port map( A1 => n637, A2 => n70, B1 => n635, B2 => n92, C1 
                           => n644, C2 => n80, ZN => n224);
   U27 : OAI222_X1 port map( A1 => n637, A2 => n67, B1 => n635, B2 => n96, C1 
                           => n644, C2 => n83, ZN => n212);
   U28 : NOR2_X1 port map( A1 => n40, A2 => n642, ZN => n493);
   U29 : OAI22_X1 port map( A1 => n115, A2 => n642, B1 => n126, B2 => n638, ZN 
                           => n383);
   U30 : INV_X1 port map( A => n454, ZN => n636);
   U31 : AOI21_X1 port map( B1 => n134, B2 => n2, A => n519, ZN => n286);
   U32 : AOI21_X1 port map( B1 => n129, B2 => n3, A => n519, ZN => n312);
   U33 : BUF_X1 port map( A => n138, Z => n33);
   U34 : BUF_X1 port map( A => n138, Z => n32);
   U35 : NOR2_X1 port map( A1 => n383, A2 => n359, ZN => n197);
   U36 : NOR2_X1 port map( A1 => n118, A2 => n359, ZN => n181);
   U37 : BUF_X1 port map( A => n138, Z => n34);
   U38 : NAND2_X1 port map( A1 => n488, A2 => n5, ZN => n505);
   U39 : INV_X1 port map( A => n182, ZN => n118);
   U40 : INV_X1 port map( A => n172, ZN => n54);
   U41 : INV_X1 port map( A => n139, ZN => n58);
   U42 : INV_X1 port map( A => n348, ZN => n52);
   U43 : INV_X1 port map( A => n337, ZN => n44);
   U44 : INV_X1 port map( A => n480, ZN => n88);
   U45 : INV_X1 port map( A => n314, ZN => n56);
   U46 : INV_X1 port map( A => n290, ZN => n50);
   U47 : INV_X1 port map( A => n271, ZN => n46);
   U48 : INV_X1 port map( A => n257, ZN => n101);
   U49 : INV_X1 port map( A => n440, ZN => n93);
   U50 : INV_X1 port map( A => n302, ZN => n97);
   U51 : NOR2_X1 port map( A1 => n612, A2 => n148, ZN => n150);
   U52 : NOR2_X1 port map( A1 => n639, A2 => n646, ZN => n454);
   U53 : NAND2_X1 port map( A1 => n484, A2 => n630, ZN => n281);
   U54 : AOI222_X1 port map( A1 => n370, A2 => n262, B1 => n320, B2 => n260, C1
                           => n185, C2 => n3, ZN => n238);
   U55 : INV_X1 port map( A => n356, ZN => n642);
   U56 : AOI222_X1 port map( A1 => n168, A2 => n262, B1 => n355, B2 => n260, C1
                           => n170, C2 => n3, ZN => n471);
   U57 : AOI222_X1 port map( A1 => n402, A2 => n262, B1 => n403, B2 => n260, C1
                           => n464, C2 => n2, ZN => n461);
   U58 : NAND2_X1 port map( A1 => n488, A2 => n262, ZN => n157);
   U59 : NAND2_X1 port map( A1 => n488, A2 => n260, ZN => n158);
   U60 : OAI222_X1 port map( A1 => n374, A2 => n638, B1 => n645, B2 => n375, C1
                           => n376, C2 => n642, ZN => n172);
   U61 : OAI222_X1 port map( A1 => n131, A2 => n638, B1 => n362, B2 => n645, C1
                           => n363, C2 => n642, ZN => n139);
   U62 : OAI222_X1 port map( A1 => n613, A2 => n638, B1 => n293, B2 => n645, C1
                           => n405, C2 => n642, ZN => n348);
   U63 : OAI222_X1 port map( A1 => n615, A2 => n638, B1 => n45, B2 => n645, C1 
                           => n387, C2 => n642, ZN => n337);
   U64 : AOI221_X1 port map( B1 => n129, B2 => n262, C1 => n355, C2 => n2, A =>
                           n359, ZN => n159);
   U65 : AOI221_X1 port map( B1 => n134, B2 => n262, C1 => n403, C2 => n3, A =>
                           n359, ZN => n347);
   U66 : OAI221_X1 port map( B1 => n105, B2 => n638, C1 => n89, C2 => n642, A 
                           => n607, ZN => n480);
   U67 : AOI22_X1 port map( A1 => n454, A2 => n320, B1 => n260, B2 => n370, ZN 
                           => n607);
   U68 : AOI222_X1 port map( A1 => n169, A2 => n185, B1 => n493, B2 => n320, C1
                           => n167, C2 => n370, ZN => n550);
   U69 : AOI222_X1 port map( A1 => n165, A2 => n166, B1 => n167, B2 => n168, C1
                           => n169, C2 => n170, ZN => n164);
   U70 : AOI222_X1 port map( A1 => n165, A2 => n516, B1 => n167, B2 => n402, C1
                           => n169, C2 => n464, ZN => n581);
   U71 : AOI222_X1 port map( A1 => n165, A2 => n184, B1 => n167, B2 => n185, C1
                           => n169, C2 => n186, ZN => n183);
   U72 : AOI222_X1 port map( A1 => n165, A2 => n178, B1 => n167, B2 => n186, C1
                           => n169, C2 => n184, ZN => n239);
   U73 : AOI222_X1 port map( A1 => n169, A2 => n168, B1 => n493, B2 => n128, C1
                           => n167, C2 => n355, ZN => n534);
   U74 : AOI222_X1 port map( A1 => n169, A2 => n402, B1 => n493, B2 => n133, C1
                           => n167, C2 => n403, ZN => n520);
   U75 : AOI222_X1 port map( A1 => n169, A2 => n453, B1 => n493, B2 => n382, C1
                           => n167, C2 => n506, ZN => n507);
   U76 : OAI222_X1 port map( A1 => n637, A2 => n74, B1 => n635, B2 => n100, C1 
                           => n644, C2 => n196, ZN => n200);
   U77 : INV_X1 port map( A => n260, ZN => n645);
   U78 : NOR2_X1 port map( A1 => n647, A2 => B(4), ZN => n488);
   U79 : INV_X1 port map( A => n262, ZN => n638);
   U80 : OAI222_X1 port map( A1 => n132, A2 => n14, B1 => n27, B2 => n614, C1 
                           => n1, C2 => n102, ZN => n602);
   U81 : OAI221_X1 port map( B1 => n363, B2 => n638, C1 => n61, C2 => n642, A 
                           => n522, ZN => n314);
   U82 : AOI22_X1 port map( A1 => n454, A2 => n57, B1 => n260, B2 => n420, ZN 
                           => n522);
   U83 : OAI221_X1 port map( B1 => n405, B2 => n638, C1 => n72, C2 => n642, A 
                           => n509, ZN => n290);
   U84 : AOI22_X1 port map( A1 => n454, A2 => n51, B1 => n260, B2 => n407, ZN 
                           => n509);
   U85 : OAI221_X1 port map( B1 => n387, B2 => n638, C1 => n75, C2 => n642, A 
                           => n496, ZN => n271);
   U86 : AOI22_X1 port map( A1 => n454, A2 => n390, B1 => n260, B2 => n389, ZN 
                           => n496);
   U87 : INV_X1 port map( A => n228, ZN => n625);
   U88 : OAI21_X1 port map( B1 => n612, B2 => n630, A => n486, ZN => n253);
   U89 : AOI221_X1 port map( B1 => n199, B2 => n361, C1 => B(4), C2 => n55, A 
                           => n418, ZN => n409);
   U90 : INV_X1 port map( A => n214, ZN => n55);
   U91 : OAI222_X1 port map( A1 => n61, A2 => n644, B1 => n363, B2 => n635, C1 
                           => n81, C2 => n637, ZN => n418);
   U92 : AOI221_X1 port map( B1 => n199, B2 => n350, C1 => B(4), C2 => n49, A 
                           => n404, ZN => n392);
   U93 : INV_X1 port map( A => n202, ZN => n49);
   U94 : OAI222_X1 port map( A1 => n72, A2 => n644, B1 => n405, B2 => n635, C1 
                           => n84, C2 => n637, ZN => n404);
   U95 : AOI221_X1 port map( B1 => n199, B2 => n339, C1 => B(4), C2 => n47, A 
                           => n386, ZN => n378);
   U96 : INV_X1 port map( A => n188, ZN => n47);
   U97 : OAI222_X1 port map( A1 => n75, A2 => n644, B1 => n387, B2 => n635, C1 
                           => n86, C2 => n637, ZN => n386);
   U98 : AOI221_X1 port map( B1 => n199, B2 => n324, C1 => n38, C2 => n172, A 
                           => n371, ZN => n365);
   U99 : OAI222_X1 port map( A1 => n78, A2 => n644, B1 => n62, B2 => n635, C1 
                           => n90, C2 => n637, ZN => n371);
   U100 : AOI221_X1 port map( B1 => n199, B2 => n313, C1 => n38, C2 => n139, A 
                           => n360, ZN => n352);
   U101 : OAI222_X1 port map( A1 => n81, A2 => n644, B1 => n61, B2 => n635, C1 
                           => n94, C2 => n637, ZN => n360);
   U102 : AOI221_X1 port map( B1 => n199, B2 => n289, C1 => n38, C2 => n348, A 
                           => n349, ZN => n341);
   U103 : OAI222_X1 port map( A1 => n84, A2 => n644, B1 => n72, B2 => n635, C1 
                           => n98, C2 => n637, ZN => n349);
   U104 : AOI221_X1 port map( B1 => n199, B2 => n270, C1 => n38, C2 => n337, A 
                           => n338, ZN => n328);
   U105 : OAI222_X1 port map( A1 => n86, A2 => n644, B1 => n75, B2 => n635, C1 
                           => n103, C2 => n637, ZN => n338);
   U106 : NOR2_X1 port map( A1 => n612, A2 => n646, ZN => n359);
   U107 : AOI221_X1 port map( B1 => n276, B2 => n479, C1 => n627, C2 => n480, A
                           => n279, ZN => n478);
   U108 : OAI21_X1 port map( B1 => n482, B2 => n281, A => n282, ZN => n479);
   U109 : AOI21_X1 port map( B1 => n283, B2 => n485, A => n285, ZN => n482);
   U110 : OAI21_X1 port map( B1 => n88, B2 => n287, A => n288, ZN => n485);
   U111 : AOI221_X1 port map( B1 => n276, B2 => n470, C1 => n627, C2 => n434, A
                           => n279, ZN => n469);
   U112 : OAI21_X1 port map( B1 => n472, B2 => n281, A => n282, ZN => n470);
   U113 : AOI21_X1 port map( B1 => n283, B2 => n473, A => n285, ZN => n472);
   U114 : OAI21_X1 port map( B1 => n93, B2 => n287, A => n288, ZN => n473);
   U115 : AOI221_X1 port map( B1 => n276, B2 => n460, C1 => n627, C2 => n297, A
                           => n279, ZN => n459);
   U116 : OAI21_X1 port map( B1 => n462, B2 => n281, A => n282, ZN => n460);
   U117 : AOI21_X1 port map( B1 => n283, B2 => n463, A => n285, ZN => n462);
   U118 : OAI21_X1 port map( B1 => n97, B2 => n287, A => n288, ZN => n463);
   U119 : AOI221_X1 port map( B1 => n276, B2 => n448, C1 => n627, C2 => n246, A
                           => n279, ZN => n447);
   U120 : OAI21_X1 port map( B1 => n450, B2 => n281, A => n282, ZN => n448);
   U121 : AOI21_X1 port map( B1 => n283, B2 => n451, A => n285, ZN => n450);
   U122 : OAI21_X1 port map( B1 => n101, B2 => n287, A => n288, ZN => n451);
   U123 : AOI221_X1 port map( B1 => n276, B2 => n424, C1 => n627, C2 => n106, A
                           => n279, ZN => n423);
   U124 : INV_X1 port map( A => n238, ZN => n106);
   U125 : OAI21_X1 port map( B1 => n425, B2 => n281, A => n282, ZN => n424);
   U126 : AOI21_X1 port map( B1 => n283, B2 => n426, A => n285, ZN => n425);
   U127 : AOI221_X1 port map( B1 => n276, B2 => n411, C1 => n627, C2 => n223, A
                           => n279, ZN => n410);
   U128 : OAI21_X1 port map( B1 => n414, B2 => n281, A => n282, ZN => n411);
   U129 : AOI21_X1 port map( B1 => n283, B2 => n415, A => n285, ZN => n414);
   U130 : OAI21_X1 port map( B1 => n109, B2 => n287, A => n288, ZN => n415);
   U131 : AOI221_X1 port map( B1 => n276, B2 => n394, C1 => n627, C2 => n211, A
                           => n279, ZN => n393);
   U132 : OAI21_X1 port map( B1 => n397, B2 => n281, A => n282, ZN => n394);
   U133 : AOI21_X1 port map( B1 => n283, B2 => n398, A => n285, ZN => n397);
   U134 : OAI21_X1 port map( B1 => n112, B2 => n287, A => n288, ZN => n398);
   U135 : AOI221_X1 port map( B1 => n276, B2 => n380, C1 => n627, C2 => n114, A
                           => n279, ZN => n379);
   U136 : OAI21_X1 port map( B1 => n384, B2 => n281, A => n282, ZN => n380);
   U137 : AOI21_X1 port map( B1 => n283, B2 => n385, A => n285, ZN => n384);
   U138 : OAI21_X1 port map( B1 => n197, B2 => n287, A => n288, ZN => n385);
   U139 : AOI221_X1 port map( B1 => n276, B2 => n367, C1 => n627, C2 => n118, A
                           => n279, ZN => n366);
   U140 : OAI21_X1 port map( B1 => n368, B2 => n281, A => n282, ZN => n367);
   U141 : AOI21_X1 port map( B1 => n283, B2 => n369, A => n285, ZN => n368);
   U142 : OAI21_X1 port map( B1 => n181, B2 => n287, A => n288, ZN => n369);
   U143 : AOI221_X1 port map( B1 => n276, B2 => n354, C1 => n627, C2 => n121, A
                           => n279, ZN => n353);
   U144 : INV_X1 port map( A => n163, ZN => n121);
   U145 : OAI21_X1 port map( B1 => n357, B2 => n281, A => n282, ZN => n354);
   U146 : AOI21_X1 port map( B1 => n283, B2 => n358, A => n285, ZN => n357);
   U147 : AOI221_X1 port map( B1 => n276, B2 => n343, C1 => n627, C2 => n124, A
                           => n279, ZN => n342);
   U148 : INV_X1 port map( A => n344, ZN => n124);
   U149 : OAI21_X1 port map( B1 => n345, B2 => n281, A => n282, ZN => n343);
   U150 : AOI21_X1 port map( B1 => n283, B2 => n346, A => n285, ZN => n345);
   U151 : NOR2_X1 port map( A1 => n612, A2 => n2, ZN => n519);
   U152 : AOI221_X1 port map( B1 => n165, B2 => n429, C1 => n199, C2 => n373, A
                           => n492, ZN => n477);
   U153 : OAI222_X1 port map( A1 => n374, A2 => n635, B1 => n375, B2 => n640, 
                           C1 => n376, C2 => n644, ZN => n492);
   U154 : AOI221_X1 port map( B1 => n165, B2 => n474, C1 => n199, C2 => n419, A
                           => n475, ZN => n468);
   U155 : OAI222_X1 port map( A1 => n131, A2 => n635, B1 => n362, B2 => n640, 
                           C1 => n363, C2 => n644, ZN => n475);
   U156 : AOI221_X1 port map( B1 => n165, B2 => n465, C1 => n199, C2 => n406, A
                           => n466, ZN => n458);
   U157 : OAI222_X1 port map( A1 => n613, A2 => n635, B1 => n293, B2 => n640, 
                           C1 => n405, C2 => n644, ZN => n466);
   U158 : AOI221_X1 port map( B1 => n165, B2 => n455, C1 => n199, C2 => n388, A
                           => n456, ZN => n446);
   U159 : OAI222_X1 port map( A1 => n615, A2 => n635, B1 => n45, B2 => n640, C1
                           => n387, C2 => n644, ZN => n456);
   U160 : AOI221_X1 port map( B1 => n165, B2 => n373, C1 => n199, C2 => n372, A
                           => n427, ZN => n422);
   U161 : OAI221_X1 port map( B1 => n376, B2 => n635, C1 => n62, C2 => n644, A 
                           => n428, ZN => n427);
   U162 : OAI22_X1 port map( A1 => n8, A2 => n130, B1 => n1, B2 => n135, ZN => 
                           n533);
   U163 : NOR2_X1 port map( A1 => n612, A2 => n8, ZN => n382);
   U164 : OAI221_X1 port map( B1 => n109, B2 => n160, C1 => n92, C2 => n161, A 
                           => n162, ZN => n220);
   U165 : OAI221_X1 port map( B1 => n112, B2 => n160, C1 => n96, C2 => n161, A 
                           => n162, ZN => n208);
   U166 : OAI221_X1 port map( B1 => n197, B2 => n160, C1 => n100, C2 => n161, A
                           => n162, ZN => n194);
   U167 : AOI22_X1 port map( A1 => n480, A2 => n38, B1 => n42, B2 => n63, ZN =>
                           n587);
   U168 : INV_X1 port map( A => n601, ZN => n63);
   U169 : AOI221_X1 port map( B1 => n4, B2 => n602, C1 => n454, C2 => n184, A 
                           => n603, ZN => n601);
   U170 : OAI22_X1 port map( A1 => n617, A2 => n638, B1 => n64, B2 => n645, ZN 
                           => n603);
   U171 : AOI22_X1 port map( A1 => n420, A2 => n2, B1 => n57, B2 => n262, ZN =>
                           n214);
   U172 : AOI22_X1 port map( A1 => n407, A2 => n5, B1 => n51, B2 => n262, ZN =>
                           n202);
   U173 : AOI22_X1 port map( A1 => n389, A2 => n3, B1 => n390, B2 => n262, ZN 
                           => n188);
   U174 : AOI22_X1 port map( A1 => n452, A2 => n4, B1 => n453, B2 => n262, ZN 
                           => n449);
   U175 : AOI22_X1 port map( A1 => n168, A2 => n3, B1 => n355, B2 => n262, ZN 
                           => n413);
   U176 : AOI22_X1 port map( A1 => n402, A2 => n5, B1 => n403, B2 => n262, ZN 
                           => n396);
   U177 : AOI22_X1 port map( A1 => n370, A2 => n4, B1 => n320, B2 => n262, ZN 
                           => n182);
   U178 : AOI22_X1 port map( A1 => n355, A2 => n2, B1 => n128, B2 => n262, ZN 
                           => n163);
   U179 : AOI22_X1 port map( A1 => n403, A2 => n4, B1 => n133, B2 => n262, ZN 
                           => n344);
   U180 : AOI21_X1 port map( B1 => n148, B2 => n217, A => n150, ZN => n216);
   U181 : OAI21_X1 port map( B1 => n218, B2 => n152, A => n153, ZN => n217);
   U182 : AOI211_X1 port map( C1 => n643, C2 => n219, A => n220, B => n221, ZN 
                           => n218);
   U183 : OAI22_X1 port map( A1 => n70, A2 => n157, B1 => n80, B2 => n158, ZN 
                           => n221);
   U184 : AOI21_X1 port map( B1 => n148, B2 => n205, A => n150, ZN => n204);
   U185 : OAI21_X1 port map( B1 => n206, B2 => n152, A => n153, ZN => n205);
   U186 : AOI211_X1 port map( C1 => n643, C2 => n207, A => n208, B => n209, ZN 
                           => n206);
   U187 : OAI22_X1 port map( A1 => n67, A2 => n157, B1 => n83, B2 => n158, ZN 
                           => n209);
   U188 : AOI21_X1 port map( B1 => n148, B2 => n191, A => n150, ZN => n190);
   U189 : OAI21_X1 port map( B1 => n192, B2 => n152, A => n153, ZN => n191);
   U190 : AOI211_X1 port map( C1 => n643, C2 => n193, A => n194, B => n195, ZN 
                           => n192);
   U191 : OAI22_X1 port map( A1 => n74, A2 => n157, B1 => n196, B2 => n158, ZN 
                           => n195);
   U192 : OAI211_X1 port map( C1 => n126, C2 => n645, A => n401, B => n449, ZN 
                           => n257);
   U193 : AOI21_X1 port map( B1 => n320, B2 => n4, A => n519, ZN => n323);
   U194 : AOI21_X1 port map( B1 => n506, B2 => n5, A => n519, ZN => n336);
   U195 : NAND2_X1 port map( A1 => n484, A2 => n632, ZN => n249);
   U196 : OAI21_X1 port map( B1 => n417, B2 => n636, A => n471, ZN => n440);
   U197 : OAI21_X1 port map( B1 => n400, B2 => n636, A => n461, ZN => n302);
   U198 : OAI21_X1 port map( B1 => n412, B2 => n636, A => n471, ZN => n434);
   U199 : OAI21_X1 port map( B1 => n395, B2 => n636, A => n461, ZN => n297);
   U200 : OAI21_X1 port map( B1 => n412, B2 => n645, A => n413, ZN => n223);
   U201 : OAI21_X1 port map( B1 => n395, B2 => n645, A => n396, ZN => n211);
   U202 : OAI21_X1 port map( B1 => n333, B2 => n646, A => n449, ZN => n246);
   U203 : NOR2_X1 port map( A1 => n612, A2 => n484, ZN => n483);
   U204 : OAI21_X1 port map( B1 => n237, B2 => n287, A => n288, ZN => n426);
   U205 : OAI21_X1 port map( B1 => n159, B2 => n287, A => n288, ZN => n358);
   U206 : OAI21_X1 port map( B1 => n347, B2 => n287, A => n288, ZN => n346);
   U207 : OAI21_X1 port map( B1 => n336, B2 => n287, A => n288, ZN => n335);
   U208 : BUF_X1 port map( A => n137, Z => n35);
   U209 : BUF_X1 port map( A => n137, Z => n36);
   U210 : OAI21_X1 port map( B1 => n233, B2 => n152, A => n153, ZN => n232);
   U211 : AOI211_X1 port map( C1 => n643, C2 => n234, A => n235, B => n236, ZN 
                           => n233);
   U212 : OAI22_X1 port map( A1 => n64, A2 => n157, B1 => n77, B2 => n158, ZN 
                           => n236);
   U213 : OAI221_X1 port map( B1 => n237, B2 => n160, C1 => n89, C2 => n161, A 
                           => n162, ZN => n235);
   U214 : OAI21_X1 port map( B1 => n177, B2 => n152, A => n153, ZN => n176);
   U215 : AOI211_X1 port map( C1 => n643, C2 => n178, A => n179, B => n180, ZN 
                           => n177);
   U216 : OAI22_X1 port map( A1 => n77, A2 => n157, B1 => n89, B2 => n158, ZN 
                           => n180);
   U217 : OAI221_X1 port map( B1 => n181, B2 => n160, C1 => n105, C2 => n161, A
                           => n162, ZN => n179);
   U218 : OAI21_X1 port map( B1 => n151, B2 => n152, A => n153, ZN => n149);
   U219 : AOI211_X1 port map( C1 => n643, C2 => n154, A => n155, B => n156, ZN 
                           => n151);
   U220 : OAI22_X1 port map( A1 => n80, A2 => n157, B1 => n92, B2 => n158, ZN 
                           => n156);
   U221 : OAI221_X1 port map( B1 => n159, B2 => n160, C1 => n108, C2 => n161, A
                           => n162, ZN => n155);
   U222 : OAI21_X1 port map( B1 => n576, B2 => n152, A => n153, ZN => n575);
   U223 : AOI211_X1 port map( C1 => n643, C2 => n305, A => n577, B => n578, ZN 
                           => n576);
   U224 : OAI22_X1 port map( A1 => n83, A2 => n157, B1 => n96, B2 => n158, ZN 
                           => n578);
   U225 : OAI221_X1 port map( B1 => n347, B2 => n160, C1 => n111, C2 => n161, A
                           => n162, ZN => n577);
   U226 : OAI21_X1 port map( B1 => n559, B2 => n152, A => n153, ZN => n558);
   U227 : AOI211_X1 port map( C1 => n643, C2 => n261, A => n560, B => n561, ZN 
                           => n559);
   U228 : OAI22_X1 port map( A1 => n196, A2 => n157, B1 => n100, B2 => n158, ZN
                           => n561);
   U229 : OAI221_X1 port map( B1 => n336, B2 => n160, C1 => n115, C2 => n161, A
                           => n162, ZN => n560);
   U230 : OAI21_X1 port map( B1 => n547, B2 => n152, A => n153, ZN => n546);
   U231 : AOI211_X1 port map( C1 => n643, C2 => n184, A => n548, B => n549, ZN 
                           => n547);
   U232 : OAI22_X1 port map( A1 => n89, A2 => n157, B1 => n105, B2 => n158, ZN 
                           => n549);
   U233 : OAI221_X1 port map( B1 => n323, B2 => n160, C1 => n117, C2 => n161, A
                           => n162, ZN => n548);
   U234 : OAI21_X1 port map( B1 => n530, B2 => n152, A => n153, ZN => n529);
   U235 : AOI211_X1 port map( C1 => n643, C2 => n166, A => n531, B => n532, ZN 
                           => n530);
   U236 : OAI22_X1 port map( A1 => n92, A2 => n157, B1 => n108, B2 => n158, ZN 
                           => n532);
   U237 : OAI221_X1 port map( B1 => n312, B2 => n160, C1 => n120, C2 => n161, A
                           => n162, ZN => n531);
   U238 : OAI21_X1 port map( B1 => n515, B2 => n152, A => n153, ZN => n514);
   U239 : AOI211_X1 port map( C1 => n643, C2 => n516, A => n517, B => n518, ZN 
                           => n515);
   U240 : OAI22_X1 port map( A1 => n96, A2 => n157, B1 => n111, B2 => n158, ZN 
                           => n518);
   U241 : OAI221_X1 port map( B1 => n286, B2 => n160, C1 => n123, C2 => n161, A
                           => n162, ZN => n517);
   U242 : INV_X1 port map( A => n452, ZN => n100);
   U243 : INV_X1 port map( A => n170, ZN => n92);
   U244 : INV_X1 port map( A => n464, ZN => n96);
   U245 : INV_X1 port map( A => n186, ZN => n89);
   U246 : INV_X1 port map( A => n166, ZN => n80);
   U247 : INV_X1 port map( A => n516, ZN => n83);
   U248 : NOR2_X1 port map( A1 => n135, A2 => n8, ZN => n580);
   U249 : OAI21_X1 port map( B1 => n587, B2 => n255, A => n256, ZN => n595);
   U250 : AOI21_X1 port map( B1 => n251, B2 => n438, A => n253, ZN => n437);
   U251 : OAI21_X1 port map( B1 => n439, B2 => n255, A => n256, ZN => n438);
   U252 : AOI22_X1 port map( A1 => n435, A2 => n39, B1 => B(4), B2 => n440, ZN 
                           => n439);
   U253 : AOI21_X1 port map( B1 => n251, B2 => n300, A => n253, ZN => n299);
   U254 : OAI21_X1 port map( B1 => n301, B2 => n255, A => n256, ZN => n300);
   U255 : AOI22_X1 port map( A1 => n298, A2 => n39, B1 => B(4), B2 => n302, ZN 
                           => n301);
   U256 : AOI21_X1 port map( B1 => n251, B2 => n252, A => n253, ZN => n248);
   U257 : OAI21_X1 port map( B1 => n254, B2 => n255, A => n256, ZN => n252);
   U258 : AOI22_X1 port map( A1 => n247, A2 => n39, B1 => B(4), B2 => n257, ZN 
                           => n254);
   U259 : BUF_X1 port map( A => n356, Z => n2);
   U260 : BUF_X1 port map( A => n356, Z => n3);
   U261 : INV_X1 port map( A => n293, ZN => n51);
   U262 : INV_X1 port map( A => n184, ZN => n77);
   U263 : INV_X1 port map( A => n506, ZN => n126);
   U265 : INV_X1 port map( A => n185, ZN => n105);
   U266 : INV_X1 port map( A => n390, ZN => n45);
   U268 : BUF_X1 port map( A => n356, Z => n4);
   U270 : BUF_X1 port map( A => n356, Z => n5);
   U271 : INV_X1 port map( A => n453, ZN => n115);
   U272 : INV_X1 port map( A => n412, ZN => n128);
   U273 : INV_X1 port map( A => n395, ZN => n133);
   U274 : INV_X1 port map( A => n154, ZN => n70);
   U275 : INV_X1 port map( A => n305, ZN => n67);
   U276 : INV_X1 port map( A => n178, ZN => n64);
   U277 : INV_X1 port map( A => n168, ZN => n108);
   U278 : INV_X1 port map( A => n402, ZN => n111);
   U279 : INV_X1 port map( A => n261, ZN => n74);
   U280 : INV_X1 port map( A => n419, ZN => n81);
   U281 : INV_X1 port map( A => n406, ZN => n84);
   U282 : INV_X1 port map( A => n388, ZN => n86);
   U283 : BUF_X1 port map( A => n43, Z => n41);
   U284 : INV_X1 port map( A => n362, ZN => n57);
   U285 : INV_X1 port map( A => n474, ZN => n61);
   U286 : INV_X1 port map( A => n465, ZN => n72);
   U287 : INV_X1 port map( A => n455, ZN => n75);
   U288 : INV_X1 port map( A => n267, ZN => n8);
   U289 : INV_X1 port map( A => n355, ZN => n120);
   U290 : INV_X1 port map( A => n403, ZN => n123);
   U291 : BUF_X1 port map( A => n43, Z => n42);
   U292 : BUF_X1 port map( A => n43, Z => n39);
   U293 : BUF_X1 port map( A => n43, Z => n40);
   U294 : INV_X1 port map( A => n370, ZN => n117);
   U295 : INV_X1 port map( A => n373, ZN => n78);
   U296 : INV_X1 port map( A => n420, ZN => n131);
   U297 : INV_X1 port map( A => n407, ZN => n613);
   U298 : INV_X1 port map( A => n389, ZN => n615);
   U299 : INV_X1 port map( A => n417, ZN => n129);
   U300 : INV_X1 port map( A => n400, ZN => n134);
   U301 : INV_X1 port map( A => n429, ZN => n62);
   U302 : INV_X1 port map( A => n372, ZN => n90);
   U303 : INV_X1 port map( A => n361, ZN => n94);
   U304 : INV_X1 port map( A => n350, ZN => n98);
   U305 : INV_X1 port map( A => n339, ZN => n103);
   U306 : AND2_X1 port map( A1 => n238, A2 => n401, ZN => n237);
   U307 : INV_X1 port map( A => n234, ZN => n617);
   U308 : INV_X1 port map( A => n416, ZN => n109);
   U309 : OAI211_X1 port map( C1 => n417, C2 => n645, A => n401, B => n413, ZN 
                           => n416);
   U310 : INV_X1 port map( A => n399, ZN => n112);
   U311 : OAI211_X1 port map( C1 => n400, C2 => n645, A => n401, B => n396, ZN 
                           => n399);
   U312 : INV_X1 port map( A => n381, ZN => n114);
   U313 : AOI21_X1 port map( B1 => n260, B2 => n382, A => n383, ZN => n381);
   U314 : BUF_X1 port map( A => n137, Z => n37);
   U315 : OR4_X1 port map( A1 => B(21), A2 => B(20), A3 => B(19), A4 => B(18), 
                           ZN => n598);
   U316 : OAI22_X1 port map( A1 => n87, A2 => n1, B1 => n85, B2 => n8, ZN => 
                           n568);
   U317 : OAI22_X1 port map( A1 => n622, A2 => n1, B1 => n623, B2 => n8, ZN => 
                           n525);
   U318 : OAI22_X1 port map( A1 => n623, A2 => n1, B1 => n65, B2 => n8, ZN => 
                           n570);
   U319 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n73, B2 => n8, ZN => 
                           n552);
   U320 : AOI221_X1 port map( B1 => n31, B2 => A(5), C1 => n20, C2 => A(6), A 
                           => n541, ZN => n376);
   U321 : OAI22_X1 port map( A1 => n621, A2 => n1, B1 => n622, B2 => n8, ZN => 
                           n541);
   U322 : OAI221_X1 port map( B1 => n27, B2 => n612, C1 => n17, C2 => n135, A 
                           => n609, ZN => n320);
   U323 : AOI22_X1 port map( A1 => A(29), A2 => n10, B1 => A(28), B2 => n7, ZN 
                           => n609);
   U324 : OAI221_X1 port map( B1 => n25, B2 => n127, C1 => n15, C2 => n125, A 
                           => n535, ZN => n355);
   U325 : AOI22_X1 port map( A1 => A(26), A2 => n9, B1 => A(25), B2 => n267, ZN
                           => n535);
   U326 : OAI221_X1 port map( B1 => n26, B2 => n130, C1 => n16, C2 => n127, A 
                           => n585, ZN => n403);
   U327 : AOI22_X1 port map( A1 => A(27), A2 => n10, B1 => A(26), B2 => n7, ZN 
                           => n585);
   U328 : OR3_X1 port map( A1 => B(22), A2 => B(24), A3 => B(23), ZN => n594);
   U329 : NAND3_X1 port map( A1 => n489, A2 => n628, A3 => n600, ZN => n152);
   U330 : NOR3_X1 port map( A1 => B(12), A2 => B(14), A3 => B(13), ZN => n600);
   U331 : NAND3_X1 port map( A1 => n592, A2 => n631, A3 => n599, ZN => n146);
   U332 : INV_X1 port map( A => B(22), ZN => n631);
   U333 : NOR3_X1 port map( A1 => B(23), A2 => B(25), A3 => B(24), ZN => n599);
   U334 : OAI221_X1 port map( B1 => n27, B2 => n85, C1 => n17, C2 => n82, A => 
                           n606, ZN => n184);
   U335 : AOI22_X1 port map( A1 => A(13), A2 => n11, B1 => A(12), B2 => n7, ZN 
                           => n606);
   U336 : OAI221_X1 port map( B1 => n27, B2 => n125, C1 => n17, C2 => n122, A 
                           => n608, ZN => n370);
   U337 : AOI22_X1 port map( A1 => A(25), A2 => n9, B1 => A(24), B2 => n7, ZN 
                           => n608);
   U338 : NAND2_X1 port map( A1 => n488, A2 => n489, ZN => n287);
   U339 : OAI221_X1 port map( B1 => n25, B2 => n116, C1 => n15, C2 => n113, A 
                           => n536, ZN => n168);
   U340 : AOI22_X1 port map( A1 => A(22), A2 => n9, B1 => A(21), B2 => n267, ZN
                           => n536);
   U341 : OAI221_X1 port map( B1 => n26, B2 => n119, C1 => n16, C2 => n116, A 
                           => n583, ZN => n402);
   U342 : AOI22_X1 port map( A1 => A(23), A2 => n10, B1 => A(22), B2 => n7, ZN 
                           => n583);
   U343 : NOR2_X2 port map( A1 => n490, A2 => B(11), ZN => n283);
   U344 : NAND2_X1 port map( A1 => A(31), A2 => n647, ZN => n162);
   U345 : AOI221_X1 port map( B1 => A(1), B2 => n31, C1 => A(2), C2 => n21, A 
                           => n540, ZN => n374);
   U346 : OAI22_X1 port map( A1 => n614, A2 => n1, B1 => n616, B2 => n8, ZN => 
                           n540);
   U347 : NOR2_X2 port map( A1 => n266, A2 => n591, ZN => n144);
   U348 : NAND2_X1 port map( A1 => A(31), A2 => n152, ZN => n153);
   U349 : NAND2_X1 port map( A1 => A(31), A2 => n146, ZN => n147);
   U350 : OAI221_X1 port map( B1 => n26, B2 => n135, C1 => n16, C2 => n130, A 
                           => n564, ZN => n506);
   U351 : AOI22_X1 port map( A1 => A(28), A2 => n10, B1 => A(27), B2 => n6, ZN 
                           => n564);
   U352 : OAI221_X1 port map( B1 => n26, B2 => n122, C1 => n16, C2 => n119, A 
                           => n565, ZN => n453);
   U353 : AOI22_X1 port map( A1 => A(24), A2 => n10, B1 => A(23), B2 => n6, ZN 
                           => n565);
   U354 : NOR2_X2 port map( A1 => n646, A2 => B(2), ZN => n260);
   U355 : OAI221_X1 port map( B1 => n24, B2 => n113, C1 => n14, C2 => n110, A 
                           => n611, ZN => n185);
   U356 : AOI22_X1 port map( A1 => A(21), A2 => n11, B1 => A(20), B2 => n6, ZN 
                           => n611);
   U357 : AOI222_X1 port map( A1 => n429, A2 => n5, B1 => n619, B2 => n262, C1 
                           => n227, C2 => B(3), ZN => n327);
   U358 : INV_X1 port map( A => n376, ZN => n619);
   U359 : OAI221_X1 port map( B1 => n24, B2 => n76, C1 => n15, C2 => n73, A => 
                           n444, ZN => n154);
   U360 : AOI22_X1 port map( A1 => A(10), A2 => n11, B1 => A(9), B2 => n267, ZN
                           => n444);
   U361 : OAI221_X1 port map( B1 => n27, B2 => n79, C1 => n16, C2 => n76, A => 
                           n586, ZN => n305);
   U362 : AOI22_X1 port map( A1 => A(11), A2 => n10, B1 => A(10), B2 => n7, ZN 
                           => n586);
   U363 : OAI221_X1 port map( B1 => n26, B2 => n82, C1 => n16, C2 => n79, A => 
                           n567, ZN => n261);
   U364 : AOI22_X1 port map( A1 => A(12), A2 => n10, B1 => A(11), B2 => n6, ZN 
                           => n567);
   U365 : OAI221_X1 port map( B1 => n24, B2 => n622, C1 => n14, C2 => n621, A 
                           => n443, ZN => n219);
   U366 : AOI22_X1 port map( A1 => A(6), A2 => n11, B1 => A(5), B2 => n267, ZN 
                           => n443);
   U367 : OAI221_X1 port map( B1 => n24, B2 => n623, C1 => n14, C2 => n622, A 
                           => n306, ZN => n207);
   U368 : AOI22_X1 port map( A1 => A(7), A2 => n11, B1 => A(6), B2 => n7, ZN =>
                           n306);
   U369 : OAI221_X1 port map( B1 => n25, B2 => n65, C1 => n15, C2 => n623, A =>
                           n265, ZN => n193);
   U370 : AOI22_X1 port map( A1 => A(8), A2 => n9, B1 => A(7), B2 => n6, ZN => 
                           n265);
   U371 : OAI221_X1 port map( B1 => n27, B2 => n99, C1 => n17, C2 => n95, A => 
                           n610, ZN => n186);
   U372 : AOI22_X1 port map( A1 => A(17), A2 => n11, B1 => A(16), B2 => n7, ZN 
                           => n610);
   U373 : OAI221_X1 port map( B1 => n27, B2 => n73, C1 => n17, C2 => n65, A => 
                           n604, ZN => n178);
   U374 : AOI22_X1 port map( A1 => A(9), A2 => n9, B1 => A(8), B2 => n7, ZN => 
                           n604);
   U375 : OAI221_X1 port map( B1 => n25, B2 => n87, C1 => n15, C2 => n85, A => 
                           n537, ZN => n166);
   U376 : AOI22_X1 port map( A1 => A(14), A2 => n9, B1 => A(13), B2 => n6, ZN 
                           => n537);
   U377 : OAI221_X1 port map( B1 => n26, B2 => n91, C1 => n16, C2 => n87, A => 
                           n584, ZN => n516);
   U378 : AOI22_X1 port map( A1 => A(15), A2 => n10, B1 => A(14), B2 => n6, ZN 
                           => n584);
   U379 : OAI221_X1 port map( B1 => n25, B2 => n79, C1 => n15, C2 => n82, A => 
                           n494, ZN => n373);
   U380 : AOI22_X1 port map( A1 => A(15), A2 => n9, B1 => A(16), B2 => n267, ZN
                           => n494);
   U381 : OAI221_X1 port map( B1 => n25, B2 => n132, C1 => n15, C2 => n614, A 
                           => n523, ZN => n420);
   U382 : AOI22_X1 port map( A1 => A(4), A2 => n9, B1 => A(5), B2 => n267, ZN 
                           => n523);
   U383 : OAI221_X1 port map( B1 => n26, B2 => n614, C1 => n16, C2 => n616, A 
                           => n571, ZN => n407);
   U384 : AOI22_X1 port map( A1 => A(5), A2 => n10, B1 => A(6), B2 => n6, ZN =>
                           n571);
   U385 : OAI221_X1 port map( B1 => n26, B2 => n616, C1 => n16, C2 => n618, A 
                           => n554, ZN => n389);
   U386 : AOI22_X1 port map( A1 => A(6), A2 => n10, B1 => A(7), B2 => n6, ZN =>
                           n554);
   U387 : OAI221_X1 port map( B1 => n48, B2 => n27, C1 => n102, C2 => n14, A =>
                           n553, ZN => n390);
   U389 : AOI22_X1 port map( A1 => A(2), A2 => n10, B1 => A(3), B2 => n6, ZN =>
                           n553);
   U390 : OAI221_X1 port map( B1 => n26, B2 => n623, C1 => n16, C2 => n65, A =>
                           n542, ZN => n429);
   U391 : AOI22_X1 port map( A1 => A(11), A2 => n10, B1 => A(12), B2 => n6, ZN 
                           => n542);
   U392 : OAI221_X1 port map( B1 => n26, B2 => n110, C1 => n16, C2 => n107, A 
                           => n566, ZN => n452);
   U393 : AOI22_X1 port map( A1 => A(20), A2 => n10, B1 => A(19), B2 => n6, ZN 
                           => n566);
   U394 : OAI221_X1 port map( B1 => n26, B2 => n104, C1 => n16, C2 => n99, A =>
                           n538, ZN => n170);
   U395 : AOI22_X1 port map( A1 => A(18), A2 => n10, B1 => A(17), B2 => n6, ZN 
                           => n538);
   U396 : OAI221_X1 port map( B1 => n26, B2 => n107, C1 => n16, C2 => n104, A 
                           => n582, ZN => n464);
   U397 : AOI22_X1 port map( A1 => A(19), A2 => n10, B1 => A(18), B2 => n6, ZN 
                           => n582);
   U398 : AOI22_X1 port map( A1 => n7, A2 => A(1), B1 => n11, B2 => A(0), ZN =>
                           n362);
   U399 : NAND2_X1 port map( A1 => B(4), A2 => n579, ZN => n160);
   U400 : INV_X1 port map( A => A(31), ZN => n612);
   U401 : INV_X1 port map( A => n332, ZN => n627);
   U402 : AOI21_X1 port map( B1 => A(31), B2 => B(11), A => n487, ZN => n256);
   U403 : AOI21_X1 port map( B1 => A(31), B2 => B(25), A => n483, ZN => n250);
   U404 : OAI221_X1 port map( B1 => n24, B2 => n91, C1 => n14, C2 => n95, A => 
                           n430, ZN => n372);
   U405 : AOI22_X1 port map( A1 => A(19), A2 => n11, B1 => A(20), B2 => n7, ZN 
                           => n430);
   U406 : OAI221_X1 port map( B1 => n25, B2 => n82, C1 => n15, C2 => n85, A => 
                           n476, ZN => n419);
   U407 : AOI22_X1 port map( A1 => A(16), A2 => n9, B1 => A(17), B2 => n267, ZN
                           => n476);
   U408 : OAI221_X1 port map( B1 => n25, B2 => n85, C1 => n15, C2 => n87, A => 
                           n467, ZN => n406);
   U409 : AOI22_X1 port map( A1 => A(17), A2 => n9, B1 => A(18), B2 => n267, ZN
                           => n467);
   U410 : OAI221_X1 port map( B1 => n25, B2 => n87, C1 => n15, C2 => n91, A => 
                           n457, ZN => n388);
   U411 : AOI22_X1 port map( A1 => A(18), A2 => n9, B1 => A(19), B2 => n267, ZN
                           => n457);
   U412 : OAI221_X1 port map( B1 => n27, B2 => n621, C1 => n17, C2 => n620, A 
                           => n605, ZN => n234);
   U413 : AOI22_X1 port map( A1 => A(5), A2 => n11, B1 => A(4), B2 => n7, ZN =>
                           n605);
   U414 : OAI221_X1 port map( B1 => n258, B2 => n642, C1 => n196, C2 => n636, A
                           => n259, ZN => n247);
   U415 : AOI22_X1 port map( A1 => n260, A2 => n261, B1 => n262, B2 => n193, ZN
                           => n259);
   U416 : AOI222_X1 port map( A1 => A(4), A2 => n11, B1 => A(6), B2 => n29, C1 
                           => A(5), C2 => n18, ZN => n258);
   U417 : OAI221_X1 port map( B1 => n303, B2 => n642, C1 => n83, C2 => n636, A 
                           => n304, ZN => n298);
   U418 : AOI22_X1 port map( A1 => n260, A2 => n305, B1 => n262, B2 => n207, ZN
                           => n304);
   U419 : AOI222_X1 port map( A1 => A(3), A2 => n11, B1 => A(5), B2 => n28, C1 
                           => A(4), C2 => n19, ZN => n303);
   U420 : OAI221_X1 port map( B1 => n441, B2 => n642, C1 => n80, C2 => n636, A 
                           => n442, ZN => n435);
   U421 : AOI22_X1 port map( A1 => n260, A2 => n154, B1 => n262, B2 => n219, ZN
                           => n442);
   U422 : AOI222_X1 port map( A1 => A(2), A2 => n9, B1 => A(4), B2 => n28, C1 
                           => A(3), C2 => n18, ZN => n441);
   U423 : OAI221_X1 port map( B1 => n24, B2 => n95, C1 => n14, C2 => n99, A => 
                           n421, ZN => n361);
   U424 : AOI22_X1 port map( A1 => A(20), A2 => n11, B1 => A(21), B2 => n6, ZN 
                           => n421);
   U425 : OAI221_X1 port map( B1 => n25, B2 => n65, C1 => n15, C2 => n73, A => 
                           n524, ZN => n474);
   U426 : AOI22_X1 port map( A1 => A(12), A2 => n9, B1 => A(13), B2 => n267, ZN
                           => n524);
   U427 : OAI221_X1 port map( B1 => n24, B2 => n99, C1 => n14, C2 => n104, A =>
                           n408, ZN => n350);
   U429 : AOI22_X1 port map( A1 => A(21), A2 => n9, B1 => A(22), B2 => n7, ZN 
                           => n408);
   U430 : OAI221_X1 port map( B1 => n25, B2 => n73, C1 => n15, C2 => n76, A => 
                           n510, ZN => n465);
   U431 : AOI22_X1 port map( A1 => A(13), A2 => n9, B1 => A(14), B2 => n267, ZN
                           => n510);
   U432 : OAI221_X1 port map( B1 => n24, B2 => n104, C1 => n14, C2 => n107, A 
                           => n391, ZN => n339);
   U433 : AOI22_X1 port map( A1 => A(22), A2 => n10, B1 => A(23), B2 => n6, ZN 
                           => n391);
   U434 : OAI221_X1 port map( B1 => n25, B2 => n76, C1 => n15, C2 => n79, A => 
                           n497, ZN => n455);
   U435 : AOI22_X1 port map( A1 => A(14), A2 => n9, B1 => A(15), B2 => n6, ZN 
                           => n497);
   U436 : OAI221_X1 port map( B1 => n24, B2 => n107, C1 => n14, C2 => n110, A 
                           => n377, ZN => n324);
   U437 : AOI22_X1 port map( A1 => A(23), A2 => n9, B1 => A(24), B2 => n7, ZN 
                           => n377);
   U438 : OAI221_X1 port map( B1 => n24, B2 => n110, C1 => n14, C2 => n113, A 
                           => n364, ZN => n313);
   U439 : AOI22_X1 port map( A1 => A(24), A2 => n11, B1 => A(25), B2 => n6, ZN 
                           => n364);
   U440 : OAI221_X1 port map( B1 => n24, B2 => n113, C1 => n14, C2 => n116, A 
                           => n351, ZN => n289);
   U441 : AOI22_X1 port map( A1 => A(25), A2 => n9, B1 => A(26), B2 => n7, ZN 
                           => n351);
   U442 : OAI221_X1 port map( B1 => n24, B2 => n116, C1 => n14, C2 => n119, A 
                           => n340, ZN => n270);
   U443 : AOI22_X1 port map( A1 => A(26), A2 => n10, B1 => A(27), B2 => n6, ZN 
                           => n340);
   U444 : AOI221_X1 port map( B1 => n169, B2 => n452, C1 => n167, C2 => n453, A
                           => n563, ZN => n562);
   U445 : NOR3_X1 port map( A1 => n40, A2 => B(3), A3 => n333, ZN => n563);
   U446 : AOI221_X1 port map( B1 => n242, B2 => n432, C1 => n626, C2 => n71, A 
                           => n244, ZN => n431);
   U447 : INV_X1 port map( A => n433, ZN => n71);
   U448 : OAI21_X1 port map( B1 => n437, B2 => n249, A => n250, ZN => n432);
   U449 : AOI22_X1 port map( A1 => n434, A2 => n38, B1 => n41, B2 => n435, ZN 
                           => n433);
   U450 : AOI221_X1 port map( B1 => n242, B2 => n295, C1 => n626, C2 => n68, A 
                           => n244, ZN => n294);
   U451 : INV_X1 port map( A => n296, ZN => n68);
   U452 : OAI21_X1 port map( B1 => n299, B2 => n249, A => n250, ZN => n295);
   U453 : AOI22_X1 port map( A1 => n297, A2 => n38, B1 => n41, B2 => n298, ZN 
                           => n296);
   U454 : AOI221_X1 port map( B1 => n242, B2 => n243, C1 => n626, C2 => n59, A 
                           => n244, ZN => n241);
   U455 : INV_X1 port map( A => n245, ZN => n59);
   U456 : OAI21_X1 port map( B1 => n248, B2 => n249, A => n250, ZN => n243);
   U457 : AOI22_X1 port map( A1 => n246, A2 => n38, B1 => n42, B2 => n247, ZN 
                           => n245);
   U458 : AOI22_X1 port map( A1 => n639, A2 => n506, B1 => B(2), B2 => n382, ZN
                           => n333);
   U459 : AOI221_X1 port map( B1 => n276, B2 => n319, C1 => n278, C2 => n320, A
                           => n279, ZN => n318);
   U460 : OAI21_X1 port map( B1 => n321, B2 => n281, A => n282, ZN => n319);
   U462 : AOI21_X1 port map( B1 => n283, B2 => n322, A => n285, ZN => n321);
   U463 : OAI21_X1 port map( B1 => n323, B2 => n287, A => n288, ZN => n322);
   U464 : AOI221_X1 port map( B1 => n276, B2 => n309, C1 => n278, C2 => n128, A
                           => n279, ZN => n308);
   U465 : OAI21_X1 port map( B1 => n310, B2 => n281, A => n282, ZN => n309);
   U466 : AOI21_X1 port map( B1 => n283, B2 => n311, A => n285, ZN => n310);
   U467 : OAI21_X1 port map( B1 => n312, B2 => n287, A => n288, ZN => n311);
   U468 : AOI221_X1 port map( B1 => n276, B2 => n277, C1 => n278, C2 => n133, A
                           => n279, ZN => n275);
   U469 : OAI21_X1 port map( B1 => n280, B2 => n281, A => n282, ZN => n277);
   U470 : AOI21_X1 port map( B1 => n283, B2 => n284, A => n285, ZN => n280);
   U471 : OAI21_X1 port map( B1 => n286, B2 => n287, A => n288, ZN => n284);
   U472 : AOI221_X1 port map( B1 => n165, B2 => n324, C1 => n38, C2 => n53, A 
                           => n325, ZN => n317);
   U473 : INV_X1 port map( A => n327, ZN => n53);
   U474 : OAI222_X1 port map( A1 => n78, A2 => n635, B1 => n326, B2 => n641, C1
                           => n90, C2 => n644, ZN => n325);
   U475 : AOI222_X1 port map( A1 => A(27), A2 => n10, B1 => A(25), B2 => n28, 
                           C1 => A(26), C2 => n19, ZN => n326);
   U476 : AOI221_X1 port map( B1 => n165, B2 => n313, C1 => n38, C2 => n314, A 
                           => n315, ZN => n307);
   U477 : OAI222_X1 port map( A1 => n81, A2 => n635, B1 => n316, B2 => n641, C1
                           => n94, C2 => n644, ZN => n315);
   U478 : AOI222_X1 port map( A1 => A(28), A2 => n11, B1 => A(26), B2 => n28, 
                           C1 => A(27), C2 => n18, ZN => n316);
   U479 : AOI221_X1 port map( B1 => n165, B2 => n289, C1 => n38, C2 => n290, A 
                           => n291, ZN => n274);
   U480 : OAI222_X1 port map( A1 => n84, A2 => n635, B1 => n292, B2 => n641, C1
                           => n98, C2 => n644, ZN => n291);
   U481 : AOI222_X1 port map( A1 => A(29), A2 => n11, B1 => A(27), B2 => n31, 
                           C1 => A(28), C2 => n18, ZN => n292);
   U482 : AOI221_X1 port map( B1 => n165, B2 => n270, C1 => n38, C2 => n271, A 
                           => n272, ZN => n268);
   U483 : OAI222_X1 port map( A1 => n86, A2 => n635, B1 => n273, B2 => n641, C1
                           => n103, C2 => n644, ZN => n272);
   U484 : AOI222_X1 port map( A1 => A(30), A2 => n11, B1 => A(28), B2 => n30, 
                           C1 => A(29), C2 => n20, ZN => n273);
   U485 : NOR2_X1 port map( A1 => n490, A2 => B(18), ZN => n251);
   U486 : OAI22_X1 port map( A1 => B(2), A2 => n374, B1 => n639, B2 => n375, ZN
                           => n227);
   U487 : AOI21_X1 port map( B1 => n20, B2 => A(31), A => n533, ZN => n412);
   U488 : AOI21_X1 port map( B1 => n11, B2 => A(31), A => n580, ZN => n395);
   U489 : AOI21_X1 port map( B1 => B(1), B2 => A(31), A => n533, ZN => n417);
   U490 : AOI21_X1 port map( B1 => n8, B2 => A(31), A => n580, ZN => n400);
   U491 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n267);
   U492 : AOI211_X1 port map( C1 => n276, C2 => n330, A => n279, B => n331, ZN 
                           => n329);
   U493 : OAI21_X1 port map( B1 => n334, B2 => n281, A => n282, ZN => n330);
   U494 : NOR3_X1 port map( A1 => n332, A2 => B(3), A3 => n333, ZN => n331);
   U495 : AOI21_X1 port map( B1 => n283, B2 => n335, A => n285, ZN => n334);
   U496 : OAI221_X1 port map( B1 => n587, B2 => n436, C1 => n48, C2 => n32, A 
                           => n588, ZN => RES(0));
   U497 : AOI21_X1 port map( B1 => n242, B2 => n589, A => n244, ZN => n588);
   U498 : OAI21_X1 port map( B1 => n593, B2 => n249, A => n250, ZN => n589);
   U499 : AOI21_X1 port map( B1 => n251, B2 => n595, A => n253, ZN => n593);
   U500 : AND2_X1 port map( A1 => n491, A2 => n632, ZN => n276);
   U501 : NAND2_X1 port map( A1 => A(31), A2 => n490, ZN => n486);
   U502 : NOR2_X1 port map( A1 => B(2), A2 => B(3), ZN => n356);
   U503 : INV_X1 port map( A => A(10), ZN => n65);
   U504 : NAND2_X1 port map( A1 => n454, A2 => A(31), ZN => n401);
   U505 : OAI21_X1 port map( B1 => n489, B2 => n612, A => n162, ZN => n487);
   U506 : INV_X1 port map( A => B(3), ZN => n646);
   U507 : INV_X1 port map( A => A(11), ZN => n73);
   U508 : INV_X1 port map( A => A(15), ZN => n85);
   U509 : INV_X1 port map( A => A(16), ZN => n87);
   U510 : INV_X1 port map( A => A(9), ZN => n623);
   U511 : OAI21_X1 port map( B1 => n502, B2 => n152, A => n153, ZN => n501);
   U512 : AOI211_X1 port map( C1 => B(4), C2 => A(31), A => n503, B => n504, ZN
                           => n502);
   U513 : OAI22_X1 port map( A1 => n196, A2 => n505, B1 => n100, B2 => n157, ZN
                           => n504);
   U514 : OAI221_X1 port map( B1 => n126, B2 => n161, C1 => n115, C2 => n158, A
                           => n162, ZN => n503);
   U515 : NAND2_X1 port map( A1 => A(0), A2 => n7, ZN => n375);
   U516 : NOR2_X1 port map( A1 => n269, A2 => n38, ZN => n228);
   U517 : INV_X1 port map( A => A(30), ZN => n135);
   U518 : INV_X1 port map( A => A(12), ZN => n76);
   U519 : INV_X1 port map( A => A(13), ZN => n79);
   U520 : INV_X1 port map( A => A(14), ZN => n82);
   U521 : INV_X1 port map( A => A(19), ZN => n99);
   U522 : INV_X1 port map( A => A(20), ZN => n104);
   U523 : INV_X1 port map( A => A(21), ZN => n107);
   U524 : INV_X1 port map( A => A(22), ZN => n110);
   U525 : INV_X1 port map( A => A(23), ZN => n113);
   U526 : INV_X1 port map( A => A(24), ZN => n116);
   U527 : OR4_X1 port map( A1 => B(13), A2 => B(14), A3 => B(12), A4 => n596, 
                           ZN => n490);
   U528 : OR3_X1 port map( A1 => B(15), A2 => B(17), A3 => B(16), ZN => n596);
   U529 : INV_X1 port map( A => B(2), ZN => n639);
   U530 : INV_X1 port map( A => A(8), ZN => n622);
   U531 : INV_X1 port map( A => A(3), ZN => n614);
   U532 : AND3_X1 port map( A1 => n579, A2 => n591, A3 => n597, ZN => n445);
   U533 : NOR3_X1 port map( A1 => n152, A2 => n146, A3 => n629, ZN => n597);
   U534 : INV_X1 port map( A => n148, ZN => n629);
   U535 : AND2_X1 port map( A1 => n491, A2 => n648, ZN => n242);
   U536 : INV_X1 port map( A => A(17), ZN => n91);
   U537 : INV_X1 port map( A => A(7), ZN => n621);
   U538 : INV_X1 port map( A => A(18), ZN => n95);
   U539 : INV_X1 port map( A => A(25), ZN => n119);
   U540 : INV_X1 port map( A => A(29), ZN => n130);
   U541 : INV_X1 port map( A => B(25), ZN => n632);
   U542 : INV_X1 port map( A => A(4), ZN => n616);
   U543 : INV_X1 port map( A => A(27), ZN => n125);
   U544 : INV_X1 port map( A => A(26), ZN => n122);
   U545 : INV_X1 port map( A => A(6), ZN => n620);
   U546 : INV_X1 port map( A => A(5), ZN => n618);
   U547 : INV_X1 port map( A => A(28), ZN => n127);
   U548 : NAND2_X1 port map( A1 => n34, A2 => n648, ZN => n137);
   U549 : INV_X1 port map( A => A(2), ZN => n132);
   U550 : INV_X1 port map( A => n579, ZN => n647);
   U551 : OR2_X1 port map( A1 => n624, A2 => B(1), ZN => n1);
   U552 : INV_X1 port map( A => n436, ZN => n626);
   U553 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n263);
   U554 : NAND2_X1 port map( A1 => B(1), A2 => n624, ZN => n264);
   U555 : INV_X1 port map( A => A(1), ZN => n102);
   U556 : INV_X1 port map( A => B(11), ZN => n628);
   U557 : INV_X1 port map( A => A(0), ZN => n48);
   U558 : INV_X1 port map( A => B(18), ZN => n630);
   U559 : INV_X1 port map( A => B(0), ZN => n624);
   U560 : INV_X1 port map( A => B(4), ZN => n43);
   U561 : NOR3_X1 port map( A1 => B(9), A2 => B(8), A3 => B(10), ZN => n489);
   U562 : NOR3_X1 port map( A1 => B(7), A2 => B(6), A3 => B(5), ZN => n579);
   U563 : NOR3_X1 port map( A1 => B(28), A2 => B(27), A3 => B(26), ZN => n592);
   U564 : NAND3_X1 port map( A1 => n445, A2 => n34, A3 => LEFT_RIGHT, ZN => 
                           n269);
   U565 : NOR2_X1 port map( A1 => n481, A2 => LEFT_RIGHT, ZN => n244);
   U566 : AOI221_X1 port map( B1 => n140, B2 => n229, C1 => n142, C2 => n230, A
                           => n144, ZN => n225);
   U567 : OAI21_X1 port map( B1 => n231, B2 => n146, A => n147, ZN => n230);
   U568 : OAI221_X1 port map( B1 => n617, B2 => n641, C1 => n238, C2 => n40, A 
                           => n239, ZN => n229);
   U569 : AOI21_X1 port map( B1 => n148, B2 => n232, A => n150, ZN => n231);
   U570 : AOI221_X1 port map( B1 => n140, B2 => n498, C1 => n142, C2 => n499, A
                           => n144, ZN => n495);
   U571 : OAI21_X1 port map( B1 => n500, B2 => n146, A => n147, ZN => n499);
   U572 : OAI221_X1 port map( B1 => n100, B2 => n637, C1 => n196, C2 => n641, A
                           => n507, ZN => n498);
   U573 : AOI21_X1 port map( B1 => n148, B2 => n501, A => n150, ZN => n500);
   U574 : AOI221_X1 port map( B1 => n140, B2 => n69, C1 => n142, C2 => n215, A 
                           => n144, ZN => n213);
   U575 : INV_X1 port map( A => n222, ZN => n69);
   U576 : OAI21_X1 port map( B1 => n216, B2 => n146, A => n147, ZN => n215);
   U577 : AOI221_X1 port map( B1 => n219, B2 => n199, C1 => n223, C2 => n38, A 
                           => n224, ZN => n222);
   U578 : AOI221_X1 port map( B1 => n140, B2 => n66, C1 => n142, C2 => n203, A 
                           => n144, ZN => n201);
   U579 : INV_X1 port map( A => n210, ZN => n66);
   U580 : OAI21_X1 port map( B1 => n204, B2 => n146, A => n147, ZN => n203);
   U581 : AOI221_X1 port map( B1 => n207, B2 => n199, C1 => n211, C2 => n38, A 
                           => n212, ZN => n210);
   U582 : AOI221_X1 port map( B1 => n140, B2 => n60, C1 => n142, C2 => n189, A 
                           => n144, ZN => n187);
   U583 : INV_X1 port map( A => n198, ZN => n60);
   U584 : OAI21_X1 port map( B1 => n190, B2 => n146, A => n147, ZN => n189);
   U585 : AOI221_X1 port map( B1 => n193, B2 => n199, C1 => n114, C2 => n38, A 
                           => n200, ZN => n198);
   U586 : AOI221_X1 port map( B1 => n140, B2 => n173, C1 => n142, C2 => n174, A
                           => n144, ZN => n171);
   U587 : OAI21_X1 port map( B1 => n175, B2 => n146, A => n147, ZN => n174);
   U588 : OAI221_X1 port map( B1 => n64, B2 => n641, C1 => n182, C2 => n40, A 
                           => n183, ZN => n173);
   U589 : AOI21_X1 port map( B1 => n148, B2 => n176, A => n150, ZN => n175);
   U590 : AOI221_X1 port map( B1 => n140, B2 => n141, C1 => n142, C2 => n143, A
                           => n144, ZN => n136);
   U591 : OAI21_X1 port map( B1 => n145, B2 => n146, A => n147, ZN => n143);
   U592 : OAI221_X1 port map( B1 => n70, B2 => n641, C1 => n163, C2 => n41, A 
                           => n164, ZN => n141);
   U593 : AOI21_X1 port map( B1 => n148, B2 => n149, A => n150, ZN => n145);
   U594 : AOI221_X1 port map( B1 => n140, B2 => n572, C1 => n142, C2 => n573, A
                           => n144, ZN => n569);
   U595 : OAI21_X1 port map( B1 => n574, B2 => n146, A => n147, ZN => n573);
   U596 : OAI221_X1 port map( B1 => n67, B2 => n641, C1 => n344, C2 => n41, A 
                           => n581, ZN => n572);
   U597 : AOI21_X1 port map( B1 => n148, B2 => n575, A => n150, ZN => n574);
   U598 : AOI221_X1 port map( B1 => n140, B2 => n555, C1 => n142, C2 => n556, A
                           => n144, ZN => n551);
   U599 : OAI21_X1 port map( B1 => n557, B2 => n146, A => n147, ZN => n556);
   U600 : OAI221_X1 port map( B1 => n196, B2 => n637, C1 => n74, C2 => n641, A 
                           => n562, ZN => n555);
   U601 : AOI21_X1 port map( B1 => n148, B2 => n558, A => n150, ZN => n557);
   U602 : AOI221_X1 port map( B1 => n140, B2 => n543, C1 => n142, C2 => n544, A
                           => n144, ZN => n539);
   U603 : OAI21_X1 port map( B1 => n545, B2 => n146, A => n147, ZN => n544);
   U604 : OAI221_X1 port map( B1 => n89, B2 => n637, C1 => n77, C2 => n641, A 
                           => n550, ZN => n543);
   U605 : AOI21_X1 port map( B1 => n148, B2 => n546, A => n150, ZN => n545);
   U606 : AOI221_X1 port map( B1 => n140, B2 => n526, C1 => n142, C2 => n527, A
                           => n144, ZN => n521);
   U607 : OAI21_X1 port map( B1 => n528, B2 => n146, A => n147, ZN => n527);
   U608 : OAI221_X1 port map( B1 => n92, B2 => n637, C1 => n80, C2 => n641, A 
                           => n534, ZN => n526);
   U609 : AOI21_X1 port map( B1 => n148, B2 => n529, A => n150, ZN => n528);
   U610 : AOI221_X1 port map( B1 => n140, B2 => n511, C1 => n142, C2 => n512, A
                           => n144, ZN => n508);
   U611 : OAI21_X1 port map( B1 => n513, B2 => n146, A => n147, ZN => n512);
   U612 : OAI221_X1 port map( B1 => n96, B2 => n637, C1 => n83, C2 => n641, A 
                           => n520, ZN => n511);
   U613 : AOI21_X1 port map( B1 => n148, B2 => n514, A => n150, ZN => n513);
   U614 : AOI21_X1 port map( B1 => n633, B2 => n590, A => n144, ZN => n481);
   U615 : INV_X1 port map( A => n592, ZN => n633);
   U616 : NOR2_X1 port map( A1 => B(29), A2 => B(30), ZN => n591);
   U617 : INV_X1 port map( A => n590, ZN => n266);
   U618 : AND2_X1 port map( A1 => n140, A2 => n199, ZN => n278);
   U619 : NAND2_X1 port map( A1 => n140, A2 => n39, ZN => n332);
   U620 : NAND2_X1 port map( A1 => n140, A2 => n648, ZN => n436);
   U621 : INV_X1 port map( A => LEFT_RIGHT, ZN => n648);
   U622 : AND2_X1 port map( A1 => n142, A2 => n592, ZN => n491);
   U623 : NOR2_X2 port map( A1 => n634, A2 => LOGIC_ARITH, ZN => n142);
   U624 : INV_X1 port map( A => n591, ZN => n634);
   U625 : AND2_X1 port map( A1 => LOGIC_ARITH, A2 => n445, ZN => n140);
   U626 : NOR2_X1 port map( A1 => n612, A2 => LOGIC_ARITH, ZN => n590);
   U627 : OAI222_X1 port map( A1 => n268, A2 => n269, B1 => LEFT_RIGHT, B2 => 
                           n266, C1 => n612, C2 => n33, ZN => RES(31));
   U628 : OAI222_X1 port map( A1 => n187, A2 => n35, B1 => n188, B2 => n625, C1
                           => n621, C2 => n32, ZN => RES(7));
   U629 : OAI222_X1 port map( A1 => n171, A2 => n35, B1 => n54, B2 => n625, C1 
                           => n622, C2 => n32, ZN => RES(8));
   U630 : OAI222_X1 port map( A1 => n136, A2 => n35, B1 => n58, B2 => n625, C1 
                           => n623, C2 => n32, ZN => RES(9));
   U631 : OAI222_X1 port map( A1 => n551, A2 => n35, B1 => n44, B2 => n625, C1 
                           => n73, C2 => n34, ZN => RES(11));
   U632 : OAI222_X1 port map( A1 => n539, A2 => n35, B1 => n327, B2 => n625, C1
                           => n76, C2 => n34, ZN => RES(12));
   U633 : OAI222_X1 port map( A1 => n521, A2 => n35, B1 => n56, B2 => n625, C1 
                           => n79, C2 => n34, ZN => RES(13));
   U634 : OAI222_X1 port map( A1 => n508, A2 => n35, B1 => n50, B2 => n625, C1 
                           => n82, C2 => n34, ZN => RES(14));
   U635 : OAI222_X1 port map( A1 => n468, A2 => n269, B1 => n469, B2 => n36, C1
                           => n91, C2 => n33, ZN => RES(17));
   U636 : OAI222_X1 port map( A1 => n495, A2 => n35, B1 => n46, B2 => n625, C1 
                           => n85, C2 => n34, ZN => RES(15));
   U640 : OAI222_X1 port map( A1 => n458, A2 => n269, B1 => n459, B2 => n37, C1
                           => n95, C2 => n33, ZN => RES(18));
   U643 : OAI222_X1 port map( A1 => n446, A2 => n269, B1 => n447, B2 => n36, C1
                           => n99, C2 => n33, ZN => RES(19));
   U644 : OAI222_X1 port map( A1 => n422, A2 => n269, B1 => n423, B2 => n36, C1
                           => n104, C2 => n33, ZN => RES(20));
   U645 : OAI222_X1 port map( A1 => n409, A2 => n269, B1 => n410, B2 => n36, C1
                           => n107, C2 => n33, ZN => RES(21));
   U646 : OAI222_X1 port map( A1 => n392, A2 => n269, B1 => n393, B2 => n36, C1
                           => n110, C2 => n33, ZN => RES(22));
   U647 : OAI222_X1 port map( A1 => n378, A2 => n269, B1 => n379, B2 => n36, C1
                           => n113, C2 => n33, ZN => RES(23));
   U648 : OAI222_X1 port map( A1 => n365, A2 => n269, B1 => n366, B2 => n36, C1
                           => n116, C2 => n33, ZN => RES(24));
   U649 : OAI222_X1 port map( A1 => n352, A2 => n269, B1 => n353, B2 => n36, C1
                           => n119, C2 => n33, ZN => RES(25));
   U650 : OAI222_X1 port map( A1 => n213, A2 => n35, B1 => n214, B2 => n625, C1
                           => n618, C2 => n32, ZN => RES(5));
   U651 : OAI222_X1 port map( A1 => n201, A2 => n35, B1 => n202, B2 => n625, C1
                           => n620, C2 => n32, ZN => RES(6));
   U652 : OAI222_X1 port map( A1 => n569, A2 => n35, B1 => n52, B2 => n625, C1 
                           => n65, C2 => n34, ZN => RES(10));
   U653 : OAI222_X1 port map( A1 => n477, A2 => n269, B1 => n478, B2 => n37, C1
                           => n87, C2 => n34, ZN => RES(16));
   U654 : OAI222_X1 port map( A1 => n341, A2 => n269, B1 => n342, B2 => n36, C1
                           => n122, C2 => n33, ZN => RES(26));
   U655 : OAI222_X1 port map( A1 => n328, A2 => n269, B1 => n329, B2 => n36, C1
                           => n125, C2 => n33, ZN => RES(27));
   U656 : OAI222_X1 port map( A1 => n317, A2 => n269, B1 => n318, B2 => n36, C1
                           => n127, C2 => n33, ZN => RES(28));
   U657 : OAI222_X1 port map( A1 => n307, A2 => n269, B1 => n308, B2 => n36, C1
                           => n130, C2 => n32, ZN => RES(29));
   U658 : OAI222_X1 port map( A1 => n274, A2 => n269, B1 => n275, B2 => n37, C1
                           => n135, C2 => n32, ZN => RES(30));
   U659 : OAI221_X1 port map( B1 => n293, B2 => n240, C1 => n132, C2 => n32, A 
                           => n294, ZN => RES(2));
   U660 : OAI221_X1 port map( B1 => n362, B2 => n240, C1 => n102, C2 => n32, A 
                           => n431, ZN => RES(1));
   U661 : OAI221_X1 port map( B1 => n45, B2 => n240, C1 => n614, C2 => n32, A 
                           => n241, ZN => RES(3));
   U662 : OAI221_X1 port map( B1 => n225, B2 => n35, C1 => n616, C2 => n32, A 
                           => n226, ZN => RES(4));
   U663 : NOR4_X4 port map( A1 => B(16), A2 => B(17), A3 => B(15), A4 => n598, 
                           ZN => n148);
   U664 : INV_X1 port map( A => n8, ZN => n6);
   U665 : INV_X1 port map( A => n8, ZN => n7);
   U666 : INV_X1 port map( A => n1, ZN => n9);
   U667 : INV_X1 port map( A => n1, ZN => n10);
   U668 : INV_X1 port map( A => n1, ZN => n11);
   U669 : CLKBUF_X1 port map( A => n264, Z => n12);
   U670 : CLKBUF_X1 port map( A => n264, Z => n13);
   U671 : INV_X1 port map( A => n20, ZN => n17);
   U672 : INV_X1 port map( A => n12, ZN => n18);
   U673 : INV_X1 port map( A => n12, ZN => n19);
   U674 : INV_X1 port map( A => n12, ZN => n20);
   U675 : INV_X1 port map( A => n13, ZN => n21);
   U676 : CLKBUF_X1 port map( A => n263, Z => n22);
   U677 : CLKBUF_X1 port map( A => n263, Z => n23);
   U678 : INV_X1 port map( A => n22, ZN => n28);
   U679 : INV_X1 port map( A => n23, ZN => n29);
   U680 : INV_X1 port map( A => n23, ZN => n30);
   U681 : INV_X1 port map( A => n263, ZN => n31);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity comparator_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  OPSel : in std_logic_vector
         (0 to 2);  RES : out std_logic_vector (31 downto 0));

end comparator_NBIT32;

architecture SYN_bhv of comparator_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component comparator_NBIT32_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   signal X_Logic0_port, N26, N27, N28, N29, N30, N31, n10, n15, n16, n17, n18,
      n19, n20, RES_0_port, n2, n3, n4 : std_logic;

begin
   RES <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, RES_0_port 
      );
   
   X_Logic0_port <= '0';
   n10 <= '0';
   r57 : comparator_NBIT32_DW01_cmp6_0 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), TC => n10, LT => N30, GT => N28,
                           EQ => N26, LE => N31, GE => N29, NE => N27);
   U3 : INV_X1 port map( A => n15, ZN => RES_0_port);
   U4 : AOI21_X1 port map( B1 => n16, B2 => n4, A => n17, ZN => n15);
   U5 : NOR3_X1 port map( A1 => n4, A2 => OPSel(1), A3 => n18, ZN => n17);
   U6 : OAI22_X1 port map( A1 => n19, A2 => n3, B1 => OPSel(1), B2 => n20, ZN 
                           => n16);
   U7 : INV_X1 port map( A => OPSel(1), ZN => n3);
   U8 : AOI22_X1 port map( A1 => N28, A2 => n2, B1 => N29, B2 => OPSel(2), ZN 
                           => n19);
   U9 : INV_X1 port map( A => OPSel(2), ZN => n2);
   U10 : AOI22_X1 port map( A1 => N30, A2 => n2, B1 => OPSel(2), B2 => N31, ZN 
                           => n18);
   U11 : AOI22_X1 port map( A1 => N26, A2 => n2, B1 => N27, B2 => OPSel(2), ZN 
                           => n20);
   U12 : INV_X1 port map( A => OPSel(0), ZN => n4);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_NBIT32 is

   port( OP1, OP2 : in std_logic_vector (31 downto 0);  ALU_OPC : in 
         std_logic_vector (0 to 3);  ALU_RES : out std_logic_vector (31 downto 
         0));

end ALU_NBIT32;

architecture SYN_struct of ALU_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux21_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux41_NBIT32_1
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component P4Adder_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component shifter_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  LOGIC_ARITH, LEFT_RIGHT 
            : in std_logic;  RES : out std_logic_vector (31 downto 0));
   end component;
   
   component comparator_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  OPSel : in 
            std_logic_vector (0 to 2);  RES : out std_logic_vector (31 downto 
            0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, select_type_sig_1_port, select_type_sig_0_port, 
      select_zero_sig, A_SHF_31_port, A_SHF_30_port, A_SHF_29_port, 
      A_SHF_28_port, A_SHF_27_port, A_SHF_26_port, A_SHF_25_port, A_SHF_24_port
      , A_SHF_23_port, A_SHF_22_port, A_SHF_21_port, A_SHF_20_port, 
      A_SHF_19_port, A_SHF_18_port, A_SHF_17_port, A_SHF_16_port, A_SHF_15_port
      , A_SHF_14_port, A_SHF_13_port, A_SHF_12_port, A_SHF_11_port, 
      A_SHF_10_port, A_SHF_9_port, A_SHF_8_port, A_SHF_7_port, A_SHF_6_port, 
      A_SHF_5_port, A_SHF_4_port, A_SHF_3_port, A_SHF_2_port, A_SHF_1_port, 
      A_SHF_0_port, B_SHF_31_port, B_SHF_30_port, B_SHF_29_port, B_SHF_28_port,
      B_SHF_27_port, B_SHF_26_port, B_SHF_25_port, B_SHF_24_port, B_SHF_23_port
      , B_SHF_22_port, B_SHF_21_port, B_SHF_20_port, B_SHF_19_port, 
      B_SHF_18_port, B_SHF_17_port, B_SHF_16_port, B_SHF_15_port, B_SHF_14_port
      , B_SHF_13_port, B_SHF_12_port, B_SHF_11_port, B_SHF_10_port, 
      B_SHF_9_port, B_SHF_8_port, B_SHF_7_port, B_SHF_6_port, B_SHF_5_port, 
      B_SHF_4_port, B_SHF_3_port, B_SHF_2_port, B_SHF_1_port, B_SHF_0_port, 
      A_ADD_31_port, A_ADD_30_port, A_ADD_29_port, A_ADD_28_port, A_ADD_27_port
      , A_ADD_26_port, A_ADD_25_port, A_ADD_24_port, A_ADD_23_port, 
      A_ADD_22_port, A_ADD_21_port, A_ADD_20_port, A_ADD_19_port, A_ADD_18_port
      , A_ADD_17_port, A_ADD_16_port, A_ADD_15_port, A_ADD_14_port, 
      A_ADD_13_port, A_ADD_12_port, A_ADD_11_port, A_ADD_10_port, A_ADD_9_port,
      A_ADD_8_port, A_ADD_7_port, A_ADD_6_port, A_ADD_5_port, A_ADD_4_port, 
      A_ADD_3_port, A_ADD_2_port, A_ADD_1_port, A_ADD_0_port, B_ADD_31_port, 
      B_ADD_30_port, B_ADD_29_port, B_ADD_28_port, B_ADD_27_port, B_ADD_26_port
      , B_ADD_25_port, B_ADD_24_port, B_ADD_23_port, B_ADD_22_port, 
      B_ADD_21_port, B_ADD_20_port, B_ADD_19_port, B_ADD_18_port, B_ADD_17_port
      , B_ADD_16_port, B_ADD_15_port, B_ADD_14_port, B_ADD_13_port, 
      B_ADD_12_port, B_ADD_11_port, B_ADD_10_port, B_ADD_9_port, B_ADD_8_port, 
      B_ADD_7_port, B_ADD_6_port, B_ADD_5_port, B_ADD_4_port, B_ADD_3_port, 
      B_ADD_2_port, B_ADD_1_port, B_ADD_0_port, LOGIC_ARITH, OPSel_0_port, 
      LOGIC_RES_31_port, LOGIC_RES_30_port, LOGIC_RES_29_port, 
      LOGIC_RES_28_port, LOGIC_RES_27_port, LOGIC_RES_26_port, 
      LOGIC_RES_25_port, LOGIC_RES_24_port, LOGIC_RES_23_port, 
      LOGIC_RES_22_port, LOGIC_RES_21_port, LOGIC_RES_20_port, 
      LOGIC_RES_19_port, LOGIC_RES_18_port, LOGIC_RES_17_port, 
      LOGIC_RES_16_port, LOGIC_RES_15_port, LOGIC_RES_14_port, 
      LOGIC_RES_13_port, LOGIC_RES_12_port, LOGIC_RES_11_port, 
      LOGIC_RES_10_port, LOGIC_RES_9_port, LOGIC_RES_8_port, LOGIC_RES_7_port, 
      LOGIC_RES_6_port, LOGIC_RES_5_port, LOGIC_RES_4_port, LOGIC_RES_3_port, 
      LOGIC_RES_2_port, LOGIC_RES_1_port, LOGIC_RES_0_port, COMP_RES_31_port, 
      COMP_RES_30_port, COMP_RES_29_port, COMP_RES_28_port, COMP_RES_27_port, 
      COMP_RES_26_port, COMP_RES_25_port, COMP_RES_24_port, COMP_RES_23_port, 
      COMP_RES_22_port, COMP_RES_21_port, COMP_RES_20_port, COMP_RES_19_port, 
      COMP_RES_18_port, COMP_RES_17_port, COMP_RES_16_port, COMP_RES_15_port, 
      COMP_RES_14_port, COMP_RES_13_port, COMP_RES_12_port, COMP_RES_11_port, 
      COMP_RES_10_port, COMP_RES_9_port, COMP_RES_8_port, COMP_RES_7_port, 
      COMP_RES_6_port, COMP_RES_5_port, COMP_RES_4_port, COMP_RES_3_port, 
      COMP_RES_2_port, COMP_RES_1_port, COMP_RES_0_port, SHIFT_RES_31_port, 
      SHIFT_RES_30_port, SHIFT_RES_29_port, SHIFT_RES_28_port, 
      SHIFT_RES_27_port, SHIFT_RES_26_port, SHIFT_RES_25_port, 
      SHIFT_RES_24_port, SHIFT_RES_23_port, SHIFT_RES_22_port, 
      SHIFT_RES_21_port, SHIFT_RES_20_port, SHIFT_RES_19_port, 
      SHIFT_RES_18_port, SHIFT_RES_17_port, SHIFT_RES_16_port, 
      SHIFT_RES_15_port, SHIFT_RES_14_port, SHIFT_RES_13_port, 
      SHIFT_RES_12_port, SHIFT_RES_11_port, SHIFT_RES_10_port, SHIFT_RES_9_port
      , SHIFT_RES_8_port, SHIFT_RES_7_port, SHIFT_RES_6_port, SHIFT_RES_5_port,
      SHIFT_RES_4_port, SHIFT_RES_3_port, SHIFT_RES_2_port, SHIFT_RES_1_port, 
      SHIFT_RES_0_port, ADD_SUB_RES_31_port, ADD_SUB_RES_30_port, 
      ADD_SUB_RES_29_port, ADD_SUB_RES_28_port, ADD_SUB_RES_27_port, 
      ADD_SUB_RES_26_port, ADD_SUB_RES_25_port, ADD_SUB_RES_24_port, 
      ADD_SUB_RES_23_port, ADD_SUB_RES_22_port, ADD_SUB_RES_21_port, 
      ADD_SUB_RES_20_port, ADD_SUB_RES_19_port, ADD_SUB_RES_18_port, 
      ADD_SUB_RES_17_port, ADD_SUB_RES_16_port, ADD_SUB_RES_15_port, 
      ADD_SUB_RES_14_port, ADD_SUB_RES_13_port, ADD_SUB_RES_12_port, 
      ADD_SUB_RES_11_port, ADD_SUB_RES_10_port, ADD_SUB_RES_9_port, 
      ADD_SUB_RES_8_port, ADD_SUB_RES_7_port, ADD_SUB_RES_6_port, 
      ADD_SUB_RES_5_port, ADD_SUB_RES_4_port, ADD_SUB_RES_3_port, 
      ADD_SUB_RES_2_port, ADD_SUB_RES_1_port, ADD_SUB_RES_0_port, 
      sig_intraMux_31_port, sig_intraMux_30_port, sig_intraMux_29_port, 
      sig_intraMux_28_port, sig_intraMux_27_port, sig_intraMux_26_port, 
      sig_intraMux_25_port, sig_intraMux_24_port, sig_intraMux_23_port, 
      sig_intraMux_22_port, sig_intraMux_21_port, sig_intraMux_20_port, 
      sig_intraMux_19_port, sig_intraMux_18_port, sig_intraMux_17_port, 
      sig_intraMux_16_port, sig_intraMux_15_port, sig_intraMux_14_port, 
      sig_intraMux_13_port, sig_intraMux_12_port, sig_intraMux_11_port, 
      sig_intraMux_10_port, sig_intraMux_9_port, sig_intraMux_8_port, 
      sig_intraMux_7_port, sig_intraMux_6_port, sig_intraMux_5_port, 
      sig_intraMux_4_port, sig_intraMux_3_port, sig_intraMux_2_port, 
      sig_intraMux_1_port, sig_intraMux_0_port, n78, n79, n80, n81, n82, n83, 
      n84, n85, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99
      , n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n1, n2,
      n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n77, n86, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n_1371, n_1372, n_1373, n_1374, 
      n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, 
      n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, 
      n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, 
      n_1402 : std_logic;

begin
   
   X_Logic0_port <= '0';
   U177 : NOR2_X2 port map( A1 => n13, A2 => n55, ZN => A_SHF_31_port);
   U317 : NAND3_X1 port map( A1 => n185, A2 => n184, A3 => n186, ZN => n79);
   U318 : NAND3_X1 port map( A1 => n84, A2 => n83, A3 => n87, ZN => 
                           OPSel_0_port);
   U319 : NAND3_X1 port map( A1 => ALU_OPC(0), A2 => n186, A3 => n88, ZN => n87
                           );
   U320 : NAND3_X1 port map( A1 => ALU_OPC(0), A2 => n186, A3 => n89, ZN => n83
                           );
   U321 : NAND3_X1 port map( A1 => ALU_OPC(0), A2 => ALU_OPC(3), A3 => n89, ZN 
                           => n84);
   U322 : NAND3_X1 port map( A1 => ALU_OPC(1), A2 => ALU_OPC(2), A3 => n155, ZN
                           => n157);
   U323 : NAND3_X1 port map( A1 => ALU_OPC(1), A2 => ALU_OPC(2), A3 => n154, ZN
                           => n85);
   U324 : NAND3_X1 port map( A1 => n185, A2 => n184, A3 => n155, ZN => n156);
   Comp : comparator_NBIT32 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, OPSel(0) => n183, OPSel(1) => n182, 
                           OPSel(2) => OPSel_0_port, RES(31) => n_1371, RES(30)
                           => n_1372, RES(29) => n_1373, RES(28) => n_1374, 
                           RES(27) => n_1375, RES(26) => n_1376, RES(25) => 
                           n_1377, RES(24) => n_1378, RES(23) => n_1379, 
                           RES(22) => n_1380, RES(21) => n_1381, RES(20) => 
                           n_1382, RES(19) => n_1383, RES(18) => n_1384, 
                           RES(17) => n_1385, RES(16) => n_1386, RES(15) => 
                           n_1387, RES(14) => n_1388, RES(13) => n_1389, 
                           RES(12) => n_1390, RES(11) => n_1391, RES(10) => 
                           n_1392, RES(9) => n_1393, RES(8) => n_1394, RES(7) 
                           => n_1395, RES(6) => n_1396, RES(5) => n_1397, 
                           RES(4) => n_1398, RES(3) => n_1399, RES(2) => n_1400
                           , RES(1) => n_1401, RES(0) => COMP_RES_0_port);
   Shift : shifter_NBIT32 port map( A(31) => A_SHF_31_port, A(30) => 
                           A_SHF_30_port, A(29) => A_SHF_29_port, A(28) => 
                           A_SHF_28_port, A(27) => A_SHF_27_port, A(26) => 
                           A_SHF_26_port, A(25) => A_SHF_25_port, A(24) => 
                           A_SHF_24_port, A(23) => A_SHF_23_port, A(22) => 
                           A_SHF_22_port, A(21) => A_SHF_21_port, A(20) => 
                           A_SHF_20_port, A(19) => A_SHF_19_port, A(18) => 
                           A_SHF_18_port, A(17) => A_SHF_17_port, A(16) => 
                           A_SHF_16_port, A(15) => A_SHF_15_port, A(14) => 
                           A_SHF_14_port, A(13) => A_SHF_13_port, A(12) => 
                           A_SHF_12_port, A(11) => A_SHF_11_port, A(10) => 
                           A_SHF_10_port, A(9) => A_SHF_9_port, A(8) => 
                           A_SHF_8_port, A(7) => A_SHF_7_port, A(6) => 
                           A_SHF_6_port, A(5) => A_SHF_5_port, A(4) => 
                           A_SHF_4_port, A(3) => A_SHF_3_port, A(2) => 
                           A_SHF_2_port, A(1) => A_SHF_1_port, A(0) => 
                           A_SHF_0_port, B(31) => B_SHF_31_port, B(30) => 
                           B_SHF_30_port, B(29) => B_SHF_29_port, B(28) => 
                           B_SHF_28_port, B(27) => B_SHF_27_port, B(26) => 
                           B_SHF_26_port, B(25) => B_SHF_25_port, B(24) => 
                           B_SHF_24_port, B(23) => B_SHF_23_port, B(22) => 
                           B_SHF_22_port, B(21) => B_SHF_21_port, B(20) => 
                           B_SHF_20_port, B(19) => B_SHF_19_port, B(18) => 
                           B_SHF_18_port, B(17) => B_SHF_17_port, B(16) => 
                           B_SHF_16_port, B(15) => B_SHF_15_port, B(14) => 
                           B_SHF_14_port, B(13) => B_SHF_13_port, B(12) => 
                           B_SHF_12_port, B(11) => B_SHF_11_port, B(10) => 
                           B_SHF_10_port, B(9) => B_SHF_9_port, B(8) => 
                           B_SHF_8_port, B(7) => B_SHF_7_port, B(6) => 
                           B_SHF_6_port, B(5) => B_SHF_5_port, B(4) => 
                           B_SHF_4_port, B(3) => B_SHF_3_port, B(2) => 
                           B_SHF_2_port, B(1) => B_SHF_1_port, B(0) => 
                           B_SHF_0_port, LOGIC_ARITH => LOGIC_ARITH, LEFT_RIGHT
                           => n180, RES(31) => SHIFT_RES_31_port, RES(30) => 
                           SHIFT_RES_30_port, RES(29) => SHIFT_RES_29_port, 
                           RES(28) => SHIFT_RES_28_port, RES(27) => 
                           SHIFT_RES_27_port, RES(26) => SHIFT_RES_26_port, 
                           RES(25) => SHIFT_RES_25_port, RES(24) => 
                           SHIFT_RES_24_port, RES(23) => SHIFT_RES_23_port, 
                           RES(22) => SHIFT_RES_22_port, RES(21) => 
                           SHIFT_RES_21_port, RES(20) => SHIFT_RES_20_port, 
                           RES(19) => SHIFT_RES_19_port, RES(18) => 
                           SHIFT_RES_18_port, RES(17) => SHIFT_RES_17_port, 
                           RES(16) => SHIFT_RES_16_port, RES(15) => 
                           SHIFT_RES_15_port, RES(14) => SHIFT_RES_14_port, 
                           RES(13) => SHIFT_RES_13_port, RES(12) => 
                           SHIFT_RES_12_port, RES(11) => SHIFT_RES_11_port, 
                           RES(10) => SHIFT_RES_10_port, RES(9) => 
                           SHIFT_RES_9_port, RES(8) => SHIFT_RES_8_port, RES(7)
                           => SHIFT_RES_7_port, RES(6) => SHIFT_RES_6_port, 
                           RES(5) => SHIFT_RES_5_port, RES(4) => 
                           SHIFT_RES_4_port, RES(3) => SHIFT_RES_3_port, RES(2)
                           => SHIFT_RES_2_port, RES(1) => SHIFT_RES_1_port, 
                           RES(0) => SHIFT_RES_0_port);
   Add_Sub_unit : P4Adder_NBIT32 port map( A(31) => A_ADD_31_port, A(30) => 
                           A_ADD_30_port, A(29) => A_ADD_29_port, A(28) => 
                           A_ADD_28_port, A(27) => A_ADD_27_port, A(26) => 
                           A_ADD_26_port, A(25) => A_ADD_25_port, A(24) => 
                           A_ADD_24_port, A(23) => A_ADD_23_port, A(22) => 
                           A_ADD_22_port, A(21) => A_ADD_21_port, A(20) => 
                           A_ADD_20_port, A(19) => A_ADD_19_port, A(18) => 
                           A_ADD_18_port, A(17) => A_ADD_17_port, A(16) => 
                           A_ADD_16_port, A(15) => A_ADD_15_port, A(14) => 
                           A_ADD_14_port, A(13) => A_ADD_13_port, A(12) => 
                           A_ADD_12_port, A(11) => A_ADD_11_port, A(10) => 
                           A_ADD_10_port, A(9) => A_ADD_9_port, A(8) => 
                           A_ADD_8_port, A(7) => A_ADD_7_port, A(6) => 
                           A_ADD_6_port, A(5) => A_ADD_5_port, A(4) => 
                           A_ADD_4_port, A(3) => A_ADD_3_port, A(2) => 
                           A_ADD_2_port, A(1) => A_ADD_1_port, A(0) => 
                           A_ADD_0_port, B(31) => B_ADD_31_port, B(30) => 
                           B_ADD_30_port, B(29) => B_ADD_29_port, B(28) => 
                           B_ADD_28_port, B(27) => B_ADD_27_port, B(26) => 
                           B_ADD_26_port, B(25) => B_ADD_25_port, B(24) => 
                           B_ADD_24_port, B(23) => B_ADD_23_port, B(22) => 
                           B_ADD_22_port, B(21) => B_ADD_21_port, B(20) => 
                           B_ADD_20_port, B(19) => B_ADD_19_port, B(18) => 
                           B_ADD_18_port, B(17) => B_ADD_17_port, B(16) => 
                           B_ADD_16_port, B(15) => B_ADD_15_port, B(14) => 
                           B_ADD_14_port, B(13) => B_ADD_13_port, B(12) => 
                           B_ADD_12_port, B(11) => B_ADD_11_port, B(10) => 
                           B_ADD_10_port, B(9) => B_ADD_9_port, B(8) => 
                           B_ADD_8_port, B(7) => B_ADD_7_port, B(6) => 
                           B_ADD_6_port, B(5) => B_ADD_5_port, B(4) => 
                           B_ADD_4_port, B(3) => B_ADD_3_port, B(2) => 
                           B_ADD_2_port, B(1) => B_ADD_1_port, B(0) => 
                           B_ADD_0_port, Cin => n1, S(31) => 
                           ADD_SUB_RES_31_port, S(30) => ADD_SUB_RES_30_port, 
                           S(29) => ADD_SUB_RES_29_port, S(28) => 
                           ADD_SUB_RES_28_port, S(27) => ADD_SUB_RES_27_port, 
                           S(26) => ADD_SUB_RES_26_port, S(25) => 
                           ADD_SUB_RES_25_port, S(24) => ADD_SUB_RES_24_port, 
                           S(23) => ADD_SUB_RES_23_port, S(22) => 
                           ADD_SUB_RES_22_port, S(21) => ADD_SUB_RES_21_port, 
                           S(20) => ADD_SUB_RES_20_port, S(19) => 
                           ADD_SUB_RES_19_port, S(18) => ADD_SUB_RES_18_port, 
                           S(17) => ADD_SUB_RES_17_port, S(16) => 
                           ADD_SUB_RES_16_port, S(15) => ADD_SUB_RES_15_port, 
                           S(14) => ADD_SUB_RES_14_port, S(13) => 
                           ADD_SUB_RES_13_port, S(12) => ADD_SUB_RES_12_port, 
                           S(11) => ADD_SUB_RES_11_port, S(10) => 
                           ADD_SUB_RES_10_port, S(9) => ADD_SUB_RES_9_port, 
                           S(8) => ADD_SUB_RES_8_port, S(7) => 
                           ADD_SUB_RES_7_port, S(6) => ADD_SUB_RES_6_port, S(5)
                           => ADD_SUB_RES_5_port, S(4) => ADD_SUB_RES_4_port, 
                           S(3) => ADD_SUB_RES_3_port, S(2) => 
                           ADD_SUB_RES_2_port, S(1) => ADD_SUB_RES_1_port, S(0)
                           => ADD_SUB_RES_0_port, Cout => n_1402);
   Res_mux : mux41_NBIT32_1 port map( A(31) => ADD_SUB_RES_31_port, A(30) => 
                           ADD_SUB_RES_30_port, A(29) => ADD_SUB_RES_29_port, 
                           A(28) => ADD_SUB_RES_28_port, A(27) => 
                           ADD_SUB_RES_27_port, A(26) => ADD_SUB_RES_26_port, 
                           A(25) => ADD_SUB_RES_25_port, A(24) => 
                           ADD_SUB_RES_24_port, A(23) => ADD_SUB_RES_23_port, 
                           A(22) => ADD_SUB_RES_22_port, A(21) => 
                           ADD_SUB_RES_21_port, A(20) => ADD_SUB_RES_20_port, 
                           A(19) => ADD_SUB_RES_19_port, A(18) => 
                           ADD_SUB_RES_18_port, A(17) => ADD_SUB_RES_17_port, 
                           A(16) => ADD_SUB_RES_16_port, A(15) => 
                           ADD_SUB_RES_15_port, A(14) => ADD_SUB_RES_14_port, 
                           A(13) => ADD_SUB_RES_13_port, A(12) => 
                           ADD_SUB_RES_12_port, A(11) => ADD_SUB_RES_11_port, 
                           A(10) => ADD_SUB_RES_10_port, A(9) => 
                           ADD_SUB_RES_9_port, A(8) => ADD_SUB_RES_8_port, A(7)
                           => ADD_SUB_RES_7_port, A(6) => ADD_SUB_RES_6_port, 
                           A(5) => ADD_SUB_RES_5_port, A(4) => 
                           ADD_SUB_RES_4_port, A(3) => ADD_SUB_RES_3_port, A(2)
                           => ADD_SUB_RES_2_port, A(1) => ADD_SUB_RES_1_port, 
                           A(0) => ADD_SUB_RES_0_port, B(31) => 
                           LOGIC_RES_31_port, B(30) => LOGIC_RES_30_port, B(29)
                           => LOGIC_RES_29_port, B(28) => LOGIC_RES_28_port, 
                           B(27) => LOGIC_RES_27_port, B(26) => 
                           LOGIC_RES_26_port, B(25) => LOGIC_RES_25_port, B(24)
                           => LOGIC_RES_24_port, B(23) => LOGIC_RES_23_port, 
                           B(22) => LOGIC_RES_22_port, B(21) => 
                           LOGIC_RES_21_port, B(20) => LOGIC_RES_20_port, B(19)
                           => LOGIC_RES_19_port, B(18) => LOGIC_RES_18_port, 
                           B(17) => LOGIC_RES_17_port, B(16) => 
                           LOGIC_RES_16_port, B(15) => LOGIC_RES_15_port, B(14)
                           => LOGIC_RES_14_port, B(13) => LOGIC_RES_13_port, 
                           B(12) => LOGIC_RES_12_port, B(11) => 
                           LOGIC_RES_11_port, B(10) => LOGIC_RES_10_port, B(9) 
                           => LOGIC_RES_9_port, B(8) => LOGIC_RES_8_port, B(7) 
                           => LOGIC_RES_7_port, B(6) => LOGIC_RES_6_port, B(5) 
                           => LOGIC_RES_5_port, B(4) => LOGIC_RES_4_port, B(3) 
                           => LOGIC_RES_3_port, B(2) => LOGIC_RES_2_port, B(1) 
                           => LOGIC_RES_1_port, B(0) => LOGIC_RES_0_port, C(31)
                           => SHIFT_RES_31_port, C(30) => SHIFT_RES_30_port, 
                           C(29) => SHIFT_RES_29_port, C(28) => 
                           SHIFT_RES_28_port, C(27) => SHIFT_RES_27_port, C(26)
                           => SHIFT_RES_26_port, C(25) => SHIFT_RES_25_port, 
                           C(24) => SHIFT_RES_24_port, C(23) => 
                           SHIFT_RES_23_port, C(22) => SHIFT_RES_22_port, C(21)
                           => SHIFT_RES_21_port, C(20) => SHIFT_RES_20_port, 
                           C(19) => SHIFT_RES_19_port, C(18) => 
                           SHIFT_RES_18_port, C(17) => SHIFT_RES_17_port, C(16)
                           => SHIFT_RES_16_port, C(15) => SHIFT_RES_15_port, 
                           C(14) => SHIFT_RES_14_port, C(13) => 
                           SHIFT_RES_13_port, C(12) => SHIFT_RES_12_port, C(11)
                           => SHIFT_RES_11_port, C(10) => SHIFT_RES_10_port, 
                           C(9) => SHIFT_RES_9_port, C(8) => SHIFT_RES_8_port, 
                           C(7) => SHIFT_RES_7_port, C(6) => SHIFT_RES_6_port, 
                           C(5) => SHIFT_RES_5_port, C(4) => SHIFT_RES_4_port, 
                           C(3) => SHIFT_RES_3_port, C(2) => SHIFT_RES_2_port, 
                           C(1) => SHIFT_RES_1_port, C(0) => SHIFT_RES_0_port, 
                           D(31) => COMP_RES_31_port, D(30) => COMP_RES_30_port
                           , D(29) => COMP_RES_29_port, D(28) => 
                           COMP_RES_28_port, D(27) => COMP_RES_27_port, D(26) 
                           => COMP_RES_26_port, D(25) => COMP_RES_25_port, 
                           D(24) => COMP_RES_24_port, D(23) => COMP_RES_23_port
                           , D(22) => COMP_RES_22_port, D(21) => 
                           COMP_RES_21_port, D(20) => COMP_RES_20_port, D(19) 
                           => COMP_RES_19_port, D(18) => COMP_RES_18_port, 
                           D(17) => COMP_RES_17_port, D(16) => COMP_RES_16_port
                           , D(15) => COMP_RES_15_port, D(14) => 
                           COMP_RES_14_port, D(13) => COMP_RES_13_port, D(12) 
                           => COMP_RES_12_port, D(11) => COMP_RES_11_port, 
                           D(10) => COMP_RES_10_port, D(9) => COMP_RES_9_port, 
                           D(8) => COMP_RES_8_port, D(7) => COMP_RES_7_port, 
                           D(6) => COMP_RES_6_port, D(5) => COMP_RES_5_port, 
                           D(4) => COMP_RES_4_port, D(3) => COMP_RES_3_port, 
                           D(2) => COMP_RES_2_port, D(1) => COMP_RES_1_port, 
                           D(0) => COMP_RES_0_port, S(1) => 
                           select_type_sig_1_port, S(0) => 
                           select_type_sig_0_port, Z(31) => 
                           sig_intraMux_31_port, Z(30) => sig_intraMux_30_port,
                           Z(29) => sig_intraMux_29_port, Z(28) => 
                           sig_intraMux_28_port, Z(27) => sig_intraMux_27_port,
                           Z(26) => sig_intraMux_26_port, Z(25) => 
                           sig_intraMux_25_port, Z(24) => sig_intraMux_24_port,
                           Z(23) => sig_intraMux_23_port, Z(22) => 
                           sig_intraMux_22_port, Z(21) => sig_intraMux_21_port,
                           Z(20) => sig_intraMux_20_port, Z(19) => 
                           sig_intraMux_19_port, Z(18) => sig_intraMux_18_port,
                           Z(17) => sig_intraMux_17_port, Z(16) => 
                           sig_intraMux_16_port, Z(15) => sig_intraMux_15_port,
                           Z(14) => sig_intraMux_14_port, Z(13) => 
                           sig_intraMux_13_port, Z(12) => sig_intraMux_12_port,
                           Z(11) => sig_intraMux_11_port, Z(10) => 
                           sig_intraMux_10_port, Z(9) => sig_intraMux_9_port, 
                           Z(8) => sig_intraMux_8_port, Z(7) => 
                           sig_intraMux_7_port, Z(6) => sig_intraMux_6_port, 
                           Z(5) => sig_intraMux_5_port, Z(4) => 
                           sig_intraMux_4_port, Z(3) => sig_intraMux_3_port, 
                           Z(2) => sig_intraMux_2_port, Z(1) => 
                           sig_intraMux_1_port, Z(0) => sig_intraMux_0_port);
   Zeros_mux : mux21_NBIT32_1 port map( A(31) => sig_intraMux_31_port, A(30) =>
                           sig_intraMux_30_port, A(29) => sig_intraMux_29_port,
                           A(28) => sig_intraMux_28_port, A(27) => 
                           sig_intraMux_27_port, A(26) => sig_intraMux_26_port,
                           A(25) => sig_intraMux_25_port, A(24) => 
                           sig_intraMux_24_port, A(23) => sig_intraMux_23_port,
                           A(22) => sig_intraMux_22_port, A(21) => 
                           sig_intraMux_21_port, A(20) => sig_intraMux_20_port,
                           A(19) => sig_intraMux_19_port, A(18) => 
                           sig_intraMux_18_port, A(17) => sig_intraMux_17_port,
                           A(16) => sig_intraMux_16_port, A(15) => 
                           sig_intraMux_15_port, A(14) => sig_intraMux_14_port,
                           A(13) => sig_intraMux_13_port, A(12) => 
                           sig_intraMux_12_port, A(11) => sig_intraMux_11_port,
                           A(10) => sig_intraMux_10_port, A(9) => 
                           sig_intraMux_9_port, A(8) => sig_intraMux_8_port, 
                           A(7) => sig_intraMux_7_port, A(6) => 
                           sig_intraMux_6_port, A(5) => sig_intraMux_5_port, 
                           A(4) => sig_intraMux_4_port, A(3) => 
                           sig_intraMux_3_port, A(2) => sig_intraMux_2_port, 
                           A(1) => sig_intraMux_1_port, A(0) => 
                           sig_intraMux_0_port, B(31) => X_Logic0_port, B(30) 
                           => X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, S => select_zero_sig, Z(31) => 
                           ALU_RES(31), Z(30) => ALU_RES(30), Z(29) => 
                           ALU_RES(29), Z(28) => ALU_RES(28), Z(27) => 
                           ALU_RES(27), Z(26) => ALU_RES(26), Z(25) => 
                           ALU_RES(25), Z(24) => ALU_RES(24), Z(23) => 
                           ALU_RES(23), Z(22) => ALU_RES(22), Z(21) => 
                           ALU_RES(21), Z(20) => ALU_RES(20), Z(19) => 
                           ALU_RES(19), Z(18) => ALU_RES(18), Z(17) => 
                           ALU_RES(17), Z(16) => ALU_RES(16), Z(15) => 
                           ALU_RES(15), Z(14) => ALU_RES(14), Z(13) => 
                           ALU_RES(13), Z(12) => ALU_RES(12), Z(11) => 
                           ALU_RES(11), Z(10) => ALU_RES(10), Z(9) => 
                           ALU_RES(9), Z(8) => ALU_RES(8), Z(7) => ALU_RES(7), 
                           Z(6) => ALU_RES(6), Z(5) => ALU_RES(5), Z(4) => 
                           ALU_RES(4), Z(3) => ALU_RES(3), Z(2) => ALU_RES(2), 
                           Z(1) => ALU_RES(1), Z(0) => ALU_RES(0));
   U2 : NOR2_X1 port map( A1 => n13, A2 => n58, ZN => A_SHF_5_port);
   U3 : NOR2_X1 port map( A1 => n13, A2 => n59, ZN => A_SHF_6_port);
   U4 : BUF_X1 port map( A => n158, Z => n23);
   U5 : BUF_X1 port map( A => n158, Z => n24);
   U6 : BUF_X1 port map( A => n158, Z => n25);
   U7 : BUF_X1 port map( A => n177, Z => n5);
   U8 : BUF_X1 port map( A => n177, Z => n6);
   U9 : BUF_X1 port map( A => n177, Z => n7);
   U10 : BUF_X1 port map( A => n177, Z => n9);
   U11 : BUF_X1 port map( A => n177, Z => n8);
   U12 : BUF_X1 port map( A => n179, Z => n17);
   U13 : BUF_X1 port map( A => n179, Z => n18);
   U14 : BUF_X1 port map( A => n179, Z => n21);
   U15 : BUF_X1 port map( A => n179, Z => n20);
   U16 : BUF_X1 port map( A => n179, Z => n19);
   U17 : BUF_X1 port map( A => n176, Z => n2);
   U18 : BUF_X1 port map( A => n176, Z => n3);
   U19 : BUF_X1 port map( A => n176, Z => n4);
   U20 : AND2_X1 port map( A1 => n28, A2 => n29, ZN => n158);
   U21 : NOR2_X1 port map( A1 => n15, A2 => n168, ZN => B_SHF_3_port);
   U22 : NOR2_X1 port map( A1 => n12, A2 => n50, ZN => A_SHF_27_port);
   U23 : NOR2_X1 port map( A1 => n12, A2 => n49, ZN => A_SHF_26_port);
   U24 : NOR2_X1 port map( A1 => n13, A2 => n64, ZN => B_SHF_10_port);
   U25 : NOR2_X1 port map( A1 => n16, A2 => n174, ZN => B_SHF_9_port);
   U26 : NOR2_X1 port map( A1 => n16, A2 => n173, ZN => B_SHF_8_port);
   U27 : NOR2_X1 port map( A1 => n11, A2 => n39, ZN => A_SHF_17_port);
   U28 : NOR2_X1 port map( A1 => n13, A2 => n60, ZN => A_SHF_7_port);
   U29 : NOR2_X1 port map( A1 => n15, A2 => n165, ZN => B_SHF_2_port);
   U30 : NOR2_X1 port map( A1 => n11, A2 => n40, ZN => A_SHF_18_port);
   U31 : NOR2_X1 port map( A1 => n12, A2 => n48, ZN => A_SHF_25_port);
   U32 : NOR2_X1 port map( A1 => n13, A2 => n57, ZN => A_SHF_4_port);
   U33 : NOR2_X1 port map( A1 => n12, A2 => n51, ZN => A_SHF_28_port);
   U34 : NOR2_X1 port map( A1 => n15, A2 => n170, ZN => B_SHF_5_port);
   U35 : NOR2_X1 port map( A1 => n16, A2 => n172, ZN => B_SHF_7_port);
   U36 : NOR2_X1 port map( A1 => n16, A2 => n171, ZN => B_SHF_6_port);
   U37 : NOR2_X1 port map( A1 => n23, A2 => n31, ZN => A_ADD_0_port);
   U38 : NOR2_X1 port map( A1 => n13, A2 => n61, ZN => A_SHF_8_port);
   U39 : NOR2_X1 port map( A1 => n12, A2 => n53, ZN => A_SHF_2_port);
   U40 : NOR2_X1 port map( A1 => n25, A2 => n57, ZN => A_ADD_4_port);
   U41 : NOR2_X1 port map( A1 => n25, A2 => n58, ZN => A_ADD_5_port);
   U42 : NOR2_X1 port map( A1 => n25, A2 => n59, ZN => A_ADD_6_port);
   U43 : NOR2_X1 port map( A1 => n25, A2 => n61, ZN => A_ADD_8_port);
   U44 : NOR2_X1 port map( A1 => n25, A2 => n62, ZN => A_ADD_9_port);
   U45 : NOR2_X1 port map( A1 => n25, A2 => n56, ZN => A_ADD_3_port);
   U46 : NOR2_X1 port map( A1 => n25, A2 => n60, ZN => A_ADD_7_port);
   U47 : NOR2_X1 port map( A1 => n25, A2 => n55, ZN => A_ADD_31_port);
   U48 : NOR2_X1 port map( A1 => n23, A2 => n42, ZN => A_ADD_1_port);
   U49 : NOR2_X1 port map( A1 => n24, A2 => n53, ZN => A_ADD_2_port);
   U50 : NOR2_X1 port map( A1 => n23, A2 => n32, ZN => A_ADD_10_port);
   U51 : NOR2_X1 port map( A1 => n23, A2 => n34, ZN => A_ADD_12_port);
   U52 : NOR2_X1 port map( A1 => n23, A2 => n35, ZN => A_ADD_13_port);
   U53 : NOR2_X1 port map( A1 => n23, A2 => n36, ZN => A_ADD_14_port);
   U54 : NOR2_X1 port map( A1 => n23, A2 => n38, ZN => A_ADD_16_port);
   U55 : NOR2_X1 port map( A1 => n23, A2 => n39, ZN => A_ADD_17_port);
   U56 : NOR2_X1 port map( A1 => n23, A2 => n40, ZN => A_ADD_18_port);
   U57 : NOR2_X1 port map( A1 => n24, A2 => n43, ZN => A_ADD_20_port);
   U58 : NOR2_X1 port map( A1 => n24, A2 => n44, ZN => A_ADD_21_port);
   U59 : NOR2_X1 port map( A1 => n24, A2 => n45, ZN => A_ADD_22_port);
   U60 : NOR2_X1 port map( A1 => n24, A2 => n47, ZN => A_ADD_24_port);
   U61 : NOR2_X1 port map( A1 => n24, A2 => n48, ZN => A_ADD_25_port);
   U62 : NOR2_X1 port map( A1 => n24, A2 => n49, ZN => A_ADD_26_port);
   U63 : NOR2_X1 port map( A1 => n24, A2 => n51, ZN => A_ADD_28_port);
   U64 : NOR2_X1 port map( A1 => n24, A2 => n52, ZN => A_ADD_29_port);
   U65 : NOR2_X1 port map( A1 => n24, A2 => n54, ZN => A_ADD_30_port);
   U66 : NOR2_X1 port map( A1 => n23, A2 => n33, ZN => A_ADD_11_port);
   U67 : NOR2_X1 port map( A1 => n23, A2 => n37, ZN => A_ADD_15_port);
   U68 : NOR2_X1 port map( A1 => n23, A2 => n41, ZN => A_ADD_19_port);
   U69 : NOR2_X1 port map( A1 => n24, A2 => n46, ZN => A_ADD_23_port);
   U70 : NOR2_X1 port map( A1 => n24, A2 => n50, ZN => A_ADD_27_port);
   U71 : NOR2_X1 port map( A1 => n14, A2 => n74, ZN => B_SHF_1_port);
   U72 : NOR2_X1 port map( A1 => n12, A2 => n43, ZN => A_SHF_20_port);
   U73 : NOR2_X1 port map( A1 => n11, A2 => n34, ZN => A_SHF_12_port);
   U74 : NOR2_X1 port map( A1 => n12, A2 => n44, ZN => A_SHF_21_port);
   U75 : NOR2_X1 port map( A1 => n11, A2 => n35, ZN => A_SHF_13_port);
   U76 : NOR2_X1 port map( A1 => n11, A2 => n41, ZN => A_SHF_19_port);
   U77 : NOR2_X1 port map( A1 => n12, A2 => n45, ZN => A_SHF_22_port);
   U78 : NOR2_X1 port map( A1 => n11, A2 => n36, ZN => A_SHF_14_port);
   U79 : NOR2_X1 port map( A1 => n12, A2 => n46, ZN => A_SHF_23_port);
   U80 : NOR2_X1 port map( A1 => n12, A2 => n47, ZN => A_SHF_24_port);
   U81 : NOR2_X1 port map( A1 => n15, A2 => n163, ZN => B_SHF_28_port);
   U82 : NOR2_X1 port map( A1 => n15, A2 => n162, ZN => B_SHF_27_port);
   U83 : NOR2_X1 port map( A1 => n15, A2 => n161, ZN => B_SHF_26_port);
   U84 : NOR2_X1 port map( A1 => n11, A2 => n42, ZN => A_SHF_1_port);
   U85 : NOR2_X1 port map( A1 => n13, A2 => n65, ZN => B_SHF_11_port);
   U86 : NOR2_X1 port map( A1 => n13, A2 => n62, ZN => A_SHF_9_port);
   U87 : NOR2_X1 port map( A1 => n11, A2 => n31, ZN => A_SHF_0_port);
   U88 : NOR2_X1 port map( A1 => n11, A2 => n33, ZN => A_SHF_11_port);
   U89 : NOR2_X1 port map( A1 => n11, A2 => n37, ZN => A_SHF_15_port);
   U90 : NOR2_X1 port map( A1 => n12, A2 => n52, ZN => A_SHF_29_port);
   U91 : NOR2_X1 port map( A1 => n11, A2 => n38, ZN => A_SHF_16_port);
   U92 : NOR2_X1 port map( A1 => n13, A2 => n56, ZN => A_SHF_3_port);
   U93 : NOR2_X1 port map( A1 => n14, A2 => n72, ZN => B_SHF_18_port);
   U94 : BUF_X1 port map( A => n178, Z => n13);
   U95 : BUF_X1 port map( A => n178, Z => n14);
   U96 : BUF_X1 port map( A => n178, Z => n11);
   U97 : BUF_X1 port map( A => n178, Z => n12);
   U98 : BUF_X1 port map( A => n178, Z => n15);
   U99 : NOR2_X1 port map( A1 => n15, A2 => n164, ZN => B_SHF_29_port);
   U100 : NOR2_X1 port map( A1 => n15, A2 => n166, ZN => B_SHF_30_port);
   U101 : NOR2_X1 port map( A1 => n15, A2 => n160, ZN => B_SHF_25_port);
   U102 : NOR2_X1 port map( A1 => n13, A2 => n63, ZN => B_SHF_0_port);
   U103 : NOR2_X1 port map( A1 => n14, A2 => n70, ZN => B_SHF_16_port);
   U104 : NOR2_X1 port map( A1 => n11, A2 => n32, ZN => A_SHF_10_port);
   U105 : NOR2_X1 port map( A1 => n14, A2 => n71, ZN => B_SHF_17_port);
   U106 : NOR2_X1 port map( A1 => n14, A2 => n69, ZN => B_SHF_15_port);
   U107 : BUF_X1 port map( A => n156, Z => n27);
   U108 : BUF_X1 port map( A => n156, Z => n26);
   U109 : NOR2_X1 port map( A1 => n15, A2 => n159, ZN => B_SHF_24_port);
   U110 : NOR2_X1 port map( A1 => n14, A2 => n86, ZN => B_SHF_23_port);
   U111 : NOR2_X1 port map( A1 => n14, A2 => n77, ZN => B_SHF_22_port);
   U112 : NOR2_X1 port map( A1 => n15, A2 => n169, ZN => B_SHF_4_port);
   U113 : NAND4_X1 port map( A1 => n80, A2 => n81, A3 => n82, A4 => n181, ZN =>
                           select_type_sig_0_port);
   U114 : NOR2_X1 port map( A1 => n12, A2 => n54, ZN => A_SHF_30_port);
   U115 : INV_X1 port map( A => n81, ZN => n179);
   U116 : NOR2_X1 port map( A1 => n14, A2 => n73, ZN => B_SHF_19_port);
   U117 : NOR2_X1 port map( A1 => n14, A2 => n67, ZN => B_SHF_13_port);
   U118 : NOR2_X1 port map( A1 => n14, A2 => n76, ZN => B_SHF_21_port);
   U119 : NOR2_X1 port map( A1 => n14, A2 => n68, ZN => B_SHF_14_port);
   U120 : NOR2_X1 port map( A1 => n14, A2 => n75, ZN => B_SHF_20_port);
   U121 : NOR2_X1 port map( A1 => n13, A2 => n66, ZN => B_SHF_12_port);
   U122 : NAND2_X1 port map( A1 => n16, A2 => n181, ZN => 
                           select_type_sig_1_port);
   U123 : BUF_X1 port map( A => n156, Z => n28);
   U124 : INV_X1 port map( A => n80, ZN => n177);
   U125 : INV_X1 port map( A => n82, ZN => n176);
   U126 : NOR2_X1 port map( A1 => n15, A2 => n167, ZN => B_SHF_31_port);
   U127 : OAI22_X1 port map( A1 => n63, A2 => n28, B1 => OP2(0), B2 => n29, ZN 
                           => B_ADD_0_port);
   U128 : OAI22_X1 port map( A1 => n74, A2 => n27, B1 => OP2(1), B2 => n30, ZN 
                           => B_ADD_1_port);
   U129 : OAI22_X1 port map( A1 => n165, A2 => n26, B1 => OP2(2), B2 => n29, ZN
                           => B_ADD_2_port);
   U130 : OAI22_X1 port map( A1 => n169, A2 => n26, B1 => OP2(4), B2 => n29, ZN
                           => B_ADD_4_port);
   U131 : OAI22_X1 port map( A1 => n170, A2 => n26, B1 => OP2(5), B2 => n29, ZN
                           => B_ADD_5_port);
   U132 : OAI22_X1 port map( A1 => n171, A2 => n26, B1 => OP2(6), B2 => n29, ZN
                           => B_ADD_6_port);
   U133 : OAI22_X1 port map( A1 => n173, A2 => n26, B1 => OP2(8), B2 => n29, ZN
                           => B_ADD_8_port);
   U134 : OAI22_X1 port map( A1 => n174, A2 => n26, B1 => OP2(9), B2 => n29, ZN
                           => B_ADD_9_port);
   U135 : OAI22_X1 port map( A1 => n71, A2 => n27, B1 => OP2(17), B2 => n30, ZN
                           => B_ADD_17_port);
   U136 : OAI22_X1 port map( A1 => n72, A2 => n27, B1 => OP2(18), B2 => n30, ZN
                           => B_ADD_18_port);
   U137 : OAI22_X1 port map( A1 => n75, A2 => n27, B1 => OP2(20), B2 => n30, ZN
                           => B_ADD_20_port);
   U138 : OAI22_X1 port map( A1 => n76, A2 => n27, B1 => OP2(21), B2 => n30, ZN
                           => B_ADD_21_port);
   U139 : OAI22_X1 port map( A1 => n77, A2 => n27, B1 => OP2(22), B2 => n30, ZN
                           => B_ADD_22_port);
   U140 : OAI22_X1 port map( A1 => n159, A2 => n27, B1 => OP2(24), B2 => n30, 
                           ZN => B_ADD_24_port);
   U141 : OAI22_X1 port map( A1 => n160, A2 => n27, B1 => OP2(25), B2 => n30, 
                           ZN => B_ADD_25_port);
   U142 : OAI22_X1 port map( A1 => n161, A2 => n27, B1 => OP2(26), B2 => n30, 
                           ZN => B_ADD_26_port);
   U143 : OAI22_X1 port map( A1 => n163, A2 => n26, B1 => OP2(28), B2 => n29, 
                           ZN => B_ADD_28_port);
   U144 : OAI22_X1 port map( A1 => n164, A2 => n26, B1 => OP2(29), B2 => n29, 
                           ZN => B_ADD_29_port);
   U145 : OAI22_X1 port map( A1 => n166, A2 => n26, B1 => OP2(30), B2 => n29, 
                           ZN => B_ADD_30_port);
   U146 : OAI22_X1 port map( A1 => n168, A2 => n26, B1 => OP2(3), B2 => n29, ZN
                           => B_ADD_3_port);
   U147 : OAI22_X1 port map( A1 => n172, A2 => n26, B1 => OP2(7), B2 => n29, ZN
                           => B_ADD_7_port);
   U148 : OAI22_X1 port map( A1 => n73, A2 => n27, B1 => OP2(19), B2 => n30, ZN
                           => B_ADD_19_port);
   U149 : OAI22_X1 port map( A1 => n86, A2 => n27, B1 => OP2(23), B2 => n30, ZN
                           => B_ADD_23_port);
   U150 : OAI22_X1 port map( A1 => n162, A2 => n27, B1 => OP2(27), B2 => n30, 
                           ZN => B_ADD_27_port);
   U151 : OAI22_X1 port map( A1 => n167, A2 => n26, B1 => OP2(31), B2 => n29, 
                           ZN => B_ADD_31_port);
   U152 : OAI22_X1 port map( A1 => n64, A2 => n28, B1 => OP2(10), B2 => n30, ZN
                           => B_ADD_10_port);
   U153 : OAI22_X1 port map( A1 => n66, A2 => n28, B1 => OP2(12), B2 => n29, ZN
                           => B_ADD_12_port);
   U154 : OAI22_X1 port map( A1 => n67, A2 => n28, B1 => OP2(13), B2 => n30, ZN
                           => B_ADD_13_port);
   U155 : OAI22_X1 port map( A1 => n68, A2 => n28, B1 => OP2(14), B2 => n29, ZN
                           => B_ADD_14_port);
   U156 : OAI22_X1 port map( A1 => n70, A2 => n28, B1 => OP2(16), B2 => n30, ZN
                           => B_ADD_16_port);
   U157 : OAI22_X1 port map( A1 => n65, A2 => n28, B1 => OP2(11), B2 => n29, ZN
                           => B_ADD_11_port);
   U158 : OAI22_X1 port map( A1 => n69, A2 => n28, B1 => OP2(15), B2 => n30, ZN
                           => B_ADD_15_port);
   U159 : OAI22_X1 port map( A1 => n152, A2 => n63, B1 => n153, B2 => n31, ZN 
                           => LOGIC_RES_0_port);
   U160 : AOI21_X1 port map( B1 => n7, B2 => n63, A => n19, ZN => n153);
   U161 : AOI221_X1 port map( B1 => OP1(0), B2 => n4, C1 => n5, C2 => n31, A =>
                           n17, ZN => n152);
   U162 : OAI22_X1 port map( A1 => n130, A2 => n74, B1 => n131, B2 => n42, ZN 
                           => LOGIC_RES_1_port);
   U163 : AOI21_X1 port map( B1 => n9, B2 => n74, A => n21, ZN => n131);
   U164 : AOI221_X1 port map( B1 => OP1(1), B2 => n3, C1 => n6, C2 => n42, A =>
                           n18, ZN => n130);
   U165 : OAI22_X1 port map( A1 => n108, A2 => n165, B1 => n109, B2 => n53, ZN 
                           => LOGIC_RES_2_port);
   U166 : AOI21_X1 port map( B1 => n8, B2 => n165, A => n20, ZN => n109);
   U167 : AOI221_X1 port map( B1 => OP1(2), B2 => n2, C1 => n7, C2 => n53, A =>
                           n19, ZN => n108);
   U168 : OAI22_X1 port map( A1 => n102, A2 => n168, B1 => n103, B2 => n56, ZN 
                           => LOGIC_RES_3_port);
   U169 : AOI21_X1 port map( B1 => n8, B2 => n168, A => n20, ZN => n103);
   U170 : AOI221_X1 port map( B1 => OP1(3), B2 => n2, C1 => n6, C2 => n56, A =>
                           n18, ZN => n102);
   U171 : OAI22_X1 port map( A1 => n100, A2 => n169, B1 => n101, B2 => n57, ZN 
                           => LOGIC_RES_4_port);
   U172 : AOI21_X1 port map( B1 => n8, B2 => n169, A => n20, ZN => n101);
   U173 : AOI221_X1 port map( B1 => OP1(4), B2 => n2, C1 => n6, C2 => n57, A =>
                           n18, ZN => n100);
   U174 : OAI22_X1 port map( A1 => n98, A2 => n170, B1 => n99, B2 => n58, ZN =>
                           LOGIC_RES_5_port);
   U175 : AOI21_X1 port map( B1 => n7, B2 => n170, A => n19, ZN => n99);
   U176 : AOI221_X1 port map( B1 => OP1(5), B2 => n2, C1 => n6, C2 => n58, A =>
                           n18, ZN => n98);
   U178 : OAI22_X1 port map( A1 => n96, A2 => n171, B1 => n97, B2 => n59, ZN =>
                           LOGIC_RES_6_port);
   U179 : AOI21_X1 port map( B1 => n7, B2 => n171, A => n19, ZN => n97);
   U180 : AOI221_X1 port map( B1 => OP1(6), B2 => n2, C1 => n5, C2 => n59, A =>
                           n17, ZN => n96);
   U181 : OAI22_X1 port map( A1 => n94, A2 => n172, B1 => n95, B2 => n60, ZN =>
                           LOGIC_RES_7_port);
   U182 : AOI21_X1 port map( B1 => n8, B2 => n172, A => n20, ZN => n95);
   U183 : AOI221_X1 port map( B1 => OP1(7), B2 => n2, C1 => n5, C2 => n60, A =>
                           n17, ZN => n94);
   U184 : OAI22_X1 port map( A1 => n92, A2 => n173, B1 => n93, B2 => n61, ZN =>
                           LOGIC_RES_8_port);
   U185 : AOI21_X1 port map( B1 => n7, B2 => n173, A => n19, ZN => n93);
   U186 : AOI221_X1 port map( B1 => OP1(8), B2 => n2, C1 => n5, C2 => n61, A =>
                           n17, ZN => n92);
   U187 : OAI22_X1 port map( A1 => n90, A2 => n174, B1 => n91, B2 => n62, ZN =>
                           LOGIC_RES_9_port);
   U188 : AOI21_X1 port map( B1 => n8, B2 => n174, A => n20, ZN => n91);
   U189 : AOI221_X1 port map( B1 => n2, B2 => OP1(9), C1 => n5, C2 => n62, A =>
                           n17, ZN => n90);
   U190 : OAI22_X1 port map( A1 => n150, A2 => n64, B1 => n151, B2 => n32, ZN 
                           => LOGIC_RES_10_port);
   U191 : AOI21_X1 port map( B1 => n10, B2 => n64, A => n22, ZN => n151);
   U192 : AOI221_X1 port map( B1 => OP1(10), B2 => n4, C1 => n5, C2 => n32, A 
                           => n17, ZN => n150);
   U193 : OAI22_X1 port map( A1 => n148, A2 => n65, B1 => n149, B2 => n33, ZN 
                           => LOGIC_RES_11_port);
   U194 : AOI21_X1 port map( B1 => n10, B2 => n65, A => n22, ZN => n149);
   U195 : AOI221_X1 port map( B1 => OP1(11), B2 => n4, C1 => n5, C2 => n33, A 
                           => n17, ZN => n148);
   U196 : OAI22_X1 port map( A1 => n146, A2 => n66, B1 => n147, B2 => n34, ZN 
                           => LOGIC_RES_12_port);
   U197 : AOI21_X1 port map( B1 => n10, B2 => n66, A => n21, ZN => n147);
   U198 : AOI221_X1 port map( B1 => OP1(12), B2 => n4, C1 => n5, C2 => n34, A 
                           => n17, ZN => n146);
   U199 : OAI22_X1 port map( A1 => n144, A2 => n67, B1 => n145, B2 => n35, ZN 
                           => LOGIC_RES_13_port);
   U200 : AOI21_X1 port map( B1 => n10, B2 => n67, A => n21, ZN => n145);
   U201 : AOI221_X1 port map( B1 => OP1(13), B2 => n4, C1 => n5, C2 => n35, A 
                           => n17, ZN => n144);
   U202 : OAI22_X1 port map( A1 => n142, A2 => n68, B1 => n143, B2 => n36, ZN 
                           => LOGIC_RES_14_port);
   U203 : AOI21_X1 port map( B1 => n9, B2 => n68, A => n21, ZN => n143);
   U204 : AOI221_X1 port map( B1 => OP1(14), B2 => n4, C1 => n5, C2 => n36, A 
                           => n17, ZN => n142);
   U205 : OAI22_X1 port map( A1 => n140, A2 => n69, B1 => n141, B2 => n37, ZN 
                           => LOGIC_RES_15_port);
   U206 : AOI21_X1 port map( B1 => n9, B2 => n69, A => n21, ZN => n141);
   U207 : AOI221_X1 port map( B1 => OP1(15), B2 => n4, C1 => n5, C2 => n37, A 
                           => n17, ZN => n140);
   U208 : OAI22_X1 port map( A1 => n138, A2 => n70, B1 => n139, B2 => n38, ZN 
                           => LOGIC_RES_16_port);
   U209 : AOI21_X1 port map( B1 => n9, B2 => n70, A => n21, ZN => n139);
   U210 : AOI221_X1 port map( B1 => OP1(16), B2 => n4, C1 => n5, C2 => n38, A 
                           => n17, ZN => n138);
   U211 : OAI22_X1 port map( A1 => n136, A2 => n71, B1 => n137, B2 => n39, ZN 
                           => LOGIC_RES_17_port);
   U212 : AOI21_X1 port map( B1 => n9, B2 => n71, A => n21, ZN => n137);
   U213 : AOI221_X1 port map( B1 => OP1(17), B2 => n3, C1 => n6, C2 => n39, A 
                           => n18, ZN => n136);
   U214 : OAI22_X1 port map( A1 => n134, A2 => n72, B1 => n135, B2 => n40, ZN 
                           => LOGIC_RES_18_port);
   U215 : AOI21_X1 port map( B1 => n9, B2 => n72, A => n21, ZN => n135);
   U216 : AOI221_X1 port map( B1 => OP1(18), B2 => n3, C1 => n6, C2 => n40, A 
                           => n18, ZN => n134);
   U217 : OAI22_X1 port map( A1 => n132, A2 => n73, B1 => n133, B2 => n41, ZN 
                           => LOGIC_RES_19_port);
   U218 : AOI21_X1 port map( B1 => n9, B2 => n73, A => n21, ZN => n133);
   U219 : AOI221_X1 port map( B1 => OP1(19), B2 => n3, C1 => n6, C2 => n41, A 
                           => n18, ZN => n132);
   U220 : OAI22_X1 port map( A1 => n128, A2 => n75, B1 => n129, B2 => n43, ZN 
                           => LOGIC_RES_20_port);
   U221 : AOI21_X1 port map( B1 => n9, B2 => n75, A => n21, ZN => n129);
   U222 : AOI221_X1 port map( B1 => OP1(20), B2 => n3, C1 => n6, C2 => n43, A 
                           => n18, ZN => n128);
   U223 : OAI22_X1 port map( A1 => n126, A2 => n76, B1 => n127, B2 => n44, ZN 
                           => LOGIC_RES_21_port);
   U224 : AOI21_X1 port map( B1 => n9, B2 => n76, A => n21, ZN => n127);
   U225 : AOI221_X1 port map( B1 => OP1(21), B2 => n3, C1 => n6, C2 => n44, A 
                           => n18, ZN => n126);
   U226 : OAI22_X1 port map( A1 => n124, A2 => n77, B1 => n125, B2 => n45, ZN 
                           => LOGIC_RES_22_port);
   U227 : AOI21_X1 port map( B1 => n9, B2 => n77, A => n21, ZN => n125);
   U228 : AOI221_X1 port map( B1 => OP1(22), B2 => n3, C1 => n6, C2 => n45, A 
                           => n18, ZN => n124);
   U229 : OAI22_X1 port map( A1 => n122, A2 => n86, B1 => n123, B2 => n46, ZN 
                           => LOGIC_RES_23_port);
   U230 : AOI21_X1 port map( B1 => n9, B2 => n86, A => n21, ZN => n123);
   U231 : AOI221_X1 port map( B1 => OP1(23), B2 => n3, C1 => n6, C2 => n46, A 
                           => n18, ZN => n122);
   U232 : OAI22_X1 port map( A1 => n120, A2 => n159, B1 => n121, B2 => n47, ZN 
                           => LOGIC_RES_24_port);
   U233 : AOI21_X1 port map( B1 => n9, B2 => n159, A => n20, ZN => n121);
   U234 : AOI221_X1 port map( B1 => OP1(24), B2 => n3, C1 => n7, C2 => n47, A 
                           => n19, ZN => n120);
   U235 : OAI22_X1 port map( A1 => n118, A2 => n160, B1 => n119, B2 => n48, ZN 
                           => LOGIC_RES_25_port);
   U236 : AOI21_X1 port map( B1 => n8, B2 => n160, A => n20, ZN => n119);
   U237 : AOI221_X1 port map( B1 => OP1(25), B2 => n3, C1 => n7, C2 => n48, A 
                           => n19, ZN => n118);
   U238 : OAI22_X1 port map( A1 => n116, A2 => n161, B1 => n117, B2 => n49, ZN 
                           => LOGIC_RES_26_port);
   U239 : AOI21_X1 port map( B1 => n8, B2 => n161, A => n20, ZN => n117);
   U240 : AOI221_X1 port map( B1 => OP1(26), B2 => n3, C1 => n6, C2 => n49, A 
                           => n18, ZN => n116);
   U241 : OAI22_X1 port map( A1 => n114, A2 => n162, B1 => n115, B2 => n50, ZN 
                           => LOGIC_RES_27_port);
   U242 : AOI21_X1 port map( B1 => n8, B2 => n162, A => n20, ZN => n115);
   U243 : AOI221_X1 port map( B1 => OP1(27), B2 => n3, C1 => n7, C2 => n50, A 
                           => n19, ZN => n114);
   U244 : OAI22_X1 port map( A1 => n112, A2 => n163, B1 => n113, B2 => n51, ZN 
                           => LOGIC_RES_28_port);
   U245 : AOI21_X1 port map( B1 => n8, B2 => n163, A => n20, ZN => n113);
   U246 : AOI221_X1 port map( B1 => OP1(28), B2 => n2, C1 => n7, C2 => n51, A 
                           => n19, ZN => n112);
   U247 : OAI22_X1 port map( A1 => n110, A2 => n164, B1 => n111, B2 => n52, ZN 
                           => LOGIC_RES_29_port);
   U248 : AOI21_X1 port map( B1 => n8, B2 => n164, A => n20, ZN => n111);
   U249 : AOI221_X1 port map( B1 => OP1(29), B2 => n2, C1 => n7, C2 => n52, A 
                           => n19, ZN => n110);
   U250 : OAI22_X1 port map( A1 => n106, A2 => n166, B1 => n107, B2 => n54, ZN 
                           => LOGIC_RES_30_port);
   U251 : AOI21_X1 port map( B1 => n8, B2 => n166, A => n20, ZN => n107);
   U252 : AOI221_X1 port map( B1 => OP1(30), B2 => n2, C1 => n7, C2 => n54, A 
                           => n19, ZN => n106);
   U253 : OAI22_X1 port map( A1 => n104, A2 => n167, B1 => n105, B2 => n55, ZN 
                           => LOGIC_RES_31_port);
   U254 : AOI21_X1 port map( B1 => n8, B2 => n167, A => n20, ZN => n105);
   U255 : AOI221_X1 port map( B1 => OP1(31), B2 => n2, C1 => n7, C2 => n55, A 
                           => n19, ZN => n104);
   U256 : INV_X1 port map( A => n85, ZN => n180);
   U257 : INV_X1 port map( A => OPSel_0_port, ZN => n181);
   U258 : INV_X1 port map( A => OP1(10), ZN => n32);
   U259 : INV_X1 port map( A => OP1(16), ZN => n38);
   U260 : INV_X1 port map( A => OP1(20), ZN => n43);
   U261 : INV_X1 port map( A => OP1(4), ZN => n57);
   U262 : INV_X1 port map( A => OP1(12), ZN => n34);
   U263 : INV_X1 port map( A => OP1(21), ZN => n44);
   U264 : INV_X1 port map( A => OP1(13), ZN => n35);
   U265 : INV_X1 port map( A => OP1(22), ZN => n45);
   U266 : INV_X1 port map( A => OP1(14), ZN => n36);
   U267 : INV_X1 port map( A => OP1(0), ZN => n31);
   U268 : INV_X1 port map( A => OP1(1), ZN => n42);
   U269 : INV_X1 port map( A => OP1(2), ZN => n53);
   U270 : INV_X1 port map( A => OP1(17), ZN => n39);
   U271 : INV_X1 port map( A => OP1(18), ZN => n40);
   U272 : INV_X1 port map( A => OP1(5), ZN => n58);
   U273 : INV_X1 port map( A => OP1(6), ZN => n59);
   U274 : INV_X1 port map( A => OP1(24), ZN => n47);
   U275 : INV_X1 port map( A => OP1(25), ZN => n48);
   U276 : INV_X1 port map( A => OP1(28), ZN => n51);
   U277 : INV_X1 port map( A => OP1(29), ZN => n52);
   U278 : INV_X1 port map( A => OP1(30), ZN => n54);
   U279 : INV_X1 port map( A => OP1(8), ZN => n61);
   U280 : INV_X1 port map( A => OP1(9), ZN => n62);
   U281 : INV_X1 port map( A => OP1(26), ZN => n49);
   U282 : INV_X1 port map( A => OP1(3), ZN => n56);
   U283 : INV_X1 port map( A => OP1(7), ZN => n60);
   U284 : INV_X1 port map( A => OP1(11), ZN => n33);
   U285 : INV_X1 port map( A => OP1(15), ZN => n37);
   U286 : INV_X1 port map( A => OP1(19), ZN => n41);
   U287 : INV_X1 port map( A => OP1(23), ZN => n46);
   U288 : INV_X1 port map( A => OP1(27), ZN => n50);
   U289 : INV_X1 port map( A => OP1(31), ZN => n55);
   U290 : INV_X1 port map( A => OP2(1), ZN => n74);
   U291 : INV_X1 port map( A => OP2(0), ZN => n63);
   U292 : INV_X1 port map( A => OP2(2), ZN => n165);
   U293 : INV_X1 port map( A => OP2(6), ZN => n171);
   U294 : INV_X1 port map( A => OP2(5), ZN => n170);
   U295 : INV_X1 port map( A => OP2(4), ZN => n169);
   U296 : INV_X1 port map( A => OP2(13), ZN => n67);
   U297 : INV_X1 port map( A => OP2(14), ZN => n68);
   U298 : INV_X1 port map( A => OP2(12), ZN => n66);
   U299 : INV_X1 port map( A => OP2(16), ZN => n70);
   U300 : INV_X1 port map( A => OP2(17), ZN => n71);
   U301 : INV_X1 port map( A => OP2(8), ZN => n173);
   U302 : INV_X1 port map( A => OP2(9), ZN => n174);
   U303 : INV_X1 port map( A => OP2(10), ZN => n64);
   U304 : INV_X1 port map( A => OP2(18), ZN => n72);
   U305 : INV_X1 port map( A => OP2(21), ZN => n76);
   U306 : INV_X1 port map( A => OP2(20), ZN => n75);
   U307 : INV_X1 port map( A => OP2(30), ZN => n166);
   U308 : INV_X1 port map( A => OP2(29), ZN => n164);
   U309 : INV_X1 port map( A => OP2(24), ZN => n159);
   U310 : INV_X1 port map( A => OP2(22), ZN => n77);
   U311 : INV_X1 port map( A => OP2(25), ZN => n160);
   U312 : INV_X1 port map( A => OP2(26), ZN => n161);
   U313 : INV_X1 port map( A => OP2(28), ZN => n163);
   U314 : INV_X1 port map( A => OP2(3), ZN => n168);
   U315 : INV_X1 port map( A => OP2(7), ZN => n172);
   U316 : INV_X1 port map( A => OP2(11), ZN => n65);
   U325 : INV_X1 port map( A => OP2(15), ZN => n69);
   U326 : INV_X1 port map( A => OP2(19), ZN => n73);
   U327 : INV_X1 port map( A => OP2(23), ZN => n86);
   U328 : INV_X1 port map( A => OP2(27), ZN => n162);
   U329 : INV_X1 port map( A => OP2(31), ZN => n167);
   U330 : AND2_X1 port map( A1 => n154, A2 => n89, ZN => n1);
   U331 : INV_X1 port map( A => n83, ZN => n182);
   U332 : INV_X1 port map( A => LOGIC_ARITH, ZN => n178);
   U333 : NAND2_X1 port map( A1 => n155, A2 => n89, ZN => n82);
   U334 : NAND2_X1 port map( A1 => n155, A2 => n88, ZN => n80);
   U335 : NAND2_X1 port map( A1 => n154, A2 => n88, ZN => n81);
   U336 : INV_X1 port map( A => n84, ZN => n183);
   U337 : NOR2_X1 port map( A1 => n185, A2 => ALU_OPC(1), ZN => n89);
   U338 : NOR2_X1 port map( A1 => n186, A2 => ALU_OPC(0), ZN => n155);
   U339 : NOR2_X1 port map( A1 => n184, A2 => ALU_OPC(2), ZN => n88);
   U340 : NOR2_X1 port map( A1 => ALU_OPC(0), A2 => ALU_OPC(3), ZN => n154);
   U341 : NAND2_X1 port map( A1 => n85, A2 => n157, ZN => LOGIC_ARITH);
   U342 : OAI21_X1 port map( B1 => n78, B2 => n175, A => n79, ZN => 
                           select_zero_sig);
   U343 : INV_X1 port map( A => ALU_OPC(0), ZN => n175);
   U344 : AOI22_X1 port map( A1 => ALU_OPC(3), A2 => n185, B1 => ALU_OPC(1), B2
                           => ALU_OPC(2), ZN => n78);
   U345 : INV_X1 port map( A => ALU_OPC(2), ZN => n185);
   U346 : INV_X1 port map( A => ALU_OPC(3), ZN => n186);
   U347 : INV_X1 port map( A => ALU_OPC(1), ZN => n184);
   U348 : CLKBUF_X1 port map( A => n177, Z => n10);
   U349 : CLKBUF_X1 port map( A => n178, Z => n16);
   U350 : CLKBUF_X1 port map( A => n179, Z => n22);
   U351 : INV_X1 port map( A => n1, ZN => n29);
   U352 : INV_X1 port map( A => n1, ZN => n30);
   COMP_RES_1_port <= '0';
   COMP_RES_2_port <= '0';
   COMP_RES_3_port <= '0';
   COMP_RES_4_port <= '0';
   COMP_RES_5_port <= '0';
   COMP_RES_6_port <= '0';
   COMP_RES_7_port <= '0';
   COMP_RES_8_port <= '0';
   COMP_RES_9_port <= '0';
   COMP_RES_10_port <= '0';
   COMP_RES_11_port <= '0';
   COMP_RES_12_port <= '0';
   COMP_RES_13_port <= '0';
   COMP_RES_14_port <= '0';
   COMP_RES_15_port <= '0';
   COMP_RES_16_port <= '0';
   COMP_RES_17_port <= '0';
   COMP_RES_18_port <= '0';
   COMP_RES_19_port <= '0';
   COMP_RES_20_port <= '0';
   COMP_RES_21_port <= '0';
   COMP_RES_22_port <= '0';
   COMP_RES_23_port <= '0';
   COMP_RES_24_port <= '0';
   COMP_RES_25_port <= '0';
   COMP_RES_26_port <= '0';
   COMP_RES_27_port <= '0';
   COMP_RES_28_port <= '0';
   COMP_RES_29_port <= '0';
   COMP_RES_30_port <= '0';
   COMP_RES_31_port <= '0';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_0 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_0;

architecture SYN_bhv of mux41_NBIT32_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n1, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n6, Z => n72);
   U2 : BUF_X1 port map( A => n6, Z => n73);
   U3 : BUF_X1 port map( A => n4, Z => n78);
   U4 : BUF_X1 port map( A => n4, Z => n79);
   U5 : BUF_X1 port map( A => n7, Z => n1);
   U6 : BUF_X1 port map( A => n7, Z => n70);
   U7 : BUF_X1 port map( A => n5, Z => n75);
   U8 : BUF_X1 port map( A => n5, Z => n76);
   U9 : BUF_X1 port map( A => n6, Z => n74);
   U10 : BUF_X1 port map( A => n4, Z => n80);
   U11 : BUF_X1 port map( A => n7, Z => n71);
   U12 : BUF_X1 port map( A => n5, Z => n77);
   U13 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n6);
   U14 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n7);
   U15 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n4);
   U16 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n5);
   U17 : INV_X1 port map( A => S(0), ZN => n81);
   U18 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => Z(20));
   U19 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN 
                           => n45);
   U20 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN 
                           => n44);
   U21 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => Z(17));
   U22 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n53);
   U23 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n52);
   U24 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => Z(13));
   U25 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN 
                           => n61);
   U26 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n60);
   U27 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => Z(0));
   U28 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n69);
   U29 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n68);
   U30 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => Z(6));
   U31 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n13);
   U32 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n12);
   U33 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => Z(31));
   U34 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN 
                           => n21);
   U35 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN 
                           => n20);
   U36 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => Z(28));
   U37 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n29);
   U38 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n28);
   U39 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => Z(24));
   U40 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN 
                           => n37);
   U41 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN 
                           => n36);
   U42 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => Z(21));
   U43 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n43);
   U44 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n42);
   U45 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => Z(18));
   U46 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n51);
   U47 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n50);
   U48 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => Z(14));
   U49 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN 
                           => n59);
   U50 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n58);
   U51 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => Z(10));
   U52 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN 
                           => n67);
   U53 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n66);
   U54 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => Z(7));
   U55 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n11);
   U56 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n10);
   U57 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => Z(3));
   U58 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN =>
                           n19);
   U59 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN =>
                           n18);
   U60 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => Z(29));
   U61 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n27);
   U62 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n26);
   U63 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => Z(25));
   U64 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n35);
   U65 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n34);
   U66 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => Z(22));
   U67 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n41);
   U68 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n40);
   U69 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => Z(19));
   U70 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN 
                           => n49);
   U71 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n48);
   U72 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => Z(15));
   U73 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN 
                           => n57);
   U74 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n56);
   U75 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => Z(11));
   U76 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN 
                           => n65);
   U77 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n64);
   U78 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => Z(8));
   U79 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n9);
   U80 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n8);
   U81 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => Z(4));
   U82 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN =>
                           n17);
   U83 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN =>
                           n16);
   U84 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => Z(2));
   U85 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN =>
                           n25);
   U86 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN =>
                           n24);
   U87 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => Z(26));
   U88 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n33);
   U89 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n32);
   U90 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => Z(23));
   U91 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN 
                           => n39);
   U92 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN 
                           => n38);
   U93 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => Z(1));
   U94 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN =>
                           n47);
   U95 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN => 
                           n46);
   U96 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => Z(16));
   U97 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n55);
   U98 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n54);
   U99 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => Z(12));
   U100 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN
                           => n63);
   U101 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n62);
   U102 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Z(9));
   U103 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN 
                           => n3);
   U104 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN 
                           => n2);
   U105 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => Z(5));
   U106 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN 
                           => n15);
   U107 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN 
                           => n14);
   U108 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => Z(30));
   U109 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN
                           => n23);
   U110 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN
                           => n22);
   U111 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => Z(27));
   U112 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN
                           => n31);
   U113 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN
                           => n30);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FWD_Unit is

   port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB : in 
         std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;  
         FWDA, FWDB : out std_logic_vector (1 downto 0));

end FWD_Unit;

architecture SYN_bhv of FWD_Unit is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42 : std_logic;

begin
   
   U3 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => FWDB(1));
   U4 : AOI21_X1 port map( B1 => n3, B2 => n4, A => n5, ZN => n1);
   U5 : INV_X1 port map( A => n6, ZN => n3);
   U6 : NOR2_X1 port map( A1 => n2, A2 => n7, ZN => FWDB(0));
   U7 : MUX2_X1 port map( A => n6, B => n8, S => n5, Z => n7);
   U8 : AND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => n5);
   U9 : NOR2_X1 port map( A1 => n13, A2 => n14, ZN => n12);
   U10 : XOR2_X1 port map( A => ADD_WR_MEM(4), B => ADD_RS2(4), Z => n14);
   U11 : XOR2_X1 port map( A => ADD_WR_MEM(3), B => ADD_RS2(3), Z => n13);
   U12 : XNOR2_X1 port map( A => ADD_RS2(1), B => ADD_WR_MEM(1), ZN => n11);
   U13 : XNOR2_X1 port map( A => ADD_RS2(2), B => ADD_WR_MEM(2), ZN => n10);
   U14 : XNOR2_X1 port map( A => ADD_RS2(0), B => ADD_WR_MEM(0), ZN => n9);
   U15 : NAND4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           n6);
   U16 : NOR2_X1 port map( A1 => n19, A2 => n20, ZN => n18);
   U17 : XOR2_X1 port map( A => ADD_WR_WB(3), B => ADD_RS2(3), Z => n20);
   U18 : XOR2_X1 port map( A => ADD_WR_WB(2), B => ADD_RS2(2), Z => n19);
   U19 : XNOR2_X1 port map( A => ADD_RS2(4), B => ADD_WR_WB(4), ZN => n17);
   U20 : XNOR2_X1 port map( A => ADD_RS2(1), B => ADD_WR_WB(1), ZN => n16);
   U21 : XNOR2_X1 port map( A => ADD_RS2(0), B => ADD_WR_WB(0), ZN => n15);
   U22 : NOR2_X1 port map( A1 => n21, A2 => n2, ZN => FWDA(1));
   U23 : AOI21_X1 port map( B1 => n22, B2 => n4, A => n23, ZN => n21);
   U24 : OAI21_X1 port map( B1 => n24, B2 => n25, A => RF_WE_WB, ZN => n4);
   U25 : OR2_X1 port map( A1 => ADD_WR_WB(0), A2 => ADD_WR_WB(1), ZN => n25);
   U26 : OR3_X1 port map( A1 => ADD_WR_WB(3), A2 => ADD_WR_WB(4), A3 => 
                           ADD_WR_WB(2), ZN => n24);
   U27 : INV_X1 port map( A => n26, ZN => n22);
   U28 : NOR2_X1 port map( A1 => n2, A2 => n27, ZN => FWDA(0));
   U29 : MUX2_X1 port map( A => n26, B => n8, S => n23, Z => n27);
   U30 : AND4_X1 port map( A1 => n28, A2 => n29, A3 => n30, A4 => n31, ZN => 
                           n23);
   U31 : NOR2_X1 port map( A1 => n32, A2 => n33, ZN => n31);
   U32 : XOR2_X1 port map( A => ADD_WR_MEM(4), B => ADD_RS1(4), Z => n33);
   U33 : XOR2_X1 port map( A => ADD_WR_MEM(3), B => ADD_RS1(3), Z => n32);
   U34 : XNOR2_X1 port map( A => ADD_RS1(1), B => ADD_WR_MEM(1), ZN => n30);
   U35 : XNOR2_X1 port map( A => ADD_RS1(2), B => ADD_WR_MEM(2), ZN => n29);
   U36 : XNOR2_X1 port map( A => ADD_RS1(0), B => ADD_WR_MEM(0), ZN => n28);
   U37 : INV_X1 port map( A => n34, ZN => n8);
   U38 : OAI21_X1 port map( B1 => n35, B2 => n36, A => RF_WE_MEM, ZN => n34);
   U39 : OR2_X1 port map( A1 => ADD_WR_MEM(0), A2 => ADD_WR_MEM(1), ZN => n36);
   U40 : OR3_X1 port map( A1 => ADD_WR_MEM(3), A2 => ADD_WR_MEM(4), A3 => 
                           ADD_WR_MEM(2), ZN => n35);
   U41 : NAND4_X1 port map( A1 => n37, A2 => n38, A3 => n39, A4 => n40, ZN => 
                           n26);
   U42 : NOR2_X1 port map( A1 => n41, A2 => n42, ZN => n40);
   U43 : XOR2_X1 port map( A => ADD_WR_WB(3), B => ADD_RS1(3), Z => n42);
   U44 : XOR2_X1 port map( A => ADD_WR_WB(2), B => ADD_RS1(2), Z => n41);
   U45 : XNOR2_X1 port map( A => ADD_RS1(4), B => ADD_WR_WB(4), ZN => n39);
   U46 : XNOR2_X1 port map( A => ADD_RS1(1), B => ADD_WR_WB(1), ZN => n38);
   U47 : XNOR2_X1 port map( A => ADD_RS1(0), B => ADD_WR_WB(0), ZN => n37);
   U48 : INV_X1 port map( A => RST, ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N2 is

   port( DIN : in std_logic_vector (1 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (1 downto 0));

end regn_N2;

architecture SYN_bhv of regn_N2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   DOUT_reg_1_inst : DFFR_X1 port map( D => n6, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n4);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n5, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n3);
   U2 : OAI21_X1 port map( B1 => n3, B2 => EN, A => n1, ZN => n5);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n1);
   U4 : OAI21_X1 port map( B1 => n4, B2 => EN, A => n2, ZN => n6);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Branch_Cond_Unit_NBIT32 is

   port( RST : in std_logic;  A : in std_logic_vector (31 downto 0);  ALU_OPC :
         in std_logic_vector (0 to 3);  JUMP_TYPE : in std_logic_vector (1 
         downto 0);  PC_SEL : out std_logic_vector (1 downto 0);  ZERO : out 
         std_logic);

end Branch_Cond_Unit_NBIT32;

architecture SYN_bhv of Branch_Cond_Unit_NBIT32 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n1, n2 : std_logic;

begin
   
   U3 : NOR4_X1 port map( A1 => A(23), A2 => A(22), A3 => A(21), A4 => A(20), 
                           ZN => n15);
   U4 : NOR4_X1 port map( A1 => A(9), A2 => A(8), A3 => A(7), A4 => A(6), ZN =>
                           n19);
   U5 : NAND4_X1 port map( A1 => n12, A2 => n13, A3 => n14, A4 => n15, ZN => 
                           n11);
   U6 : NOR4_X1 port map( A1 => A(12), A2 => A(11), A3 => A(10), A4 => A(0), ZN
                           => n12);
   U7 : NOR4_X1 port map( A1 => A(16), A2 => A(15), A3 => A(14), A4 => A(13), 
                           ZN => n13);
   U8 : NOR4_X1 port map( A1 => A(1), A2 => A(19), A3 => A(18), A4 => A(17), ZN
                           => n14);
   U9 : NAND4_X1 port map( A1 => n16, A2 => n17, A3 => n18, A4 => n19, ZN => 
                           n10);
   U10 : NOR4_X1 port map( A1 => A(27), A2 => A(26), A3 => A(25), A4 => A(24), 
                           ZN => n16);
   U11 : NOR4_X1 port map( A1 => A(30), A2 => A(2), A3 => A(29), A4 => A(28), 
                           ZN => n17);
   U12 : NOR4_X1 port map( A1 => A(5), A2 => A(4), A3 => A(3), A4 => A(31), ZN 
                           => n18);
   U13 : NOR4_X1 port map( A1 => ALU_OPC(3), A2 => n1, A3 => ALU_OPC(1), A4 => 
                           ALU_OPC(2), ZN => n7);
   U14 : OAI211_X1 port map( C1 => n5, C2 => n6, A => JUMP_TYPE(0), B => RST, 
                           ZN => n4);
   U15 : AND2_X1 port map( A1 => n7, A2 => n8, ZN => n6);
   U16 : NOR4_X1 port map( A1 => n8, A2 => n9, A3 => n7, A4 => n1, ZN => n5);
   U17 : NOR2_X1 port map( A1 => n10, A2 => n11, ZN => n8);
   U18 : NAND2_X1 port map( A1 => JUMP_TYPE(1), A2 => RST, ZN => n3);
   U19 : INV_X1 port map( A => ALU_OPC(0), ZN => n1);
   U20 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => ZERO);
   U21 : OAI22_X1 port map( A1 => JUMP_TYPE(0), A2 => n3, B1 => JUMP_TYPE(1), 
                           B2 => n4, ZN => PC_SEL(0));
   U22 : NOR2_X1 port map( A1 => n2, A2 => n3, ZN => PC_SEL(1));
   U23 : INV_X1 port map( A => JUMP_TYPE(0), ZN => n2);
   U24 : OR2_X1 port map( A1 => ALU_OPC(2), A2 => ALU_OPC(1), ZN => n9);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity register_file_NBIT_ADD5_NBIT_DATA32 is

   port( CLK, RST, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RS1, 
         ADD_RS2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_NBIT_ADD5_NBIT_DATA32;

architecture SYN_bhv of register_file_NBIT_ADD5_NBIT_DATA32 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
      n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, 
      n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, 
      n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, 
      n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, 
      n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, 
      n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, 
      n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, 
      n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, 
      n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, 
      n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, 
      n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, 
      n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, 
      n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, 
      n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, 
      n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, 
      n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, 
      n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, 
      n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, 
      n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, 
      n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, 
      n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, 
      n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, 
      n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
      n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, 
      n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, 
      n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, 
      n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, 
      n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, 
      n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, 
      n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, 
      n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, 
      n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, 
      n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, 
      n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, 
      n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, 
      n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, 
      n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, 
      n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, 
      n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, 
      n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, 
      n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, 
      n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, 
      n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, 
      n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, 
      n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, 
      n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, 
      n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, 
      n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, 
      n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, 
      n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, 
      n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
      n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, 
      n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, 
      n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, 
      n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, 
      n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, 
      n3553, n3554, n3555, n3556, n3557, n3558, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
      n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
      n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
      n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
      n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
      n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
      n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
      n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
      n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, 
      n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, 
      n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, 
      n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, 
      n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, 
      n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, 
      n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, 
      n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, 
      n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, 
      n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, 
      n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, 
      n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, 
      n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, 
      n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
      n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, 
      n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, 
      n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, 
      n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, 
      n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, 
      n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, 
      n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, 
      n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, 
      n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, 
      n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, 
      n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, 
      n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, 
      n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, 
      n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, 
      n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, 
      n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, 
      n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, 
      n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, 
      n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, 
      n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, 
      n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, 
      n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, 
      n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, 
      n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, 
      n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, 
      n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, 
      n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, 
      n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, 
      n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, 
      n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, 
      n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, 
      n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, 
      n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, 
      n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, 
      n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, 
      n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, 
      n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, 
      n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, 
      n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, 
      n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, 
      n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, 
      n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
      n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
      n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, 
      n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, 
      n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, 
      n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, 
      n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, 
      n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, 
      n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, 
      n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, 
      n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, 
      n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, 
      n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, 
      n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, 
      n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, 
      n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, 
      n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, 
      n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, 
      n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, 
      n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, 
      n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, 
      n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, 
      n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
      n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, 
      n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, 
      n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, 
      n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, 
      n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, 
      n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, 
      n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, 
      n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, 
      n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, 
      n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, 
      n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, 
      n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, 
      n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, 
      n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, 
      n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, 
      n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, 
      n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, 
      n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, 
      n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, 
      n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, 
      n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, 
      n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, 
      n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, 
      n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, 
      n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, 
      n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, 
      n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, 
      n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, 
      n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, 
      n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, 
      n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, 
      n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, 
      n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, 
      n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, 
      n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, 
      n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, 
      n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, 
      n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, 
      n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, 
      n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, 
      n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, 
      n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, 
      n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, 
      n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, 
      n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, 
      n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, 
      n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, 
      n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, 
      n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, 
      n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, 
      n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, 
      n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, 
      n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, 
      n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, 
      n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, 
      n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, 
      n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, 
      n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, 
      n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, 
      n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, 
      n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, 
      n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, 
      n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, 
      n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, 
      n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, 
      n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, 
      n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, 
      n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, 
      n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, 
      n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, 
      n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, 
      n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, 
      n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, 
      n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
      n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
      n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
      n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, 
      n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
      n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
      n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, 
      n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, 
      n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, 
      n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, 
      n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
      n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, 
      n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, 
      n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, 
      n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
      n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, 
      n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, 
      n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, 
      n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, 
      n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, 
      n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, 
      n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, 
      n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, 
      n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, 
      n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, 
      n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, 
      n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, 
      n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, 
      n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, 
      n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, 
      n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, 
      n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, 
      n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, 
      n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, 
      n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, 
      n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, 
      n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, 
      n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, 
      n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, 
      n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, 
      n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, 
      n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, 
      n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, 
      n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, 
      n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, 
      n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, 
      n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, 
      n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, 
      n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, 
      n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, 
      n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, 
      n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, 
      n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, 
      n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, 
      n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, 
      n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, 
      n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, 
      n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, 
      n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, 
      n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, 
      n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, 
      n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, 
      n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, 
      n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, 
      n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, 
      n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, 
      n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, 
      n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, 
      n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, 
      n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, 
      n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, 
      n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, 
      n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, 
      n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, 
      n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, 
      n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, 
      n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, 
      n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, 
      n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, 
      n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, 
      n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, 
      n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, 
      n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, 
      n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, 
      n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, 
      n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, 
      n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, 
      n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, 
      n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, 
      n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, 
      n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, 
      n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, 
      n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, 
      n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, 
      n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, 
      n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, 
      n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, 
      n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, 
      n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, 
      n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, 
      n2978, n2979, n2980, n2981, n2982, n3559, n3560, n3561, n3562, n3563, 
      n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, 
      n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, 
      n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, 
      n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, 
      n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, 
      n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, 
      n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, 
      n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, 
      n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, 
      n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, 
      n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, 
      n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, 
      n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, 
      n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, 
      n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, 
      n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, 
      n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, 
      n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, 
      n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, 
      n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, 
      n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, 
      n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, 
      n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, 
      n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, 
      n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, 
      n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, 
      n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, 
      n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, 
      n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, 
      n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, 
      n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, 
      n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, 
      n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, 
      n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, 
      n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, 
      n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, 
      n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, 
      n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, 
      n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, 
      n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, 
      n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, 
      n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, 
      n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, 
      n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, 
      n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, 
      n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, 
      n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, 
      n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, 
      n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, 
      n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, 
      n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, 
      n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, 
      n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, 
      n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, 
      n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, 
      n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, 
      n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, 
      n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, 
      n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, 
      n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, 
      n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, 
      n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, 
      n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, 
      n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, 
      n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, 
      n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, 
      n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, 
      n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, 
      n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, 
      n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, 
      n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, 
      n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, 
      n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, 
      n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, 
      n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, 
      n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, 
      n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, 
      n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, 
      n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, 
      n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, 
      n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, 
      n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, 
      n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, 
      n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, 
      n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, 
      n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, 
      n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, 
      n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, 
      n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, 
      n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, 
      n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, 
      n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, 
      n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, 
      n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, 
      n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, 
      n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, 
      n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, 
      n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, 
      n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, 
      n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, 
      n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, 
      n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, 
      n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, 
      n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, 
      n4604, n4605, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, 
      n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, 
      n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, 
      n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, 
      n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, 
      n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, 
      n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, 
      n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, 
      n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, 
      n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, 
      n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, 
      n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, 
      n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, 
      n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, 
      n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, 
      n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, 
      n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, 
      n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, 
      n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, 
      n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, 
      n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, 
      n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, 
      n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, 
      n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, 
      n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, 
      n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, 
      n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, 
      n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, 
      n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, 
      n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, 
      n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, 
      n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, 
      n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, 
      n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, 
      n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, 
      n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, 
      n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, 
      n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, 
      n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, 
      n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, 
      n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, 
      n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, 
      n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, 
      n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, 
      n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, 
      n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, 
      n_1815, n_1816, n_1817, n_1818 : std_logic;

begin
   
   REGISTERS_reg_10_31_inst : DFFR_X1 port map( D => n3430, CK => CLK, RN => 
                           n434, Q => n2662, QN => n_1403);
   REGISTERS_reg_10_30_inst : DFFR_X1 port map( D => n3429, CK => CLK, RN => 
                           n434, Q => n2685, QN => n_1404);
   REGISTERS_reg_10_29_inst : DFFR_X1 port map( D => n3428, CK => CLK, RN => 
                           n434, Q => n2708, QN => n_1405);
   REGISTERS_reg_10_28_inst : DFFR_X1 port map( D => n3427, CK => CLK, RN => 
                           n434, Q => n2731, QN => n_1406);
   REGISTERS_reg_10_27_inst : DFFR_X1 port map( D => n3426, CK => CLK, RN => 
                           n434, Q => n2754, QN => n_1407);
   REGISTERS_reg_10_26_inst : DFFR_X1 port map( D => n3425, CK => CLK, RN => 
                           n434, Q => n2777, QN => n_1408);
   REGISTERS_reg_10_25_inst : DFFR_X1 port map( D => n3424, CK => CLK, RN => 
                           n434, Q => n2800, QN => n_1409);
   REGISTERS_reg_10_24_inst : DFFR_X1 port map( D => n3423, CK => CLK, RN => 
                           n434, Q => n2823, QN => n_1410);
   REGISTERS_reg_10_23_inst : DFFR_X1 port map( D => n3422, CK => CLK, RN => 
                           n434, Q => n2846, QN => n_1411);
   REGISTERS_reg_10_22_inst : DFFR_X1 port map( D => n3421, CK => CLK, RN => 
                           n434, Q => n2869, QN => n_1412);
   REGISTERS_reg_10_21_inst : DFFR_X1 port map( D => n3420, CK => CLK, RN => 
                           n434, Q => n2892, QN => n_1413);
   REGISTERS_reg_10_20_inst : DFFR_X1 port map( D => n3419, CK => CLK, RN => 
                           n434, Q => n2915, QN => n_1414);
   REGISTERS_reg_10_19_inst : DFFR_X1 port map( D => n3418, CK => CLK, RN => 
                           n435, Q => n2938, QN => n_1415);
   REGISTERS_reg_10_18_inst : DFFR_X1 port map( D => n3417, CK => CLK, RN => 
                           n435, Q => n2961, QN => n_1416);
   REGISTERS_reg_10_17_inst : DFFR_X1 port map( D => n3416, CK => CLK, RN => 
                           n435, Q => n3560, QN => n_1417);
   REGISTERS_reg_10_16_inst : DFFR_X1 port map( D => n3415, CK => CLK, RN => 
                           n435, Q => n3583, QN => n_1418);
   REGISTERS_reg_10_15_inst : DFFR_X1 port map( D => n3414, CK => CLK, RN => 
                           n435, Q => n3606, QN => n_1419);
   REGISTERS_reg_10_14_inst : DFFR_X1 port map( D => n3413, CK => CLK, RN => 
                           n435, Q => n3629, QN => n_1420);
   REGISTERS_reg_10_13_inst : DFFR_X1 port map( D => n3412, CK => CLK, RN => 
                           n435, Q => n3652, QN => n_1421);
   REGISTERS_reg_10_12_inst : DFFR_X1 port map( D => n3411, CK => CLK, RN => 
                           n435, Q => n3675, QN => n_1422);
   REGISTERS_reg_10_11_inst : DFFR_X1 port map( D => n3410, CK => CLK, RN => 
                           n435, Q => n3698, QN => n_1423);
   REGISTERS_reg_10_10_inst : DFFR_X1 port map( D => n3409, CK => CLK, RN => 
                           n435, Q => n3721, QN => n_1424);
   REGISTERS_reg_10_9_inst : DFFR_X1 port map( D => n3408, CK => CLK, RN => 
                           n435, Q => n3744, QN => n_1425);
   REGISTERS_reg_10_8_inst : DFFR_X1 port map( D => n3407, CK => CLK, RN => 
                           n435, Q => n3767, QN => n_1426);
   REGISTERS_reg_10_7_inst : DFFR_X1 port map( D => n3406, CK => CLK, RN => 
                           n436, Q => n3790, QN => n_1427);
   REGISTERS_reg_10_6_inst : DFFR_X1 port map( D => n3405, CK => CLK, RN => 
                           n436, Q => n3813, QN => n_1428);
   REGISTERS_reg_10_5_inst : DFFR_X1 port map( D => n3404, CK => CLK, RN => 
                           n436, Q => n3836, QN => n_1429);
   REGISTERS_reg_10_4_inst : DFFR_X1 port map( D => n3403, CK => CLK, RN => 
                           n436, Q => n3859, QN => n_1430);
   REGISTERS_reg_10_3_inst : DFFR_X1 port map( D => n3402, CK => CLK, RN => 
                           n436, Q => n3882, QN => n_1431);
   REGISTERS_reg_10_2_inst : DFFR_X1 port map( D => n3401, CK => CLK, RN => 
                           n436, Q => n3905, QN => n_1432);
   REGISTERS_reg_10_1_inst : DFFR_X1 port map( D => n3400, CK => CLK, RN => 
                           n436, Q => n3928, QN => n_1433);
   REGISTERS_reg_10_0_inst : DFFR_X1 port map( D => n3399, CK => CLK, RN => 
                           n436, Q => n3951, QN => n_1434);
   REGISTERS_reg_11_31_inst : DFFR_X1 port map( D => n3398, CK => CLK, RN => 
                           n436, Q => n2661, QN => n_1435);
   REGISTERS_reg_11_30_inst : DFFR_X1 port map( D => n3397, CK => CLK, RN => 
                           n436, Q => n2684, QN => n_1436);
   REGISTERS_reg_11_29_inst : DFFR_X1 port map( D => n3396, CK => CLK, RN => 
                           n436, Q => n2707, QN => n_1437);
   REGISTERS_reg_11_28_inst : DFFR_X1 port map( D => n3395, CK => CLK, RN => 
                           n436, Q => n2730, QN => n_1438);
   REGISTERS_reg_11_27_inst : DFFR_X1 port map( D => n3394, CK => CLK, RN => 
                           n437, Q => n2753, QN => n_1439);
   REGISTERS_reg_11_26_inst : DFFR_X1 port map( D => n3393, CK => CLK, RN => 
                           n437, Q => n2776, QN => n_1440);
   REGISTERS_reg_11_25_inst : DFFR_X1 port map( D => n3392, CK => CLK, RN => 
                           n437, Q => n2799, QN => n_1441);
   REGISTERS_reg_11_24_inst : DFFR_X1 port map( D => n3391, CK => CLK, RN => 
                           n437, Q => n2822, QN => n_1442);
   REGISTERS_reg_11_23_inst : DFFR_X1 port map( D => n3390, CK => CLK, RN => 
                           n437, Q => n2845, QN => n_1443);
   REGISTERS_reg_11_22_inst : DFFR_X1 port map( D => n3389, CK => CLK, RN => 
                           n437, Q => n2868, QN => n_1444);
   REGISTERS_reg_11_21_inst : DFFR_X1 port map( D => n3388, CK => CLK, RN => 
                           n437, Q => n2891, QN => n_1445);
   REGISTERS_reg_11_20_inst : DFFR_X1 port map( D => n3387, CK => CLK, RN => 
                           n437, Q => n2914, QN => n_1446);
   REGISTERS_reg_11_19_inst : DFFR_X1 port map( D => n3386, CK => CLK, RN => 
                           n437, Q => n2937, QN => n_1447);
   REGISTERS_reg_11_18_inst : DFFR_X1 port map( D => n3385, CK => CLK, RN => 
                           n437, Q => n2960, QN => n_1448);
   REGISTERS_reg_11_17_inst : DFFR_X1 port map( D => n3384, CK => CLK, RN => 
                           n437, Q => n3559, QN => n_1449);
   REGISTERS_reg_11_16_inst : DFFR_X1 port map( D => n3383, CK => CLK, RN => 
                           n437, Q => n3582, QN => n_1450);
   REGISTERS_reg_11_15_inst : DFFR_X1 port map( D => n3382, CK => CLK, RN => 
                           n438, Q => n3605, QN => n_1451);
   REGISTERS_reg_11_14_inst : DFFR_X1 port map( D => n3381, CK => CLK, RN => 
                           n438, Q => n3628, QN => n_1452);
   REGISTERS_reg_11_13_inst : DFFR_X1 port map( D => n3380, CK => CLK, RN => 
                           n438, Q => n3651, QN => n_1453);
   REGISTERS_reg_11_12_inst : DFFR_X1 port map( D => n3379, CK => CLK, RN => 
                           n438, Q => n3674, QN => n_1454);
   REGISTERS_reg_11_11_inst : DFFR_X1 port map( D => n3378, CK => CLK, RN => 
                           n438, Q => n3697, QN => n_1455);
   REGISTERS_reg_11_10_inst : DFFR_X1 port map( D => n3377, CK => CLK, RN => 
                           n438, Q => n3720, QN => n_1456);
   REGISTERS_reg_11_9_inst : DFFR_X1 port map( D => n3376, CK => CLK, RN => 
                           n438, Q => n3743, QN => n_1457);
   REGISTERS_reg_11_8_inst : DFFR_X1 port map( D => n3375, CK => CLK, RN => 
                           n438, Q => n3766, QN => n_1458);
   REGISTERS_reg_11_7_inst : DFFR_X1 port map( D => n3374, CK => CLK, RN => 
                           n438, Q => n3789, QN => n_1459);
   REGISTERS_reg_11_6_inst : DFFR_X1 port map( D => n3373, CK => CLK, RN => 
                           n438, Q => n3812, QN => n_1460);
   REGISTERS_reg_11_5_inst : DFFR_X1 port map( D => n3372, CK => CLK, RN => 
                           n438, Q => n3835, QN => n_1461);
   REGISTERS_reg_11_4_inst : DFFR_X1 port map( D => n3371, CK => CLK, RN => 
                           n438, Q => n3858, QN => n_1462);
   REGISTERS_reg_11_3_inst : DFFR_X1 port map( D => n3370, CK => CLK, RN => 
                           n439, Q => n3881, QN => n_1463);
   REGISTERS_reg_11_2_inst : DFFR_X1 port map( D => n3369, CK => CLK, RN => 
                           n439, Q => n3904, QN => n_1464);
   REGISTERS_reg_11_1_inst : DFFR_X1 port map( D => n3368, CK => CLK, RN => 
                           n439, Q => n3927, QN => n_1465);
   REGISTERS_reg_11_0_inst : DFFR_X1 port map( D => n3367, CK => CLK, RN => 
                           n439, Q => n3950, QN => n_1466);
   REGISTERS_reg_14_31_inst : DFFR_X1 port map( D => n3366, CK => CLK, RN => 
                           n444, Q => n2658, QN => n_1467);
   REGISTERS_reg_14_30_inst : DFFR_X1 port map( D => n3365, CK => CLK, RN => 
                           n444, Q => n2681, QN => n_1468);
   REGISTERS_reg_14_29_inst : DFFR_X1 port map( D => n3364, CK => CLK, RN => 
                           n444, Q => n2704, QN => n_1469);
   REGISTERS_reg_14_28_inst : DFFR_X1 port map( D => n3363, CK => CLK, RN => 
                           n444, Q => n2727, QN => n_1470);
   REGISTERS_reg_14_27_inst : DFFR_X1 port map( D => n3362, CK => CLK, RN => 
                           n445, Q => n2750, QN => n_1471);
   REGISTERS_reg_14_26_inst : DFFR_X1 port map( D => n3361, CK => CLK, RN => 
                           n445, Q => n2773, QN => n_1472);
   REGISTERS_reg_14_25_inst : DFFR_X1 port map( D => n3360, CK => CLK, RN => 
                           n445, Q => n2796, QN => n_1473);
   REGISTERS_reg_14_24_inst : DFFR_X1 port map( D => n3359, CK => CLK, RN => 
                           n445, Q => n2819, QN => n_1474);
   REGISTERS_reg_14_23_inst : DFFR_X1 port map( D => n3358, CK => CLK, RN => 
                           n445, Q => n2842, QN => n_1475);
   REGISTERS_reg_14_22_inst : DFFR_X1 port map( D => n3357, CK => CLK, RN => 
                           n445, Q => n2865, QN => n_1476);
   REGISTERS_reg_14_21_inst : DFFR_X1 port map( D => n3356, CK => CLK, RN => 
                           n445, Q => n2888, QN => n_1477);
   REGISTERS_reg_14_20_inst : DFFR_X1 port map( D => n3355, CK => CLK, RN => 
                           n445, Q => n2911, QN => n_1478);
   REGISTERS_reg_14_19_inst : DFFR_X1 port map( D => n3354, CK => CLK, RN => 
                           n445, Q => n2934, QN => n_1479);
   REGISTERS_reg_14_18_inst : DFFR_X1 port map( D => n3353, CK => CLK, RN => 
                           n445, Q => n2957, QN => n_1480);
   REGISTERS_reg_14_17_inst : DFFR_X1 port map( D => n3352, CK => CLK, RN => 
                           n445, Q => n2980, QN => n_1481);
   REGISTERS_reg_14_16_inst : DFFR_X1 port map( D => n3351, CK => CLK, RN => 
                           n445, Q => n3579, QN => n_1482);
   REGISTERS_reg_14_15_inst : DFFR_X1 port map( D => n3350, CK => CLK, RN => 
                           n446, Q => n3602, QN => n_1483);
   REGISTERS_reg_14_14_inst : DFFR_X1 port map( D => n3349, CK => CLK, RN => 
                           n446, Q => n3625, QN => n_1484);
   REGISTERS_reg_14_13_inst : DFFR_X1 port map( D => n3348, CK => CLK, RN => 
                           n446, Q => n3648, QN => n_1485);
   REGISTERS_reg_14_12_inst : DFFR_X1 port map( D => n3347, CK => CLK, RN => 
                           n446, Q => n3671, QN => n_1486);
   REGISTERS_reg_14_11_inst : DFFR_X1 port map( D => n3346, CK => CLK, RN => 
                           n446, Q => n3694, QN => n_1487);
   REGISTERS_reg_14_10_inst : DFFR_X1 port map( D => n3345, CK => CLK, RN => 
                           n446, Q => n3717, QN => n_1488);
   REGISTERS_reg_14_9_inst : DFFR_X1 port map( D => n3344, CK => CLK, RN => 
                           n446, Q => n3740, QN => n_1489);
   REGISTERS_reg_14_8_inst : DFFR_X1 port map( D => n3343, CK => CLK, RN => 
                           n446, Q => n3763, QN => n_1490);
   REGISTERS_reg_14_7_inst : DFFR_X1 port map( D => n3342, CK => CLK, RN => 
                           n446, Q => n3786, QN => n_1491);
   REGISTERS_reg_14_6_inst : DFFR_X1 port map( D => n3341, CK => CLK, RN => 
                           n446, Q => n3809, QN => n_1492);
   REGISTERS_reg_14_5_inst : DFFR_X1 port map( D => n3340, CK => CLK, RN => 
                           n446, Q => n3832, QN => n_1493);
   REGISTERS_reg_14_4_inst : DFFR_X1 port map( D => n3339, CK => CLK, RN => 
                           n446, Q => n3855, QN => n_1494);
   REGISTERS_reg_14_3_inst : DFFR_X1 port map( D => n3338, CK => CLK, RN => 
                           n447, Q => n3878, QN => n_1495);
   REGISTERS_reg_14_2_inst : DFFR_X1 port map( D => n3337, CK => CLK, RN => 
                           n447, Q => n3901, QN => n_1496);
   REGISTERS_reg_14_1_inst : DFFR_X1 port map( D => n3336, CK => CLK, RN => 
                           n447, Q => n3924, QN => n_1497);
   REGISTERS_reg_14_0_inst : DFFR_X1 port map( D => n3335, CK => CLK, RN => 
                           n447, Q => n3947, QN => n_1498);
   REGISTERS_reg_15_31_inst : DFFR_X1 port map( D => n3334, CK => CLK, RN => 
                           n447, Q => n2657, QN => n_1499);
   REGISTERS_reg_15_30_inst : DFFR_X1 port map( D => n3333, CK => CLK, RN => 
                           n447, Q => n2680, QN => n_1500);
   REGISTERS_reg_15_29_inst : DFFR_X1 port map( D => n3332, CK => CLK, RN => 
                           n447, Q => n2703, QN => n_1501);
   REGISTERS_reg_15_28_inst : DFFR_X1 port map( D => n3331, CK => CLK, RN => 
                           n447, Q => n2726, QN => n_1502);
   REGISTERS_reg_15_27_inst : DFFR_X1 port map( D => n3330, CK => CLK, RN => 
                           n447, Q => n2749, QN => n_1503);
   REGISTERS_reg_15_26_inst : DFFR_X1 port map( D => n3329, CK => CLK, RN => 
                           n447, Q => n2772, QN => n_1504);
   REGISTERS_reg_15_25_inst : DFFR_X1 port map( D => n3328, CK => CLK, RN => 
                           n447, Q => n2795, QN => n_1505);
   REGISTERS_reg_15_24_inst : DFFR_X1 port map( D => n3327, CK => CLK, RN => 
                           n447, Q => n2818, QN => n_1506);
   REGISTERS_reg_15_23_inst : DFFR_X1 port map( D => n3326, CK => CLK, RN => 
                           n448, Q => n2841, QN => n_1507);
   REGISTERS_reg_15_22_inst : DFFR_X1 port map( D => n3325, CK => CLK, RN => 
                           n448, Q => n2864, QN => n_1508);
   REGISTERS_reg_15_21_inst : DFFR_X1 port map( D => n3324, CK => CLK, RN => 
                           n448, Q => n2887, QN => n_1509);
   REGISTERS_reg_15_20_inst : DFFR_X1 port map( D => n3323, CK => CLK, RN => 
                           n448, Q => n2910, QN => n_1510);
   REGISTERS_reg_15_19_inst : DFFR_X1 port map( D => n3322, CK => CLK, RN => 
                           n448, Q => n2933, QN => n_1511);
   REGISTERS_reg_15_18_inst : DFFR_X1 port map( D => n3321, CK => CLK, RN => 
                           n448, Q => n2956, QN => n_1512);
   REGISTERS_reg_15_17_inst : DFFR_X1 port map( D => n3320, CK => CLK, RN => 
                           n448, Q => n2979, QN => n_1513);
   REGISTERS_reg_15_16_inst : DFFR_X1 port map( D => n3319, CK => CLK, RN => 
                           n448, Q => n3578, QN => n_1514);
   REGISTERS_reg_15_15_inst : DFFR_X1 port map( D => n3318, CK => CLK, RN => 
                           n448, Q => n3601, QN => n_1515);
   REGISTERS_reg_15_14_inst : DFFR_X1 port map( D => n3317, CK => CLK, RN => 
                           n448, Q => n3624, QN => n_1516);
   REGISTERS_reg_15_13_inst : DFFR_X1 port map( D => n3316, CK => CLK, RN => 
                           n448, Q => n3647, QN => n_1517);
   REGISTERS_reg_15_12_inst : DFFR_X1 port map( D => n3315, CK => CLK, RN => 
                           n448, Q => n3670, QN => n_1518);
   REGISTERS_reg_15_11_inst : DFFR_X1 port map( D => n3314, CK => CLK, RN => 
                           n449, Q => n3693, QN => n_1519);
   REGISTERS_reg_15_10_inst : DFFR_X1 port map( D => n3313, CK => CLK, RN => 
                           n449, Q => n3716, QN => n_1520);
   REGISTERS_reg_15_9_inst : DFFR_X1 port map( D => n3312, CK => CLK, RN => 
                           n449, Q => n3739, QN => n_1521);
   REGISTERS_reg_15_8_inst : DFFR_X1 port map( D => n3311, CK => CLK, RN => 
                           n449, Q => n3762, QN => n_1522);
   REGISTERS_reg_15_7_inst : DFFR_X1 port map( D => n3310, CK => CLK, RN => 
                           n449, Q => n3785, QN => n_1523);
   REGISTERS_reg_15_6_inst : DFFR_X1 port map( D => n3309, CK => CLK, RN => 
                           n449, Q => n3808, QN => n_1524);
   REGISTERS_reg_15_5_inst : DFFR_X1 port map( D => n3308, CK => CLK, RN => 
                           n449, Q => n3831, QN => n_1525);
   REGISTERS_reg_15_4_inst : DFFR_X1 port map( D => n3307, CK => CLK, RN => 
                           n449, Q => n3854, QN => n_1526);
   REGISTERS_reg_15_3_inst : DFFR_X1 port map( D => n3306, CK => CLK, RN => 
                           n449, Q => n3877, QN => n_1527);
   REGISTERS_reg_15_2_inst : DFFR_X1 port map( D => n3305, CK => CLK, RN => 
                           n449, Q => n3900, QN => n_1528);
   REGISTERS_reg_15_1_inst : DFFR_X1 port map( D => n3304, CK => CLK, RN => 
                           n449, Q => n3923, QN => n_1529);
   REGISTERS_reg_15_0_inst : DFFR_X1 port map( D => n3303, CK => CLK, RN => 
                           n449, Q => n3946, QN => n_1530);
   REGISTERS_reg_18_30_inst : DFFR_X1 port map( D => n3301, CK => CLK, RN => 
                           n455, Q => n2699, QN => n_1531);
   REGISTERS_reg_18_29_inst : DFFR_X1 port map( D => n3300, CK => CLK, RN => 
                           n455, Q => n2722, QN => n_1532);
   REGISTERS_reg_18_28_inst : DFFR_X1 port map( D => n3299, CK => CLK, RN => 
                           n455, Q => n2745, QN => n_1533);
   REGISTERS_reg_18_27_inst : DFFR_X1 port map( D => n3298, CK => CLK, RN => 
                           n455, Q => n2768, QN => n_1534);
   REGISTERS_reg_18_26_inst : DFFR_X1 port map( D => n3297, CK => CLK, RN => 
                           n455, Q => n2791, QN => n_1535);
   REGISTERS_reg_18_25_inst : DFFR_X1 port map( D => n3296, CK => CLK, RN => 
                           n455, Q => n2814, QN => n_1536);
   REGISTERS_reg_18_24_inst : DFFR_X1 port map( D => n3295, CK => CLK, RN => 
                           n455, Q => n2837, QN => n_1537);
   REGISTERS_reg_18_23_inst : DFFR_X1 port map( D => n3294, CK => CLK, RN => 
                           n456, Q => n2860, QN => n_1538);
   REGISTERS_reg_18_22_inst : DFFR_X1 port map( D => n3293, CK => CLK, RN => 
                           n456, Q => n2883, QN => n_1539);
   REGISTERS_reg_18_21_inst : DFFR_X1 port map( D => n3292, CK => CLK, RN => 
                           n456, Q => n2906, QN => n_1540);
   REGISTERS_reg_18_20_inst : DFFR_X1 port map( D => n3291, CK => CLK, RN => 
                           n456, Q => n2929, QN => n_1541);
   REGISTERS_reg_18_19_inst : DFFR_X1 port map( D => n3290, CK => CLK, RN => 
                           n456, Q => n2952, QN => n_1542);
   REGISTERS_reg_18_18_inst : DFFR_X1 port map( D => n3289, CK => CLK, RN => 
                           n456, Q => n2975, QN => n_1543);
   REGISTERS_reg_18_17_inst : DFFR_X1 port map( D => n3288, CK => CLK, RN => 
                           n456, Q => n3574, QN => n_1544);
   REGISTERS_reg_18_16_inst : DFFR_X1 port map( D => n3287, CK => CLK, RN => 
                           n456, Q => n3597, QN => n_1545);
   REGISTERS_reg_18_15_inst : DFFR_X1 port map( D => n3286, CK => CLK, RN => 
                           n456, Q => n3620, QN => n_1546);
   REGISTERS_reg_18_14_inst : DFFR_X1 port map( D => n3285, CK => CLK, RN => 
                           n456, Q => n3643, QN => n_1547);
   REGISTERS_reg_18_13_inst : DFFR_X1 port map( D => n3284, CK => CLK, RN => 
                           n456, Q => n3666, QN => n_1548);
   REGISTERS_reg_18_12_inst : DFFR_X1 port map( D => n3283, CK => CLK, RN => 
                           n456, Q => n3689, QN => n_1549);
   REGISTERS_reg_18_11_inst : DFFR_X1 port map( D => n3282, CK => CLK, RN => 
                           n457, Q => n3712, QN => n_1550);
   REGISTERS_reg_18_10_inst : DFFR_X1 port map( D => n3281, CK => CLK, RN => 
                           n457, Q => n3735, QN => n_1551);
   REGISTERS_reg_18_9_inst : DFFR_X1 port map( D => n3280, CK => CLK, RN => 
                           n457, Q => n3758, QN => n_1552);
   REGISTERS_reg_18_8_inst : DFFR_X1 port map( D => n3279, CK => CLK, RN => 
                           n457, Q => n3781, QN => n_1553);
   REGISTERS_reg_18_7_inst : DFFR_X1 port map( D => n3278, CK => CLK, RN => 
                           n457, Q => n3804, QN => n_1554);
   REGISTERS_reg_18_6_inst : DFFR_X1 port map( D => n3277, CK => CLK, RN => 
                           n457, Q => n3827, QN => n_1555);
   REGISTERS_reg_18_5_inst : DFFR_X1 port map( D => n3276, CK => CLK, RN => 
                           n457, Q => n3850, QN => n_1556);
   REGISTERS_reg_18_4_inst : DFFR_X1 port map( D => n3275, CK => CLK, RN => 
                           n457, Q => n3873, QN => n_1557);
   REGISTERS_reg_18_3_inst : DFFR_X1 port map( D => n3274, CK => CLK, RN => 
                           n457, Q => n3896, QN => n_1558);
   REGISTERS_reg_18_2_inst : DFFR_X1 port map( D => n3273, CK => CLK, RN => 
                           n457, Q => n3919, QN => n_1559);
   REGISTERS_reg_18_1_inst : DFFR_X1 port map( D => n3272, CK => CLK, RN => 
                           n457, Q => n3942, QN => n_1560);
   REGISTERS_reg_18_0_inst : DFFR_X1 port map( D => n3271, CK => CLK, RN => 
                           n457, Q => n3965, QN => n_1561);
   REGISTERS_reg_19_31_inst : DFFR_X1 port map( D => n3270, CK => CLK, RN => 
                           n458, Q => n2675, QN => n_1562);
   REGISTERS_reg_19_30_inst : DFFR_X1 port map( D => n3269, CK => CLK, RN => 
                           n458, Q => n2698, QN => n_1563);
   REGISTERS_reg_19_29_inst : DFFR_X1 port map( D => n3268, CK => CLK, RN => 
                           n458, Q => n2721, QN => n_1564);
   REGISTERS_reg_19_28_inst : DFFR_X1 port map( D => n3267, CK => CLK, RN => 
                           n458, Q => n2744, QN => n_1565);
   REGISTERS_reg_19_27_inst : DFFR_X1 port map( D => n3266, CK => CLK, RN => 
                           n458, Q => n2767, QN => n_1566);
   REGISTERS_reg_19_26_inst : DFFR_X1 port map( D => n3265, CK => CLK, RN => 
                           n458, Q => n2790, QN => n_1567);
   REGISTERS_reg_19_25_inst : DFFR_X1 port map( D => n3264, CK => CLK, RN => 
                           n458, Q => n2813, QN => n_1568);
   REGISTERS_reg_19_24_inst : DFFR_X1 port map( D => n3263, CK => CLK, RN => 
                           n458, Q => n2836, QN => n_1569);
   REGISTERS_reg_19_23_inst : DFFR_X1 port map( D => n3262, CK => CLK, RN => 
                           n458, Q => n2859, QN => n_1570);
   REGISTERS_reg_19_22_inst : DFFR_X1 port map( D => n3261, CK => CLK, RN => 
                           n458, Q => n2882, QN => n_1571);
   REGISTERS_reg_19_21_inst : DFFR_X1 port map( D => n3260, CK => CLK, RN => 
                           n458, Q => n2905, QN => n_1572);
   REGISTERS_reg_19_20_inst : DFFR_X1 port map( D => n3259, CK => CLK, RN => 
                           n458, Q => n2928, QN => n_1573);
   REGISTERS_reg_19_19_inst : DFFR_X1 port map( D => n3258, CK => CLK, RN => 
                           n459, Q => n2951, QN => n_1574);
   REGISTERS_reg_19_18_inst : DFFR_X1 port map( D => n3257, CK => CLK, RN => 
                           n459, Q => n2974, QN => n_1575);
   REGISTERS_reg_19_17_inst : DFFR_X1 port map( D => n3256, CK => CLK, RN => 
                           n459, Q => n3573, QN => n_1576);
   REGISTERS_reg_19_16_inst : DFFR_X1 port map( D => n3255, CK => CLK, RN => 
                           n459, Q => n3596, QN => n_1577);
   REGISTERS_reg_19_15_inst : DFFR_X1 port map( D => n3254, CK => CLK, RN => 
                           n459, Q => n3619, QN => n_1578);
   REGISTERS_reg_19_14_inst : DFFR_X1 port map( D => n3253, CK => CLK, RN => 
                           n459, Q => n3642, QN => n_1579);
   REGISTERS_reg_19_13_inst : DFFR_X1 port map( D => n3252, CK => CLK, RN => 
                           n459, Q => n3665, QN => n_1580);
   REGISTERS_reg_19_12_inst : DFFR_X1 port map( D => n3251, CK => CLK, RN => 
                           n459, Q => n3688, QN => n_1581);
   REGISTERS_reg_19_11_inst : DFFR_X1 port map( D => n3250, CK => CLK, RN => 
                           n459, Q => n3711, QN => n_1582);
   REGISTERS_reg_19_10_inst : DFFR_X1 port map( D => n3249, CK => CLK, RN => 
                           n459, Q => n3734, QN => n_1583);
   REGISTERS_reg_19_9_inst : DFFR_X1 port map( D => n3248, CK => CLK, RN => 
                           n459, Q => n3757, QN => n_1584);
   REGISTERS_reg_19_8_inst : DFFR_X1 port map( D => n3247, CK => CLK, RN => 
                           n459, Q => n3780, QN => n_1585);
   REGISTERS_reg_19_7_inst : DFFR_X1 port map( D => n3246, CK => CLK, RN => 
                           n460, Q => n3803, QN => n_1586);
   REGISTERS_reg_19_6_inst : DFFR_X1 port map( D => n3245, CK => CLK, RN => 
                           n460, Q => n3826, QN => n_1587);
   REGISTERS_reg_19_5_inst : DFFR_X1 port map( D => n3244, CK => CLK, RN => 
                           n460, Q => n3849, QN => n_1588);
   REGISTERS_reg_19_4_inst : DFFR_X1 port map( D => n3243, CK => CLK, RN => 
                           n460, Q => n3872, QN => n_1589);
   REGISTERS_reg_19_3_inst : DFFR_X1 port map( D => n3242, CK => CLK, RN => 
                           n460, Q => n3895, QN => n_1590);
   REGISTERS_reg_19_2_inst : DFFR_X1 port map( D => n3241, CK => CLK, RN => 
                           n460, Q => n3918, QN => n_1591);
   REGISTERS_reg_19_1_inst : DFFR_X1 port map( D => n3240, CK => CLK, RN => 
                           n460, Q => n3941, QN => n_1592);
   REGISTERS_reg_19_0_inst : DFFR_X1 port map( D => n3239, CK => CLK, RN => 
                           n460, Q => n3964, QN => n_1593);
   REGISTERS_reg_25_31_inst : DFFR_X1 port map( D => n3142, CK => CLK, RN => 
                           n474, Q => n2668, QN => n_1594);
   REGISTERS_reg_25_30_inst : DFFR_X1 port map( D => n3141, CK => CLK, RN => 
                           n474, Q => n2691, QN => n_1595);
   REGISTERS_reg_25_29_inst : DFFR_X1 port map( D => n3140, CK => CLK, RN => 
                           n474, Q => n2714, QN => n_1596);
   REGISTERS_reg_25_28_inst : DFFR_X1 port map( D => n3139, CK => CLK, RN => 
                           n474, Q => n2737, QN => n_1597);
   REGISTERS_reg_25_27_inst : DFFR_X1 port map( D => n3138, CK => CLK, RN => 
                           n474, Q => n2760, QN => n_1598);
   REGISTERS_reg_25_26_inst : DFFR_X1 port map( D => n3137, CK => CLK, RN => 
                           n474, Q => n2783, QN => n_1599);
   REGISTERS_reg_25_25_inst : DFFR_X1 port map( D => n3136, CK => CLK, RN => 
                           n474, Q => n2806, QN => n_1600);
   REGISTERS_reg_25_24_inst : DFFR_X1 port map( D => n3135, CK => CLK, RN => 
                           n474, Q => n2829, QN => n_1601);
   REGISTERS_reg_25_23_inst : DFFR_X1 port map( D => n3134, CK => CLK, RN => 
                           n474, Q => n2852, QN => n_1602);
   REGISTERS_reg_25_22_inst : DFFR_X1 port map( D => n3133, CK => CLK, RN => 
                           n474, Q => n2875, QN => n_1603);
   REGISTERS_reg_25_21_inst : DFFR_X1 port map( D => n3132, CK => CLK, RN => 
                           n474, Q => n2898, QN => n_1604);
   REGISTERS_reg_25_20_inst : DFFR_X1 port map( D => n3131, CK => CLK, RN => 
                           n474, Q => n2921, QN => n_1605);
   REGISTERS_reg_25_19_inst : DFFR_X1 port map( D => n3130, CK => CLK, RN => 
                           n475, Q => n2944, QN => n_1606);
   REGISTERS_reg_25_18_inst : DFFR_X1 port map( D => n3129, CK => CLK, RN => 
                           n475, Q => n2967, QN => n_1607);
   REGISTERS_reg_25_17_inst : DFFR_X1 port map( D => n3128, CK => CLK, RN => 
                           n475, Q => n3566, QN => n_1608);
   REGISTERS_reg_25_16_inst : DFFR_X1 port map( D => n3127, CK => CLK, RN => 
                           n475, Q => n3589, QN => n_1609);
   REGISTERS_reg_25_15_inst : DFFR_X1 port map( D => n3126, CK => CLK, RN => 
                           n475, Q => n3612, QN => n_1610);
   REGISTERS_reg_25_14_inst : DFFR_X1 port map( D => n3125, CK => CLK, RN => 
                           n475, Q => n3635, QN => n_1611);
   REGISTERS_reg_25_13_inst : DFFR_X1 port map( D => n3124, CK => CLK, RN => 
                           n475, Q => n3658, QN => n_1612);
   REGISTERS_reg_25_12_inst : DFFR_X1 port map( D => n3123, CK => CLK, RN => 
                           n475, Q => n3681, QN => n_1613);
   REGISTERS_reg_25_11_inst : DFFR_X1 port map( D => n3122, CK => CLK, RN => 
                           n475, Q => n3704, QN => n_1614);
   REGISTERS_reg_25_10_inst : DFFR_X1 port map( D => n3121, CK => CLK, RN => 
                           n475, Q => n3727, QN => n_1615);
   REGISTERS_reg_25_9_inst : DFFR_X1 port map( D => n3120, CK => CLK, RN => 
                           n475, Q => n3750, QN => n_1616);
   REGISTERS_reg_25_8_inst : DFFR_X1 port map( D => n3119, CK => CLK, RN => 
                           n475, Q => n3773, QN => n_1617);
   REGISTERS_reg_25_7_inst : DFFR_X1 port map( D => n3118, CK => CLK, RN => 
                           n476, Q => n3796, QN => n_1618);
   REGISTERS_reg_25_6_inst : DFFR_X1 port map( D => n3117, CK => CLK, RN => 
                           n476, Q => n3819, QN => n_1619);
   REGISTERS_reg_25_5_inst : DFFR_X1 port map( D => n3116, CK => CLK, RN => 
                           n476, Q => n3842, QN => n_1620);
   REGISTERS_reg_25_4_inst : DFFR_X1 port map( D => n3115, CK => CLK, RN => 
                           n476, Q => n3865, QN => n_1621);
   REGISTERS_reg_25_3_inst : DFFR_X1 port map( D => n3114, CK => CLK, RN => 
                           n476, Q => n3888, QN => n_1622);
   REGISTERS_reg_25_2_inst : DFFR_X1 port map( D => n3113, CK => CLK, RN => 
                           n476, Q => n3911, QN => n_1623);
   REGISTERS_reg_25_1_inst : DFFR_X1 port map( D => n3112, CK => CLK, RN => 
                           n476, Q => n3934, QN => n_1624);
   REGISTERS_reg_25_0_inst : DFFR_X1 port map( D => n3111, CK => CLK, RN => 
                           n476, Q => n3957, QN => n_1625);
   REGISTERS_reg_29_31_inst : DFFR_X1 port map( D => n3078, CK => CLK, RN => 
                           n484, Q => n4061, QN => n_1626);
   REGISTERS_reg_29_30_inst : DFFR_X1 port map( D => n3077, CK => CLK, RN => 
                           n484, Q => n4060, QN => n_1627);
   REGISTERS_reg_29_29_inst : DFFR_X1 port map( D => n3076, CK => CLK, RN => 
                           n484, Q => n4059, QN => n_1628);
   REGISTERS_reg_29_28_inst : DFFR_X1 port map( D => n3075, CK => CLK, RN => 
                           n484, Q => n4058, QN => n_1629);
   REGISTERS_reg_29_27_inst : DFFR_X1 port map( D => n3074, CK => CLK, RN => 
                           n485, Q => n4057, QN => n_1630);
   REGISTERS_reg_29_26_inst : DFFR_X1 port map( D => n3073, CK => CLK, RN => 
                           n485, Q => n4056, QN => n_1631);
   REGISTERS_reg_29_25_inst : DFFR_X1 port map( D => n3072, CK => CLK, RN => 
                           n485, Q => n4055, QN => n_1632);
   REGISTERS_reg_29_24_inst : DFFR_X1 port map( D => n3071, CK => CLK, RN => 
                           n485, Q => n4054, QN => n_1633);
   REGISTERS_reg_29_23_inst : DFFR_X1 port map( D => n3070, CK => CLK, RN => 
                           n485, Q => n4053, QN => n_1634);
   REGISTERS_reg_29_22_inst : DFFR_X1 port map( D => n3069, CK => CLK, RN => 
                           n485, Q => n4052, QN => n_1635);
   REGISTERS_reg_29_21_inst : DFFR_X1 port map( D => n3068, CK => CLK, RN => 
                           n485, Q => n4051, QN => n_1636);
   REGISTERS_reg_29_20_inst : DFFR_X1 port map( D => n3067, CK => CLK, RN => 
                           n485, Q => n4050, QN => n_1637);
   REGISTERS_reg_29_19_inst : DFFR_X1 port map( D => n3066, CK => CLK, RN => 
                           n485, Q => n4049, QN => n_1638);
   REGISTERS_reg_29_18_inst : DFFR_X1 port map( D => n3065, CK => CLK, RN => 
                           n485, Q => n4048, QN => n_1639);
   REGISTERS_reg_29_17_inst : DFFR_X1 port map( D => n3064, CK => CLK, RN => 
                           n485, Q => n4047, QN => n_1640);
   REGISTERS_reg_29_16_inst : DFFR_X1 port map( D => n3063, CK => CLK, RN => 
                           n485, Q => n4046, QN => n_1641);
   REGISTERS_reg_29_15_inst : DFFR_X1 port map( D => n3062, CK => CLK, RN => 
                           n486, Q => n4045, QN => n_1642);
   REGISTERS_reg_29_14_inst : DFFR_X1 port map( D => n3061, CK => CLK, RN => 
                           n486, Q => n4044, QN => n_1643);
   REGISTERS_reg_29_13_inst : DFFR_X1 port map( D => n3060, CK => CLK, RN => 
                           n486, Q => n4043, QN => n_1644);
   REGISTERS_reg_29_12_inst : DFFR_X1 port map( D => n3059, CK => CLK, RN => 
                           n486, Q => n4042, QN => n_1645);
   REGISTERS_reg_29_11_inst : DFFR_X1 port map( D => n3058, CK => CLK, RN => 
                           n486, Q => n4041, QN => n_1646);
   REGISTERS_reg_29_10_inst : DFFR_X1 port map( D => n3057, CK => CLK, RN => 
                           n486, Q => n4040, QN => n_1647);
   REGISTERS_reg_29_9_inst : DFFR_X1 port map( D => n3056, CK => CLK, RN => 
                           n486, Q => n4039, QN => n_1648);
   REGISTERS_reg_29_8_inst : DFFR_X1 port map( D => n3055, CK => CLK, RN => 
                           n486, Q => n4038, QN => n_1649);
   REGISTERS_reg_29_7_inst : DFFR_X1 port map( D => n3054, CK => CLK, RN => 
                           n486, Q => n4037, QN => n_1650);
   REGISTERS_reg_29_6_inst : DFFR_X1 port map( D => n3053, CK => CLK, RN => 
                           n486, Q => n4036, QN => n_1651);
   REGISTERS_reg_29_5_inst : DFFR_X1 port map( D => n3052, CK => CLK, RN => 
                           n486, Q => n4035, QN => n_1652);
   REGISTERS_reg_29_4_inst : DFFR_X1 port map( D => n3051, CK => CLK, RN => 
                           n486, Q => n4034, QN => n_1653);
   REGISTERS_reg_29_3_inst : DFFR_X1 port map( D => n3050, CK => CLK, RN => 
                           n487, Q => n4033, QN => n_1654);
   REGISTERS_reg_29_2_inst : DFFR_X1 port map( D => n3049, CK => CLK, RN => 
                           n487, Q => n4032, QN => n_1655);
   REGISTERS_reg_29_1_inst : DFFR_X1 port map( D => n3048, CK => CLK, RN => 
                           n487, Q => n4031, QN => n_1656);
   REGISTERS_reg_29_0_inst : DFFR_X1 port map( D => n3047, CK => CLK, RN => 
                           n487, Q => n4030, QN => n_1657);
   OUT2_reg_31_inst : DFF_X1 port map( D => n3015, CK => CLK, Q => OUT2(31), QN
                           => n2654);
   OUT2_reg_30_inst : DFF_X1 port map( D => n3016, CK => CLK, Q => OUT2(30), QN
                           => n2677);
   OUT2_reg_29_inst : DFF_X1 port map( D => n3017, CK => CLK, Q => OUT2(29), QN
                           => n2700);
   OUT2_reg_28_inst : DFF_X1 port map( D => n3018, CK => CLK, Q => OUT2(28), QN
                           => n2723);
   OUT2_reg_27_inst : DFF_X1 port map( D => n3019, CK => CLK, Q => OUT2(27), QN
                           => n2746);
   OUT2_reg_26_inst : DFF_X1 port map( D => n3020, CK => CLK, Q => OUT2(26), QN
                           => n2769);
   OUT2_reg_25_inst : DFF_X1 port map( D => n3021, CK => CLK, Q => OUT2(25), QN
                           => n2792);
   OUT2_reg_24_inst : DFF_X1 port map( D => n3022, CK => CLK, Q => OUT2(24), QN
                           => n2815);
   OUT2_reg_23_inst : DFF_X1 port map( D => n3023, CK => CLK, Q => OUT2(23), QN
                           => n2838);
   OUT2_reg_22_inst : DFF_X1 port map( D => n3024, CK => CLK, Q => OUT2(22), QN
                           => n2861);
   OUT2_reg_21_inst : DFF_X1 port map( D => n3025, CK => CLK, Q => OUT2(21), QN
                           => n2884);
   OUT2_reg_20_inst : DFF_X1 port map( D => n3026, CK => CLK, Q => OUT2(20), QN
                           => n2907);
   OUT2_reg_19_inst : DFF_X1 port map( D => n3027, CK => CLK, Q => OUT2(19), QN
                           => n2930);
   OUT2_reg_18_inst : DFF_X1 port map( D => n3028, CK => CLK, Q => OUT2(18), QN
                           => n2953);
   OUT2_reg_17_inst : DFF_X1 port map( D => n3029, CK => CLK, Q => OUT2(17), QN
                           => n2976);
   OUT2_reg_16_inst : DFF_X1 port map( D => n3030, CK => CLK, Q => OUT2(16), QN
                           => n3575);
   OUT2_reg_15_inst : DFF_X1 port map( D => n3031, CK => CLK, Q => OUT2(15), QN
                           => n3598);
   OUT2_reg_14_inst : DFF_X1 port map( D => n3032, CK => CLK, Q => OUT2(14), QN
                           => n3621);
   OUT2_reg_13_inst : DFF_X1 port map( D => n3033, CK => CLK, Q => OUT2(13), QN
                           => n3644);
   OUT2_reg_12_inst : DFF_X1 port map( D => n3034, CK => CLK, Q => OUT2(12), QN
                           => n3667);
   OUT2_reg_11_inst : DFF_X1 port map( D => n3035, CK => CLK, Q => OUT2(11), QN
                           => n3690);
   OUT2_reg_10_inst : DFF_X1 port map( D => n3036, CK => CLK, Q => OUT2(10), QN
                           => n3713);
   OUT2_reg_9_inst : DFF_X1 port map( D => n3037, CK => CLK, Q => OUT2(9), QN 
                           => n3736);
   OUT2_reg_8_inst : DFF_X1 port map( D => n3038, CK => CLK, Q => OUT2(8), QN 
                           => n3759);
   OUT2_reg_7_inst : DFF_X1 port map( D => n3039, CK => CLK, Q => OUT2(7), QN 
                           => n3782);
   OUT2_reg_6_inst : DFF_X1 port map( D => n3040, CK => CLK, Q => OUT2(6), QN 
                           => n3805);
   OUT2_reg_5_inst : DFF_X1 port map( D => n3041, CK => CLK, Q => OUT2(5), QN 
                           => n3828);
   OUT2_reg_4_inst : DFF_X1 port map( D => n3042, CK => CLK, Q => OUT2(4), QN 
                           => n3851);
   OUT2_reg_3_inst : DFF_X1 port map( D => n3043, CK => CLK, Q => OUT2(3), QN 
                           => n3874);
   OUT2_reg_2_inst : DFF_X1 port map( D => n3044, CK => CLK, Q => OUT2(2), QN 
                           => n3897);
   OUT2_reg_1_inst : DFF_X1 port map( D => n3045, CK => CLK, Q => OUT2(1), QN 
                           => n3920);
   OUT2_reg_0_inst : DFF_X1 port map( D => n3046, CK => CLK, Q => OUT2(0), QN 
                           => n3943);
   OUT1_reg_31_inst : DFF_X1 port map( D => n3014, CK => CLK, Q => OUT1(31), QN
                           => n2653);
   OUT1_reg_30_inst : DFF_X1 port map( D => n3013, CK => CLK, Q => OUT1(30), QN
                           => n2652);
   OUT1_reg_29_inst : DFF_X1 port map( D => n3012, CK => CLK, Q => OUT1(29), QN
                           => n2651);
   OUT1_reg_28_inst : DFF_X1 port map( D => n3011, CK => CLK, Q => OUT1(28), QN
                           => n2650);
   OUT1_reg_27_inst : DFF_X1 port map( D => n3010, CK => CLK, Q => OUT1(27), QN
                           => n2649);
   OUT1_reg_26_inst : DFF_X1 port map( D => n3009, CK => CLK, Q => OUT1(26), QN
                           => n2648);
   OUT1_reg_25_inst : DFF_X1 port map( D => n3008, CK => CLK, Q => OUT1(25), QN
                           => n2647);
   OUT1_reg_24_inst : DFF_X1 port map( D => n3007, CK => CLK, Q => OUT1(24), QN
                           => n2646);
   OUT1_reg_23_inst : DFF_X1 port map( D => n3006, CK => CLK, Q => OUT1(23), QN
                           => n2645);
   OUT1_reg_22_inst : DFF_X1 port map( D => n3005, CK => CLK, Q => OUT1(22), QN
                           => n2644);
   OUT1_reg_21_inst : DFF_X1 port map( D => n3004, CK => CLK, Q => OUT1(21), QN
                           => n2643);
   OUT1_reg_20_inst : DFF_X1 port map( D => n3003, CK => CLK, Q => OUT1(20), QN
                           => n2642);
   OUT1_reg_19_inst : DFF_X1 port map( D => n3002, CK => CLK, Q => OUT1(19), QN
                           => n2641);
   OUT1_reg_18_inst : DFF_X1 port map( D => n3001, CK => CLK, Q => OUT1(18), QN
                           => n2640);
   OUT1_reg_17_inst : DFF_X1 port map( D => n3000, CK => CLK, Q => OUT1(17), QN
                           => n2639);
   OUT1_reg_16_inst : DFF_X1 port map( D => n2999, CK => CLK, Q => OUT1(16), QN
                           => n2638);
   OUT1_reg_15_inst : DFF_X1 port map( D => n2998, CK => CLK, Q => OUT1(15), QN
                           => n2637);
   OUT1_reg_14_inst : DFF_X1 port map( D => n2997, CK => CLK, Q => OUT1(14), QN
                           => n2636);
   OUT1_reg_13_inst : DFF_X1 port map( D => n2996, CK => CLK, Q => OUT1(13), QN
                           => n2635);
   OUT1_reg_12_inst : DFF_X1 port map( D => n2995, CK => CLK, Q => OUT1(12), QN
                           => n2634);
   OUT1_reg_11_inst : DFF_X1 port map( D => n2994, CK => CLK, Q => OUT1(11), QN
                           => n2633);
   OUT1_reg_10_inst : DFF_X1 port map( D => n2993, CK => CLK, Q => OUT1(10), QN
                           => n2632);
   OUT1_reg_9_inst : DFF_X1 port map( D => n2992, CK => CLK, Q => OUT1(9), QN 
                           => n2631);
   OUT1_reg_8_inst : DFF_X1 port map( D => n2991, CK => CLK, Q => OUT1(8), QN 
                           => n2630);
   OUT1_reg_7_inst : DFF_X1 port map( D => n2990, CK => CLK, Q => OUT1(7), QN 
                           => n2629);
   OUT1_reg_6_inst : DFF_X1 port map( D => n2989, CK => CLK, Q => OUT1(6), QN 
                           => n2628);
   OUT1_reg_5_inst : DFF_X1 port map( D => n2988, CK => CLK, Q => OUT1(5), QN 
                           => n2627);
   OUT1_reg_4_inst : DFF_X1 port map( D => n2987, CK => CLK, Q => OUT1(4), QN 
                           => n2626);
   OUT1_reg_3_inst : DFF_X1 port map( D => n2986, CK => CLK, Q => OUT1(3), QN 
                           => n2625);
   OUT1_reg_2_inst : DFF_X1 port map( D => n2985, CK => CLK, Q => OUT1(2), QN 
                           => n2624);
   OUT1_reg_1_inst : DFF_X1 port map( D => n2984, CK => CLK, Q => OUT1(1), QN 
                           => n2623);
   OUT1_reg_0_inst : DFF_X1 port map( D => n2983, CK => CLK, Q => OUT1(0), QN 
                           => n2622);
   REGISTERS_reg_24_31_inst : DFFR_X1 port map( D => n3174, CK => CLK, RN => 
                           RST, Q => n2669, QN => n1435);
   REGISTERS_reg_24_30_inst : DFFR_X1 port map( D => n3173, CK => CLK, RN => 
                           n471, Q => n2692, QN => n1419);
   REGISTERS_reg_24_29_inst : DFFR_X1 port map( D => n3172, CK => CLK, RN => 
                           n471, Q => n2715, QN => n1403);
   REGISTERS_reg_24_28_inst : DFFR_X1 port map( D => n3171, CK => CLK, RN => 
                           n471, Q => n2738, QN => n1387);
   REGISTERS_reg_24_27_inst : DFFR_X1 port map( D => n3170, CK => CLK, RN => 
                           n471, Q => n2761, QN => n1371);
   REGISTERS_reg_24_26_inst : DFFR_X1 port map( D => n3169, CK => CLK, RN => 
                           n471, Q => n2784, QN => n1355);
   REGISTERS_reg_24_25_inst : DFFR_X1 port map( D => n3168, CK => CLK, RN => 
                           n471, Q => n2807, QN => n1339);
   REGISTERS_reg_24_24_inst : DFFR_X1 port map( D => n3167, CK => CLK, RN => 
                           n471, Q => n2830, QN => n1323);
   REGISTERS_reg_24_23_inst : DFFR_X1 port map( D => n3166, CK => CLK, RN => 
                           n472, Q => n2853, QN => n1307);
   REGISTERS_reg_24_22_inst : DFFR_X1 port map( D => n3165, CK => CLK, RN => 
                           n472, Q => n2876, QN => n1291);
   REGISTERS_reg_24_21_inst : DFFR_X1 port map( D => n3164, CK => CLK, RN => 
                           n472, Q => n2899, QN => n1275);
   REGISTERS_reg_24_20_inst : DFFR_X1 port map( D => n3163, CK => CLK, RN => 
                           n472, Q => n2922, QN => n1259);
   REGISTERS_reg_24_19_inst : DFFR_X1 port map( D => n3162, CK => CLK, RN => 
                           n472, Q => n2945, QN => n1243);
   REGISTERS_reg_24_18_inst : DFFR_X1 port map( D => n3161, CK => CLK, RN => 
                           n472, Q => n2968, QN => n1227);
   REGISTERS_reg_24_17_inst : DFFR_X1 port map( D => n3160, CK => CLK, RN => 
                           n472, Q => n3567, QN => n1211);
   REGISTERS_reg_24_16_inst : DFFR_X1 port map( D => n3159, CK => CLK, RN => 
                           n472, Q => n3590, QN => n1195);
   REGISTERS_reg_24_15_inst : DFFR_X1 port map( D => n3158, CK => CLK, RN => 
                           n472, Q => n3613, QN => n1179);
   REGISTERS_reg_24_14_inst : DFFR_X1 port map( D => n3157, CK => CLK, RN => 
                           n472, Q => n3636, QN => n1163);
   REGISTERS_reg_24_13_inst : DFFR_X1 port map( D => n3156, CK => CLK, RN => 
                           n472, Q => n3659, QN => n1147);
   REGISTERS_reg_24_12_inst : DFFR_X1 port map( D => n3155, CK => CLK, RN => 
                           n472, Q => n3682, QN => n1131);
   REGISTERS_reg_24_11_inst : DFFR_X1 port map( D => n3154, CK => CLK, RN => 
                           n473, Q => n3705, QN => n1115);
   REGISTERS_reg_24_10_inst : DFFR_X1 port map( D => n3153, CK => CLK, RN => 
                           n473, Q => n3728, QN => n1099);
   REGISTERS_reg_24_9_inst : DFFR_X1 port map( D => n3152, CK => CLK, RN => 
                           n473, Q => n3751, QN => n1083);
   REGISTERS_reg_24_8_inst : DFFR_X1 port map( D => n3151, CK => CLK, RN => 
                           n473, Q => n3774, QN => n1067);
   REGISTERS_reg_24_7_inst : DFFR_X1 port map( D => n3150, CK => CLK, RN => 
                           n473, Q => n3797, QN => n1051);
   REGISTERS_reg_24_6_inst : DFFR_X1 port map( D => n3149, CK => CLK, RN => 
                           n473, Q => n3820, QN => n1035);
   REGISTERS_reg_24_5_inst : DFFR_X1 port map( D => n3148, CK => CLK, RN => 
                           n473, Q => n3843, QN => n1019);
   REGISTERS_reg_24_4_inst : DFFR_X1 port map( D => n3147, CK => CLK, RN => 
                           n473, Q => n3866, QN => n1003);
   REGISTERS_reg_24_3_inst : DFFR_X1 port map( D => n3146, CK => CLK, RN => 
                           n473, Q => n3889, QN => n987);
   REGISTERS_reg_24_2_inst : DFFR_X1 port map( D => n3145, CK => CLK, RN => 
                           n473, Q => n3912, QN => n971);
   REGISTERS_reg_24_1_inst : DFFR_X1 port map( D => n3144, CK => CLK, RN => 
                           n473, Q => n3935, QN => n955);
   REGISTERS_reg_24_0_inst : DFFR_X1 port map( D => n3143, CK => CLK, RN => 
                           n473, Q => n3958, QN => n938);
   REGISTERS_reg_23_31_inst : DFFR_X1 port map( D => n3206, CK => CLK, RN => 
                           n468, Q => n2672, QN => n1437);
   REGISTERS_reg_23_30_inst : DFFR_X1 port map( D => n3205, CK => CLK, RN => 
                           n468, Q => n2695, QN => n1420);
   REGISTERS_reg_23_29_inst : DFFR_X1 port map( D => n3204, CK => CLK, RN => 
                           n468, Q => n2718, QN => n1404);
   REGISTERS_reg_23_28_inst : DFFR_X1 port map( D => n3203, CK => CLK, RN => 
                           n468, Q => n2741, QN => n1388);
   REGISTERS_reg_23_27_inst : DFFR_X1 port map( D => n3202, CK => CLK, RN => 
                           n469, Q => n2764, QN => n1372);
   REGISTERS_reg_23_26_inst : DFFR_X1 port map( D => n3201, CK => CLK, RN => 
                           n469, Q => n2787, QN => n1356);
   REGISTERS_reg_23_25_inst : DFFR_X1 port map( D => n3200, CK => CLK, RN => 
                           n469, Q => n2810, QN => n1340);
   REGISTERS_reg_23_24_inst : DFFR_X1 port map( D => n3199, CK => CLK, RN => 
                           n469, Q => n2833, QN => n1324);
   REGISTERS_reg_23_23_inst : DFFR_X1 port map( D => n3198, CK => CLK, RN => 
                           n469, Q => n2856, QN => n1308);
   REGISTERS_reg_23_22_inst : DFFR_X1 port map( D => n3197, CK => CLK, RN => 
                           n469, Q => n2879, QN => n1292);
   REGISTERS_reg_23_21_inst : DFFR_X1 port map( D => n3196, CK => CLK, RN => 
                           n469, Q => n2902, QN => n1276);
   REGISTERS_reg_23_20_inst : DFFR_X1 port map( D => n3195, CK => CLK, RN => 
                           n469, Q => n2925, QN => n1260);
   REGISTERS_reg_23_19_inst : DFFR_X1 port map( D => n3194, CK => CLK, RN => 
                           n469, Q => n2948, QN => n1244);
   REGISTERS_reg_23_18_inst : DFFR_X1 port map( D => n3193, CK => CLK, RN => 
                           n469, Q => n2971, QN => n1228);
   REGISTERS_reg_23_17_inst : DFFR_X1 port map( D => n3192, CK => CLK, RN => 
                           n469, Q => n3570, QN => n1212);
   REGISTERS_reg_23_16_inst : DFFR_X1 port map( D => n3191, CK => CLK, RN => 
                           n469, Q => n3593, QN => n1196);
   REGISTERS_reg_23_15_inst : DFFR_X1 port map( D => n3190, CK => CLK, RN => 
                           n470, Q => n3616, QN => n1180);
   REGISTERS_reg_23_14_inst : DFFR_X1 port map( D => n3189, CK => CLK, RN => 
                           n470, Q => n3639, QN => n1164);
   REGISTERS_reg_23_13_inst : DFFR_X1 port map( D => n3188, CK => CLK, RN => 
                           n470, Q => n3662, QN => n1148);
   REGISTERS_reg_23_12_inst : DFFR_X1 port map( D => n3187, CK => CLK, RN => 
                           n470, Q => n3685, QN => n1132);
   REGISTERS_reg_23_11_inst : DFFR_X1 port map( D => n3186, CK => CLK, RN => 
                           n470, Q => n3708, QN => n1116);
   REGISTERS_reg_23_10_inst : DFFR_X1 port map( D => n3185, CK => CLK, RN => 
                           n470, Q => n3731, QN => n1100);
   REGISTERS_reg_23_9_inst : DFFR_X1 port map( D => n3184, CK => CLK, RN => 
                           n470, Q => n3754, QN => n1084);
   REGISTERS_reg_23_8_inst : DFFR_X1 port map( D => n3183, CK => CLK, RN => 
                           n470, Q => n3777, QN => n1068);
   REGISTERS_reg_23_7_inst : DFFR_X1 port map( D => n3182, CK => CLK, RN => 
                           n470, Q => n3800, QN => n1052);
   REGISTERS_reg_23_6_inst : DFFR_X1 port map( D => n3181, CK => CLK, RN => 
                           n470, Q => n3823, QN => n1036);
   REGISTERS_reg_23_5_inst : DFFR_X1 port map( D => n3180, CK => CLK, RN => 
                           n470, Q => n3846, QN => n1020);
   REGISTERS_reg_23_4_inst : DFFR_X1 port map( D => n3179, CK => CLK, RN => 
                           n470, Q => n3869, QN => n1004);
   REGISTERS_reg_23_3_inst : DFFR_X1 port map( D => n3178, CK => CLK, RN => 
                           n471, Q => n3892, QN => n988);
   REGISTERS_reg_23_2_inst : DFFR_X1 port map( D => n3177, CK => CLK, RN => 
                           n471, Q => n3915, QN => n972);
   REGISTERS_reg_23_1_inst : DFFR_X1 port map( D => n3176, CK => CLK, RN => 
                           n471, Q => n3938, QN => n956);
   REGISTERS_reg_23_0_inst : DFFR_X1 port map( D => n3175, CK => CLK, RN => 
                           n471, Q => n3961, QN => n939);
   REGISTERS_reg_22_31_inst : DFFR_X1 port map( D => n3238, CK => CLK, RN => 
                           n466, Q => n2673, QN => n2320);
   REGISTERS_reg_22_30_inst : DFFR_X1 port map( D => n3237, CK => CLK, RN => 
                           n466, Q => n2696, QN => n2299);
   REGISTERS_reg_22_29_inst : DFFR_X1 port map( D => n3236, CK => CLK, RN => 
                           n466, Q => n2719, QN => n2287);
   REGISTERS_reg_22_28_inst : DFFR_X1 port map( D => n3235, CK => CLK, RN => 
                           n466, Q => n2742, QN => n2275);
   REGISTERS_reg_22_27_inst : DFFR_X1 port map( D => n3234, CK => CLK, RN => 
                           n466, Q => n2765, QN => n2263);
   REGISTERS_reg_22_26_inst : DFFR_X1 port map( D => n3233, CK => CLK, RN => 
                           n466, Q => n2788, QN => n2251);
   REGISTERS_reg_22_25_inst : DFFR_X1 port map( D => n3232, CK => CLK, RN => 
                           n466, Q => n2811, QN => n2239);
   REGISTERS_reg_22_24_inst : DFFR_X1 port map( D => n3231, CK => CLK, RN => 
                           n466, Q => n2834, QN => n2227);
   REGISTERS_reg_22_23_inst : DFFR_X1 port map( D => n3230, CK => CLK, RN => 
                           n466, Q => n2857, QN => n2215);
   REGISTERS_reg_22_22_inst : DFFR_X1 port map( D => n3229, CK => CLK, RN => 
                           n466, Q => n2880, QN => n2203);
   REGISTERS_reg_22_21_inst : DFFR_X1 port map( D => n3228, CK => CLK, RN => 
                           n466, Q => n2903, QN => n2191);
   REGISTERS_reg_22_20_inst : DFFR_X1 port map( D => n3227, CK => CLK, RN => 
                           n466, Q => n2926, QN => n2179);
   REGISTERS_reg_22_19_inst : DFFR_X1 port map( D => n3226, CK => CLK, RN => 
                           n467, Q => n2949, QN => n2167);
   REGISTERS_reg_22_18_inst : DFFR_X1 port map( D => n3225, CK => CLK, RN => 
                           n467, Q => n2972, QN => n2155);
   REGISTERS_reg_22_17_inst : DFFR_X1 port map( D => n3224, CK => CLK, RN => 
                           n467, Q => n3571, QN => n2143);
   REGISTERS_reg_22_16_inst : DFFR_X1 port map( D => n3223, CK => CLK, RN => 
                           n467, Q => n3594, QN => n2131);
   REGISTERS_reg_22_15_inst : DFFR_X1 port map( D => n3222, CK => CLK, RN => 
                           n467, Q => n3617, QN => n2119);
   REGISTERS_reg_22_14_inst : DFFR_X1 port map( D => n3221, CK => CLK, RN => 
                           n467, Q => n3640, QN => n2107);
   REGISTERS_reg_22_13_inst : DFFR_X1 port map( D => n3220, CK => CLK, RN => 
                           n467, Q => n3663, QN => n2095);
   REGISTERS_reg_22_12_inst : DFFR_X1 port map( D => n3219, CK => CLK, RN => 
                           n467, Q => n3686, QN => n2083);
   REGISTERS_reg_22_11_inst : DFFR_X1 port map( D => n3218, CK => CLK, RN => 
                           n467, Q => n3709, QN => n2071);
   REGISTERS_reg_22_10_inst : DFFR_X1 port map( D => n3217, CK => CLK, RN => 
                           n467, Q => n3732, QN => n2059);
   REGISTERS_reg_22_9_inst : DFFR_X1 port map( D => n3216, CK => CLK, RN => 
                           n467, Q => n3755, QN => n2047);
   REGISTERS_reg_22_8_inst : DFFR_X1 port map( D => n3215, CK => CLK, RN => 
                           n467, Q => n3778, QN => n2035);
   REGISTERS_reg_22_7_inst : DFFR_X1 port map( D => n3214, CK => CLK, RN => 
                           n468, Q => n3801, QN => n2023);
   REGISTERS_reg_22_6_inst : DFFR_X1 port map( D => n3213, CK => CLK, RN => 
                           n468, Q => n3824, QN => n2011);
   REGISTERS_reg_22_5_inst : DFFR_X1 port map( D => n3212, CK => CLK, RN => 
                           n468, Q => n3847, QN => n1999);
   REGISTERS_reg_22_4_inst : DFFR_X1 port map( D => n3211, CK => CLK, RN => 
                           n468, Q => n3870, QN => n1987);
   REGISTERS_reg_22_3_inst : DFFR_X1 port map( D => n3210, CK => CLK, RN => 
                           n468, Q => n3893, QN => n1975);
   REGISTERS_reg_22_2_inst : DFFR_X1 port map( D => n3209, CK => CLK, RN => 
                           n468, Q => n3916, QN => n1963);
   REGISTERS_reg_22_1_inst : DFFR_X1 port map( D => n3208, CK => CLK, RN => 
                           n468, Q => n3939, QN => n1951);
   REGISTERS_reg_22_0_inst : DFFR_X1 port map( D => n3207, CK => CLK, RN => 
                           n468, Q => n3962, QN => n1922);
   REGISTERS_reg_7_31_inst : DFFR_X1 port map( D => n3462, CK => CLK, RN => 
                           n426, Q => n2664, QN => n2331);
   REGISTERS_reg_7_30_inst : DFFR_X1 port map( D => n3461, CK => CLK, RN => 
                           n426, Q => n2687, QN => n2306);
   REGISTERS_reg_7_29_inst : DFFR_X1 port map( D => n3460, CK => CLK, RN => 
                           n426, Q => n2710, QN => n2294);
   REGISTERS_reg_7_28_inst : DFFR_X1 port map( D => n3459, CK => CLK, RN => 
                           n426, Q => n2733, QN => n2282);
   REGISTERS_reg_7_27_inst : DFFR_X1 port map( D => n3458, CK => CLK, RN => 
                           n426, Q => n2756, QN => n2270);
   REGISTERS_reg_7_26_inst : DFFR_X1 port map( D => n3457, CK => CLK, RN => 
                           n426, Q => n2779, QN => n2258);
   REGISTERS_reg_7_25_inst : DFFR_X1 port map( D => n3456, CK => CLK, RN => 
                           n426, Q => n2802, QN => n2246);
   REGISTERS_reg_7_24_inst : DFFR_X1 port map( D => n3455, CK => CLK, RN => 
                           n426, Q => n2825, QN => n2234);
   REGISTERS_reg_7_23_inst : DFFR_X1 port map( D => n3454, CK => CLK, RN => 
                           n426, Q => n2848, QN => n2222);
   REGISTERS_reg_7_22_inst : DFFR_X1 port map( D => n3453, CK => CLK, RN => 
                           n426, Q => n2871, QN => n2210);
   REGISTERS_reg_7_21_inst : DFFR_X1 port map( D => n3452, CK => CLK, RN => 
                           n426, Q => n2894, QN => n2198);
   REGISTERS_reg_7_20_inst : DFFR_X1 port map( D => n3451, CK => CLK, RN => 
                           n426, Q => n2917, QN => n2186);
   REGISTERS_reg_7_19_inst : DFFR_X1 port map( D => n3450, CK => CLK, RN => 
                           n427, Q => n2940, QN => n2174);
   REGISTERS_reg_7_18_inst : DFFR_X1 port map( D => n3449, CK => CLK, RN => 
                           n427, Q => n2963, QN => n2162);
   REGISTERS_reg_7_17_inst : DFFR_X1 port map( D => n3448, CK => CLK, RN => 
                           n427, Q => n3562, QN => n2150);
   REGISTERS_reg_7_16_inst : DFFR_X1 port map( D => n3447, CK => CLK, RN => 
                           n427, Q => n3585, QN => n2138);
   REGISTERS_reg_7_15_inst : DFFR_X1 port map( D => n3446, CK => CLK, RN => 
                           n427, Q => n3608, QN => n2126);
   REGISTERS_reg_7_14_inst : DFFR_X1 port map( D => n3445, CK => CLK, RN => 
                           n427, Q => n3631, QN => n2114);
   REGISTERS_reg_7_13_inst : DFFR_X1 port map( D => n3444, CK => CLK, RN => 
                           n427, Q => n3654, QN => n2102);
   REGISTERS_reg_7_12_inst : DFFR_X1 port map( D => n3443, CK => CLK, RN => 
                           n427, Q => n3677, QN => n2090);
   REGISTERS_reg_7_11_inst : DFFR_X1 port map( D => n3442, CK => CLK, RN => 
                           n427, Q => n3700, QN => n2078);
   REGISTERS_reg_7_10_inst : DFFR_X1 port map( D => n3441, CK => CLK, RN => 
                           n427, Q => n3723, QN => n2066);
   REGISTERS_reg_7_9_inst : DFFR_X1 port map( D => n3440, CK => CLK, RN => n427
                           , Q => n3746, QN => n2054);
   REGISTERS_reg_7_8_inst : DFFR_X1 port map( D => n3439, CK => CLK, RN => n427
                           , Q => n3769, QN => n2042);
   REGISTERS_reg_7_7_inst : DFFR_X1 port map( D => n3438, CK => CLK, RN => n428
                           , Q => n3792, QN => n2030);
   REGISTERS_reg_7_6_inst : DFFR_X1 port map( D => n3437, CK => CLK, RN => n428
                           , Q => n3815, QN => n2018);
   REGISTERS_reg_7_5_inst : DFFR_X1 port map( D => n3436, CK => CLK, RN => n428
                           , Q => n3838, QN => n2006);
   REGISTERS_reg_7_4_inst : DFFR_X1 port map( D => n3435, CK => CLK, RN => n428
                           , Q => n3861, QN => n1994);
   REGISTERS_reg_7_3_inst : DFFR_X1 port map( D => n3434, CK => CLK, RN => n428
                           , Q => n3884, QN => n1982);
   REGISTERS_reg_7_2_inst : DFFR_X1 port map( D => n3433, CK => CLK, RN => n428
                           , Q => n3907, QN => n1970);
   REGISTERS_reg_7_1_inst : DFFR_X1 port map( D => n3432, CK => CLK, RN => n428
                           , Q => n3930, QN => n1958);
   REGISTERS_reg_7_0_inst : DFFR_X1 port map( D => n3431, CK => CLK, RN => n428
                           , Q => n3953, QN => n1942);
   REGISTERS_reg_6_31_inst : DFFR_X1 port map( D => n3494, CK => CLK, RN => 
                           n423, Q => n2665, QN => n2330);
   REGISTERS_reg_6_30_inst : DFFR_X1 port map( D => n3493, CK => CLK, RN => 
                           n423, Q => n2688, QN => n2305);
   REGISTERS_reg_6_29_inst : DFFR_X1 port map( D => n3492, CK => CLK, RN => 
                           n423, Q => n2711, QN => n2293);
   REGISTERS_reg_6_28_inst : DFFR_X1 port map( D => n3491, CK => CLK, RN => 
                           n423, Q => n2734, QN => n2281);
   REGISTERS_reg_6_27_inst : DFFR_X1 port map( D => n3490, CK => CLK, RN => 
                           n423, Q => n2757, QN => n2269);
   REGISTERS_reg_6_26_inst : DFFR_X1 port map( D => n3489, CK => CLK, RN => 
                           n423, Q => n2780, QN => n2257);
   REGISTERS_reg_6_25_inst : DFFR_X1 port map( D => n3488, CK => CLK, RN => 
                           n423, Q => n2803, QN => n2245);
   REGISTERS_reg_6_24_inst : DFFR_X1 port map( D => n3487, CK => CLK, RN => 
                           n423, Q => n2826, QN => n2233);
   REGISTERS_reg_6_23_inst : DFFR_X1 port map( D => n3486, CK => CLK, RN => 
                           n424, Q => n2849, QN => n2221);
   REGISTERS_reg_6_22_inst : DFFR_X1 port map( D => n3485, CK => CLK, RN => 
                           n424, Q => n2872, QN => n2209);
   REGISTERS_reg_6_21_inst : DFFR_X1 port map( D => n3484, CK => CLK, RN => 
                           n424, Q => n2895, QN => n2197);
   REGISTERS_reg_6_20_inst : DFFR_X1 port map( D => n3483, CK => CLK, RN => 
                           n424, Q => n2918, QN => n2185);
   REGISTERS_reg_6_19_inst : DFFR_X1 port map( D => n3482, CK => CLK, RN => 
                           n424, Q => n2941, QN => n2173);
   REGISTERS_reg_6_18_inst : DFFR_X1 port map( D => n3481, CK => CLK, RN => 
                           n424, Q => n2964, QN => n2161);
   REGISTERS_reg_6_17_inst : DFFR_X1 port map( D => n3480, CK => CLK, RN => 
                           n424, Q => n3563, QN => n2149);
   REGISTERS_reg_6_16_inst : DFFR_X1 port map( D => n3479, CK => CLK, RN => 
                           n424, Q => n3586, QN => n2137);
   REGISTERS_reg_6_15_inst : DFFR_X1 port map( D => n3478, CK => CLK, RN => 
                           n424, Q => n3609, QN => n2125);
   REGISTERS_reg_6_14_inst : DFFR_X1 port map( D => n3477, CK => CLK, RN => 
                           n424, Q => n3632, QN => n2113);
   REGISTERS_reg_6_13_inst : DFFR_X1 port map( D => n3476, CK => CLK, RN => 
                           n424, Q => n3655, QN => n2101);
   REGISTERS_reg_6_12_inst : DFFR_X1 port map( D => n3475, CK => CLK, RN => 
                           n424, Q => n3678, QN => n2089);
   REGISTERS_reg_6_11_inst : DFFR_X1 port map( D => n3474, CK => CLK, RN => 
                           n425, Q => n3701, QN => n2077);
   REGISTERS_reg_6_10_inst : DFFR_X1 port map( D => n3473, CK => CLK, RN => 
                           n425, Q => n3724, QN => n2065);
   REGISTERS_reg_6_9_inst : DFFR_X1 port map( D => n3472, CK => CLK, RN => n425
                           , Q => n3747, QN => n2053);
   REGISTERS_reg_6_8_inst : DFFR_X1 port map( D => n3471, CK => CLK, RN => n425
                           , Q => n3770, QN => n2041);
   REGISTERS_reg_6_7_inst : DFFR_X1 port map( D => n3470, CK => CLK, RN => n425
                           , Q => n3793, QN => n2029);
   REGISTERS_reg_6_6_inst : DFFR_X1 port map( D => n3469, CK => CLK, RN => n425
                           , Q => n3816, QN => n2017);
   REGISTERS_reg_6_5_inst : DFFR_X1 port map( D => n3468, CK => CLK, RN => n425
                           , Q => n3839, QN => n2005);
   REGISTERS_reg_6_4_inst : DFFR_X1 port map( D => n3467, CK => CLK, RN => n425
                           , Q => n3862, QN => n1993);
   REGISTERS_reg_6_3_inst : DFFR_X1 port map( D => n3466, CK => CLK, RN => n425
                           , Q => n3885, QN => n1981);
   REGISTERS_reg_6_2_inst : DFFR_X1 port map( D => n3465, CK => CLK, RN => n425
                           , Q => n3908, QN => n1969);
   REGISTERS_reg_6_1_inst : DFFR_X1 port map( D => n3464, CK => CLK, RN => n425
                           , Q => n3931, QN => n1957);
   REGISTERS_reg_6_0_inst : DFFR_X1 port map( D => n3463, CK => CLK, RN => n425
                           , Q => n3954, QN => n1940);
   REGISTERS_reg_3_31_inst : DFFR_X1 port map( D => n3526, CK => CLK, RN => 
                           n415, Q => n2666, QN => n2338);
   REGISTERS_reg_3_30_inst : DFFR_X1 port map( D => n3525, CK => CLK, RN => 
                           n415, Q => n2689, QN => n2309);
   REGISTERS_reg_3_29_inst : DFFR_X1 port map( D => n3524, CK => CLK, RN => 
                           n415, Q => n2712, QN => n2297);
   REGISTERS_reg_3_28_inst : DFFR_X1 port map( D => n3523, CK => CLK, RN => 
                           n415, Q => n2735, QN => n2285);
   REGISTERS_reg_3_27_inst : DFFR_X1 port map( D => n3522, CK => CLK, RN => 
                           n415, Q => n2758, QN => n2273);
   REGISTERS_reg_3_26_inst : DFFR_X1 port map( D => n3521, CK => CLK, RN => 
                           n415, Q => n2781, QN => n2261);
   REGISTERS_reg_3_25_inst : DFFR_X1 port map( D => n3520, CK => CLK, RN => 
                           n415, Q => n2804, QN => n2249);
   REGISTERS_reg_3_24_inst : DFFR_X1 port map( D => n3519, CK => CLK, RN => 
                           n415, Q => n2827, QN => n2237);
   REGISTERS_reg_3_23_inst : DFFR_X1 port map( D => n3518, CK => CLK, RN => 
                           n416, Q => n2850, QN => n2225);
   REGISTERS_reg_3_22_inst : DFFR_X1 port map( D => n3517, CK => CLK, RN => 
                           n416, Q => n2873, QN => n2213);
   REGISTERS_reg_3_21_inst : DFFR_X1 port map( D => n3516, CK => CLK, RN => 
                           n416, Q => n2896, QN => n2201);
   REGISTERS_reg_3_20_inst : DFFR_X1 port map( D => n3515, CK => CLK, RN => 
                           n416, Q => n2919, QN => n2189);
   REGISTERS_reg_3_19_inst : DFFR_X1 port map( D => n3514, CK => CLK, RN => 
                           n416, Q => n2942, QN => n2177);
   REGISTERS_reg_3_18_inst : DFFR_X1 port map( D => n3513, CK => CLK, RN => 
                           n416, Q => n2965, QN => n2165);
   REGISTERS_reg_3_17_inst : DFFR_X1 port map( D => n3512, CK => CLK, RN => 
                           n416, Q => n3564, QN => n2153);
   REGISTERS_reg_3_16_inst : DFFR_X1 port map( D => n3511, CK => CLK, RN => 
                           n416, Q => n3587, QN => n2141);
   REGISTERS_reg_3_15_inst : DFFR_X1 port map( D => n3510, CK => CLK, RN => 
                           n416, Q => n3610, QN => n2129);
   REGISTERS_reg_3_14_inst : DFFR_X1 port map( D => n3509, CK => CLK, RN => 
                           n416, Q => n3633, QN => n2117);
   REGISTERS_reg_3_13_inst : DFFR_X1 port map( D => n3508, CK => CLK, RN => 
                           n416, Q => n3656, QN => n2105);
   REGISTERS_reg_3_12_inst : DFFR_X1 port map( D => n3507, CK => CLK, RN => 
                           n416, Q => n3679, QN => n2093);
   REGISTERS_reg_3_11_inst : DFFR_X1 port map( D => n3506, CK => CLK, RN => 
                           n417, Q => n3702, QN => n2081);
   REGISTERS_reg_3_10_inst : DFFR_X1 port map( D => n3505, CK => CLK, RN => 
                           n417, Q => n3725, QN => n2069);
   REGISTERS_reg_3_9_inst : DFFR_X1 port map( D => n3504, CK => CLK, RN => n417
                           , Q => n3748, QN => n2057);
   REGISTERS_reg_3_8_inst : DFFR_X1 port map( D => n3503, CK => CLK, RN => n417
                           , Q => n3771, QN => n2045);
   REGISTERS_reg_3_7_inst : DFFR_X1 port map( D => n3502, CK => CLK, RN => n417
                           , Q => n3794, QN => n2033);
   REGISTERS_reg_3_6_inst : DFFR_X1 port map( D => n3501, CK => CLK, RN => n417
                           , Q => n3817, QN => n2021);
   REGISTERS_reg_3_5_inst : DFFR_X1 port map( D => n3500, CK => CLK, RN => n417
                           , Q => n3840, QN => n2009);
   REGISTERS_reg_3_4_inst : DFFR_X1 port map( D => n3499, CK => CLK, RN => n417
                           , Q => n3863, QN => n1997);
   REGISTERS_reg_3_3_inst : DFFR_X1 port map( D => n3498, CK => CLK, RN => n417
                           , Q => n3886, QN => n1985);
   REGISTERS_reg_3_2_inst : DFFR_X1 port map( D => n3497, CK => CLK, RN => n417
                           , Q => n3909, QN => n1973);
   REGISTERS_reg_3_1_inst : DFFR_X1 port map( D => n3496, CK => CLK, RN => n417
                           , Q => n3932, QN => n1961);
   REGISTERS_reg_3_0_inst : DFFR_X1 port map( D => n3495, CK => CLK, RN => n417
                           , Q => n3955, QN => n1948);
   REGISTERS_reg_2_31_inst : DFFR_X1 port map( D => n3558, CK => CLK, RN => 
                           n412, Q => n2667, QN => n2337);
   REGISTERS_reg_2_30_inst : DFFR_X1 port map( D => n3557, CK => CLK, RN => 
                           n412, Q => n2690, QN => n2308);
   REGISTERS_reg_2_29_inst : DFFR_X1 port map( D => n3556, CK => CLK, RN => 
                           n412, Q => n2713, QN => n2296);
   REGISTERS_reg_2_28_inst : DFFR_X1 port map( D => n3555, CK => CLK, RN => 
                           n412, Q => n2736, QN => n2284);
   REGISTERS_reg_2_27_inst : DFFR_X1 port map( D => n3554, CK => CLK, RN => 
                           n413, Q => n2759, QN => n2272);
   REGISTERS_reg_2_26_inst : DFFR_X1 port map( D => n3553, CK => CLK, RN => 
                           n413, Q => n2782, QN => n2260);
   REGISTERS_reg_2_25_inst : DFFR_X1 port map( D => n3552, CK => CLK, RN => 
                           n413, Q => n2805, QN => n2248);
   REGISTERS_reg_2_24_inst : DFFR_X1 port map( D => n3551, CK => CLK, RN => 
                           n413, Q => n2828, QN => n2236);
   REGISTERS_reg_2_23_inst : DFFR_X1 port map( D => n3550, CK => CLK, RN => 
                           n413, Q => n2851, QN => n2224);
   REGISTERS_reg_2_22_inst : DFFR_X1 port map( D => n3549, CK => CLK, RN => 
                           n413, Q => n2874, QN => n2212);
   REGISTERS_reg_2_21_inst : DFFR_X1 port map( D => n3548, CK => CLK, RN => 
                           n413, Q => n2897, QN => n2200);
   REGISTERS_reg_2_20_inst : DFFR_X1 port map( D => n3547, CK => CLK, RN => 
                           n413, Q => n2920, QN => n2188);
   REGISTERS_reg_2_19_inst : DFFR_X1 port map( D => n3546, CK => CLK, RN => 
                           n413, Q => n2943, QN => n2176);
   REGISTERS_reg_2_18_inst : DFFR_X1 port map( D => n3545, CK => CLK, RN => 
                           n413, Q => n2966, QN => n2164);
   REGISTERS_reg_2_17_inst : DFFR_X1 port map( D => n3544, CK => CLK, RN => 
                           n413, Q => n3565, QN => n2152);
   REGISTERS_reg_2_16_inst : DFFR_X1 port map( D => n3543, CK => CLK, RN => 
                           n413, Q => n3588, QN => n2140);
   REGISTERS_reg_2_15_inst : DFFR_X1 port map( D => n3542, CK => CLK, RN => 
                           n414, Q => n3611, QN => n2128);
   REGISTERS_reg_2_14_inst : DFFR_X1 port map( D => n3541, CK => CLK, RN => 
                           n414, Q => n3634, QN => n2116);
   REGISTERS_reg_2_13_inst : DFFR_X1 port map( D => n3540, CK => CLK, RN => 
                           n414, Q => n3657, QN => n2104);
   REGISTERS_reg_2_12_inst : DFFR_X1 port map( D => n3539, CK => CLK, RN => 
                           n414, Q => n3680, QN => n2092);
   REGISTERS_reg_2_11_inst : DFFR_X1 port map( D => n3538, CK => CLK, RN => 
                           n414, Q => n3703, QN => n2080);
   REGISTERS_reg_2_10_inst : DFFR_X1 port map( D => n3537, CK => CLK, RN => 
                           n414, Q => n3726, QN => n2068);
   REGISTERS_reg_2_9_inst : DFFR_X1 port map( D => n3536, CK => CLK, RN => n414
                           , Q => n3749, QN => n2056);
   REGISTERS_reg_2_8_inst : DFFR_X1 port map( D => n3535, CK => CLK, RN => n414
                           , Q => n3772, QN => n2044);
   REGISTERS_reg_2_7_inst : DFFR_X1 port map( D => n3534, CK => CLK, RN => n414
                           , Q => n3795, QN => n2032);
   REGISTERS_reg_2_6_inst : DFFR_X1 port map( D => n3533, CK => CLK, RN => n414
                           , Q => n3818, QN => n2020);
   REGISTERS_reg_2_5_inst : DFFR_X1 port map( D => n3532, CK => CLK, RN => n414
                           , Q => n3841, QN => n2008);
   REGISTERS_reg_2_4_inst : DFFR_X1 port map( D => n3531, CK => CLK, RN => n414
                           , Q => n3864, QN => n1996);
   REGISTERS_reg_2_3_inst : DFFR_X1 port map( D => n3530, CK => CLK, RN => n415
                           , Q => n3887, QN => n1984);
   REGISTERS_reg_2_2_inst : DFFR_X1 port map( D => n3529, CK => CLK, RN => n415
                           , Q => n3910, QN => n1972);
   REGISTERS_reg_2_1_inst : DFFR_X1 port map( D => n3528, CK => CLK, RN => n415
                           , Q => n3933, QN => n1960);
   REGISTERS_reg_2_0_inst : DFFR_X1 port map( D => n3527, CK => CLK, RN => n415
                           , Q => n3956, QN => n1946);
   REGISTERS_reg_28_31_inst : DFFR_X1 port map( D => n3110, CK => CLK, RN => 
                           n482, Q => n4093, QN => n_1658);
   REGISTERS_reg_28_30_inst : DFFR_X1 port map( D => n3109, CK => CLK, RN => 
                           n482, Q => n4092, QN => n_1659);
   REGISTERS_reg_28_29_inst : DFFR_X1 port map( D => n3108, CK => CLK, RN => 
                           n482, Q => n4091, QN => n_1660);
   REGISTERS_reg_28_28_inst : DFFR_X1 port map( D => n3107, CK => CLK, RN => 
                           n482, Q => n4090, QN => n_1661);
   REGISTERS_reg_28_27_inst : DFFR_X1 port map( D => n3106, CK => CLK, RN => 
                           n482, Q => n4089, QN => n_1662);
   REGISTERS_reg_28_26_inst : DFFR_X1 port map( D => n3105, CK => CLK, RN => 
                           n482, Q => n4088, QN => n_1663);
   REGISTERS_reg_28_25_inst : DFFR_X1 port map( D => n3104, CK => CLK, RN => 
                           n482, Q => n4087, QN => n_1664);
   REGISTERS_reg_28_24_inst : DFFR_X1 port map( D => n3103, CK => CLK, RN => 
                           n482, Q => n4086, QN => n_1665);
   REGISTERS_reg_28_23_inst : DFFR_X1 port map( D => n3102, CK => CLK, RN => 
                           n482, Q => n4085, QN => n_1666);
   REGISTERS_reg_28_22_inst : DFFR_X1 port map( D => n3101, CK => CLK, RN => 
                           n482, Q => n4084, QN => n_1667);
   REGISTERS_reg_28_21_inst : DFFR_X1 port map( D => n3100, CK => CLK, RN => 
                           n482, Q => n4083, QN => n_1668);
   REGISTERS_reg_28_20_inst : DFFR_X1 port map( D => n3099, CK => CLK, RN => 
                           n482, Q => n4082, QN => n_1669);
   REGISTERS_reg_28_19_inst : DFFR_X1 port map( D => n3098, CK => CLK, RN => 
                           n483, Q => n4081, QN => n_1670);
   REGISTERS_reg_28_18_inst : DFFR_X1 port map( D => n3097, CK => CLK, RN => 
                           n483, Q => n4080, QN => n_1671);
   REGISTERS_reg_28_17_inst : DFFR_X1 port map( D => n3096, CK => CLK, RN => 
                           n483, Q => n4079, QN => n_1672);
   REGISTERS_reg_28_16_inst : DFFR_X1 port map( D => n3095, CK => CLK, RN => 
                           n483, Q => n4078, QN => n_1673);
   REGISTERS_reg_28_15_inst : DFFR_X1 port map( D => n3094, CK => CLK, RN => 
                           n483, Q => n4077, QN => n_1674);
   REGISTERS_reg_28_14_inst : DFFR_X1 port map( D => n3093, CK => CLK, RN => 
                           n483, Q => n4076, QN => n_1675);
   REGISTERS_reg_28_13_inst : DFFR_X1 port map( D => n3092, CK => CLK, RN => 
                           n483, Q => n4075, QN => n_1676);
   REGISTERS_reg_28_12_inst : DFFR_X1 port map( D => n3091, CK => CLK, RN => 
                           n483, Q => n4074, QN => n_1677);
   REGISTERS_reg_28_11_inst : DFFR_X1 port map( D => n3090, CK => CLK, RN => 
                           n483, Q => n4073, QN => n_1678);
   REGISTERS_reg_28_10_inst : DFFR_X1 port map( D => n3089, CK => CLK, RN => 
                           n483, Q => n4072, QN => n_1679);
   REGISTERS_reg_28_9_inst : DFFR_X1 port map( D => n3088, CK => CLK, RN => 
                           n483, Q => n4071, QN => n_1680);
   REGISTERS_reg_28_8_inst : DFFR_X1 port map( D => n3087, CK => CLK, RN => 
                           n483, Q => n4070, QN => n_1681);
   REGISTERS_reg_28_7_inst : DFFR_X1 port map( D => n3086, CK => CLK, RN => 
                           n484, Q => n4069, QN => n_1682);
   REGISTERS_reg_28_6_inst : DFFR_X1 port map( D => n3085, CK => CLK, RN => 
                           n484, Q => n4068, QN => n_1683);
   REGISTERS_reg_28_5_inst : DFFR_X1 port map( D => n3084, CK => CLK, RN => 
                           n484, Q => n4067, QN => n_1684);
   REGISTERS_reg_28_4_inst : DFFR_X1 port map( D => n3083, CK => CLK, RN => 
                           n484, Q => n4066, QN => n_1685);
   REGISTERS_reg_28_3_inst : DFFR_X1 port map( D => n3082, CK => CLK, RN => 
                           n484, Q => n4065, QN => n_1686);
   REGISTERS_reg_28_2_inst : DFFR_X1 port map( D => n3081, CK => CLK, RN => 
                           n484, Q => n4064, QN => n_1687);
   REGISTERS_reg_28_1_inst : DFFR_X1 port map( D => n3080, CK => CLK, RN => 
                           n484, Q => n4063, QN => n_1688);
   REGISTERS_reg_28_0_inst : DFFR_X1 port map( D => n3079, CK => CLK, RN => 
                           n484, Q => n4062, QN => n_1689);
   REGISTERS_reg_18_31_inst : DFFR_X1 port map( D => n3302, CK => CLK, RN => 
                           n455, Q => n2676, QN => n_1690);
   REGISTERS_reg_27_31_inst : DFFR_X1 port map( D => n4413, CK => CLK, RN => 
                           RST, Q => n1518, QN => n_1691);
   REGISTERS_reg_27_30_inst : DFFR_X1 port map( D => n4412, CK => CLK, RN => 
                           n479, Q => n1517, QN => n_1692);
   REGISTERS_reg_27_29_inst : DFFR_X1 port map( D => n4411, CK => CLK, RN => 
                           n479, Q => n1516, QN => n_1693);
   REGISTERS_reg_27_28_inst : DFFR_X1 port map( D => n4410, CK => CLK, RN => 
                           n479, Q => n1515, QN => n_1694);
   REGISTERS_reg_27_27_inst : DFFR_X1 port map( D => n4409, CK => CLK, RN => 
                           n479, Q => n1514, QN => n_1695);
   REGISTERS_reg_27_26_inst : DFFR_X1 port map( D => n4408, CK => CLK, RN => 
                           n479, Q => n1513, QN => n_1696);
   REGISTERS_reg_27_25_inst : DFFR_X1 port map( D => n4407, CK => CLK, RN => 
                           n479, Q => n1512, QN => n_1697);
   REGISTERS_reg_27_24_inst : DFFR_X1 port map( D => n4406, CK => CLK, RN => 
                           n479, Q => n1511, QN => n_1698);
   REGISTERS_reg_27_23_inst : DFFR_X1 port map( D => n4405, CK => CLK, RN => 
                           n480, Q => n1510, QN => n_1699);
   REGISTERS_reg_27_22_inst : DFFR_X1 port map( D => n4404, CK => CLK, RN => 
                           n480, Q => n1509, QN => n_1700);
   REGISTERS_reg_27_21_inst : DFFR_X1 port map( D => n4403, CK => CLK, RN => 
                           n480, Q => n1508, QN => n_1701);
   REGISTERS_reg_27_20_inst : DFFR_X1 port map( D => n4402, CK => CLK, RN => 
                           n480, Q => n1507, QN => n_1702);
   REGISTERS_reg_27_19_inst : DFFR_X1 port map( D => n4401, CK => CLK, RN => 
                           n480, Q => n1506, QN => n_1703);
   REGISTERS_reg_27_18_inst : DFFR_X1 port map( D => n4400, CK => CLK, RN => 
                           n480, Q => n1505, QN => n_1704);
   REGISTERS_reg_27_17_inst : DFFR_X1 port map( D => n4399, CK => CLK, RN => 
                           n480, Q => n1504, QN => n_1705);
   REGISTERS_reg_27_16_inst : DFFR_X1 port map( D => n4398, CK => CLK, RN => 
                           n480, Q => n1503, QN => n_1706);
   REGISTERS_reg_27_15_inst : DFFR_X1 port map( D => n4397, CK => CLK, RN => 
                           n480, Q => n1502, QN => n_1707);
   REGISTERS_reg_27_14_inst : DFFR_X1 port map( D => n4396, CK => CLK, RN => 
                           n480, Q => n1501, QN => n_1708);
   REGISTERS_reg_27_13_inst : DFFR_X1 port map( D => n4395, CK => CLK, RN => 
                           n480, Q => n1500, QN => n_1709);
   REGISTERS_reg_27_12_inst : DFFR_X1 port map( D => n4394, CK => CLK, RN => 
                           n480, Q => n1499, QN => n_1710);
   REGISTERS_reg_27_11_inst : DFFR_X1 port map( D => n4393, CK => CLK, RN => 
                           n481, Q => n1498, QN => n_1711);
   REGISTERS_reg_27_10_inst : DFFR_X1 port map( D => n4392, CK => CLK, RN => 
                           n481, Q => n1497, QN => n_1712);
   REGISTERS_reg_27_9_inst : DFFR_X1 port map( D => n4391, CK => CLK, RN => 
                           n481, Q => n1496, QN => n_1713);
   REGISTERS_reg_27_8_inst : DFFR_X1 port map( D => n4390, CK => CLK, RN => 
                           n481, Q => n1495, QN => n_1714);
   REGISTERS_reg_27_7_inst : DFFR_X1 port map( D => n4389, CK => CLK, RN => 
                           n481, Q => n1494, QN => n_1715);
   REGISTERS_reg_27_6_inst : DFFR_X1 port map( D => n4388, CK => CLK, RN => 
                           n481, Q => n1493, QN => n_1716);
   REGISTERS_reg_27_5_inst : DFFR_X1 port map( D => n4387, CK => CLK, RN => 
                           n481, Q => n1492, QN => n_1717);
   REGISTERS_reg_27_4_inst : DFFR_X1 port map( D => n4386, CK => CLK, RN => 
                           n481, Q => n1491, QN => n_1718);
   REGISTERS_reg_27_3_inst : DFFR_X1 port map( D => n4385, CK => CLK, RN => 
                           n481, Q => n1490, QN => n_1719);
   REGISTERS_reg_27_2_inst : DFFR_X1 port map( D => n4384, CK => CLK, RN => 
                           n481, Q => n1489, QN => n_1720);
   REGISTERS_reg_27_1_inst : DFFR_X1 port map( D => n4383, CK => CLK, RN => 
                           n481, Q => n1488, QN => n_1721);
   REGISTERS_reg_27_0_inst : DFFR_X1 port map( D => n4382, CK => CLK, RN => 
                           n481, Q => n1487, QN => n_1722);
   REGISTERS_reg_4_31_inst : DFFR_X1 port map( D => n4317, CK => CLK, RN => 
                           n418, Q => n1874, QN => n_1723);
   REGISTERS_reg_4_30_inst : DFFR_X1 port map( D => n4316, CK => CLK, RN => 
                           n418, Q => n1873, QN => n_1724);
   REGISTERS_reg_4_29_inst : DFFR_X1 port map( D => n4315, CK => CLK, RN => 
                           n418, Q => n1872, QN => n_1725);
   REGISTERS_reg_4_28_inst : DFFR_X1 port map( D => n4314, CK => CLK, RN => 
                           n418, Q => n1871, QN => n_1726);
   REGISTERS_reg_4_27_inst : DFFR_X1 port map( D => n4313, CK => CLK, RN => 
                           n418, Q => n1870, QN => n_1727);
   REGISTERS_reg_4_26_inst : DFFR_X1 port map( D => n4312, CK => CLK, RN => 
                           n418, Q => n1869, QN => n_1728);
   REGISTERS_reg_4_25_inst : DFFR_X1 port map( D => n4311, CK => CLK, RN => 
                           n418, Q => n1868, QN => n_1729);
   REGISTERS_reg_4_24_inst : DFFR_X1 port map( D => n4310, CK => CLK, RN => 
                           n418, Q => n1867, QN => n_1730);
   REGISTERS_reg_4_23_inst : DFFR_X1 port map( D => n4309, CK => CLK, RN => 
                           n418, Q => n1866, QN => n_1731);
   REGISTERS_reg_4_22_inst : DFFR_X1 port map( D => n4308, CK => CLK, RN => 
                           n418, Q => n1865, QN => n_1732);
   REGISTERS_reg_4_21_inst : DFFR_X1 port map( D => n4307, CK => CLK, RN => 
                           n418, Q => n1864, QN => n_1733);
   REGISTERS_reg_4_20_inst : DFFR_X1 port map( D => n4306, CK => CLK, RN => 
                           n418, Q => n1863, QN => n_1734);
   REGISTERS_reg_4_19_inst : DFFR_X1 port map( D => n4305, CK => CLK, RN => 
                           n419, Q => n1862, QN => n_1735);
   REGISTERS_reg_4_18_inst : DFFR_X1 port map( D => n4304, CK => CLK, RN => 
                           n419, Q => n1861, QN => n_1736);
   REGISTERS_reg_4_17_inst : DFFR_X1 port map( D => n4303, CK => CLK, RN => 
                           n419, Q => n1860, QN => n_1737);
   REGISTERS_reg_4_16_inst : DFFR_X1 port map( D => n4302, CK => CLK, RN => 
                           n419, Q => n1859, QN => n_1738);
   REGISTERS_reg_4_15_inst : DFFR_X1 port map( D => n4301, CK => CLK, RN => 
                           n419, Q => n1858, QN => n_1739);
   REGISTERS_reg_4_14_inst : DFFR_X1 port map( D => n4300, CK => CLK, RN => 
                           n419, Q => n1857, QN => n_1740);
   REGISTERS_reg_4_13_inst : DFFR_X1 port map( D => n4299, CK => CLK, RN => 
                           n419, Q => n1856, QN => n_1741);
   REGISTERS_reg_4_12_inst : DFFR_X1 port map( D => n4298, CK => CLK, RN => 
                           n419, Q => n1855, QN => n_1742);
   REGISTERS_reg_4_11_inst : DFFR_X1 port map( D => n4297, CK => CLK, RN => 
                           n419, Q => n1854, QN => n_1743);
   REGISTERS_reg_4_10_inst : DFFR_X1 port map( D => n4296, CK => CLK, RN => 
                           n419, Q => n1853, QN => n_1744);
   REGISTERS_reg_4_9_inst : DFFR_X1 port map( D => n4295, CK => CLK, RN => n419
                           , Q => n1852, QN => n_1745);
   REGISTERS_reg_4_8_inst : DFFR_X1 port map( D => n4294, CK => CLK, RN => n419
                           , Q => n1851, QN => n_1746);
   REGISTERS_reg_4_7_inst : DFFR_X1 port map( D => n4293, CK => CLK, RN => n420
                           , Q => n1850, QN => n_1747);
   REGISTERS_reg_4_6_inst : DFFR_X1 port map( D => n4292, CK => CLK, RN => n420
                           , Q => n1849, QN => n_1748);
   REGISTERS_reg_4_5_inst : DFFR_X1 port map( D => n4291, CK => CLK, RN => n420
                           , Q => n1848, QN => n_1749);
   REGISTERS_reg_4_4_inst : DFFR_X1 port map( D => n4290, CK => CLK, RN => n420
                           , Q => n1847, QN => n_1750);
   REGISTERS_reg_4_3_inst : DFFR_X1 port map( D => n4289, CK => CLK, RN => n420
                           , Q => n1846, QN => n_1751);
   REGISTERS_reg_4_2_inst : DFFR_X1 port map( D => n4288, CK => CLK, RN => n420
                           , Q => n1845, QN => n_1752);
   REGISTERS_reg_4_1_inst : DFFR_X1 port map( D => n4287, CK => CLK, RN => n420
                           , Q => n1844, QN => n_1753);
   REGISTERS_reg_4_0_inst : DFFR_X1 port map( D => n4286, CK => CLK, RN => n420
                           , Q => n1843, QN => n_1754);
   REGISTERS_reg_26_31_inst : DFFR_X1 port map( D => n4350, CK => CLK, RN => 
                           n476, Q => n1550, QN => n_1755);
   REGISTERS_reg_26_30_inst : DFFR_X1 port map( D => n4381, CK => CLK, RN => 
                           n476, Q => n1549, QN => n_1756);
   REGISTERS_reg_26_29_inst : DFFR_X1 port map( D => n4380, CK => CLK, RN => 
                           n476, Q => n1548, QN => n_1757);
   REGISTERS_reg_26_28_inst : DFFR_X1 port map( D => n4379, CK => CLK, RN => 
                           n476, Q => n1547, QN => n_1758);
   REGISTERS_reg_26_27_inst : DFFR_X1 port map( D => n4378, CK => CLK, RN => 
                           n477, Q => n1546, QN => n_1759);
   REGISTERS_reg_26_26_inst : DFFR_X1 port map( D => n4377, CK => CLK, RN => 
                           n477, Q => n1545, QN => n_1760);
   REGISTERS_reg_26_25_inst : DFFR_X1 port map( D => n4376, CK => CLK, RN => 
                           n477, Q => n1544, QN => n_1761);
   REGISTERS_reg_26_24_inst : DFFR_X1 port map( D => n4375, CK => CLK, RN => 
                           n477, Q => n1543, QN => n_1762);
   REGISTERS_reg_26_23_inst : DFFR_X1 port map( D => n4374, CK => CLK, RN => 
                           n477, Q => n1542, QN => n_1763);
   REGISTERS_reg_26_22_inst : DFFR_X1 port map( D => n4373, CK => CLK, RN => 
                           n477, Q => n1541, QN => n_1764);
   REGISTERS_reg_26_21_inst : DFFR_X1 port map( D => n4372, CK => CLK, RN => 
                           n477, Q => n1540, QN => n_1765);
   REGISTERS_reg_26_20_inst : DFFR_X1 port map( D => n4371, CK => CLK, RN => 
                           n477, Q => n1539, QN => n_1766);
   REGISTERS_reg_26_19_inst : DFFR_X1 port map( D => n4370, CK => CLK, RN => 
                           n477, Q => n1538, QN => n_1767);
   REGISTERS_reg_26_18_inst : DFFR_X1 port map( D => n4369, CK => CLK, RN => 
                           n477, Q => n1537, QN => n_1768);
   REGISTERS_reg_26_17_inst : DFFR_X1 port map( D => n4368, CK => CLK, RN => 
                           n477, Q => n1536, QN => n_1769);
   REGISTERS_reg_26_16_inst : DFFR_X1 port map( D => n4367, CK => CLK, RN => 
                           n477, Q => n1535, QN => n_1770);
   REGISTERS_reg_26_15_inst : DFFR_X1 port map( D => n4366, CK => CLK, RN => 
                           n478, Q => n1534, QN => n_1771);
   REGISTERS_reg_26_14_inst : DFFR_X1 port map( D => n4365, CK => CLK, RN => 
                           n478, Q => n1533, QN => n_1772);
   REGISTERS_reg_26_13_inst : DFFR_X1 port map( D => n4364, CK => CLK, RN => 
                           n478, Q => n1532, QN => n_1773);
   REGISTERS_reg_26_12_inst : DFFR_X1 port map( D => n4363, CK => CLK, RN => 
                           n478, Q => n1531, QN => n_1774);
   REGISTERS_reg_26_11_inst : DFFR_X1 port map( D => n4362, CK => CLK, RN => 
                           n478, Q => n1530, QN => n_1775);
   REGISTERS_reg_26_10_inst : DFFR_X1 port map( D => n4361, CK => CLK, RN => 
                           n478, Q => n1529, QN => n_1776);
   REGISTERS_reg_26_9_inst : DFFR_X1 port map( D => n4360, CK => CLK, RN => 
                           n478, Q => n1528, QN => n_1777);
   REGISTERS_reg_26_8_inst : DFFR_X1 port map( D => n4359, CK => CLK, RN => 
                           n478, Q => n1527, QN => n_1778);
   REGISTERS_reg_26_7_inst : DFFR_X1 port map( D => n4358, CK => CLK, RN => 
                           n478, Q => n1526, QN => n_1779);
   REGISTERS_reg_26_6_inst : DFFR_X1 port map( D => n4357, CK => CLK, RN => 
                           n478, Q => n1525, QN => n_1780);
   REGISTERS_reg_26_5_inst : DFFR_X1 port map( D => n4356, CK => CLK, RN => 
                           n478, Q => n1524, QN => n_1781);
   REGISTERS_reg_26_4_inst : DFFR_X1 port map( D => n4355, CK => CLK, RN => 
                           n478, Q => n1523, QN => n_1782);
   REGISTERS_reg_26_3_inst : DFFR_X1 port map( D => n4354, CK => CLK, RN => 
                           n479, Q => n1522, QN => n_1783);
   REGISTERS_reg_26_2_inst : DFFR_X1 port map( D => n4353, CK => CLK, RN => 
                           n479, Q => n1521, QN => n_1784);
   REGISTERS_reg_26_1_inst : DFFR_X1 port map( D => n4352, CK => CLK, RN => 
                           n479, Q => n1520, QN => n_1785);
   REGISTERS_reg_26_0_inst : DFFR_X1 port map( D => n4351, CK => CLK, RN => 
                           n479, Q => n1519, QN => n_1786);
   REGISTERS_reg_17_31_inst : DFFR_X1 port map( D => n4541, CK => CLK, RN => 
                           n452, Q => n1648, QN => n_1787);
   REGISTERS_reg_17_30_inst : DFFR_X1 port map( D => n4540, CK => CLK, RN => 
                           n452, Q => n1647, QN => n_1788);
   REGISTERS_reg_17_29_inst : DFFR_X1 port map( D => n4539, CK => CLK, RN => 
                           n452, Q => n1646, QN => n_1789);
   REGISTERS_reg_17_28_inst : DFFR_X1 port map( D => n4538, CK => CLK, RN => 
                           n452, Q => n1645, QN => n_1790);
   REGISTERS_reg_17_27_inst : DFFR_X1 port map( D => n4537, CK => CLK, RN => 
                           n453, Q => n1644, QN => n_1791);
   REGISTERS_reg_17_26_inst : DFFR_X1 port map( D => n4536, CK => CLK, RN => 
                           n453, Q => n1643, QN => n_1792);
   REGISTERS_reg_17_25_inst : DFFR_X1 port map( D => n4535, CK => CLK, RN => 
                           n453, Q => n1642, QN => n_1793);
   REGISTERS_reg_17_24_inst : DFFR_X1 port map( D => n4534, CK => CLK, RN => 
                           n453, Q => n1641, QN => n_1794);
   REGISTERS_reg_17_23_inst : DFFR_X1 port map( D => n4533, CK => CLK, RN => 
                           n453, Q => n1640, QN => n_1795);
   REGISTERS_reg_17_22_inst : DFFR_X1 port map( D => n4532, CK => CLK, RN => 
                           n453, Q => n1639, QN => n_1796);
   REGISTERS_reg_17_21_inst : DFFR_X1 port map( D => n4531, CK => CLK, RN => 
                           n453, Q => n1638, QN => n_1797);
   REGISTERS_reg_17_20_inst : DFFR_X1 port map( D => n4530, CK => CLK, RN => 
                           n453, Q => n1637, QN => n_1798);
   REGISTERS_reg_17_19_inst : DFFR_X1 port map( D => n4529, CK => CLK, RN => 
                           n453, Q => n1636, QN => n_1799);
   REGISTERS_reg_17_18_inst : DFFR_X1 port map( D => n4528, CK => CLK, RN => 
                           n453, Q => n1635, QN => n_1800);
   REGISTERS_reg_17_17_inst : DFFR_X1 port map( D => n4527, CK => CLK, RN => 
                           n453, Q => n1634, QN => n_1801);
   REGISTERS_reg_17_16_inst : DFFR_X1 port map( D => n4526, CK => CLK, RN => 
                           n453, Q => n1633, QN => n_1802);
   REGISTERS_reg_17_15_inst : DFFR_X1 port map( D => n4525, CK => CLK, RN => 
                           n454, Q => n1632, QN => n_1803);
   REGISTERS_reg_17_14_inst : DFFR_X1 port map( D => n4524, CK => CLK, RN => 
                           n454, Q => n1631, QN => n_1804);
   REGISTERS_reg_17_13_inst : DFFR_X1 port map( D => n4523, CK => CLK, RN => 
                           n454, Q => n1630, QN => n_1805);
   REGISTERS_reg_17_12_inst : DFFR_X1 port map( D => n4522, CK => CLK, RN => 
                           n454, Q => n1629, QN => n_1806);
   REGISTERS_reg_17_11_inst : DFFR_X1 port map( D => n4521, CK => CLK, RN => 
                           n454, Q => n1628, QN => n_1807);
   REGISTERS_reg_17_10_inst : DFFR_X1 port map( D => n4520, CK => CLK, RN => 
                           n454, Q => n1627, QN => n_1808);
   REGISTERS_reg_17_9_inst : DFFR_X1 port map( D => n4519, CK => CLK, RN => 
                           n454, Q => n1626, QN => n_1809);
   REGISTERS_reg_17_8_inst : DFFR_X1 port map( D => n4518, CK => CLK, RN => 
                           n454, Q => n1625, QN => n_1810);
   REGISTERS_reg_17_7_inst : DFFR_X1 port map( D => n4517, CK => CLK, RN => 
                           n454, Q => n1624, QN => n_1811);
   REGISTERS_reg_17_6_inst : DFFR_X1 port map( D => n4516, CK => CLK, RN => 
                           n454, Q => n1623, QN => n_1812);
   REGISTERS_reg_17_5_inst : DFFR_X1 port map( D => n4515, CK => CLK, RN => 
                           n454, Q => n1622, QN => n_1813);
   REGISTERS_reg_17_4_inst : DFFR_X1 port map( D => n4514, CK => CLK, RN => 
                           n454, Q => n1621, QN => n_1814);
   REGISTERS_reg_17_3_inst : DFFR_X1 port map( D => n4513, CK => CLK, RN => 
                           n455, Q => n1620, QN => n_1815);
   REGISTERS_reg_17_2_inst : DFFR_X1 port map( D => n4512, CK => CLK, RN => 
                           n455, Q => n1619, QN => n_1816);
   REGISTERS_reg_17_1_inst : DFFR_X1 port map( D => n4511, CK => CLK, RN => 
                           n455, Q => n1618, QN => n_1817);
   REGISTERS_reg_17_0_inst : DFFR_X1 port map( D => n4510, CK => CLK, RN => 
                           n455, Q => n1617, QN => n_1818);
   REGISTERS_reg_5_31_inst : DFFR_X1 port map( D => n4349, CK => CLK, RN => 
                           n420, Q => n1842, QN => n2663);
   REGISTERS_reg_5_30_inst : DFFR_X1 port map( D => n4348, CK => CLK, RN => 
                           n420, Q => n1841, QN => n2686);
   REGISTERS_reg_5_29_inst : DFFR_X1 port map( D => n4347, CK => CLK, RN => 
                           n420, Q => n1840, QN => n2709);
   REGISTERS_reg_5_28_inst : DFFR_X1 port map( D => n4346, CK => CLK, RN => 
                           n420, Q => n1839, QN => n2732);
   REGISTERS_reg_5_27_inst : DFFR_X1 port map( D => n4345, CK => CLK, RN => 
                           n421, Q => n1838, QN => n2755);
   REGISTERS_reg_5_26_inst : DFFR_X1 port map( D => n4344, CK => CLK, RN => 
                           n421, Q => n1837, QN => n2778);
   REGISTERS_reg_5_25_inst : DFFR_X1 port map( D => n4343, CK => CLK, RN => 
                           n421, Q => n1836, QN => n2801);
   REGISTERS_reg_5_24_inst : DFFR_X1 port map( D => n4342, CK => CLK, RN => 
                           n421, Q => n1835, QN => n2824);
   REGISTERS_reg_5_23_inst : DFFR_X1 port map( D => n4341, CK => CLK, RN => 
                           n421, Q => n1834, QN => n2847);
   REGISTERS_reg_5_22_inst : DFFR_X1 port map( D => n4340, CK => CLK, RN => 
                           n421, Q => n1833, QN => n2870);
   REGISTERS_reg_5_21_inst : DFFR_X1 port map( D => n4339, CK => CLK, RN => 
                           n421, Q => n1832, QN => n2893);
   REGISTERS_reg_5_20_inst : DFFR_X1 port map( D => n4338, CK => CLK, RN => 
                           n421, Q => n1831, QN => n2916);
   REGISTERS_reg_5_19_inst : DFFR_X1 port map( D => n4337, CK => CLK, RN => 
                           n421, Q => n1830, QN => n2939);
   REGISTERS_reg_5_18_inst : DFFR_X1 port map( D => n4336, CK => CLK, RN => 
                           n421, Q => n1829, QN => n2962);
   REGISTERS_reg_5_17_inst : DFFR_X1 port map( D => n4335, CK => CLK, RN => 
                           n421, Q => n1828, QN => n3561);
   REGISTERS_reg_5_16_inst : DFFR_X1 port map( D => n4334, CK => CLK, RN => 
                           n421, Q => n1827, QN => n3584);
   REGISTERS_reg_5_15_inst : DFFR_X1 port map( D => n4333, CK => CLK, RN => 
                           n422, Q => n1826, QN => n3607);
   REGISTERS_reg_5_14_inst : DFFR_X1 port map( D => n4332, CK => CLK, RN => 
                           n422, Q => n1825, QN => n3630);
   REGISTERS_reg_5_13_inst : DFFR_X1 port map( D => n4331, CK => CLK, RN => 
                           n422, Q => n1824, QN => n3653);
   REGISTERS_reg_5_12_inst : DFFR_X1 port map( D => n4330, CK => CLK, RN => 
                           n422, Q => n1823, QN => n3676);
   REGISTERS_reg_5_11_inst : DFFR_X1 port map( D => n4329, CK => CLK, RN => 
                           n422, Q => n1822, QN => n3699);
   REGISTERS_reg_5_10_inst : DFFR_X1 port map( D => n4328, CK => CLK, RN => 
                           n422, Q => n1821, QN => n3722);
   REGISTERS_reg_5_9_inst : DFFR_X1 port map( D => n4327, CK => CLK, RN => n422
                           , Q => n1820, QN => n3745);
   REGISTERS_reg_5_8_inst : DFFR_X1 port map( D => n4326, CK => CLK, RN => n422
                           , Q => n1819, QN => n3768);
   REGISTERS_reg_5_7_inst : DFFR_X1 port map( D => n4325, CK => CLK, RN => n422
                           , Q => n1818, QN => n3791);
   REGISTERS_reg_5_6_inst : DFFR_X1 port map( D => n4324, CK => CLK, RN => n422
                           , Q => n1817, QN => n3814);
   REGISTERS_reg_5_5_inst : DFFR_X1 port map( D => n4323, CK => CLK, RN => n422
                           , Q => n1816, QN => n3837);
   REGISTERS_reg_5_4_inst : DFFR_X1 port map( D => n4322, CK => CLK, RN => n422
                           , Q => n1815, QN => n3860);
   REGISTERS_reg_5_3_inst : DFFR_X1 port map( D => n4321, CK => CLK, RN => n423
                           , Q => n1814, QN => n3883);
   REGISTERS_reg_5_2_inst : DFFR_X1 port map( D => n4320, CK => CLK, RN => n423
                           , Q => n1813, QN => n3906);
   REGISTERS_reg_5_1_inst : DFFR_X1 port map( D => n4319, CK => CLK, RN => n423
                           , Q => n1812, QN => n3929);
   REGISTERS_reg_5_0_inst : DFFR_X1 port map( D => n4318, CK => CLK, RN => n423
                           , Q => n1811, QN => n3952);
   REGISTERS_reg_31_31_inst : DFFR_X1 port map( D => n4477, CK => CLK, RN => 
                           n490, Q => n1454, QN => n3997);
   REGISTERS_reg_31_30_inst : DFFR_X1 port map( D => n4476, CK => CLK, RN => 
                           n490, Q => n1430, QN => n3996);
   REGISTERS_reg_31_29_inst : DFFR_X1 port map( D => n4475, CK => CLK, RN => 
                           n490, Q => n1414, QN => n3995);
   REGISTERS_reg_31_28_inst : DFFR_X1 port map( D => n4474, CK => CLK, RN => 
                           n490, Q => n1398, QN => n3994);
   REGISTERS_reg_31_27_inst : DFFR_X1 port map( D => n4473, CK => CLK, RN => 
                           n490, Q => n1382, QN => n3993);
   REGISTERS_reg_31_26_inst : DFFR_X1 port map( D => n4472, CK => CLK, RN => 
                           n490, Q => n1366, QN => n3992);
   REGISTERS_reg_31_25_inst : DFFR_X1 port map( D => n4471, CK => CLK, RN => 
                           n490, Q => n1350, QN => n3991);
   REGISTERS_reg_31_24_inst : DFFR_X1 port map( D => n4470, CK => CLK, RN => 
                           n490, Q => n1334, QN => n3990);
   REGISTERS_reg_31_23_inst : DFFR_X1 port map( D => n4469, CK => CLK, RN => 
                           n490, Q => n1318, QN => n3989);
   REGISTERS_reg_31_22_inst : DFFR_X1 port map( D => n4468, CK => CLK, RN => 
                           n490, Q => n1302, QN => n3988);
   REGISTERS_reg_31_21_inst : DFFR_X1 port map( D => n4467, CK => CLK, RN => 
                           n490, Q => n1286, QN => n3987);
   REGISTERS_reg_31_20_inst : DFFR_X1 port map( D => n4466, CK => CLK, RN => 
                           n490, Q => n1270, QN => n3986);
   REGISTERS_reg_31_19_inst : DFFR_X1 port map( D => n4465, CK => CLK, RN => 
                           n491, Q => n1254, QN => n3985);
   REGISTERS_reg_31_18_inst : DFFR_X1 port map( D => n4464, CK => CLK, RN => 
                           n491, Q => n1238, QN => n3984);
   REGISTERS_reg_31_17_inst : DFFR_X1 port map( D => n4463, CK => CLK, RN => 
                           n491, Q => n1222, QN => n3983);
   REGISTERS_reg_31_16_inst : DFFR_X1 port map( D => n4462, CK => CLK, RN => 
                           n491, Q => n1206, QN => n3982);
   REGISTERS_reg_31_15_inst : DFFR_X1 port map( D => n4461, CK => CLK, RN => 
                           n491, Q => n1190, QN => n3981);
   REGISTERS_reg_31_14_inst : DFFR_X1 port map( D => n4460, CK => CLK, RN => 
                           n491, Q => n1174, QN => n3980);
   REGISTERS_reg_31_13_inst : DFFR_X1 port map( D => n4459, CK => CLK, RN => 
                           n491, Q => n1158, QN => n3979);
   REGISTERS_reg_31_12_inst : DFFR_X1 port map( D => n4458, CK => CLK, RN => 
                           n491, Q => n1142, QN => n3978);
   REGISTERS_reg_31_11_inst : DFFR_X1 port map( D => n4457, CK => CLK, RN => 
                           n491, Q => n1126, QN => n3977);
   REGISTERS_reg_31_10_inst : DFFR_X1 port map( D => n4456, CK => CLK, RN => 
                           n491, Q => n1110, QN => n3976);
   REGISTERS_reg_31_9_inst : DFFR_X1 port map( D => n4455, CK => CLK, RN => 
                           n491, Q => n1094, QN => n3975);
   REGISTERS_reg_31_8_inst : DFFR_X1 port map( D => n4454, CK => CLK, RN => 
                           n491, Q => n1078, QN => n3974);
   REGISTERS_reg_31_7_inst : DFFR_X1 port map( D => n4453, CK => CLK, RN => 
                           n492, Q => n1062, QN => n3973);
   REGISTERS_reg_31_6_inst : DFFR_X1 port map( D => n4452, CK => CLK, RN => 
                           n492, Q => n1046, QN => n3972);
   REGISTERS_reg_31_5_inst : DFFR_X1 port map( D => n4451, CK => CLK, RN => 
                           n492, Q => n1030, QN => n3971);
   REGISTERS_reg_31_4_inst : DFFR_X1 port map( D => n4450, CK => CLK, RN => 
                           n492, Q => n1014, QN => n3970);
   REGISTERS_reg_31_3_inst : DFFR_X1 port map( D => n4449, CK => CLK, RN => 
                           n492, Q => n998, QN => n3969);
   REGISTERS_reg_31_2_inst : DFFR_X1 port map( D => n4448, CK => CLK, RN => 
                           n492, Q => n982, QN => n3968);
   REGISTERS_reg_31_1_inst : DFFR_X1 port map( D => n4447, CK => CLK, RN => 
                           n492, Q => n966, QN => n3967);
   REGISTERS_reg_31_0_inst : DFFR_X1 port map( D => n4446, CK => CLK, RN => 
                           n492, Q => n950, QN => n3966);
   REGISTERS_reg_21_31_inst : DFFR_X1 port map( D => n4605, CK => CLK, RN => 
                           n463, Q => n1584, QN => n2671);
   REGISTERS_reg_21_30_inst : DFFR_X1 port map( D => n4604, CK => CLK, RN => 
                           n463, Q => n1583, QN => n2694);
   REGISTERS_reg_21_29_inst : DFFR_X1 port map( D => n4603, CK => CLK, RN => 
                           n463, Q => n1582, QN => n2717);
   REGISTERS_reg_21_28_inst : DFFR_X1 port map( D => n4602, CK => CLK, RN => 
                           n463, Q => n1581, QN => n2740);
   REGISTERS_reg_21_27_inst : DFFR_X1 port map( D => n4601, CK => CLK, RN => 
                           n463, Q => n1580, QN => n2763);
   REGISTERS_reg_21_26_inst : DFFR_X1 port map( D => n4600, CK => CLK, RN => 
                           n463, Q => n1579, QN => n2786);
   REGISTERS_reg_21_25_inst : DFFR_X1 port map( D => n4599, CK => CLK, RN => 
                           n463, Q => n1578, QN => n2809);
   REGISTERS_reg_21_24_inst : DFFR_X1 port map( D => n4598, CK => CLK, RN => 
                           n463, Q => n1577, QN => n2832);
   REGISTERS_reg_21_23_inst : DFFR_X1 port map( D => n4597, CK => CLK, RN => 
                           n464, Q => n1576, QN => n2855);
   REGISTERS_reg_21_22_inst : DFFR_X1 port map( D => n4596, CK => CLK, RN => 
                           n464, Q => n1575, QN => n2878);
   REGISTERS_reg_21_21_inst : DFFR_X1 port map( D => n4595, CK => CLK, RN => 
                           n464, Q => n1574, QN => n2901);
   REGISTERS_reg_21_20_inst : DFFR_X1 port map( D => n4594, CK => CLK, RN => 
                           n464, Q => n1573, QN => n2924);
   REGISTERS_reg_21_19_inst : DFFR_X1 port map( D => n4593, CK => CLK, RN => 
                           n464, Q => n1572, QN => n2947);
   REGISTERS_reg_21_18_inst : DFFR_X1 port map( D => n4592, CK => CLK, RN => 
                           n464, Q => n1571, QN => n2970);
   REGISTERS_reg_21_17_inst : DFFR_X1 port map( D => n4591, CK => CLK, RN => 
                           n464, Q => n1570, QN => n3569);
   REGISTERS_reg_21_16_inst : DFFR_X1 port map( D => n4590, CK => CLK, RN => 
                           n464, Q => n1569, QN => n3592);
   REGISTERS_reg_21_15_inst : DFFR_X1 port map( D => n4589, CK => CLK, RN => 
                           n464, Q => n1568, QN => n3615);
   REGISTERS_reg_21_14_inst : DFFR_X1 port map( D => n4588, CK => CLK, RN => 
                           n464, Q => n1567, QN => n3638);
   REGISTERS_reg_21_13_inst : DFFR_X1 port map( D => n4587, CK => CLK, RN => 
                           n464, Q => n1566, QN => n3661);
   REGISTERS_reg_21_12_inst : DFFR_X1 port map( D => n4586, CK => CLK, RN => 
                           n464, Q => n1565, QN => n3684);
   REGISTERS_reg_21_11_inst : DFFR_X1 port map( D => n4585, CK => CLK, RN => 
                           n465, Q => n1564, QN => n3707);
   REGISTERS_reg_21_10_inst : DFFR_X1 port map( D => n4584, CK => CLK, RN => 
                           n465, Q => n1563, QN => n3730);
   REGISTERS_reg_21_9_inst : DFFR_X1 port map( D => n4583, CK => CLK, RN => 
                           n465, Q => n1562, QN => n3753);
   REGISTERS_reg_21_8_inst : DFFR_X1 port map( D => n4582, CK => CLK, RN => 
                           n465, Q => n1561, QN => n3776);
   REGISTERS_reg_21_7_inst : DFFR_X1 port map( D => n4581, CK => CLK, RN => 
                           n465, Q => n1560, QN => n3799);
   REGISTERS_reg_21_6_inst : DFFR_X1 port map( D => n4580, CK => CLK, RN => 
                           n465, Q => n1559, QN => n3822);
   REGISTERS_reg_21_5_inst : DFFR_X1 port map( D => n4579, CK => CLK, RN => 
                           n465, Q => n1558, QN => n3845);
   REGISTERS_reg_21_4_inst : DFFR_X1 port map( D => n4578, CK => CLK, RN => 
                           n465, Q => n1557, QN => n3868);
   REGISTERS_reg_21_3_inst : DFFR_X1 port map( D => n4577, CK => CLK, RN => 
                           n465, Q => n1556, QN => n3891);
   REGISTERS_reg_21_2_inst : DFFR_X1 port map( D => n4576, CK => CLK, RN => 
                           n465, Q => n1555, QN => n3914);
   REGISTERS_reg_21_1_inst : DFFR_X1 port map( D => n4575, CK => CLK, RN => 
                           n465, Q => n1554, QN => n3937);
   REGISTERS_reg_21_0_inst : DFFR_X1 port map( D => n4574, CK => CLK, RN => 
                           n465, Q => n1553, QN => n3960);
   REGISTERS_reg_12_31_inst : DFFR_X1 port map( D => n4221, CK => CLK, RN => 
                           n439, Q => n1744, QN => n2655);
   REGISTERS_reg_12_30_inst : DFFR_X1 port map( D => n4220, CK => CLK, RN => 
                           n439, Q => n1743, QN => n2678);
   REGISTERS_reg_12_29_inst : DFFR_X1 port map( D => n4219, CK => CLK, RN => 
                           n439, Q => n1742, QN => n2701);
   REGISTERS_reg_12_28_inst : DFFR_X1 port map( D => n4218, CK => CLK, RN => 
                           n439, Q => n1741, QN => n2724);
   REGISTERS_reg_12_27_inst : DFFR_X1 port map( D => n4217, CK => CLK, RN => 
                           n439, Q => n1740, QN => n2747);
   REGISTERS_reg_12_26_inst : DFFR_X1 port map( D => n4216, CK => CLK, RN => 
                           n439, Q => n1739, QN => n2770);
   REGISTERS_reg_12_25_inst : DFFR_X1 port map( D => n4215, CK => CLK, RN => 
                           n439, Q => n1738, QN => n2793);
   REGISTERS_reg_12_24_inst : DFFR_X1 port map( D => n4214, CK => CLK, RN => 
                           n439, Q => n1737, QN => n2816);
   REGISTERS_reg_12_23_inst : DFFR_X1 port map( D => n4213, CK => CLK, RN => 
                           n440, Q => n1736, QN => n2839);
   REGISTERS_reg_12_22_inst : DFFR_X1 port map( D => n4212, CK => CLK, RN => 
                           n440, Q => n1735, QN => n2862);
   REGISTERS_reg_12_21_inst : DFFR_X1 port map( D => n4211, CK => CLK, RN => 
                           n440, Q => n1734, QN => n2885);
   REGISTERS_reg_12_20_inst : DFFR_X1 port map( D => n4210, CK => CLK, RN => 
                           n440, Q => n1733, QN => n2908);
   REGISTERS_reg_12_19_inst : DFFR_X1 port map( D => n4209, CK => CLK, RN => 
                           n440, Q => n1732, QN => n2931);
   REGISTERS_reg_12_18_inst : DFFR_X1 port map( D => n4208, CK => CLK, RN => 
                           n440, Q => n1731, QN => n2954);
   REGISTERS_reg_12_17_inst : DFFR_X1 port map( D => n4207, CK => CLK, RN => 
                           n440, Q => n1730, QN => n2977);
   REGISTERS_reg_12_16_inst : DFFR_X1 port map( D => n4206, CK => CLK, RN => 
                           n440, Q => n1729, QN => n3576);
   REGISTERS_reg_12_15_inst : DFFR_X1 port map( D => n4205, CK => CLK, RN => 
                           n440, Q => n1728, QN => n3599);
   REGISTERS_reg_12_14_inst : DFFR_X1 port map( D => n4204, CK => CLK, RN => 
                           n440, Q => n1727, QN => n3622);
   REGISTERS_reg_12_13_inst : DFFR_X1 port map( D => n4203, CK => CLK, RN => 
                           n440, Q => n1726, QN => n3645);
   REGISTERS_reg_12_12_inst : DFFR_X1 port map( D => n4202, CK => CLK, RN => 
                           n440, Q => n1725, QN => n3668);
   REGISTERS_reg_12_11_inst : DFFR_X1 port map( D => n4201, CK => CLK, RN => 
                           n441, Q => n1724, QN => n3691);
   REGISTERS_reg_12_10_inst : DFFR_X1 port map( D => n4200, CK => CLK, RN => 
                           n441, Q => n1723, QN => n3714);
   REGISTERS_reg_12_9_inst : DFFR_X1 port map( D => n4199, CK => CLK, RN => 
                           n441, Q => n1722, QN => n3737);
   REGISTERS_reg_12_8_inst : DFFR_X1 port map( D => n4198, CK => CLK, RN => 
                           n441, Q => n1721, QN => n3760);
   REGISTERS_reg_12_7_inst : DFFR_X1 port map( D => n4197, CK => CLK, RN => 
                           n441, Q => n1720, QN => n3783);
   REGISTERS_reg_12_6_inst : DFFR_X1 port map( D => n4196, CK => CLK, RN => 
                           n441, Q => n1719, QN => n3806);
   REGISTERS_reg_12_5_inst : DFFR_X1 port map( D => n4195, CK => CLK, RN => 
                           n441, Q => n1718, QN => n3829);
   REGISTERS_reg_12_4_inst : DFFR_X1 port map( D => n4194, CK => CLK, RN => 
                           n441, Q => n1717, QN => n3852);
   REGISTERS_reg_12_3_inst : DFFR_X1 port map( D => n4193, CK => CLK, RN => 
                           n441, Q => n1716, QN => n3875);
   REGISTERS_reg_12_2_inst : DFFR_X1 port map( D => n4192, CK => CLK, RN => 
                           n441, Q => n1715, QN => n3898);
   REGISTERS_reg_12_1_inst : DFFR_X1 port map( D => n4191, CK => CLK, RN => 
                           n441, Q => n1714, QN => n3921);
   REGISTERS_reg_12_0_inst : DFFR_X1 port map( D => n4190, CK => CLK, RN => 
                           n441, Q => n1713, QN => n3944);
   REGISTERS_reg_8_31_inst : DFFR_X1 port map( D => n4157, CK => CLK, RN => 
                           n428, Q => n1808, QN => n2659);
   REGISTERS_reg_8_30_inst : DFFR_X1 port map( D => n4156, CK => CLK, RN => 
                           n428, Q => n1807, QN => n2682);
   REGISTERS_reg_8_29_inst : DFFR_X1 port map( D => n4155, CK => CLK, RN => 
                           n428, Q => n1806, QN => n2705);
   REGISTERS_reg_8_28_inst : DFFR_X1 port map( D => n4154, CK => CLK, RN => 
                           n428, Q => n1805, QN => n2728);
   REGISTERS_reg_8_27_inst : DFFR_X1 port map( D => n4153, CK => CLK, RN => 
                           n429, Q => n1804, QN => n2751);
   REGISTERS_reg_8_26_inst : DFFR_X1 port map( D => n4152, CK => CLK, RN => 
                           n429, Q => n1803, QN => n2774);
   REGISTERS_reg_8_25_inst : DFFR_X1 port map( D => n4151, CK => CLK, RN => 
                           n429, Q => n1802, QN => n2797);
   REGISTERS_reg_8_24_inst : DFFR_X1 port map( D => n4150, CK => CLK, RN => 
                           n429, Q => n1801, QN => n2820);
   REGISTERS_reg_8_23_inst : DFFR_X1 port map( D => n4149, CK => CLK, RN => 
                           n429, Q => n1800, QN => n2843);
   REGISTERS_reg_8_22_inst : DFFR_X1 port map( D => n4148, CK => CLK, RN => 
                           n429, Q => n1799, QN => n2866);
   REGISTERS_reg_8_21_inst : DFFR_X1 port map( D => n4147, CK => CLK, RN => 
                           n429, Q => n1798, QN => n2889);
   REGISTERS_reg_8_20_inst : DFFR_X1 port map( D => n4146, CK => CLK, RN => 
                           n429, Q => n1797, QN => n2912);
   REGISTERS_reg_8_19_inst : DFFR_X1 port map( D => n4145, CK => CLK, RN => 
                           n429, Q => n1796, QN => n2935);
   REGISTERS_reg_8_18_inst : DFFR_X1 port map( D => n4144, CK => CLK, RN => 
                           n429, Q => n1795, QN => n2958);
   REGISTERS_reg_8_17_inst : DFFR_X1 port map( D => n4143, CK => CLK, RN => 
                           n429, Q => n1794, QN => n2981);
   REGISTERS_reg_8_16_inst : DFFR_X1 port map( D => n4142, CK => CLK, RN => 
                           n429, Q => n1793, QN => n3580);
   REGISTERS_reg_8_15_inst : DFFR_X1 port map( D => n4141, CK => CLK, RN => 
                           n430, Q => n1792, QN => n3603);
   REGISTERS_reg_8_14_inst : DFFR_X1 port map( D => n4140, CK => CLK, RN => 
                           n430, Q => n1791, QN => n3626);
   REGISTERS_reg_8_13_inst : DFFR_X1 port map( D => n4139, CK => CLK, RN => 
                           n430, Q => n1790, QN => n3649);
   REGISTERS_reg_8_12_inst : DFFR_X1 port map( D => n4138, CK => CLK, RN => 
                           n430, Q => n1789, QN => n3672);
   REGISTERS_reg_8_11_inst : DFFR_X1 port map( D => n4137, CK => CLK, RN => 
                           n430, Q => n1788, QN => n3695);
   REGISTERS_reg_8_10_inst : DFFR_X1 port map( D => n4136, CK => CLK, RN => 
                           n430, Q => n1787, QN => n3718);
   REGISTERS_reg_8_9_inst : DFFR_X1 port map( D => n4135, CK => CLK, RN => n430
                           , Q => n1786, QN => n3741);
   REGISTERS_reg_8_8_inst : DFFR_X1 port map( D => n4134, CK => CLK, RN => n430
                           , Q => n1785, QN => n3764);
   REGISTERS_reg_8_7_inst : DFFR_X1 port map( D => n4133, CK => CLK, RN => n430
                           , Q => n1784, QN => n3787);
   REGISTERS_reg_8_6_inst : DFFR_X1 port map( D => n4132, CK => CLK, RN => n430
                           , Q => n1783, QN => n3810);
   REGISTERS_reg_8_5_inst : DFFR_X1 port map( D => n4131, CK => CLK, RN => n430
                           , Q => n1782, QN => n3833);
   REGISTERS_reg_8_4_inst : DFFR_X1 port map( D => n4130, CK => CLK, RN => n430
                           , Q => n1781, QN => n3856);
   REGISTERS_reg_8_3_inst : DFFR_X1 port map( D => n4129, CK => CLK, RN => n431
                           , Q => n1780, QN => n3879);
   REGISTERS_reg_8_2_inst : DFFR_X1 port map( D => n4128, CK => CLK, RN => n431
                           , Q => n1779, QN => n3902);
   REGISTERS_reg_8_1_inst : DFFR_X1 port map( D => n4127, CK => CLK, RN => n431
                           , Q => n1778, QN => n3925);
   REGISTERS_reg_8_0_inst : DFFR_X1 port map( D => n4126, CK => CLK, RN => n431
                           , Q => n1777, QN => n3948);
   REGISTERS_reg_30_31_inst : DFFR_X1 port map( D => n4445, CK => CLK, RN => 
                           n487, Q => n1486, QN => n4029);
   REGISTERS_reg_30_30_inst : DFFR_X1 port map( D => n4444, CK => CLK, RN => 
                           n487, Q => n1485, QN => n4028);
   REGISTERS_reg_30_29_inst : DFFR_X1 port map( D => n4443, CK => CLK, RN => 
                           n487, Q => n1484, QN => n4027);
   REGISTERS_reg_30_28_inst : DFFR_X1 port map( D => n4442, CK => CLK, RN => 
                           n487, Q => n1483, QN => n4026);
   REGISTERS_reg_30_27_inst : DFFR_X1 port map( D => n4441, CK => CLK, RN => 
                           n487, Q => n1482, QN => n4025);
   REGISTERS_reg_30_26_inst : DFFR_X1 port map( D => n4440, CK => CLK, RN => 
                           n487, Q => n1481, QN => n4024);
   REGISTERS_reg_30_25_inst : DFFR_X1 port map( D => n4439, CK => CLK, RN => 
                           n487, Q => n1480, QN => n4023);
   REGISTERS_reg_30_24_inst : DFFR_X1 port map( D => n4438, CK => CLK, RN => 
                           n487, Q => n1479, QN => n4022);
   REGISTERS_reg_30_23_inst : DFFR_X1 port map( D => n4437, CK => CLK, RN => 
                           n488, Q => n1478, QN => n4021);
   REGISTERS_reg_30_22_inst : DFFR_X1 port map( D => n4436, CK => CLK, RN => 
                           n488, Q => n1477, QN => n4020);
   REGISTERS_reg_30_21_inst : DFFR_X1 port map( D => n4435, CK => CLK, RN => 
                           n488, Q => n1476, QN => n4019);
   REGISTERS_reg_30_20_inst : DFFR_X1 port map( D => n4434, CK => CLK, RN => 
                           n488, Q => n1475, QN => n4018);
   REGISTERS_reg_30_19_inst : DFFR_X1 port map( D => n4433, CK => CLK, RN => 
                           n488, Q => n1474, QN => n4017);
   REGISTERS_reg_30_18_inst : DFFR_X1 port map( D => n4432, CK => CLK, RN => 
                           n488, Q => n1473, QN => n4016);
   REGISTERS_reg_30_17_inst : DFFR_X1 port map( D => n4431, CK => CLK, RN => 
                           n488, Q => n1472, QN => n4015);
   REGISTERS_reg_30_16_inst : DFFR_X1 port map( D => n4430, CK => CLK, RN => 
                           n488, Q => n1471, QN => n4014);
   REGISTERS_reg_30_15_inst : DFFR_X1 port map( D => n4429, CK => CLK, RN => 
                           n488, Q => n1470, QN => n4013);
   REGISTERS_reg_30_14_inst : DFFR_X1 port map( D => n4428, CK => CLK, RN => 
                           n488, Q => n1469, QN => n4012);
   REGISTERS_reg_30_13_inst : DFFR_X1 port map( D => n4427, CK => CLK, RN => 
                           n488, Q => n1468, QN => n4011);
   REGISTERS_reg_30_12_inst : DFFR_X1 port map( D => n4426, CK => CLK, RN => 
                           n488, Q => n1467, QN => n4010);
   REGISTERS_reg_30_11_inst : DFFR_X1 port map( D => n4425, CK => CLK, RN => 
                           n489, Q => n1466, QN => n4009);
   REGISTERS_reg_30_10_inst : DFFR_X1 port map( D => n4424, CK => CLK, RN => 
                           n489, Q => n1465, QN => n4008);
   REGISTERS_reg_30_9_inst : DFFR_X1 port map( D => n4423, CK => CLK, RN => 
                           n489, Q => n1464, QN => n4007);
   REGISTERS_reg_30_8_inst : DFFR_X1 port map( D => n4422, CK => CLK, RN => 
                           n489, Q => n1463, QN => n4006);
   REGISTERS_reg_30_7_inst : DFFR_X1 port map( D => n4421, CK => CLK, RN => 
                           n489, Q => n1462, QN => n4005);
   REGISTERS_reg_30_6_inst : DFFR_X1 port map( D => n4420, CK => CLK, RN => 
                           n489, Q => n1461, QN => n4004);
   REGISTERS_reg_30_5_inst : DFFR_X1 port map( D => n4419, CK => CLK, RN => 
                           n489, Q => n1460, QN => n4003);
   REGISTERS_reg_30_4_inst : DFFR_X1 port map( D => n4418, CK => CLK, RN => 
                           n489, Q => n1459, QN => n4002);
   REGISTERS_reg_30_3_inst : DFFR_X1 port map( D => n4417, CK => CLK, RN => 
                           n489, Q => n1458, QN => n4001);
   REGISTERS_reg_30_2_inst : DFFR_X1 port map( D => n4416, CK => CLK, RN => 
                           n489, Q => n1457, QN => n4000);
   REGISTERS_reg_30_1_inst : DFFR_X1 port map( D => n4415, CK => CLK, RN => 
                           n489, Q => n1456, QN => n3999);
   REGISTERS_reg_30_0_inst : DFFR_X1 port map( D => n4414, CK => CLK, RN => 
                           n489, Q => n1455, QN => n3998);
   REGISTERS_reg_20_31_inst : DFFR_X1 port map( D => n4573, CK => CLK, RN => 
                           n460, Q => n1616, QN => n2670);
   REGISTERS_reg_20_30_inst : DFFR_X1 port map( D => n4572, CK => CLK, RN => 
                           n460, Q => n1615, QN => n2693);
   REGISTERS_reg_20_29_inst : DFFR_X1 port map( D => n4571, CK => CLK, RN => 
                           n460, Q => n1614, QN => n2716);
   REGISTERS_reg_20_28_inst : DFFR_X1 port map( D => n4570, CK => CLK, RN => 
                           n460, Q => n1613, QN => n2739);
   REGISTERS_reg_20_27_inst : DFFR_X1 port map( D => n4569, CK => CLK, RN => 
                           n461, Q => n1612, QN => n2762);
   REGISTERS_reg_20_26_inst : DFFR_X1 port map( D => n4568, CK => CLK, RN => 
                           n461, Q => n1611, QN => n2785);
   REGISTERS_reg_20_25_inst : DFFR_X1 port map( D => n4567, CK => CLK, RN => 
                           n461, Q => n1610, QN => n2808);
   REGISTERS_reg_20_24_inst : DFFR_X1 port map( D => n4566, CK => CLK, RN => 
                           n461, Q => n1609, QN => n2831);
   REGISTERS_reg_20_23_inst : DFFR_X1 port map( D => n4565, CK => CLK, RN => 
                           n461, Q => n1608, QN => n2854);
   REGISTERS_reg_20_22_inst : DFFR_X1 port map( D => n4564, CK => CLK, RN => 
                           n461, Q => n1607, QN => n2877);
   REGISTERS_reg_20_21_inst : DFFR_X1 port map( D => n4563, CK => CLK, RN => 
                           n461, Q => n1606, QN => n2900);
   REGISTERS_reg_20_20_inst : DFFR_X1 port map( D => n4562, CK => CLK, RN => 
                           n461, Q => n1605, QN => n2923);
   REGISTERS_reg_20_19_inst : DFFR_X1 port map( D => n4561, CK => CLK, RN => 
                           n461, Q => n1604, QN => n2946);
   REGISTERS_reg_20_18_inst : DFFR_X1 port map( D => n4560, CK => CLK, RN => 
                           n461, Q => n1603, QN => n2969);
   REGISTERS_reg_20_17_inst : DFFR_X1 port map( D => n4559, CK => CLK, RN => 
                           n461, Q => n1602, QN => n3568);
   REGISTERS_reg_20_16_inst : DFFR_X1 port map( D => n4558, CK => CLK, RN => 
                           n461, Q => n1601, QN => n3591);
   REGISTERS_reg_20_15_inst : DFFR_X1 port map( D => n4557, CK => CLK, RN => 
                           n462, Q => n1600, QN => n3614);
   REGISTERS_reg_20_14_inst : DFFR_X1 port map( D => n4556, CK => CLK, RN => 
                           n462, Q => n1599, QN => n3637);
   REGISTERS_reg_20_13_inst : DFFR_X1 port map( D => n4555, CK => CLK, RN => 
                           n462, Q => n1598, QN => n3660);
   REGISTERS_reg_20_12_inst : DFFR_X1 port map( D => n4554, CK => CLK, RN => 
                           n462, Q => n1597, QN => n3683);
   REGISTERS_reg_20_11_inst : DFFR_X1 port map( D => n4553, CK => CLK, RN => 
                           n462, Q => n1596, QN => n3706);
   REGISTERS_reg_20_10_inst : DFFR_X1 port map( D => n4552, CK => CLK, RN => 
                           n462, Q => n1595, QN => n3729);
   REGISTERS_reg_20_9_inst : DFFR_X1 port map( D => n4551, CK => CLK, RN => 
                           n462, Q => n1594, QN => n3752);
   REGISTERS_reg_20_8_inst : DFFR_X1 port map( D => n4550, CK => CLK, RN => 
                           n462, Q => n1593, QN => n3775);
   REGISTERS_reg_20_7_inst : DFFR_X1 port map( D => n4549, CK => CLK, RN => 
                           n462, Q => n1592, QN => n3798);
   REGISTERS_reg_20_6_inst : DFFR_X1 port map( D => n4548, CK => CLK, RN => 
                           n462, Q => n1591, QN => n3821);
   REGISTERS_reg_20_5_inst : DFFR_X1 port map( D => n4547, CK => CLK, RN => 
                           n462, Q => n1590, QN => n3844);
   REGISTERS_reg_20_4_inst : DFFR_X1 port map( D => n4546, CK => CLK, RN => 
                           n462, Q => n1589, QN => n3867);
   REGISTERS_reg_20_3_inst : DFFR_X1 port map( D => n4545, CK => CLK, RN => 
                           n463, Q => n1588, QN => n3890);
   REGISTERS_reg_20_2_inst : DFFR_X1 port map( D => n4544, CK => CLK, RN => 
                           n463, Q => n1587, QN => n3913);
   REGISTERS_reg_20_1_inst : DFFR_X1 port map( D => n4543, CK => CLK, RN => 
                           n463, Q => n1586, QN => n3936);
   REGISTERS_reg_20_0_inst : DFFR_X1 port map( D => n4542, CK => CLK, RN => 
                           n463, Q => n1585, QN => n3959);
   REGISTERS_reg_16_31_inst : DFFR_X1 port map( D => n4509, CK => CLK, RN => 
                           n450, Q => n1680, QN => n2674);
   REGISTERS_reg_16_30_inst : DFFR_X1 port map( D => n4508, CK => CLK, RN => 
                           n450, Q => n1679, QN => n2697);
   REGISTERS_reg_16_29_inst : DFFR_X1 port map( D => n4507, CK => CLK, RN => 
                           n450, Q => n1678, QN => n2720);
   REGISTERS_reg_16_28_inst : DFFR_X1 port map( D => n4506, CK => CLK, RN => 
                           n450, Q => n1677, QN => n2743);
   REGISTERS_reg_16_27_inst : DFFR_X1 port map( D => n4505, CK => CLK, RN => 
                           n450, Q => n1676, QN => n2766);
   REGISTERS_reg_16_26_inst : DFFR_X1 port map( D => n4504, CK => CLK, RN => 
                           n450, Q => n1675, QN => n2789);
   REGISTERS_reg_16_25_inst : DFFR_X1 port map( D => n4503, CK => CLK, RN => 
                           n450, Q => n1674, QN => n2812);
   REGISTERS_reg_16_24_inst : DFFR_X1 port map( D => n4502, CK => CLK, RN => 
                           n450, Q => n1673, QN => n2835);
   REGISTERS_reg_16_23_inst : DFFR_X1 port map( D => n4501, CK => CLK, RN => 
                           n450, Q => n1672, QN => n2858);
   REGISTERS_reg_16_22_inst : DFFR_X1 port map( D => n4500, CK => CLK, RN => 
                           n450, Q => n1671, QN => n2881);
   REGISTERS_reg_16_21_inst : DFFR_X1 port map( D => n4499, CK => CLK, RN => 
                           n450, Q => n1670, QN => n2904);
   REGISTERS_reg_16_20_inst : DFFR_X1 port map( D => n4498, CK => CLK, RN => 
                           n450, Q => n1669, QN => n2927);
   REGISTERS_reg_16_19_inst : DFFR_X1 port map( D => n4497, CK => CLK, RN => 
                           n451, Q => n1668, QN => n2950);
   REGISTERS_reg_16_18_inst : DFFR_X1 port map( D => n4496, CK => CLK, RN => 
                           n451, Q => n1667, QN => n2973);
   REGISTERS_reg_16_17_inst : DFFR_X1 port map( D => n4495, CK => CLK, RN => 
                           n451, Q => n1666, QN => n3572);
   REGISTERS_reg_16_16_inst : DFFR_X1 port map( D => n4494, CK => CLK, RN => 
                           n451, Q => n1665, QN => n3595);
   REGISTERS_reg_16_15_inst : DFFR_X1 port map( D => n4493, CK => CLK, RN => 
                           n451, Q => n1664, QN => n3618);
   REGISTERS_reg_16_14_inst : DFFR_X1 port map( D => n4492, CK => CLK, RN => 
                           n451, Q => n1663, QN => n3641);
   REGISTERS_reg_16_13_inst : DFFR_X1 port map( D => n4491, CK => CLK, RN => 
                           n451, Q => n1662, QN => n3664);
   REGISTERS_reg_16_12_inst : DFFR_X1 port map( D => n4490, CK => CLK, RN => 
                           n451, Q => n1661, QN => n3687);
   REGISTERS_reg_16_11_inst : DFFR_X1 port map( D => n4489, CK => CLK, RN => 
                           n451, Q => n1660, QN => n3710);
   REGISTERS_reg_16_10_inst : DFFR_X1 port map( D => n4488, CK => CLK, RN => 
                           n451, Q => n1659, QN => n3733);
   REGISTERS_reg_16_9_inst : DFFR_X1 port map( D => n4487, CK => CLK, RN => 
                           n451, Q => n1658, QN => n3756);
   REGISTERS_reg_16_8_inst : DFFR_X1 port map( D => n4486, CK => CLK, RN => 
                           n451, Q => n1657, QN => n3779);
   REGISTERS_reg_16_7_inst : DFFR_X1 port map( D => n4485, CK => CLK, RN => 
                           n452, Q => n1656, QN => n3802);
   REGISTERS_reg_16_6_inst : DFFR_X1 port map( D => n4484, CK => CLK, RN => 
                           n452, Q => n1655, QN => n3825);
   REGISTERS_reg_16_5_inst : DFFR_X1 port map( D => n4483, CK => CLK, RN => 
                           n452, Q => n1654, QN => n3848);
   REGISTERS_reg_16_4_inst : DFFR_X1 port map( D => n4482, CK => CLK, RN => 
                           n452, Q => n1653, QN => n3871);
   REGISTERS_reg_16_3_inst : DFFR_X1 port map( D => n4481, CK => CLK, RN => 
                           n452, Q => n1652, QN => n3894);
   REGISTERS_reg_16_2_inst : DFFR_X1 port map( D => n4480, CK => CLK, RN => 
                           n452, Q => n1651, QN => n3917);
   REGISTERS_reg_16_1_inst : DFFR_X1 port map( D => n4479, CK => CLK, RN => 
                           n452, Q => n1650, QN => n3940);
   REGISTERS_reg_16_0_inst : DFFR_X1 port map( D => n4478, CK => CLK, RN => 
                           n452, Q => n1649, QN => n3963);
   REGISTERS_reg_13_31_inst : DFFR_X1 port map( D => n4253, CK => CLK, RN => 
                           n442, Q => n1712, QN => n2656);
   REGISTERS_reg_13_30_inst : DFFR_X1 port map( D => n4252, CK => CLK, RN => 
                           n442, Q => n1711, QN => n2679);
   REGISTERS_reg_13_29_inst : DFFR_X1 port map( D => n4251, CK => CLK, RN => 
                           n442, Q => n1710, QN => n2702);
   REGISTERS_reg_13_28_inst : DFFR_X1 port map( D => n4250, CK => CLK, RN => 
                           n442, Q => n1709, QN => n2725);
   REGISTERS_reg_13_27_inst : DFFR_X1 port map( D => n4249, CK => CLK, RN => 
                           n442, Q => n1708, QN => n2748);
   REGISTERS_reg_13_26_inst : DFFR_X1 port map( D => n4248, CK => CLK, RN => 
                           n442, Q => n1707, QN => n2771);
   REGISTERS_reg_13_25_inst : DFFR_X1 port map( D => n4247, CK => CLK, RN => 
                           n442, Q => n1706, QN => n2794);
   REGISTERS_reg_13_24_inst : DFFR_X1 port map( D => n4246, CK => CLK, RN => 
                           n442, Q => n1705, QN => n2817);
   REGISTERS_reg_13_23_inst : DFFR_X1 port map( D => n4245, CK => CLK, RN => 
                           n442, Q => n1704, QN => n2840);
   REGISTERS_reg_13_22_inst : DFFR_X1 port map( D => n4244, CK => CLK, RN => 
                           n442, Q => n1703, QN => n2863);
   REGISTERS_reg_13_21_inst : DFFR_X1 port map( D => n4243, CK => CLK, RN => 
                           n442, Q => n1702, QN => n2886);
   REGISTERS_reg_13_20_inst : DFFR_X1 port map( D => n4242, CK => CLK, RN => 
                           n442, Q => n1701, QN => n2909);
   REGISTERS_reg_13_19_inst : DFFR_X1 port map( D => n4241, CK => CLK, RN => 
                           n443, Q => n1700, QN => n2932);
   REGISTERS_reg_13_18_inst : DFFR_X1 port map( D => n4240, CK => CLK, RN => 
                           n443, Q => n1699, QN => n2955);
   REGISTERS_reg_13_17_inst : DFFR_X1 port map( D => n4239, CK => CLK, RN => 
                           n443, Q => n1698, QN => n2978);
   REGISTERS_reg_13_16_inst : DFFR_X1 port map( D => n4238, CK => CLK, RN => 
                           n443, Q => n1697, QN => n3577);
   REGISTERS_reg_13_15_inst : DFFR_X1 port map( D => n4237, CK => CLK, RN => 
                           n443, Q => n1696, QN => n3600);
   REGISTERS_reg_13_14_inst : DFFR_X1 port map( D => n4236, CK => CLK, RN => 
                           n443, Q => n1695, QN => n3623);
   REGISTERS_reg_13_13_inst : DFFR_X1 port map( D => n4235, CK => CLK, RN => 
                           n443, Q => n1694, QN => n3646);
   REGISTERS_reg_13_12_inst : DFFR_X1 port map( D => n4234, CK => CLK, RN => 
                           n443, Q => n1693, QN => n3669);
   REGISTERS_reg_13_11_inst : DFFR_X1 port map( D => n4233, CK => CLK, RN => 
                           n443, Q => n1692, QN => n3692);
   REGISTERS_reg_13_10_inst : DFFR_X1 port map( D => n4232, CK => CLK, RN => 
                           n443, Q => n1691, QN => n3715);
   REGISTERS_reg_13_9_inst : DFFR_X1 port map( D => n4231, CK => CLK, RN => 
                           n443, Q => n1690, QN => n3738);
   REGISTERS_reg_13_8_inst : DFFR_X1 port map( D => n4230, CK => CLK, RN => 
                           n443, Q => n1689, QN => n3761);
   REGISTERS_reg_13_7_inst : DFFR_X1 port map( D => n4229, CK => CLK, RN => 
                           n444, Q => n1688, QN => n3784);
   REGISTERS_reg_13_6_inst : DFFR_X1 port map( D => n4228, CK => CLK, RN => 
                           n444, Q => n1687, QN => n3807);
   REGISTERS_reg_13_5_inst : DFFR_X1 port map( D => n4227, CK => CLK, RN => 
                           n444, Q => n1686, QN => n3830);
   REGISTERS_reg_13_4_inst : DFFR_X1 port map( D => n4226, CK => CLK, RN => 
                           n444, Q => n1685, QN => n3853);
   REGISTERS_reg_13_3_inst : DFFR_X1 port map( D => n4225, CK => CLK, RN => 
                           n444, Q => n1684, QN => n3876);
   REGISTERS_reg_13_2_inst : DFFR_X1 port map( D => n4224, CK => CLK, RN => 
                           n444, Q => n1683, QN => n3899);
   REGISTERS_reg_13_1_inst : DFFR_X1 port map( D => n4223, CK => CLK, RN => 
                           n444, Q => n1682, QN => n3922);
   REGISTERS_reg_13_0_inst : DFFR_X1 port map( D => n4222, CK => CLK, RN => 
                           n444, Q => n1681, QN => n3945);
   REGISTERS_reg_9_31_inst : DFFR_X1 port map( D => n4189, CK => CLK, RN => 
                           n431, Q => n1776, QN => n2660);
   REGISTERS_reg_9_30_inst : DFFR_X1 port map( D => n4188, CK => CLK, RN => 
                           n431, Q => n1775, QN => n2683);
   REGISTERS_reg_9_29_inst : DFFR_X1 port map( D => n4187, CK => CLK, RN => 
                           n431, Q => n1774, QN => n2706);
   REGISTERS_reg_9_28_inst : DFFR_X1 port map( D => n4186, CK => CLK, RN => 
                           n431, Q => n1773, QN => n2729);
   REGISTERS_reg_9_27_inst : DFFR_X1 port map( D => n4185, CK => CLK, RN => 
                           n431, Q => n1772, QN => n2752);
   REGISTERS_reg_9_26_inst : DFFR_X1 port map( D => n4184, CK => CLK, RN => 
                           n431, Q => n1771, QN => n2775);
   REGISTERS_reg_9_25_inst : DFFR_X1 port map( D => n4183, CK => CLK, RN => 
                           n431, Q => n1770, QN => n2798);
   REGISTERS_reg_9_24_inst : DFFR_X1 port map( D => n4182, CK => CLK, RN => 
                           n431, Q => n1769, QN => n2821);
   REGISTERS_reg_9_23_inst : DFFR_X1 port map( D => n4181, CK => CLK, RN => 
                           n432, Q => n1768, QN => n2844);
   REGISTERS_reg_9_22_inst : DFFR_X1 port map( D => n4180, CK => CLK, RN => 
                           n432, Q => n1767, QN => n2867);
   REGISTERS_reg_9_21_inst : DFFR_X1 port map( D => n4179, CK => CLK, RN => 
                           n432, Q => n1766, QN => n2890);
   REGISTERS_reg_9_20_inst : DFFR_X1 port map( D => n4178, CK => CLK, RN => 
                           n432, Q => n1765, QN => n2913);
   REGISTERS_reg_9_19_inst : DFFR_X1 port map( D => n4177, CK => CLK, RN => 
                           n432, Q => n1764, QN => n2936);
   REGISTERS_reg_9_18_inst : DFFR_X1 port map( D => n4176, CK => CLK, RN => 
                           n432, Q => n1763, QN => n2959);
   REGISTERS_reg_9_17_inst : DFFR_X1 port map( D => n4175, CK => CLK, RN => 
                           n432, Q => n1762, QN => n2982);
   REGISTERS_reg_9_16_inst : DFFR_X1 port map( D => n4174, CK => CLK, RN => 
                           n432, Q => n1761, QN => n3581);
   REGISTERS_reg_9_15_inst : DFFR_X1 port map( D => n4173, CK => CLK, RN => 
                           n432, Q => n1760, QN => n3604);
   REGISTERS_reg_9_14_inst : DFFR_X1 port map( D => n4172, CK => CLK, RN => 
                           n432, Q => n1759, QN => n3627);
   REGISTERS_reg_9_13_inst : DFFR_X1 port map( D => n4171, CK => CLK, RN => 
                           n432, Q => n1758, QN => n3650);
   REGISTERS_reg_9_12_inst : DFFR_X1 port map( D => n4170, CK => CLK, RN => 
                           n432, Q => n1757, QN => n3673);
   REGISTERS_reg_9_11_inst : DFFR_X1 port map( D => n4169, CK => CLK, RN => 
                           n433, Q => n1756, QN => n3696);
   REGISTERS_reg_9_10_inst : DFFR_X1 port map( D => n4168, CK => CLK, RN => 
                           n433, Q => n1755, QN => n3719);
   REGISTERS_reg_9_9_inst : DFFR_X1 port map( D => n4167, CK => CLK, RN => n433
                           , Q => n1754, QN => n3742);
   REGISTERS_reg_9_8_inst : DFFR_X1 port map( D => n4166, CK => CLK, RN => n433
                           , Q => n1753, QN => n3765);
   REGISTERS_reg_9_7_inst : DFFR_X1 port map( D => n4165, CK => CLK, RN => n433
                           , Q => n1752, QN => n3788);
   REGISTERS_reg_9_6_inst : DFFR_X1 port map( D => n4164, CK => CLK, RN => n433
                           , Q => n1751, QN => n3811);
   REGISTERS_reg_9_5_inst : DFFR_X1 port map( D => n4163, CK => CLK, RN => n433
                           , Q => n1750, QN => n3834);
   REGISTERS_reg_9_4_inst : DFFR_X1 port map( D => n4162, CK => CLK, RN => n433
                           , Q => n1749, QN => n3857);
   REGISTERS_reg_9_3_inst : DFFR_X1 port map( D => n4161, CK => CLK, RN => n433
                           , Q => n1748, QN => n3880);
   REGISTERS_reg_9_2_inst : DFFR_X1 port map( D => n4160, CK => CLK, RN => n433
                           , Q => n1747, QN => n3903);
   REGISTERS_reg_9_1_inst : DFFR_X1 port map( D => n4159, CK => CLK, RN => n433
                           , Q => n1746, QN => n3926);
   REGISTERS_reg_9_0_inst : DFFR_X1 port map( D => n4158, CK => CLK, RN => n433
                           , Q => n1745, QN => n3949);
   REGISTERS_reg_1_31_inst : DFFR_X1 port map( D => n4285, CK => CLK, RN => 
                           n410, Q => n1906, QN => n4094);
   REGISTERS_reg_1_30_inst : DFFR_X1 port map( D => n4284, CK => CLK, RN => 
                           n410, Q => n1905, QN => n4095);
   REGISTERS_reg_1_29_inst : DFFR_X1 port map( D => n4283, CK => CLK, RN => 
                           n410, Q => n1904, QN => n4096);
   REGISTERS_reg_1_28_inst : DFFR_X1 port map( D => n4282, CK => CLK, RN => 
                           n410, Q => n1903, QN => n4097);
   REGISTERS_reg_1_27_inst : DFFR_X1 port map( D => n4281, CK => CLK, RN => 
                           n410, Q => n1902, QN => n4098);
   REGISTERS_reg_1_26_inst : DFFR_X1 port map( D => n4280, CK => CLK, RN => 
                           n410, Q => n1901, QN => n4099);
   REGISTERS_reg_1_25_inst : DFFR_X1 port map( D => n4279, CK => CLK, RN => 
                           n410, Q => n1900, QN => n4100);
   REGISTERS_reg_1_24_inst : DFFR_X1 port map( D => n4278, CK => CLK, RN => 
                           n410, Q => n1899, QN => n4101);
   REGISTERS_reg_1_23_inst : DFFR_X1 port map( D => n4277, CK => CLK, RN => 
                           n410, Q => n1898, QN => n4102);
   REGISTERS_reg_1_22_inst : DFFR_X1 port map( D => n4276, CK => CLK, RN => 
                           n410, Q => n1897, QN => n4103);
   REGISTERS_reg_1_21_inst : DFFR_X1 port map( D => n4275, CK => CLK, RN => 
                           n410, Q => n1896, QN => n4104);
   REGISTERS_reg_1_20_inst : DFFR_X1 port map( D => n4274, CK => CLK, RN => 
                           n410, Q => n1895, QN => n4105);
   REGISTERS_reg_1_19_inst : DFFR_X1 port map( D => n4273, CK => CLK, RN => 
                           n411, Q => n1894, QN => n4106);
   REGISTERS_reg_1_18_inst : DFFR_X1 port map( D => n4272, CK => CLK, RN => 
                           n411, Q => n1893, QN => n4107);
   REGISTERS_reg_1_17_inst : DFFR_X1 port map( D => n4271, CK => CLK, RN => 
                           n411, Q => n1892, QN => n4108);
   REGISTERS_reg_1_16_inst : DFFR_X1 port map( D => n4270, CK => CLK, RN => 
                           n411, Q => n1891, QN => n4109);
   REGISTERS_reg_1_15_inst : DFFR_X1 port map( D => n4269, CK => CLK, RN => 
                           n411, Q => n1890, QN => n4110);
   REGISTERS_reg_1_14_inst : DFFR_X1 port map( D => n4268, CK => CLK, RN => 
                           n411, Q => n1889, QN => n4111);
   REGISTERS_reg_1_13_inst : DFFR_X1 port map( D => n4267, CK => CLK, RN => 
                           n411, Q => n1888, QN => n4112);
   REGISTERS_reg_1_12_inst : DFFR_X1 port map( D => n4266, CK => CLK, RN => 
                           n411, Q => n1887, QN => n4113);
   REGISTERS_reg_1_11_inst : DFFR_X1 port map( D => n4265, CK => CLK, RN => 
                           n411, Q => n1886, QN => n4114);
   REGISTERS_reg_1_10_inst : DFFR_X1 port map( D => n4264, CK => CLK, RN => 
                           n411, Q => n1885, QN => n4115);
   REGISTERS_reg_1_9_inst : DFFR_X1 port map( D => n4263, CK => CLK, RN => n411
                           , Q => n1884, QN => n4116);
   REGISTERS_reg_1_8_inst : DFFR_X1 port map( D => n4262, CK => CLK, RN => n411
                           , Q => n1883, QN => n4117);
   REGISTERS_reg_1_7_inst : DFFR_X1 port map( D => n4261, CK => CLK, RN => n412
                           , Q => n1882, QN => n4118);
   REGISTERS_reg_1_6_inst : DFFR_X1 port map( D => n4260, CK => CLK, RN => n412
                           , Q => n1881, QN => n4119);
   REGISTERS_reg_1_5_inst : DFFR_X1 port map( D => n4259, CK => CLK, RN => n412
                           , Q => n1880, QN => n4120);
   REGISTERS_reg_1_4_inst : DFFR_X1 port map( D => n4258, CK => CLK, RN => n412
                           , Q => n1879, QN => n4121);
   REGISTERS_reg_1_3_inst : DFFR_X1 port map( D => n4257, CK => CLK, RN => n412
                           , Q => n1878, QN => n4122);
   REGISTERS_reg_1_2_inst : DFFR_X1 port map( D => n4256, CK => CLK, RN => n412
                           , Q => n1877, QN => n4123);
   REGISTERS_reg_1_1_inst : DFFR_X1 port map( D => n4255, CK => CLK, RN => n412
                           , Q => n1876, QN => n4124);
   REGISTERS_reg_1_0_inst : DFFR_X1 port map( D => n4254, CK => CLK, RN => n412
                           , Q => n1875, QN => n4125);
   U2 : AND3_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), A3 => n1908, ZN => 
                           n1);
   U3 : AND3_X1 port map( A1 => ADD_WR(4), A2 => n1908, A3 => n1810, ZN => n2);
   U4 : AND3_X1 port map( A1 => ADD_WR(3), A2 => n1908, A3 => n1809, ZN => n3);
   U5 : AND3_X1 port map( A1 => n1908, A2 => n1810, A3 => n1809, ZN => n4);
   U6 : AND2_X1 port map( A1 => n45, A2 => ADD_WR(0), ZN => n5);
   U7 : AND2_X1 port map( A1 => n45, A2 => n1907, ZN => n6);
   U8 : AND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => n1551, ZN => 
                           n7);
   U9 : AND3_X1 port map( A1 => ADD_WR(1), A2 => n1907, A3 => n1551, ZN => n8);
   U10 : AND3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => n1552, ZN =>
                           n9);
   U11 : AND3_X1 port map( A1 => ADD_WR(2), A2 => n1907, A3 => n1552, ZN => n10
                           );
   U12 : AND3_X1 port map( A1 => ADD_WR(0), A2 => n1552, A3 => n1551, ZN => n11
                           );
   U13 : AND3_X1 port map( A1 => n1907, A2 => n1552, A3 => n1551, ZN => n12);
   U14 : AND2_X1 port map( A1 => n1, A2 => n5, ZN => n13);
   U15 : AND2_X1 port map( A1 => n1, A2 => n6, ZN => n14);
   U16 : AND2_X1 port map( A1 => n1, A2 => n9, ZN => n15);
   U17 : AND2_X1 port map( A1 => n1, A2 => n10, ZN => n16);
   U18 : AND2_X1 port map( A1 => n1, A2 => n7, ZN => n17);
   U19 : AND2_X1 port map( A1 => n1, A2 => n8, ZN => n18);
   U20 : AND2_X1 port map( A1 => n1, A2 => n11, ZN => n19);
   U21 : AND2_X1 port map( A1 => n1, A2 => n12, ZN => n20);
   U22 : AND2_X1 port map( A1 => n2, A2 => n5, ZN => n21);
   U23 : AND2_X1 port map( A1 => n2, A2 => n6, ZN => n22);
   U24 : AND2_X1 port map( A1 => n2, A2 => n9, ZN => n23);
   U25 : AND2_X1 port map( A1 => n2, A2 => n10, ZN => n24);
   U26 : AND2_X1 port map( A1 => n2, A2 => n7, ZN => n25);
   U27 : AND2_X1 port map( A1 => n2, A2 => n8, ZN => n26);
   U28 : AND2_X1 port map( A1 => n2, A2 => n11, ZN => n27);
   U29 : AND2_X1 port map( A1 => n2, A2 => n12, ZN => n28);
   U30 : AND2_X1 port map( A1 => n3, A2 => n5, ZN => n29);
   U31 : AND2_X1 port map( A1 => n3, A2 => n6, ZN => n30);
   U32 : AND2_X1 port map( A1 => n3, A2 => n9, ZN => n31);
   U33 : AND2_X1 port map( A1 => n3, A2 => n10, ZN => n32);
   U34 : AND2_X1 port map( A1 => n3, A2 => n7, ZN => n33);
   U35 : AND2_X1 port map( A1 => n3, A2 => n8, ZN => n34);
   U36 : AND2_X1 port map( A1 => n3, A2 => n11, ZN => n35);
   U37 : AND2_X1 port map( A1 => n3, A2 => n12, ZN => n36);
   U38 : AND2_X1 port map( A1 => n2349, A2 => n85, ZN => n37);
   U39 : AND2_X1 port map( A1 => n2353, A2 => n85, ZN => n38);
   U40 : AND2_X1 port map( A1 => n2356, A2 => n85, ZN => n39);
   U41 : AND2_X1 port map( A1 => n2360, A2 => n85, ZN => n40);
   U42 : AND2_X1 port map( A1 => n1912, A2 => n142, ZN => n41);
   U43 : AND2_X1 port map( A1 => n1916, A2 => n142, ZN => n42);
   U44 : AND2_X1 port map( A1 => n1919, A2 => n142, ZN => n43);
   U45 : AND2_X1 port map( A1 => n1924, A2 => n142, ZN => n44);
   U46 : AND2_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), ZN => n45);
   U47 : AND2_X1 port map( A1 => ENABLE, A2 => n492, ZN => n46);
   U48 : AND2_X1 port map( A1 => n5, A2 => n4, ZN => n47);
   U49 : AND2_X1 port map( A1 => n6, A2 => n4, ZN => n48);
   U50 : AND2_X1 port map( A1 => n9, A2 => n4, ZN => n49);
   U51 : AND2_X1 port map( A1 => n10, A2 => n4, ZN => n50);
   U52 : AND2_X1 port map( A1 => n7, A2 => n4, ZN => n51);
   U53 : AND2_X1 port map( A1 => n8, A2 => n4, ZN => n52);
   U54 : AND2_X1 port map( A1 => n11, A2 => n4, ZN => n53);
   U55 : NOR2_X1 port map( A1 => n2346, A2 => n516, ZN => n54);
   U56 : NOR2_X1 port map( A1 => n2350, A2 => n516, ZN => n55);
   U57 : NOR2_X1 port map( A1 => n2354, A2 => n516, ZN => n56);
   U58 : NOR2_X1 port map( A1 => n1909, A2 => n944, ZN => n57);
   U59 : NOR2_X1 port map( A1 => n1913, A2 => n944, ZN => n58);
   U60 : NOR2_X1 port map( A1 => n1917, A2 => n944, ZN => n59);
   U61 : AND2_X1 port map( A1 => RD1, A2 => n46, ZN => n60);
   U62 : AND2_X1 port map( A1 => RD2, A2 => n46, ZN => n61);
   U63 : NAND2_X1 port map( A1 => n2611, A2 => n2594, ZN => n62);
   U64 : NAND2_X1 port map( A1 => n2332, A2 => n2312, ZN => n63);
   U65 : NAND2_X1 port map( A1 => n2611, A2 => n2598, ZN => n64);
   U66 : NAND2_X1 port map( A1 => n2332, A2 => n2316, ZN => n65);
   U67 : AND2_X1 port map( A1 => n2617, A2 => n2616, ZN => n66);
   U68 : AND2_X1 port map( A1 => n2340, A2 => n2339, ZN => n67);
   U69 : BUF_X1 port map( A => n493, Z => n492);
   U70 : BUF_X1 port map( A => n1442, Z => n146);
   U71 : BUF_X1 port map( A => n1442, Z => n147);
   U72 : BUF_X1 port map( A => n1442, Z => n148);
   U73 : BUF_X1 port map( A => n1944, Z => n314);
   U74 : BUF_X1 port map( A => n1944, Z => n315);
   U75 : BUF_X1 port map( A => n43, Z => n164);
   U76 : BUF_X1 port map( A => n42, Z => n152);
   U77 : BUF_X1 port map( A => n43, Z => n165);
   U78 : BUF_X1 port map( A => n42, Z => n153);
   U79 : BUF_X1 port map( A => n1436, Z => n131);
   U80 : BUF_X1 port map( A => n1436, Z => n132);
   U81 : BUF_X1 port map( A => n63, Z => n128);
   U82 : BUF_X1 port map( A => n63, Z => n129);
   U83 : BUF_X1 port map( A => n1934, Z => n297);
   U84 : BUF_X1 port map( A => n1934, Z => n296);
   U85 : BUF_X1 port map( A => n1929, Z => n285);
   U86 : BUF_X1 port map( A => n1929, Z => n284);
   U87 : BUF_X1 port map( A => n2378, Z => n362);
   U88 : BUF_X1 port map( A => n2378, Z => n363);
   U89 : BUF_X1 port map( A => n39, Z => n107);
   U90 : BUF_X1 port map( A => n38, Z => n95);
   U91 : BUF_X1 port map( A => n37, Z => n80);
   U92 : BUF_X1 port map( A => n39, Z => n108);
   U93 : BUF_X1 port map( A => n38, Z => n96);
   U94 : BUF_X1 port map( A => n37, Z => n81);
   U95 : BUF_X1 port map( A => n41, Z => n137);
   U96 : BUF_X1 port map( A => n41, Z => n138);
   U97 : BUF_X1 port map( A => n44, Z => n179);
   U98 : BUF_X1 port map( A => n44, Z => n180);
   U99 : BUF_X1 port map( A => n1949, Z => n321);
   U100 : BUF_X1 port map( A => n1949, Z => n320);
   U101 : BUF_X1 port map( A => n1937, Z => n303);
   U102 : BUF_X1 port map( A => n1932, Z => n291);
   U103 : BUF_X1 port map( A => n1937, Z => n302);
   U104 : BUF_X1 port map( A => n1932, Z => n290);
   U105 : BUF_X1 port map( A => n2359, Z => n326);
   U106 : BUF_X1 port map( A => n2359, Z => n327);
   U107 : BUF_X1 port map( A => n1943, Z => n312);
   U108 : BUF_X1 port map( A => n1923, Z => n279);
   U109 : BUF_X1 port map( A => n1943, Z => n311);
   U110 : BUF_X1 port map( A => n1923, Z => n278);
   U111 : BUF_X1 port map( A => n924, Z => n101);
   U112 : BUF_X1 port map( A => n921, Z => n89);
   U113 : BUF_X1 port map( A => n916, Z => n74);
   U114 : BUF_X1 port map( A => n924, Z => n102);
   U115 : BUF_X1 port map( A => n921, Z => n90);
   U116 : BUF_X1 port map( A => n916, Z => n75);
   U117 : BUF_X1 port map( A => n1445, Z => n158);
   U118 : BUF_X1 port map( A => n1445, Z => n159);
   U119 : BUF_X1 port map( A => n1947, Z => n318);
   U120 : BUF_X1 port map( A => n1947, Z => n317);
   U121 : BUF_X1 port map( A => n2358, Z => n323);
   U122 : BUF_X1 port map( A => n2358, Z => n324);
   U123 : BUF_X1 port map( A => n1921, Z => n276);
   U124 : BUF_X1 port map( A => n1921, Z => n275);
   U125 : BUF_X1 port map( A => n1936, Z => n300);
   U126 : BUF_X1 port map( A => n1931, Z => n288);
   U127 : BUF_X1 port map( A => n1936, Z => n299);
   U128 : BUF_X1 port map( A => n1931, Z => n287);
   U129 : BUF_X1 port map( A => n1941, Z => n309);
   U130 : BUF_X1 port map( A => n1941, Z => n308);
   U131 : BUF_X1 port map( A => n925, Z => n104);
   U132 : BUF_X1 port map( A => n925, Z => n105);
   U133 : BUF_X1 port map( A => n1446, Z => n161);
   U134 : BUF_X1 port map( A => n1446, Z => n162);
   U135 : BUF_X1 port map( A => n1928, Z => n282);
   U136 : BUF_X1 port map( A => n1928, Z => n281);
   U137 : BUF_X1 port map( A => n1933, Z => n294);
   U138 : BUF_X1 port map( A => n1933, Z => n293);
   U139 : BUF_X1 port map( A => n1938, Z => n305);
   U140 : BUF_X1 port map( A => n1938, Z => n306);
   U141 : BUF_X1 port map( A => n40, Z => n122);
   U142 : BUF_X1 port map( A => n40, Z => n123);
   U143 : BUF_X1 port map( A => n65, Z => n125);
   U144 : BUF_X1 port map( A => n65, Z => n126);
   U145 : BUF_X1 port map( A => n83, Z => n85);
   U146 : BUF_X1 port map( A => n140, Z => n142);
   U147 : BUF_X1 port map( A => n43, Z => n166);
   U148 : BUF_X1 port map( A => n42, Z => n154);
   U149 : BUF_X1 port map( A => n1944, Z => n316);
   U150 : BUF_X1 port map( A => n83, Z => n86);
   U151 : BUF_X1 port map( A => n140, Z => n143);
   U152 : BUF_X1 port map( A => n84, Z => n87);
   U153 : BUF_X1 port map( A => n141, Z => n144);
   U154 : BUF_X1 port map( A => n1436, Z => n133);
   U155 : BUF_X1 port map( A => n63, Z => n130);
   U156 : BUF_X1 port map( A => n1934, Z => n298);
   U157 : BUF_X1 port map( A => n1929, Z => n286);
   U158 : BUF_X1 port map( A => n2378, Z => n364);
   U159 : BUF_X1 port map( A => n39, Z => n109);
   U160 : BUF_X1 port map( A => n38, Z => n97);
   U161 : BUF_X1 port map( A => n37, Z => n82);
   U162 : BUF_X1 port map( A => n41, Z => n139);
   U163 : BUF_X1 port map( A => n44, Z => n181);
   U164 : BUF_X1 port map( A => n1949, Z => n322);
   U165 : BUF_X1 port map( A => n2359, Z => n328);
   U166 : BUF_X1 port map( A => n1943, Z => n313);
   U167 : BUF_X1 port map( A => n1923, Z => n280);
   U168 : BUF_X1 port map( A => n1937, Z => n304);
   U169 : BUF_X1 port map( A => n1932, Z => n292);
   U170 : BUF_X1 port map( A => n924, Z => n103);
   U171 : BUF_X1 port map( A => n921, Z => n91);
   U172 : BUF_X1 port map( A => n916, Z => n76);
   U173 : BUF_X1 port map( A => n1445, Z => n160);
   U174 : BUF_X1 port map( A => n1947, Z => n319);
   U175 : BUF_X1 port map( A => n2358, Z => n325);
   U176 : BUF_X1 port map( A => n1921, Z => n277);
   U177 : BUF_X1 port map( A => n1941, Z => n310);
   U178 : BUF_X1 port map( A => n1936, Z => n301);
   U179 : BUF_X1 port map( A => n1931, Z => n289);
   U180 : BUF_X1 port map( A => n925, Z => n106);
   U181 : BUF_X1 port map( A => n1446, Z => n163);
   U182 : BUF_X1 port map( A => n1928, Z => n283);
   U183 : BUF_X1 port map( A => n1933, Z => n295);
   U184 : BUF_X1 port map( A => n1938, Z => n307);
   U185 : BUF_X1 port map( A => n40, Z => n124);
   U186 : BUF_X1 port map( A => n65, Z => n127);
   U187 : BUF_X1 port map( A => n403, Z => n493);
   U188 : BUF_X1 port map( A => n84, Z => n88);
   U189 : BUF_X1 port map( A => n141, Z => n145);
   U190 : BUF_X1 port map( A => n403, Z => n494);
   U191 : BUF_X1 port map( A => n403, Z => n495);
   U192 : BUF_X1 port map( A => n404, Z => n496);
   U193 : BUF_X1 port map( A => n404, Z => n497);
   U194 : BUF_X1 port map( A => n404, Z => n498);
   U195 : BUF_X1 port map( A => n405, Z => n499);
   U196 : BUF_X1 port map( A => n405, Z => n500);
   U197 : BUF_X1 port map( A => n405, Z => n501);
   U198 : BUF_X1 port map( A => n406, Z => n502);
   U199 : BUF_X1 port map( A => n406, Z => n503);
   U200 : BUF_X1 port map( A => n406, Z => n504);
   U201 : BUF_X1 port map( A => n407, Z => n505);
   U202 : BUF_X1 port map( A => n407, Z => n506);
   U203 : BUF_X1 port map( A => n48, Z => n257);
   U204 : BUF_X1 port map( A => n48, Z => n258);
   U205 : BUF_X1 port map( A => n1438, Z => n134);
   U206 : BUF_X1 port map( A => n1438, Z => n135);
   U207 : BUF_X1 port map( A => n62, Z => n71);
   U208 : BUF_X1 port map( A => n62, Z => n72);
   U209 : BUF_X1 port map( A => n2370, Z => n344);
   U210 : BUF_X1 port map( A => n2370, Z => n345);
   U211 : BUF_X1 port map( A => n2365, Z => n332);
   U212 : BUF_X1 port map( A => n2365, Z => n333);
   U213 : BUF_X1 port map( A => n56, Z => n119);
   U214 : BUF_X1 port map( A => n56, Z => n120);
   U215 : BUF_X1 port map( A => n59, Z => n176);
   U216 : BUF_X1 port map( A => n59, Z => n177);
   U217 : BUF_X1 port map( A => n58, Z => n167);
   U218 : BUF_X1 port map( A => n58, Z => n168);
   U219 : BUF_X1 port map( A => n2381, Z => n368);
   U220 : BUF_X1 port map( A => n2381, Z => n369);
   U221 : BUF_X1 port map( A => n2373, Z => n350);
   U222 : BUF_X1 port map( A => n2368, Z => n338);
   U223 : BUF_X1 port map( A => n2373, Z => n351);
   U224 : BUF_X1 port map( A => n2368, Z => n339);
   U225 : BUF_X1 port map( A => n2377, Z => n359);
   U226 : BUF_X1 port map( A => n2377, Z => n360);
   U227 : BUF_X1 port map( A => n2380, Z => n365);
   U228 : BUF_X1 port map( A => n2380, Z => n366);
   U229 : BUF_X1 port map( A => n2372, Z => n347);
   U230 : BUF_X1 port map( A => n2367, Z => n335);
   U231 : BUF_X1 port map( A => n2372, Z => n348);
   U232 : BUF_X1 port map( A => n2367, Z => n336);
   U233 : BUF_X1 port map( A => n2376, Z => n356);
   U234 : BUF_X1 port map( A => n2376, Z => n357);
   U235 : BUF_X1 port map( A => n922, Z => n92);
   U236 : BUF_X1 port map( A => n917, Z => n77);
   U237 : BUF_X1 port map( A => n922, Z => n93);
   U238 : BUF_X1 port map( A => n917, Z => n78);
   U239 : BUF_X1 port map( A => n1443, Z => n149);
   U240 : BUF_X1 port map( A => n1443, Z => n150);
   U241 : BUF_X1 port map( A => n2364, Z => n329);
   U242 : BUF_X1 port map( A => n2364, Z => n330);
   U243 : BUF_X1 port map( A => n2369, Z => n341);
   U244 : BUF_X1 port map( A => n2369, Z => n342);
   U245 : BUF_X1 port map( A => n2374, Z => n353);
   U246 : BUF_X1 port map( A => n2374, Z => n354);
   U247 : BUF_X1 port map( A => n55, Z => n110);
   U248 : BUF_X1 port map( A => n54, Z => n98);
   U249 : BUF_X1 port map( A => n55, Z => n111);
   U250 : BUF_X1 port map( A => n54, Z => n99);
   U251 : BUF_X1 port map( A => n57, Z => n155);
   U252 : BUF_X1 port map( A => n57, Z => n156);
   U253 : BUF_X1 port map( A => n64, Z => n68);
   U254 : BUF_X1 port map( A => n64, Z => n69);
   U255 : BUF_X1 port map( A => n48, Z => n259);
   U256 : BUF_X1 port map( A => n1438, Z => n136);
   U257 : BUF_X1 port map( A => n62, Z => n73);
   U258 : BUF_X1 port map( A => n2370, Z => n346);
   U259 : BUF_X1 port map( A => n2365, Z => n334);
   U260 : BUF_X1 port map( A => n56, Z => n121);
   U261 : BUF_X1 port map( A => n59, Z => n178);
   U262 : BUF_X1 port map( A => n58, Z => n169);
   U263 : BUF_X1 port map( A => n2381, Z => n370);
   U264 : BUF_X1 port map( A => n2377, Z => n361);
   U265 : BUF_X1 port map( A => n2373, Z => n352);
   U266 : BUF_X1 port map( A => n2368, Z => n340);
   U267 : BUF_X1 port map( A => n2380, Z => n367);
   U268 : BUF_X1 port map( A => n2376, Z => n358);
   U269 : BUF_X1 port map( A => n2372, Z => n349);
   U270 : BUF_X1 port map( A => n2367, Z => n337);
   U271 : BUF_X1 port map( A => n922, Z => n94);
   U272 : BUF_X1 port map( A => n917, Z => n79);
   U273 : BUF_X1 port map( A => n1443, Z => n151);
   U274 : BUF_X1 port map( A => n2364, Z => n331);
   U275 : BUF_X1 port map( A => n2369, Z => n343);
   U276 : BUF_X1 port map( A => n2374, Z => n355);
   U277 : BUF_X1 port map( A => n55, Z => n112);
   U278 : BUF_X1 port map( A => n54, Z => n100);
   U279 : BUF_X1 port map( A => n57, Z => n157);
   U280 : BUF_X1 port map( A => n64, Z => n70);
   U281 : BUF_X1 port map( A => n920, Z => n83);
   U282 : BUF_X1 port map( A => n1441, Z => n140);
   U283 : BUF_X1 port map( A => n920, Z => n84);
   U284 : BUF_X1 port map( A => n1441, Z => n141);
   U285 : BUF_X1 port map( A => n408, Z => n405);
   U286 : BUF_X1 port map( A => n408, Z => n406);
   U287 : BUF_X1 port map( A => n409, Z => n403);
   U288 : BUF_X1 port map( A => n409, Z => n404);
   U289 : BUF_X1 port map( A => n408, Z => n407);
   U290 : BUF_X1 port map( A => n13, Z => n182);
   U291 : BUF_X1 port map( A => n13, Z => n183);
   U292 : BUF_X1 port map( A => n14, Z => n185);
   U293 : BUF_X1 port map( A => n14, Z => n186);
   U294 : BUF_X1 port map( A => n15, Z => n188);
   U295 : BUF_X1 port map( A => n15, Z => n189);
   U296 : BUF_X1 port map( A => n16, Z => n191);
   U297 : BUF_X1 port map( A => n16, Z => n192);
   U298 : BUF_X1 port map( A => n17, Z => n194);
   U299 : BUF_X1 port map( A => n17, Z => n195);
   U300 : BUF_X1 port map( A => n18, Z => n197);
   U301 : BUF_X1 port map( A => n18, Z => n198);
   U302 : BUF_X1 port map( A => n19, Z => n200);
   U303 : BUF_X1 port map( A => n19, Z => n201);
   U304 : BUF_X1 port map( A => n20, Z => n203);
   U305 : BUF_X1 port map( A => n20, Z => n204);
   U306 : BUF_X1 port map( A => n21, Z => n206);
   U307 : BUF_X1 port map( A => n21, Z => n207);
   U308 : BUF_X1 port map( A => n22, Z => n209);
   U309 : BUF_X1 port map( A => n22, Z => n210);
   U310 : BUF_X1 port map( A => n23, Z => n212);
   U311 : BUF_X1 port map( A => n23, Z => n213);
   U312 : BUF_X1 port map( A => n24, Z => n215);
   U313 : BUF_X1 port map( A => n24, Z => n216);
   U314 : BUF_X1 port map( A => n25, Z => n218);
   U315 : BUF_X1 port map( A => n25, Z => n219);
   U316 : BUF_X1 port map( A => n26, Z => n221);
   U317 : BUF_X1 port map( A => n26, Z => n222);
   U318 : BUF_X1 port map( A => n27, Z => n224);
   U319 : BUF_X1 port map( A => n27, Z => n225);
   U320 : BUF_X1 port map( A => n28, Z => n227);
   U321 : BUF_X1 port map( A => n28, Z => n228);
   U322 : BUF_X1 port map( A => n29, Z => n230);
   U323 : BUF_X1 port map( A => n29, Z => n231);
   U324 : BUF_X1 port map( A => n30, Z => n233);
   U325 : BUF_X1 port map( A => n30, Z => n234);
   U326 : BUF_X1 port map( A => n31, Z => n236);
   U327 : BUF_X1 port map( A => n31, Z => n237);
   U328 : BUF_X1 port map( A => n32, Z => n239);
   U329 : BUF_X1 port map( A => n32, Z => n240);
   U330 : BUF_X1 port map( A => n33, Z => n242);
   U331 : BUF_X1 port map( A => n33, Z => n243);
   U332 : BUF_X1 port map( A => n34, Z => n245);
   U333 : BUF_X1 port map( A => n34, Z => n246);
   U334 : BUF_X1 port map( A => n35, Z => n248);
   U335 : BUF_X1 port map( A => n35, Z => n249);
   U336 : BUF_X1 port map( A => n36, Z => n251);
   U337 : BUF_X1 port map( A => n36, Z => n252);
   U338 : BUF_X1 port map( A => n47, Z => n254);
   U339 : BUF_X1 port map( A => n47, Z => n255);
   U340 : BUF_X1 port map( A => n49, Z => n260);
   U341 : BUF_X1 port map( A => n49, Z => n261);
   U342 : BUF_X1 port map( A => n50, Z => n263);
   U343 : BUF_X1 port map( A => n50, Z => n264);
   U344 : BUF_X1 port map( A => n51, Z => n266);
   U345 : BUF_X1 port map( A => n51, Z => n267);
   U346 : BUF_X1 port map( A => n52, Z => n269);
   U347 : BUF_X1 port map( A => n52, Z => n270);
   U348 : BUF_X1 port map( A => n53, Z => n272);
   U349 : BUF_X1 port map( A => n53, Z => n273);
   U350 : BUF_X1 port map( A => n1448, Z => n170);
   U351 : BUF_X1 port map( A => n1448, Z => n171);
   U352 : BUF_X1 port map( A => n927, Z => n113);
   U353 : BUF_X1 port map( A => n927, Z => n114);
   U354 : BUF_X1 port map( A => n13, Z => n184);
   U355 : BUF_X1 port map( A => n14, Z => n187);
   U356 : BUF_X1 port map( A => n15, Z => n190);
   U357 : BUF_X1 port map( A => n16, Z => n193);
   U358 : BUF_X1 port map( A => n17, Z => n196);
   U359 : BUF_X1 port map( A => n18, Z => n199);
   U360 : BUF_X1 port map( A => n19, Z => n202);
   U361 : BUF_X1 port map( A => n20, Z => n205);
   U362 : BUF_X1 port map( A => n21, Z => n208);
   U363 : BUF_X1 port map( A => n22, Z => n211);
   U364 : BUF_X1 port map( A => n23, Z => n214);
   U365 : BUF_X1 port map( A => n24, Z => n217);
   U366 : BUF_X1 port map( A => n25, Z => n220);
   U367 : BUF_X1 port map( A => n26, Z => n223);
   U368 : BUF_X1 port map( A => n27, Z => n226);
   U369 : BUF_X1 port map( A => n28, Z => n229);
   U370 : BUF_X1 port map( A => n29, Z => n232);
   U371 : BUF_X1 port map( A => n30, Z => n235);
   U372 : BUF_X1 port map( A => n31, Z => n238);
   U373 : BUF_X1 port map( A => n32, Z => n241);
   U374 : BUF_X1 port map( A => n33, Z => n244);
   U375 : BUF_X1 port map( A => n34, Z => n247);
   U376 : BUF_X1 port map( A => n35, Z => n250);
   U377 : BUF_X1 port map( A => n36, Z => n253);
   U378 : BUF_X1 port map( A => n47, Z => n256);
   U379 : BUF_X1 port map( A => n49, Z => n262);
   U380 : BUF_X1 port map( A => n50, Z => n265);
   U381 : BUF_X1 port map( A => n51, Z => n268);
   U382 : BUF_X1 port map( A => n52, Z => n271);
   U383 : BUF_X1 port map( A => n53, Z => n274);
   U384 : BUF_X1 port map( A => n1448, Z => n172);
   U385 : BUF_X1 port map( A => n927, Z => n115);
   U386 : BUF_X1 port map( A => RST, Z => n408);
   U387 : BUF_X1 port map( A => RST, Z => n409);
   U388 : BUF_X1 port map( A => n60, Z => n116);
   U389 : BUF_X1 port map( A => n61, Z => n173);
   U390 : BUF_X1 port map( A => n60, Z => n117);
   U391 : BUF_X1 port map( A => n61, Z => n174);
   U392 : BUF_X1 port map( A => n60, Z => n118);
   U393 : BUF_X1 port map( A => n61, Z => n175);
   U394 : INV_X1 port map( A => DATAIN(0), ZN => n371);
   U395 : INV_X1 port map( A => DATAIN(1), ZN => n372);
   U396 : INV_X1 port map( A => DATAIN(2), ZN => n373);
   U397 : INV_X1 port map( A => DATAIN(3), ZN => n374);
   U398 : INV_X1 port map( A => DATAIN(4), ZN => n375);
   U399 : INV_X1 port map( A => DATAIN(5), ZN => n376);
   U400 : INV_X1 port map( A => DATAIN(6), ZN => n377);
   U401 : INV_X1 port map( A => DATAIN(7), ZN => n378);
   U402 : INV_X1 port map( A => DATAIN(8), ZN => n379);
   U403 : INV_X1 port map( A => DATAIN(10), ZN => n381);
   U404 : INV_X1 port map( A => DATAIN(11), ZN => n382);
   U405 : INV_X1 port map( A => DATAIN(12), ZN => n383);
   U406 : INV_X1 port map( A => DATAIN(13), ZN => n384);
   U407 : INV_X1 port map( A => DATAIN(14), ZN => n385);
   U408 : INV_X1 port map( A => DATAIN(15), ZN => n386);
   U409 : INV_X1 port map( A => DATAIN(16), ZN => n387);
   U410 : INV_X1 port map( A => DATAIN(17), ZN => n388);
   U411 : INV_X1 port map( A => DATAIN(18), ZN => n389);
   U412 : INV_X1 port map( A => DATAIN(19), ZN => n390);
   U413 : INV_X1 port map( A => DATAIN(20), ZN => n391);
   U414 : INV_X1 port map( A => DATAIN(21), ZN => n392);
   U415 : INV_X1 port map( A => DATAIN(22), ZN => n393);
   U416 : INV_X1 port map( A => DATAIN(23), ZN => n394);
   U417 : INV_X1 port map( A => DATAIN(24), ZN => n395);
   U418 : INV_X1 port map( A => DATAIN(25), ZN => n396);
   U419 : INV_X1 port map( A => DATAIN(26), ZN => n397);
   U420 : INV_X1 port map( A => DATAIN(27), ZN => n398);
   U421 : INV_X1 port map( A => DATAIN(28), ZN => n399);
   U422 : INV_X1 port map( A => DATAIN(29), ZN => n400);
   U423 : INV_X1 port map( A => DATAIN(30), ZN => n401);
   U424 : INV_X1 port map( A => DATAIN(31), ZN => n402);
   U425 : INV_X1 port map( A => DATAIN(9), ZN => n380);
   U426 : CLKBUF_X1 port map( A => n506, Z => n410);
   U427 : CLKBUF_X1 port map( A => n506, Z => n411);
   U428 : CLKBUF_X1 port map( A => n506, Z => n412);
   U429 : CLKBUF_X1 port map( A => n506, Z => n413);
   U430 : CLKBUF_X1 port map( A => n506, Z => n414);
   U431 : CLKBUF_X1 port map( A => n505, Z => n415);
   U432 : CLKBUF_X1 port map( A => n505, Z => n416);
   U433 : CLKBUF_X1 port map( A => n505, Z => n417);
   U434 : CLKBUF_X1 port map( A => n505, Z => n418);
   U435 : CLKBUF_X1 port map( A => n505, Z => n419);
   U436 : CLKBUF_X1 port map( A => n505, Z => n420);
   U437 : CLKBUF_X1 port map( A => n504, Z => n421);
   U438 : CLKBUF_X1 port map( A => n504, Z => n422);
   U439 : CLKBUF_X1 port map( A => n504, Z => n423);
   U440 : CLKBUF_X1 port map( A => n504, Z => n424);
   U441 : CLKBUF_X1 port map( A => n504, Z => n425);
   U442 : CLKBUF_X1 port map( A => n504, Z => n426);
   U443 : CLKBUF_X1 port map( A => n503, Z => n427);
   U444 : CLKBUF_X1 port map( A => n503, Z => n428);
   U445 : CLKBUF_X1 port map( A => n503, Z => n429);
   U446 : CLKBUF_X1 port map( A => n503, Z => n430);
   U447 : CLKBUF_X1 port map( A => n503, Z => n431);
   U448 : CLKBUF_X1 port map( A => n503, Z => n432);
   U449 : CLKBUF_X1 port map( A => n502, Z => n433);
   U450 : CLKBUF_X1 port map( A => n502, Z => n434);
   U451 : CLKBUF_X1 port map( A => n502, Z => n435);
   U452 : CLKBUF_X1 port map( A => n502, Z => n436);
   U453 : CLKBUF_X1 port map( A => n502, Z => n437);
   U454 : CLKBUF_X1 port map( A => n502, Z => n438);
   U455 : CLKBUF_X1 port map( A => n501, Z => n439);
   U456 : CLKBUF_X1 port map( A => n501, Z => n440);
   U457 : CLKBUF_X1 port map( A => n501, Z => n441);
   U458 : CLKBUF_X1 port map( A => n501, Z => n442);
   U459 : CLKBUF_X1 port map( A => n501, Z => n443);
   U460 : CLKBUF_X1 port map( A => n501, Z => n444);
   U461 : CLKBUF_X1 port map( A => n500, Z => n445);
   U462 : CLKBUF_X1 port map( A => n500, Z => n446);
   U463 : CLKBUF_X1 port map( A => n500, Z => n447);
   U464 : CLKBUF_X1 port map( A => n500, Z => n448);
   U465 : CLKBUF_X1 port map( A => n500, Z => n449);
   U466 : CLKBUF_X1 port map( A => n500, Z => n450);
   U467 : CLKBUF_X1 port map( A => n499, Z => n451);
   U468 : CLKBUF_X1 port map( A => n499, Z => n452);
   U469 : CLKBUF_X1 port map( A => n499, Z => n453);
   U470 : CLKBUF_X1 port map( A => n499, Z => n454);
   U471 : CLKBUF_X1 port map( A => n499, Z => n455);
   U472 : CLKBUF_X1 port map( A => n499, Z => n456);
   U473 : CLKBUF_X1 port map( A => n498, Z => n457);
   U474 : CLKBUF_X1 port map( A => n498, Z => n458);
   U475 : CLKBUF_X1 port map( A => n498, Z => n459);
   U476 : CLKBUF_X1 port map( A => n498, Z => n460);
   U477 : CLKBUF_X1 port map( A => n498, Z => n461);
   U478 : CLKBUF_X1 port map( A => n498, Z => n462);
   U479 : CLKBUF_X1 port map( A => n497, Z => n463);
   U480 : CLKBUF_X1 port map( A => n497, Z => n464);
   U481 : CLKBUF_X1 port map( A => n497, Z => n465);
   U482 : CLKBUF_X1 port map( A => n497, Z => n466);
   U483 : CLKBUF_X1 port map( A => n497, Z => n467);
   U484 : CLKBUF_X1 port map( A => n497, Z => n468);
   U485 : CLKBUF_X1 port map( A => n496, Z => n469);
   U486 : CLKBUF_X1 port map( A => n496, Z => n470);
   U487 : CLKBUF_X1 port map( A => n496, Z => n471);
   U488 : CLKBUF_X1 port map( A => n496, Z => n472);
   U489 : CLKBUF_X1 port map( A => n496, Z => n473);
   U490 : CLKBUF_X1 port map( A => n496, Z => n474);
   U491 : CLKBUF_X1 port map( A => n495, Z => n475);
   U492 : CLKBUF_X1 port map( A => n495, Z => n476);
   U493 : CLKBUF_X1 port map( A => n495, Z => n477);
   U494 : CLKBUF_X1 port map( A => n495, Z => n478);
   U495 : CLKBUF_X1 port map( A => n495, Z => n479);
   U496 : CLKBUF_X1 port map( A => n495, Z => n480);
   U497 : CLKBUF_X1 port map( A => n494, Z => n481);
   U498 : CLKBUF_X1 port map( A => n494, Z => n482);
   U499 : CLKBUF_X1 port map( A => n494, Z => n483);
   U500 : CLKBUF_X1 port map( A => n494, Z => n484);
   U501 : CLKBUF_X1 port map( A => n494, Z => n485);
   U502 : CLKBUF_X1 port map( A => n494, Z => n486);
   U503 : CLKBUF_X1 port map( A => n493, Z => n487);
   U504 : CLKBUF_X1 port map( A => n493, Z => n488);
   U505 : CLKBUF_X1 port map( A => n493, Z => n489);
   U506 : CLKBUF_X1 port map( A => n493, Z => n490);
   U507 : CLKBUF_X1 port map( A => n493, Z => n491);
   U508 : INV_X1 port map( A => ADD_WR(0), ZN => n1907);
   U509 : NAND3_X1 port map( A1 => n2619, A2 => n2618, A3 => n66, ZN => n507);
   U510 : NAND2_X1 port map( A1 => n116, A2 => n507, ZN => n516);
   U511 : INV_X1 port map( A => n516, ZN => n920);
   U512 : OAI211_X1 port map( C1 => n3952, C2 => n68, A => n2605, B => n2604, 
                           ZN => n508);
   U513 : AOI221_X1 port map( B1 => n353, B2 => n1843, C1 => n362, C2 => n4030,
                           A => n508, ZN => n511);
   U514 : NOR2_X1 port map( A1 => n4125, A2 => n71, ZN => n509);
   U515 : NOR4_X1 port map( A1 => n2615, A2 => n2610, A3 => n2601, A4 => n509, 
                           ZN => n510);
   U516 : NAND2_X1 port map( A1 => n511, A2 => n510, ZN => n513);
   U517 : OR2_X1 port map( A1 => n2347, A2 => n516, ZN => n917);
   U518 : NAND2_X1 port map( A1 => n2348, A2 => n85, ZN => n916);
   U519 : OAI22_X1 port map( A1 => n939, A2 => n77, B1 => n938, B2 => n74, ZN 
                           => n512);
   U520 : AOI221_X1 port map( B1 => n85, B2 => n513, C1 => n80, C2 => n1519, A 
                           => n512, ZN => n521);
   U521 : OR2_X1 port map( A1 => n2351, A2 => n516, ZN => n922);
   U522 : NAND2_X1 port map( A1 => n2352, A2 => n85, ZN => n921);
   U523 : OAI22_X1 port map( A1 => n3998, A2 => n92, B1 => n3966, B2 => n89, ZN
                           => n514);
   U524 : AOI221_X1 port map( B1 => n98, B2 => n1487, C1 => n95, C2 => n3957, A
                           => n514, ZN => n520);
   U525 : NAND2_X1 port map( A1 => n2361, A2 => n85, ZN => n925);
   U526 : NAND2_X1 port map( A1 => n2355, A2 => n85, ZN => n924);
   U527 : OAI22_X1 port map( A1 => n3963, A2 => n104, B1 => n3960, B2 => n101, 
                           ZN => n515);
   U528 : AOI221_X1 port map( B1 => n110, B2 => n4062, C1 => n107, C2 => n3964,
                           A => n515, ZN => n519);
   U529 : NAND4_X1 port map( A1 => n66, A2 => n2618, A3 => n116, A4 => n2619, 
                           ZN => n927);
   U530 : OAI22_X1 port map( A1 => n2622, A2 => n116, B1 => n371, B2 => n113, 
                           ZN => n517);
   U531 : AOI221_X1 port map( B1 => n122, B2 => n3965, C1 => n119, C2 => n1617,
                           A => n517, ZN => n518);
   U532 : NAND4_X1 port map( A1 => n521, A2 => n520, A3 => n519, A4 => n518, ZN
                           => n2983);
   U533 : OAI211_X1 port map( C1 => n3929, C2 => n68, A => n2587, B => n2586, 
                           ZN => n522);
   U534 : AOI221_X1 port map( B1 => n353, B2 => n1844, C1 => n362, C2 => n4031,
                           A => n522, ZN => n525);
   U535 : NOR2_X1 port map( A1 => n4124, A2 => n71, ZN => n523);
   U536 : NOR4_X1 port map( A1 => n2591, A2 => n2590, A3 => n2585, A4 => n523, 
                           ZN => n524);
   U537 : NAND2_X1 port map( A1 => n525, A2 => n524, ZN => n527);
   U538 : OAI22_X1 port map( A1 => n956, A2 => n77, B1 => n955, B2 => n74, ZN 
                           => n526);
   U539 : AOI221_X1 port map( B1 => n88, B2 => n527, C1 => n80, C2 => n1520, A 
                           => n526, ZN => n534);
   U540 : OAI22_X1 port map( A1 => n3999, A2 => n92, B1 => n3967, B2 => n89, ZN
                           => n528);
   U541 : AOI221_X1 port map( B1 => n98, B2 => n1488, C1 => n95, C2 => n3934, A
                           => n528, ZN => n533);
   U542 : OAI22_X1 port map( A1 => n3940, A2 => n104, B1 => n3937, B2 => n101, 
                           ZN => n529);
   U543 : AOI221_X1 port map( B1 => n110, B2 => n4063, C1 => n107, C2 => n3941,
                           A => n529, ZN => n532);
   U544 : OAI22_X1 port map( A1 => n2623, A2 => n118, B1 => n372, B2 => n113, 
                           ZN => n530);
   U545 : AOI221_X1 port map( B1 => n122, B2 => n3942, C1 => n119, C2 => n1618,
                           A => n530, ZN => n531);
   U546 : NAND4_X1 port map( A1 => n534, A2 => n533, A3 => n532, A4 => n531, ZN
                           => n2984);
   U547 : OAI211_X1 port map( C1 => n3906, C2 => n68, A => n2580, B => n2579, 
                           ZN => n535);
   U548 : AOI221_X1 port map( B1 => n353, B2 => n1845, C1 => n362, C2 => n4032,
                           A => n535, ZN => n538);
   U549 : NOR2_X1 port map( A1 => n4123, A2 => n71, ZN => n536);
   U550 : NOR4_X1 port map( A1 => n2584, A2 => n2583, A3 => n2578, A4 => n536, 
                           ZN => n537);
   U551 : NAND2_X1 port map( A1 => n538, A2 => n537, ZN => n540);
   U552 : OAI22_X1 port map( A1 => n972, A2 => n77, B1 => n971, B2 => n74, ZN 
                           => n539);
   U553 : AOI221_X1 port map( B1 => n88, B2 => n540, C1 => n80, C2 => n1521, A 
                           => n539, ZN => n547);
   U554 : OAI22_X1 port map( A1 => n4000, A2 => n92, B1 => n3968, B2 => n89, ZN
                           => n541);
   U555 : AOI221_X1 port map( B1 => n98, B2 => n1489, C1 => n95, C2 => n3911, A
                           => n541, ZN => n546);
   U556 : OAI22_X1 port map( A1 => n3917, A2 => n104, B1 => n3914, B2 => n101, 
                           ZN => n542);
   U557 : AOI221_X1 port map( B1 => n110, B2 => n4064, C1 => n107, C2 => n3918,
                           A => n542, ZN => n545);
   U558 : OAI22_X1 port map( A1 => n2624, A2 => n118, B1 => n373, B2 => n113, 
                           ZN => n543);
   U559 : AOI221_X1 port map( B1 => n122, B2 => n3919, C1 => n119, C2 => n1619,
                           A => n543, ZN => n544);
   U560 : NAND4_X1 port map( A1 => n547, A2 => n546, A3 => n545, A4 => n544, ZN
                           => n2985);
   U561 : OAI211_X1 port map( C1 => n3883, C2 => n68, A => n2573, B => n2572, 
                           ZN => n548);
   U562 : AOI221_X1 port map( B1 => n353, B2 => n1846, C1 => n362, C2 => n4033,
                           A => n548, ZN => n551);
   U563 : NOR2_X1 port map( A1 => n4122, A2 => n71, ZN => n549);
   U564 : NOR4_X1 port map( A1 => n2577, A2 => n2576, A3 => n2571, A4 => n549, 
                           ZN => n550);
   U565 : NAND2_X1 port map( A1 => n551, A2 => n550, ZN => n553);
   U566 : OAI22_X1 port map( A1 => n988, A2 => n77, B1 => n987, B2 => n74, ZN 
                           => n552);
   U567 : AOI221_X1 port map( B1 => n88, B2 => n553, C1 => n80, C2 => n1522, A 
                           => n552, ZN => n560);
   U568 : OAI22_X1 port map( A1 => n4001, A2 => n92, B1 => n3969, B2 => n89, ZN
                           => n554);
   U569 : AOI221_X1 port map( B1 => n98, B2 => n1490, C1 => n95, C2 => n3888, A
                           => n554, ZN => n559);
   U570 : OAI22_X1 port map( A1 => n3894, A2 => n104, B1 => n3891, B2 => n101, 
                           ZN => n555);
   U571 : AOI221_X1 port map( B1 => n110, B2 => n4065, C1 => n107, C2 => n3895,
                           A => n555, ZN => n558);
   U572 : OAI22_X1 port map( A1 => n2625, A2 => n118, B1 => n374, B2 => n113, 
                           ZN => n556);
   U573 : AOI221_X1 port map( B1 => n122, B2 => n3896, C1 => n119, C2 => n1620,
                           A => n556, ZN => n557);
   U574 : NAND4_X1 port map( A1 => n560, A2 => n559, A3 => n558, A4 => n557, ZN
                           => n2986);
   U575 : OAI211_X1 port map( C1 => n3860, C2 => n68, A => n2566, B => n2565, 
                           ZN => n561);
   U576 : AOI221_X1 port map( B1 => n353, B2 => n1847, C1 => n362, C2 => n4034,
                           A => n561, ZN => n564);
   U577 : NOR2_X1 port map( A1 => n4121, A2 => n71, ZN => n562);
   U578 : NOR4_X1 port map( A1 => n2570, A2 => n2569, A3 => n2564, A4 => n562, 
                           ZN => n563);
   U579 : NAND2_X1 port map( A1 => n564, A2 => n563, ZN => n566);
   U580 : OAI22_X1 port map( A1 => n1004, A2 => n77, B1 => n1003, B2 => n74, ZN
                           => n565);
   U581 : AOI221_X1 port map( B1 => n88, B2 => n566, C1 => n80, C2 => n1523, A 
                           => n565, ZN => n573);
   U582 : OAI22_X1 port map( A1 => n4002, A2 => n92, B1 => n3970, B2 => n89, ZN
                           => n567);
   U583 : AOI221_X1 port map( B1 => n98, B2 => n1491, C1 => n95, C2 => n3865, A
                           => n567, ZN => n572);
   U584 : OAI22_X1 port map( A1 => n3871, A2 => n104, B1 => n3868, B2 => n101, 
                           ZN => n568);
   U585 : AOI221_X1 port map( B1 => n110, B2 => n4066, C1 => n107, C2 => n3872,
                           A => n568, ZN => n571);
   U586 : OAI22_X1 port map( A1 => n2626, A2 => n118, B1 => n375, B2 => n113, 
                           ZN => n569);
   U587 : AOI221_X1 port map( B1 => n122, B2 => n3873, C1 => n119, C2 => n1621,
                           A => n569, ZN => n570);
   U588 : NAND4_X1 port map( A1 => n573, A2 => n572, A3 => n571, A4 => n570, ZN
                           => n2987);
   U589 : OAI211_X1 port map( C1 => n3837, C2 => n68, A => n2559, B => n2558, 
                           ZN => n574);
   U590 : AOI221_X1 port map( B1 => n353, B2 => n1848, C1 => n362, C2 => n4035,
                           A => n574, ZN => n577);
   U591 : NOR2_X1 port map( A1 => n4120, A2 => n71, ZN => n575);
   U592 : NOR4_X1 port map( A1 => n2563, A2 => n2562, A3 => n2557, A4 => n575, 
                           ZN => n576);
   U593 : NAND2_X1 port map( A1 => n577, A2 => n576, ZN => n579);
   U594 : OAI22_X1 port map( A1 => n1020, A2 => n77, B1 => n1019, B2 => n74, ZN
                           => n578);
   U595 : AOI221_X1 port map( B1 => n87, B2 => n579, C1 => n80, C2 => n1524, A 
                           => n578, ZN => n586);
   U596 : OAI22_X1 port map( A1 => n4003, A2 => n92, B1 => n3971, B2 => n89, ZN
                           => n580);
   U597 : AOI221_X1 port map( B1 => n98, B2 => n1492, C1 => n95, C2 => n3842, A
                           => n580, ZN => n585);
   U598 : OAI22_X1 port map( A1 => n3848, A2 => n104, B1 => n3845, B2 => n101, 
                           ZN => n581);
   U599 : AOI221_X1 port map( B1 => n110, B2 => n4067, C1 => n107, C2 => n3849,
                           A => n581, ZN => n584);
   U600 : OAI22_X1 port map( A1 => n2627, A2 => n118, B1 => n376, B2 => n113, 
                           ZN => n582);
   U601 : AOI221_X1 port map( B1 => n122, B2 => n3850, C1 => n119, C2 => n1622,
                           A => n582, ZN => n583);
   U602 : NAND4_X1 port map( A1 => n586, A2 => n585, A3 => n584, A4 => n583, ZN
                           => n2988);
   U603 : OAI211_X1 port map( C1 => n3814, C2 => n68, A => n2552, B => n2551, 
                           ZN => n587);
   U604 : AOI221_X1 port map( B1 => n353, B2 => n1849, C1 => n362, C2 => n4036,
                           A => n587, ZN => n590);
   U605 : NOR2_X1 port map( A1 => n4119, A2 => n71, ZN => n588);
   U606 : NOR4_X1 port map( A1 => n2556, A2 => n2555, A3 => n2550, A4 => n588, 
                           ZN => n589);
   U607 : NAND2_X1 port map( A1 => n590, A2 => n589, ZN => n592);
   U608 : OAI22_X1 port map( A1 => n1036, A2 => n77, B1 => n1035, B2 => n74, ZN
                           => n591);
   U609 : AOI221_X1 port map( B1 => n87, B2 => n592, C1 => n80, C2 => n1525, A 
                           => n591, ZN => n599);
   U610 : OAI22_X1 port map( A1 => n4004, A2 => n92, B1 => n3972, B2 => n89, ZN
                           => n593);
   U611 : AOI221_X1 port map( B1 => n98, B2 => n1493, C1 => n95, C2 => n3819, A
                           => n593, ZN => n598);
   U612 : OAI22_X1 port map( A1 => n3825, A2 => n104, B1 => n3822, B2 => n101, 
                           ZN => n594);
   U613 : AOI221_X1 port map( B1 => n110, B2 => n4068, C1 => n107, C2 => n3826,
                           A => n594, ZN => n597);
   U614 : OAI22_X1 port map( A1 => n2628, A2 => n118, B1 => n377, B2 => n113, 
                           ZN => n595);
   U615 : AOI221_X1 port map( B1 => n122, B2 => n3827, C1 => n119, C2 => n1623,
                           A => n595, ZN => n596);
   U616 : NAND4_X1 port map( A1 => n599, A2 => n598, A3 => n597, A4 => n596, ZN
                           => n2989);
   U617 : OAI211_X1 port map( C1 => n3791, C2 => n68, A => n2545, B => n2544, 
                           ZN => n600);
   U618 : AOI221_X1 port map( B1 => n353, B2 => n1850, C1 => n362, C2 => n4037,
                           A => n600, ZN => n603);
   U619 : NOR2_X1 port map( A1 => n4118, A2 => n71, ZN => n601);
   U620 : NOR4_X1 port map( A1 => n2549, A2 => n2548, A3 => n2543, A4 => n601, 
                           ZN => n602);
   U621 : NAND2_X1 port map( A1 => n603, A2 => n602, ZN => n605);
   U622 : OAI22_X1 port map( A1 => n1052, A2 => n77, B1 => n1051, B2 => n74, ZN
                           => n604);
   U623 : AOI221_X1 port map( B1 => n87, B2 => n605, C1 => n80, C2 => n1526, A 
                           => n604, ZN => n612);
   U624 : OAI22_X1 port map( A1 => n4005, A2 => n92, B1 => n3973, B2 => n89, ZN
                           => n606);
   U625 : AOI221_X1 port map( B1 => n98, B2 => n1494, C1 => n95, C2 => n3796, A
                           => n606, ZN => n611);
   U626 : OAI22_X1 port map( A1 => n3802, A2 => n104, B1 => n3799, B2 => n101, 
                           ZN => n607);
   U627 : AOI221_X1 port map( B1 => n110, B2 => n4069, C1 => n107, C2 => n3803,
                           A => n607, ZN => n610);
   U628 : OAI22_X1 port map( A1 => n2629, A2 => n118, B1 => n378, B2 => n113, 
                           ZN => n608);
   U629 : AOI221_X1 port map( B1 => n122, B2 => n3804, C1 => n119, C2 => n1624,
                           A => n608, ZN => n609);
   U630 : NAND4_X1 port map( A1 => n612, A2 => n611, A3 => n610, A4 => n609, ZN
                           => n2990);
   U631 : OAI211_X1 port map( C1 => n3768, C2 => n68, A => n2538, B => n2537, 
                           ZN => n613);
   U632 : AOI221_X1 port map( B1 => n353, B2 => n1851, C1 => n362, C2 => n4038,
                           A => n613, ZN => n616);
   U633 : NOR2_X1 port map( A1 => n4117, A2 => n71, ZN => n614);
   U634 : NOR4_X1 port map( A1 => n2542, A2 => n2541, A3 => n2536, A4 => n614, 
                           ZN => n615);
   U635 : NAND2_X1 port map( A1 => n616, A2 => n615, ZN => n618);
   U636 : OAI22_X1 port map( A1 => n1068, A2 => n77, B1 => n1067, B2 => n74, ZN
                           => n617);
   U637 : AOI221_X1 port map( B1 => n87, B2 => n618, C1 => n80, C2 => n1527, A 
                           => n617, ZN => n625);
   U638 : OAI22_X1 port map( A1 => n4006, A2 => n92, B1 => n3974, B2 => n89, ZN
                           => n619);
   U639 : AOI221_X1 port map( B1 => n98, B2 => n1495, C1 => n95, C2 => n3773, A
                           => n619, ZN => n624);
   U640 : OAI22_X1 port map( A1 => n3779, A2 => n104, B1 => n3776, B2 => n101, 
                           ZN => n620);
   U641 : AOI221_X1 port map( B1 => n110, B2 => n4070, C1 => n107, C2 => n3780,
                           A => n620, ZN => n623);
   U642 : OAI22_X1 port map( A1 => n2630, A2 => n118, B1 => n379, B2 => n113, 
                           ZN => n621);
   U643 : AOI221_X1 port map( B1 => n122, B2 => n3781, C1 => n119, C2 => n1625,
                           A => n621, ZN => n622);
   U644 : NAND4_X1 port map( A1 => n625, A2 => n624, A3 => n623, A4 => n622, ZN
                           => n2991);
   U645 : OAI211_X1 port map( C1 => n3745, C2 => n68, A => n2531, B => n2530, 
                           ZN => n626);
   U646 : AOI221_X1 port map( B1 => n353, B2 => n1852, C1 => n362, C2 => n4039,
                           A => n626, ZN => n629);
   U647 : NOR2_X1 port map( A1 => n4116, A2 => n71, ZN => n627);
   U648 : NOR4_X1 port map( A1 => n2535, A2 => n2534, A3 => n2529, A4 => n627, 
                           ZN => n628);
   U649 : NAND2_X1 port map( A1 => n629, A2 => n628, ZN => n631);
   U650 : OAI22_X1 port map( A1 => n1084, A2 => n77, B1 => n1083, B2 => n74, ZN
                           => n630);
   U651 : AOI221_X1 port map( B1 => n87, B2 => n631, C1 => n80, C2 => n1528, A 
                           => n630, ZN => n638);
   U652 : OAI22_X1 port map( A1 => n4007, A2 => n92, B1 => n3975, B2 => n89, ZN
                           => n632);
   U653 : AOI221_X1 port map( B1 => n98, B2 => n1496, C1 => n95, C2 => n3750, A
                           => n632, ZN => n637);
   U654 : OAI22_X1 port map( A1 => n3756, A2 => n104, B1 => n3753, B2 => n101, 
                           ZN => n633);
   U655 : AOI221_X1 port map( B1 => n110, B2 => n4071, C1 => n107, C2 => n3757,
                           A => n633, ZN => n636);
   U656 : OAI22_X1 port map( A1 => n2631, A2 => n118, B1 => n380, B2 => n113, 
                           ZN => n634);
   U657 : AOI221_X1 port map( B1 => n122, B2 => n3758, C1 => n119, C2 => n1626,
                           A => n634, ZN => n635);
   U658 : NAND4_X1 port map( A1 => n638, A2 => n637, A3 => n636, A4 => n635, ZN
                           => n2992);
   U659 : OAI211_X1 port map( C1 => n3722, C2 => n68, A => n2524, B => n2523, 
                           ZN => n639);
   U660 : AOI221_X1 port map( B1 => n353, B2 => n1853, C1 => n362, C2 => n4040,
                           A => n639, ZN => n642);
   U661 : NOR2_X1 port map( A1 => n4115, A2 => n71, ZN => n640);
   U662 : NOR4_X1 port map( A1 => n2528, A2 => n2527, A3 => n2522, A4 => n640, 
                           ZN => n641);
   U663 : NAND2_X1 port map( A1 => n642, A2 => n641, ZN => n644);
   U664 : OAI22_X1 port map( A1 => n1100, A2 => n77, B1 => n1099, B2 => n74, ZN
                           => n643);
   U665 : AOI221_X1 port map( B1 => n87, B2 => n644, C1 => n80, C2 => n1529, A 
                           => n643, ZN => n651);
   U666 : OAI22_X1 port map( A1 => n4008, A2 => n92, B1 => n3976, B2 => n89, ZN
                           => n645);
   U667 : AOI221_X1 port map( B1 => n98, B2 => n1497, C1 => n95, C2 => n3727, A
                           => n645, ZN => n650);
   U668 : OAI22_X1 port map( A1 => n3733, A2 => n104, B1 => n3730, B2 => n101, 
                           ZN => n646);
   U669 : AOI221_X1 port map( B1 => n110, B2 => n4072, C1 => n107, C2 => n3734,
                           A => n646, ZN => n649);
   U670 : OAI22_X1 port map( A1 => n2632, A2 => n118, B1 => n381, B2 => n113, 
                           ZN => n647);
   U671 : AOI221_X1 port map( B1 => n122, B2 => n3735, C1 => n119, C2 => n1627,
                           A => n647, ZN => n648);
   U672 : NAND4_X1 port map( A1 => n651, A2 => n650, A3 => n649, A4 => n648, ZN
                           => n2993);
   U673 : OAI211_X1 port map( C1 => n3699, C2 => n68, A => n2517, B => n2516, 
                           ZN => n652);
   U674 : AOI221_X1 port map( B1 => n353, B2 => n1854, C1 => n362, C2 => n4041,
                           A => n652, ZN => n655);
   U675 : NOR2_X1 port map( A1 => n4114, A2 => n71, ZN => n653);
   U676 : NOR4_X1 port map( A1 => n2521, A2 => n2520, A3 => n2515, A4 => n653, 
                           ZN => n654);
   U677 : NAND2_X1 port map( A1 => n655, A2 => n654, ZN => n657);
   U678 : OAI22_X1 port map( A1 => n1116, A2 => n77, B1 => n1115, B2 => n74, ZN
                           => n656);
   U679 : AOI221_X1 port map( B1 => n87, B2 => n657, C1 => n80, C2 => n1530, A 
                           => n656, ZN => n664);
   U680 : OAI22_X1 port map( A1 => n4009, A2 => n92, B1 => n3977, B2 => n89, ZN
                           => n658);
   U681 : AOI221_X1 port map( B1 => n98, B2 => n1498, C1 => n95, C2 => n3704, A
                           => n658, ZN => n663);
   U682 : OAI22_X1 port map( A1 => n3710, A2 => n104, B1 => n3707, B2 => n101, 
                           ZN => n659);
   U683 : AOI221_X1 port map( B1 => n110, B2 => n4073, C1 => n107, C2 => n3711,
                           A => n659, ZN => n662);
   U684 : OAI22_X1 port map( A1 => n2633, A2 => n117, B1 => n382, B2 => n113, 
                           ZN => n660);
   U685 : AOI221_X1 port map( B1 => n122, B2 => n3712, C1 => n119, C2 => n1628,
                           A => n660, ZN => n661);
   U686 : NAND4_X1 port map( A1 => n664, A2 => n663, A3 => n662, A4 => n661, ZN
                           => n2994);
   U687 : OAI211_X1 port map( C1 => n3676, C2 => n69, A => n2510, B => n2509, 
                           ZN => n665);
   U688 : AOI221_X1 port map( B1 => n354, B2 => n1855, C1 => n363, C2 => n4042,
                           A => n665, ZN => n668);
   U689 : NOR2_X1 port map( A1 => n4113, A2 => n72, ZN => n666);
   U690 : NOR4_X1 port map( A1 => n2514, A2 => n2513, A3 => n2508, A4 => n666, 
                           ZN => n667);
   U691 : NAND2_X1 port map( A1 => n668, A2 => n667, ZN => n670);
   U692 : OAI22_X1 port map( A1 => n1132, A2 => n78, B1 => n1131, B2 => n75, ZN
                           => n669);
   U693 : AOI221_X1 port map( B1 => n87, B2 => n670, C1 => n81, C2 => n1531, A 
                           => n669, ZN => n677);
   U694 : OAI22_X1 port map( A1 => n4010, A2 => n93, B1 => n3978, B2 => n90, ZN
                           => n671);
   U695 : AOI221_X1 port map( B1 => n99, B2 => n1499, C1 => n96, C2 => n3681, A
                           => n671, ZN => n676);
   U696 : OAI22_X1 port map( A1 => n3687, A2 => n105, B1 => n3684, B2 => n102, 
                           ZN => n672);
   U697 : AOI221_X1 port map( B1 => n111, B2 => n4074, C1 => n108, C2 => n3688,
                           A => n672, ZN => n675);
   U698 : OAI22_X1 port map( A1 => n2634, A2 => n117, B1 => n383, B2 => n114, 
                           ZN => n673);
   U699 : AOI221_X1 port map( B1 => n123, B2 => n3689, C1 => n120, C2 => n1629,
                           A => n673, ZN => n674);
   U700 : NAND4_X1 port map( A1 => n677, A2 => n676, A3 => n675, A4 => n674, ZN
                           => n2995);
   U701 : OAI211_X1 port map( C1 => n3653, C2 => n69, A => n2503, B => n2502, 
                           ZN => n678);
   U702 : AOI221_X1 port map( B1 => n354, B2 => n1856, C1 => n363, C2 => n4043,
                           A => n678, ZN => n681);
   U703 : NOR2_X1 port map( A1 => n4112, A2 => n72, ZN => n679);
   U704 : NOR4_X1 port map( A1 => n2507, A2 => n2506, A3 => n2501, A4 => n679, 
                           ZN => n680);
   U705 : NAND2_X1 port map( A1 => n681, A2 => n680, ZN => n683);
   U706 : OAI22_X1 port map( A1 => n1148, A2 => n78, B1 => n1147, B2 => n75, ZN
                           => n682);
   U707 : AOI221_X1 port map( B1 => n87, B2 => n683, C1 => n81, C2 => n1532, A 
                           => n682, ZN => n690);
   U708 : OAI22_X1 port map( A1 => n4011, A2 => n93, B1 => n3979, B2 => n90, ZN
                           => n684);
   U709 : AOI221_X1 port map( B1 => n99, B2 => n1500, C1 => n96, C2 => n3658, A
                           => n684, ZN => n689);
   U710 : OAI22_X1 port map( A1 => n3664, A2 => n105, B1 => n3661, B2 => n102, 
                           ZN => n685);
   U711 : AOI221_X1 port map( B1 => n111, B2 => n4075, C1 => n108, C2 => n3665,
                           A => n685, ZN => n688);
   U712 : OAI22_X1 port map( A1 => n2635, A2 => n117, B1 => n384, B2 => n114, 
                           ZN => n686);
   U713 : AOI221_X1 port map( B1 => n123, B2 => n3666, C1 => n120, C2 => n1630,
                           A => n686, ZN => n687);
   U714 : NAND4_X1 port map( A1 => n690, A2 => n689, A3 => n688, A4 => n687, ZN
                           => n2996);
   U715 : OAI211_X1 port map( C1 => n3630, C2 => n69, A => n2496, B => n2495, 
                           ZN => n691);
   U716 : AOI221_X1 port map( B1 => n354, B2 => n1857, C1 => n363, C2 => n4044,
                           A => n691, ZN => n694);
   U717 : NOR2_X1 port map( A1 => n4111, A2 => n72, ZN => n692);
   U718 : NOR4_X1 port map( A1 => n2500, A2 => n2499, A3 => n2494, A4 => n692, 
                           ZN => n693);
   U719 : NAND2_X1 port map( A1 => n694, A2 => n693, ZN => n696);
   U720 : OAI22_X1 port map( A1 => n1164, A2 => n78, B1 => n1163, B2 => n75, ZN
                           => n695);
   U721 : AOI221_X1 port map( B1 => n87, B2 => n696, C1 => n81, C2 => n1533, A 
                           => n695, ZN => n703);
   U722 : OAI22_X1 port map( A1 => n4012, A2 => n93, B1 => n3980, B2 => n90, ZN
                           => n697);
   U723 : AOI221_X1 port map( B1 => n99, B2 => n1501, C1 => n96, C2 => n3635, A
                           => n697, ZN => n702);
   U724 : OAI22_X1 port map( A1 => n3641, A2 => n105, B1 => n3638, B2 => n102, 
                           ZN => n698);
   U725 : AOI221_X1 port map( B1 => n111, B2 => n4076, C1 => n108, C2 => n3642,
                           A => n698, ZN => n701);
   U726 : OAI22_X1 port map( A1 => n2636, A2 => n117, B1 => n385, B2 => n114, 
                           ZN => n699);
   U727 : AOI221_X1 port map( B1 => n123, B2 => n3643, C1 => n120, C2 => n1631,
                           A => n699, ZN => n700);
   U728 : NAND4_X1 port map( A1 => n703, A2 => n702, A3 => n701, A4 => n700, ZN
                           => n2997);
   U729 : OAI211_X1 port map( C1 => n3607, C2 => n69, A => n2489, B => n2488, 
                           ZN => n704);
   U730 : AOI221_X1 port map( B1 => n354, B2 => n1858, C1 => n363, C2 => n4045,
                           A => n704, ZN => n707);
   U731 : NOR2_X1 port map( A1 => n4110, A2 => n72, ZN => n705);
   U732 : NOR4_X1 port map( A1 => n2493, A2 => n2492, A3 => n2487, A4 => n705, 
                           ZN => n706);
   U733 : NAND2_X1 port map( A1 => n707, A2 => n706, ZN => n709);
   U734 : OAI22_X1 port map( A1 => n1180, A2 => n78, B1 => n1179, B2 => n75, ZN
                           => n708);
   U735 : AOI221_X1 port map( B1 => n87, B2 => n709, C1 => n81, C2 => n1534, A 
                           => n708, ZN => n716);
   U736 : OAI22_X1 port map( A1 => n4013, A2 => n93, B1 => n3981, B2 => n90, ZN
                           => n710);
   U737 : AOI221_X1 port map( B1 => n99, B2 => n1502, C1 => n96, C2 => n3612, A
                           => n710, ZN => n715);
   U738 : OAI22_X1 port map( A1 => n3618, A2 => n105, B1 => n3615, B2 => n102, 
                           ZN => n711);
   U739 : AOI221_X1 port map( B1 => n111, B2 => n4077, C1 => n108, C2 => n3619,
                           A => n711, ZN => n714);
   U740 : OAI22_X1 port map( A1 => n2637, A2 => n117, B1 => n386, B2 => n114, 
                           ZN => n712);
   U741 : AOI221_X1 port map( B1 => n123, B2 => n3620, C1 => n120, C2 => n1632,
                           A => n712, ZN => n713);
   U742 : NAND4_X1 port map( A1 => n716, A2 => n715, A3 => n714, A4 => n713, ZN
                           => n2998);
   U743 : OAI211_X1 port map( C1 => n3584, C2 => n69, A => n2482, B => n2481, 
                           ZN => n717);
   U744 : AOI221_X1 port map( B1 => n354, B2 => n1859, C1 => n363, C2 => n4046,
                           A => n717, ZN => n720);
   U745 : NOR2_X1 port map( A1 => n4109, A2 => n72, ZN => n718);
   U746 : NOR4_X1 port map( A1 => n2486, A2 => n2485, A3 => n2480, A4 => n718, 
                           ZN => n719);
   U747 : NAND2_X1 port map( A1 => n720, A2 => n719, ZN => n722);
   U748 : OAI22_X1 port map( A1 => n1196, A2 => n78, B1 => n1195, B2 => n75, ZN
                           => n721);
   U749 : AOI221_X1 port map( B1 => n86, B2 => n722, C1 => n81, C2 => n1535, A 
                           => n721, ZN => n729);
   U750 : OAI22_X1 port map( A1 => n4014, A2 => n93, B1 => n3982, B2 => n90, ZN
                           => n723);
   U751 : AOI221_X1 port map( B1 => n99, B2 => n1503, C1 => n96, C2 => n3589, A
                           => n723, ZN => n728);
   U752 : OAI22_X1 port map( A1 => n3595, A2 => n105, B1 => n3592, B2 => n102, 
                           ZN => n724);
   U753 : AOI221_X1 port map( B1 => n111, B2 => n4078, C1 => n108, C2 => n3596,
                           A => n724, ZN => n727);
   U754 : OAI22_X1 port map( A1 => n2638, A2 => n117, B1 => n387, B2 => n114, 
                           ZN => n725);
   U755 : AOI221_X1 port map( B1 => n123, B2 => n3597, C1 => n120, C2 => n1633,
                           A => n725, ZN => n726);
   U756 : NAND4_X1 port map( A1 => n729, A2 => n728, A3 => n727, A4 => n726, ZN
                           => n2999);
   U757 : OAI211_X1 port map( C1 => n3561, C2 => n69, A => n2475, B => n2474, 
                           ZN => n730);
   U758 : AOI221_X1 port map( B1 => n354, B2 => n1860, C1 => n363, C2 => n4047,
                           A => n730, ZN => n733);
   U759 : NOR2_X1 port map( A1 => n4108, A2 => n72, ZN => n731);
   U760 : NOR4_X1 port map( A1 => n2479, A2 => n2478, A3 => n2473, A4 => n731, 
                           ZN => n732);
   U761 : NAND2_X1 port map( A1 => n733, A2 => n732, ZN => n735);
   U762 : OAI22_X1 port map( A1 => n1212, A2 => n78, B1 => n1211, B2 => n75, ZN
                           => n734);
   U763 : AOI221_X1 port map( B1 => n86, B2 => n735, C1 => n81, C2 => n1536, A 
                           => n734, ZN => n742);
   U764 : OAI22_X1 port map( A1 => n4015, A2 => n93, B1 => n3983, B2 => n90, ZN
                           => n736);
   U765 : AOI221_X1 port map( B1 => n99, B2 => n1504, C1 => n96, C2 => n3566, A
                           => n736, ZN => n741);
   U766 : OAI22_X1 port map( A1 => n3572, A2 => n105, B1 => n3569, B2 => n102, 
                           ZN => n737);
   U767 : AOI221_X1 port map( B1 => n111, B2 => n4079, C1 => n108, C2 => n3573,
                           A => n737, ZN => n740);
   U768 : OAI22_X1 port map( A1 => n2639, A2 => n117, B1 => n388, B2 => n114, 
                           ZN => n738);
   U769 : AOI221_X1 port map( B1 => n123, B2 => n3574, C1 => n120, C2 => n1634,
                           A => n738, ZN => n739);
   U770 : NAND4_X1 port map( A1 => n742, A2 => n741, A3 => n740, A4 => n739, ZN
                           => n3000);
   U771 : OAI211_X1 port map( C1 => n2962, C2 => n69, A => n2468, B => n2467, 
                           ZN => n743);
   U772 : AOI221_X1 port map( B1 => n354, B2 => n1861, C1 => n363, C2 => n4048,
                           A => n743, ZN => n746);
   U773 : NOR2_X1 port map( A1 => n4107, A2 => n72, ZN => n744);
   U774 : NOR4_X1 port map( A1 => n2472, A2 => n2471, A3 => n2466, A4 => n744, 
                           ZN => n745);
   U775 : NAND2_X1 port map( A1 => n746, A2 => n745, ZN => n748);
   U776 : OAI22_X1 port map( A1 => n1228, A2 => n78, B1 => n1227, B2 => n75, ZN
                           => n747);
   U777 : AOI221_X1 port map( B1 => n86, B2 => n748, C1 => n81, C2 => n1537, A 
                           => n747, ZN => n755);
   U778 : OAI22_X1 port map( A1 => n4016, A2 => n93, B1 => n3984, B2 => n90, ZN
                           => n749);
   U779 : AOI221_X1 port map( B1 => n99, B2 => n1505, C1 => n96, C2 => n2967, A
                           => n749, ZN => n754);
   U780 : OAI22_X1 port map( A1 => n2973, A2 => n105, B1 => n2970, B2 => n102, 
                           ZN => n750);
   U781 : AOI221_X1 port map( B1 => n111, B2 => n4080, C1 => n108, C2 => n2974,
                           A => n750, ZN => n753);
   U782 : OAI22_X1 port map( A1 => n2640, A2 => n117, B1 => n389, B2 => n114, 
                           ZN => n751);
   U783 : AOI221_X1 port map( B1 => n123, B2 => n2975, C1 => n120, C2 => n1635,
                           A => n751, ZN => n752);
   U784 : NAND4_X1 port map( A1 => n755, A2 => n754, A3 => n753, A4 => n752, ZN
                           => n3001);
   U785 : OAI211_X1 port map( C1 => n2939, C2 => n69, A => n2461, B => n2460, 
                           ZN => n756);
   U786 : AOI221_X1 port map( B1 => n354, B2 => n1862, C1 => n363, C2 => n4049,
                           A => n756, ZN => n759);
   U787 : NOR2_X1 port map( A1 => n4106, A2 => n72, ZN => n757);
   U788 : NOR4_X1 port map( A1 => n2465, A2 => n2464, A3 => n2459, A4 => n757, 
                           ZN => n758);
   U789 : NAND2_X1 port map( A1 => n759, A2 => n758, ZN => n761);
   U790 : OAI22_X1 port map( A1 => n1244, A2 => n78, B1 => n1243, B2 => n75, ZN
                           => n760);
   U791 : AOI221_X1 port map( B1 => n86, B2 => n761, C1 => n81, C2 => n1538, A 
                           => n760, ZN => n768);
   U792 : OAI22_X1 port map( A1 => n4017, A2 => n93, B1 => n3985, B2 => n90, ZN
                           => n762);
   U793 : AOI221_X1 port map( B1 => n99, B2 => n1506, C1 => n96, C2 => n2944, A
                           => n762, ZN => n767);
   U794 : OAI22_X1 port map( A1 => n2950, A2 => n105, B1 => n2947, B2 => n102, 
                           ZN => n763);
   U795 : AOI221_X1 port map( B1 => n111, B2 => n4081, C1 => n108, C2 => n2951,
                           A => n763, ZN => n766);
   U796 : OAI22_X1 port map( A1 => n2641, A2 => n117, B1 => n390, B2 => n114, 
                           ZN => n764);
   U797 : AOI221_X1 port map( B1 => n123, B2 => n2952, C1 => n120, C2 => n1636,
                           A => n764, ZN => n765);
   U798 : NAND4_X1 port map( A1 => n768, A2 => n767, A3 => n766, A4 => n765, ZN
                           => n3002);
   U799 : OAI211_X1 port map( C1 => n2916, C2 => n69, A => n2454, B => n2453, 
                           ZN => n769);
   U800 : AOI221_X1 port map( B1 => n354, B2 => n1863, C1 => n363, C2 => n4050,
                           A => n769, ZN => n772);
   U801 : NOR2_X1 port map( A1 => n4105, A2 => n72, ZN => n770);
   U802 : NOR4_X1 port map( A1 => n2458, A2 => n2457, A3 => n2452, A4 => n770, 
                           ZN => n771);
   U803 : NAND2_X1 port map( A1 => n772, A2 => n771, ZN => n774);
   U804 : OAI22_X1 port map( A1 => n1260, A2 => n78, B1 => n1259, B2 => n75, ZN
                           => n773);
   U805 : AOI221_X1 port map( B1 => n86, B2 => n774, C1 => n81, C2 => n1539, A 
                           => n773, ZN => n781);
   U806 : OAI22_X1 port map( A1 => n4018, A2 => n93, B1 => n3986, B2 => n90, ZN
                           => n775);
   U807 : AOI221_X1 port map( B1 => n99, B2 => n1507, C1 => n96, C2 => n2921, A
                           => n775, ZN => n780);
   U808 : OAI22_X1 port map( A1 => n2927, A2 => n105, B1 => n2924, B2 => n102, 
                           ZN => n776);
   U809 : AOI221_X1 port map( B1 => n111, B2 => n4082, C1 => n108, C2 => n2928,
                           A => n776, ZN => n779);
   U810 : OAI22_X1 port map( A1 => n2642, A2 => n117, B1 => n391, B2 => n114, 
                           ZN => n777);
   U811 : AOI221_X1 port map( B1 => n123, B2 => n2929, C1 => n120, C2 => n1637,
                           A => n777, ZN => n778);
   U812 : NAND4_X1 port map( A1 => n781, A2 => n780, A3 => n779, A4 => n778, ZN
                           => n3003);
   U813 : OAI211_X1 port map( C1 => n2893, C2 => n69, A => n2447, B => n2446, 
                           ZN => n782);
   U814 : AOI221_X1 port map( B1 => n354, B2 => n1864, C1 => n363, C2 => n4051,
                           A => n782, ZN => n785);
   U815 : NOR2_X1 port map( A1 => n4104, A2 => n72, ZN => n783);
   U816 : NOR4_X1 port map( A1 => n2451, A2 => n2450, A3 => n2445, A4 => n783, 
                           ZN => n784);
   U817 : NAND2_X1 port map( A1 => n785, A2 => n784, ZN => n787);
   U818 : OAI22_X1 port map( A1 => n1276, A2 => n78, B1 => n1275, B2 => n75, ZN
                           => n786);
   U819 : AOI221_X1 port map( B1 => n86, B2 => n787, C1 => n81, C2 => n1540, A 
                           => n786, ZN => n794);
   U820 : OAI22_X1 port map( A1 => n4019, A2 => n93, B1 => n3987, B2 => n90, ZN
                           => n788);
   U821 : AOI221_X1 port map( B1 => n99, B2 => n1508, C1 => n96, C2 => n2898, A
                           => n788, ZN => n793);
   U822 : OAI22_X1 port map( A1 => n2904, A2 => n105, B1 => n2901, B2 => n102, 
                           ZN => n789);
   U823 : AOI221_X1 port map( B1 => n111, B2 => n4083, C1 => n108, C2 => n2905,
                           A => n789, ZN => n792);
   U824 : OAI22_X1 port map( A1 => n2643, A2 => n117, B1 => n392, B2 => n114, 
                           ZN => n790);
   U825 : AOI221_X1 port map( B1 => n123, B2 => n2906, C1 => n120, C2 => n1638,
                           A => n790, ZN => n791);
   U826 : NAND4_X1 port map( A1 => n794, A2 => n793, A3 => n792, A4 => n791, ZN
                           => n3004);
   U827 : OAI211_X1 port map( C1 => n2870, C2 => n69, A => n2440, B => n2439, 
                           ZN => n795);
   U828 : AOI221_X1 port map( B1 => n354, B2 => n1865, C1 => n363, C2 => n4052,
                           A => n795, ZN => n798);
   U829 : NOR2_X1 port map( A1 => n4103, A2 => n72, ZN => n796);
   U830 : NOR4_X1 port map( A1 => n2444, A2 => n2443, A3 => n2438, A4 => n796, 
                           ZN => n797);
   U831 : NAND2_X1 port map( A1 => n798, A2 => n797, ZN => n800);
   U832 : OAI22_X1 port map( A1 => n1292, A2 => n78, B1 => n1291, B2 => n75, ZN
                           => n799);
   U833 : AOI221_X1 port map( B1 => n86, B2 => n800, C1 => n81, C2 => n1541, A 
                           => n799, ZN => n807);
   U834 : OAI22_X1 port map( A1 => n4020, A2 => n93, B1 => n3988, B2 => n90, ZN
                           => n801);
   U835 : AOI221_X1 port map( B1 => n99, B2 => n1509, C1 => n96, C2 => n2875, A
                           => n801, ZN => n806);
   U836 : OAI22_X1 port map( A1 => n2881, A2 => n105, B1 => n2878, B2 => n102, 
                           ZN => n802);
   U837 : AOI221_X1 port map( B1 => n111, B2 => n4084, C1 => n108, C2 => n2882,
                           A => n802, ZN => n805);
   U838 : OAI22_X1 port map( A1 => n2644, A2 => n116, B1 => n393, B2 => n114, 
                           ZN => n803);
   U839 : AOI221_X1 port map( B1 => n123, B2 => n2883, C1 => n120, C2 => n1639,
                           A => n803, ZN => n804);
   U840 : NAND4_X1 port map( A1 => n807, A2 => n806, A3 => n805, A4 => n804, ZN
                           => n3005);
   U841 : OAI211_X1 port map( C1 => n2847, C2 => n69, A => n2433, B => n2432, 
                           ZN => n808);
   U842 : AOI221_X1 port map( B1 => n354, B2 => n1866, C1 => n363, C2 => n4053,
                           A => n808, ZN => n811);
   U843 : NOR2_X1 port map( A1 => n4102, A2 => n72, ZN => n809);
   U844 : NOR4_X1 port map( A1 => n2437, A2 => n2436, A3 => n2431, A4 => n809, 
                           ZN => n810);
   U845 : NAND2_X1 port map( A1 => n811, A2 => n810, ZN => n813);
   U846 : OAI22_X1 port map( A1 => n1308, A2 => n78, B1 => n1307, B2 => n75, ZN
                           => n812);
   U847 : AOI221_X1 port map( B1 => n86, B2 => n813, C1 => n81, C2 => n1542, A 
                           => n812, ZN => n820);
   U848 : OAI22_X1 port map( A1 => n4021, A2 => n93, B1 => n3989, B2 => n90, ZN
                           => n814);
   U849 : AOI221_X1 port map( B1 => n99, B2 => n1510, C1 => n96, C2 => n2852, A
                           => n814, ZN => n819);
   U850 : OAI22_X1 port map( A1 => n2858, A2 => n105, B1 => n2855, B2 => n102, 
                           ZN => n815);
   U851 : AOI221_X1 port map( B1 => n111, B2 => n4085, C1 => n108, C2 => n2859,
                           A => n815, ZN => n818);
   U852 : OAI22_X1 port map( A1 => n2645, A2 => n116, B1 => n394, B2 => n114, 
                           ZN => n816);
   U853 : AOI221_X1 port map( B1 => n123, B2 => n2860, C1 => n120, C2 => n1640,
                           A => n816, ZN => n817);
   U854 : NAND4_X1 port map( A1 => n820, A2 => n819, A3 => n818, A4 => n817, ZN
                           => n3006);
   U855 : OAI211_X1 port map( C1 => n2824, C2 => n70, A => n2426, B => n2425, 
                           ZN => n821);
   U856 : AOI221_X1 port map( B1 => n355, B2 => n1867, C1 => n364, C2 => n4054,
                           A => n821, ZN => n824);
   U857 : NOR2_X1 port map( A1 => n4101, A2 => n73, ZN => n822);
   U858 : NOR4_X1 port map( A1 => n2430, A2 => n2429, A3 => n2424, A4 => n822, 
                           ZN => n823);
   U859 : NAND2_X1 port map( A1 => n824, A2 => n823, ZN => n826);
   U860 : OAI22_X1 port map( A1 => n1324, A2 => n79, B1 => n1323, B2 => n76, ZN
                           => n825);
   U861 : AOI221_X1 port map( B1 => n86, B2 => n826, C1 => n82, C2 => n1543, A 
                           => n825, ZN => n833);
   U862 : OAI22_X1 port map( A1 => n4022, A2 => n94, B1 => n3990, B2 => n91, ZN
                           => n827);
   U863 : AOI221_X1 port map( B1 => n100, B2 => n1511, C1 => n97, C2 => n2829, 
                           A => n827, ZN => n832);
   U864 : OAI22_X1 port map( A1 => n2835, A2 => n106, B1 => n2832, B2 => n103, 
                           ZN => n828);
   U865 : AOI221_X1 port map( B1 => n112, B2 => n4086, C1 => n109, C2 => n2836,
                           A => n828, ZN => n831);
   U866 : OAI22_X1 port map( A1 => n2646, A2 => n116, B1 => n395, B2 => n115, 
                           ZN => n829);
   U867 : AOI221_X1 port map( B1 => n124, B2 => n2837, C1 => n121, C2 => n1641,
                           A => n829, ZN => n830);
   U868 : NAND4_X1 port map( A1 => n833, A2 => n832, A3 => n831, A4 => n830, ZN
                           => n3007);
   U869 : OAI211_X1 port map( C1 => n2801, C2 => n70, A => n2419, B => n2418, 
                           ZN => n834);
   U870 : AOI221_X1 port map( B1 => n355, B2 => n1868, C1 => n364, C2 => n4055,
                           A => n834, ZN => n837);
   U871 : NOR2_X1 port map( A1 => n4100, A2 => n73, ZN => n835);
   U872 : NOR4_X1 port map( A1 => n2423, A2 => n2422, A3 => n2417, A4 => n835, 
                           ZN => n836);
   U873 : NAND2_X1 port map( A1 => n837, A2 => n836, ZN => n839);
   U874 : OAI22_X1 port map( A1 => n1340, A2 => n79, B1 => n1339, B2 => n76, ZN
                           => n838);
   U875 : AOI221_X1 port map( B1 => n86, B2 => n839, C1 => n82, C2 => n1544, A 
                           => n838, ZN => n846);
   U876 : OAI22_X1 port map( A1 => n4023, A2 => n94, B1 => n3991, B2 => n91, ZN
                           => n840);
   U877 : AOI221_X1 port map( B1 => n100, B2 => n1512, C1 => n97, C2 => n2806, 
                           A => n840, ZN => n845);
   U878 : OAI22_X1 port map( A1 => n2812, A2 => n106, B1 => n2809, B2 => n103, 
                           ZN => n841);
   U879 : AOI221_X1 port map( B1 => n112, B2 => n4087, C1 => n109, C2 => n2813,
                           A => n841, ZN => n844);
   U880 : OAI22_X1 port map( A1 => n2647, A2 => n116, B1 => n396, B2 => n115, 
                           ZN => n842);
   U881 : AOI221_X1 port map( B1 => n124, B2 => n2814, C1 => n121, C2 => n1642,
                           A => n842, ZN => n843);
   U882 : NAND4_X1 port map( A1 => n846, A2 => n845, A3 => n844, A4 => n843, ZN
                           => n3008);
   U883 : OAI211_X1 port map( C1 => n2778, C2 => n70, A => n2412, B => n2411, 
                           ZN => n847);
   U884 : AOI221_X1 port map( B1 => n355, B2 => n1869, C1 => n364, C2 => n4056,
                           A => n847, ZN => n850);
   U885 : NOR2_X1 port map( A1 => n4099, A2 => n73, ZN => n848);
   U886 : NOR4_X1 port map( A1 => n2416, A2 => n2415, A3 => n2410, A4 => n848, 
                           ZN => n849);
   U887 : NAND2_X1 port map( A1 => n850, A2 => n849, ZN => n852);
   U888 : OAI22_X1 port map( A1 => n1356, A2 => n79, B1 => n1355, B2 => n76, ZN
                           => n851);
   U889 : AOI221_X1 port map( B1 => n86, B2 => n852, C1 => n82, C2 => n1545, A 
                           => n851, ZN => n859);
   U890 : OAI22_X1 port map( A1 => n4024, A2 => n94, B1 => n3992, B2 => n91, ZN
                           => n853);
   U891 : AOI221_X1 port map( B1 => n100, B2 => n1513, C1 => n97, C2 => n2783, 
                           A => n853, ZN => n858);
   U892 : OAI22_X1 port map( A1 => n2789, A2 => n106, B1 => n2786, B2 => n103, 
                           ZN => n854);
   U893 : AOI221_X1 port map( B1 => n112, B2 => n4088, C1 => n109, C2 => n2790,
                           A => n854, ZN => n857);
   U894 : OAI22_X1 port map( A1 => n2648, A2 => n116, B1 => n397, B2 => n115, 
                           ZN => n855);
   U895 : AOI221_X1 port map( B1 => n124, B2 => n2791, C1 => n121, C2 => n1643,
                           A => n855, ZN => n856);
   U896 : NAND4_X1 port map( A1 => n859, A2 => n858, A3 => n857, A4 => n856, ZN
                           => n3009);
   U897 : OAI211_X1 port map( C1 => n2755, C2 => n70, A => n2405, B => n2404, 
                           ZN => n860);
   U898 : AOI221_X1 port map( B1 => n355, B2 => n1870, C1 => n364, C2 => n4057,
                           A => n860, ZN => n863);
   U899 : NOR2_X1 port map( A1 => n4098, A2 => n73, ZN => n861);
   U900 : NOR4_X1 port map( A1 => n2409, A2 => n2408, A3 => n2403, A4 => n861, 
                           ZN => n862);
   U901 : NAND2_X1 port map( A1 => n863, A2 => n862, ZN => n865);
   U902 : OAI22_X1 port map( A1 => n1372, A2 => n79, B1 => n1371, B2 => n76, ZN
                           => n864);
   U903 : AOI221_X1 port map( B1 => n86, B2 => n865, C1 => n82, C2 => n1546, A 
                           => n864, ZN => n872);
   U904 : OAI22_X1 port map( A1 => n4025, A2 => n94, B1 => n3993, B2 => n91, ZN
                           => n866);
   U905 : AOI221_X1 port map( B1 => n100, B2 => n1514, C1 => n97, C2 => n2760, 
                           A => n866, ZN => n871);
   U906 : OAI22_X1 port map( A1 => n2766, A2 => n106, B1 => n2763, B2 => n103, 
                           ZN => n867);
   U907 : AOI221_X1 port map( B1 => n112, B2 => n4089, C1 => n109, C2 => n2767,
                           A => n867, ZN => n870);
   U908 : OAI22_X1 port map( A1 => n2649, A2 => n116, B1 => n398, B2 => n115, 
                           ZN => n868);
   U909 : AOI221_X1 port map( B1 => n124, B2 => n2768, C1 => n121, C2 => n1644,
                           A => n868, ZN => n869);
   U910 : NAND4_X1 port map( A1 => n872, A2 => n871, A3 => n870, A4 => n869, ZN
                           => n3010);
   U911 : OAI211_X1 port map( C1 => n2732, C2 => n70, A => n2398, B => n2397, 
                           ZN => n873);
   U912 : AOI221_X1 port map( B1 => n355, B2 => n1871, C1 => n364, C2 => n4058,
                           A => n873, ZN => n876);
   U913 : NOR2_X1 port map( A1 => n4097, A2 => n73, ZN => n874);
   U914 : NOR4_X1 port map( A1 => n2402, A2 => n2401, A3 => n2396, A4 => n874, 
                           ZN => n875);
   U915 : NAND2_X1 port map( A1 => n876, A2 => n875, ZN => n878);
   U916 : OAI22_X1 port map( A1 => n1388, A2 => n79, B1 => n1387, B2 => n76, ZN
                           => n877);
   U917 : AOI221_X1 port map( B1 => n85, B2 => n878, C1 => n82, C2 => n1547, A 
                           => n877, ZN => n885);
   U918 : OAI22_X1 port map( A1 => n4026, A2 => n94, B1 => n3994, B2 => n91, ZN
                           => n879);
   U919 : AOI221_X1 port map( B1 => n100, B2 => n1515, C1 => n97, C2 => n2737, 
                           A => n879, ZN => n884);
   U920 : OAI22_X1 port map( A1 => n2743, A2 => n106, B1 => n2740, B2 => n103, 
                           ZN => n880);
   U921 : AOI221_X1 port map( B1 => n112, B2 => n4090, C1 => n109, C2 => n2744,
                           A => n880, ZN => n883);
   U922 : OAI22_X1 port map( A1 => n2650, A2 => n116, B1 => n399, B2 => n115, 
                           ZN => n881);
   U923 : AOI221_X1 port map( B1 => n124, B2 => n2745, C1 => n121, C2 => n1645,
                           A => n881, ZN => n882);
   U924 : NAND4_X1 port map( A1 => n885, A2 => n884, A3 => n883, A4 => n882, ZN
                           => n3011);
   U925 : OAI211_X1 port map( C1 => n2709, C2 => n70, A => n2391, B => n2390, 
                           ZN => n886);
   U926 : AOI221_X1 port map( B1 => n355, B2 => n1872, C1 => n364, C2 => n4059,
                           A => n886, ZN => n889);
   U927 : NOR2_X1 port map( A1 => n4096, A2 => n73, ZN => n887);
   U928 : NOR4_X1 port map( A1 => n2395, A2 => n2394, A3 => n2389, A4 => n887, 
                           ZN => n888);
   U929 : NAND2_X1 port map( A1 => n889, A2 => n888, ZN => n891);
   U930 : OAI22_X1 port map( A1 => n1404, A2 => n79, B1 => n1403, B2 => n76, ZN
                           => n890);
   U931 : AOI221_X1 port map( B1 => n85, B2 => n891, C1 => n82, C2 => n1548, A 
                           => n890, ZN => n898);
   U932 : OAI22_X1 port map( A1 => n4027, A2 => n94, B1 => n3995, B2 => n91, ZN
                           => n892);
   U933 : AOI221_X1 port map( B1 => n100, B2 => n1516, C1 => n97, C2 => n2714, 
                           A => n892, ZN => n897);
   U934 : OAI22_X1 port map( A1 => n2720, A2 => n106, B1 => n2717, B2 => n103, 
                           ZN => n893);
   U935 : AOI221_X1 port map( B1 => n112, B2 => n4091, C1 => n109, C2 => n2721,
                           A => n893, ZN => n896);
   U936 : OAI22_X1 port map( A1 => n2651, A2 => n116, B1 => n400, B2 => n115, 
                           ZN => n894);
   U937 : AOI221_X1 port map( B1 => n124, B2 => n2722, C1 => n121, C2 => n1646,
                           A => n894, ZN => n895);
   U938 : NAND4_X1 port map( A1 => n898, A2 => n897, A3 => n896, A4 => n895, ZN
                           => n3012);
   U939 : OAI211_X1 port map( C1 => n2686, C2 => n70, A => n2384, B => n2383, 
                           ZN => n899);
   U940 : AOI221_X1 port map( B1 => n355, B2 => n1873, C1 => n364, C2 => n4060,
                           A => n899, ZN => n902);
   U941 : NOR2_X1 port map( A1 => n4095, A2 => n73, ZN => n900);
   U942 : NOR4_X1 port map( A1 => n2388, A2 => n2387, A3 => n2382, A4 => n900, 
                           ZN => n901);
   U943 : NAND2_X1 port map( A1 => n902, A2 => n901, ZN => n904);
   U944 : OAI22_X1 port map( A1 => n1420, A2 => n79, B1 => n1419, B2 => n76, ZN
                           => n903);
   U945 : AOI221_X1 port map( B1 => n85, B2 => n904, C1 => n82, C2 => n1549, A 
                           => n903, ZN => n911);
   U946 : OAI22_X1 port map( A1 => n4028, A2 => n94, B1 => n3996, B2 => n91, ZN
                           => n905);
   U947 : AOI221_X1 port map( B1 => n100, B2 => n1517, C1 => n97, C2 => n2691, 
                           A => n905, ZN => n910);
   U948 : OAI22_X1 port map( A1 => n2697, A2 => n106, B1 => n2694, B2 => n103, 
                           ZN => n906);
   U949 : AOI221_X1 port map( B1 => n112, B2 => n4092, C1 => n109, C2 => n2698,
                           A => n906, ZN => n909);
   U950 : OAI22_X1 port map( A1 => n2652, A2 => n116, B1 => n401, B2 => n115, 
                           ZN => n907);
   U951 : AOI221_X1 port map( B1 => n124, B2 => n2699, C1 => n121, C2 => n1647,
                           A => n907, ZN => n908);
   U952 : NAND4_X1 port map( A1 => n911, A2 => n910, A3 => n909, A4 => n908, ZN
                           => n3013);
   U953 : OAI211_X1 port map( C1 => n2663, C2 => n70, A => n2363, B => n2362, 
                           ZN => n912);
   U954 : AOI221_X1 port map( B1 => n355, B2 => n1874, C1 => n364, C2 => n4061,
                           A => n912, ZN => n915);
   U955 : NOR2_X1 port map( A1 => n4094, A2 => n73, ZN => n913);
   U956 : NOR4_X1 port map( A1 => n2379, A2 => n2375, A3 => n2357, A4 => n913, 
                           ZN => n914);
   U957 : NAND2_X1 port map( A1 => n915, A2 => n914, ZN => n919);
   U958 : OAI22_X1 port map( A1 => n1437, A2 => n79, B1 => n1435, B2 => n76, ZN
                           => n918);
   U959 : AOI221_X1 port map( B1 => n87, B2 => n919, C1 => n82, C2 => n1550, A 
                           => n918, ZN => n932);
   U960 : OAI22_X1 port map( A1 => n4029, A2 => n94, B1 => n3997, B2 => n91, ZN
                           => n923);
   U961 : AOI221_X1 port map( B1 => n100, B2 => n1518, C1 => n97, C2 => n2668, 
                           A => n923, ZN => n931);
   U962 : OAI22_X1 port map( A1 => n2674, A2 => n106, B1 => n2671, B2 => n103, 
                           ZN => n926);
   U963 : AOI221_X1 port map( B1 => n112, B2 => n4093, C1 => n109, C2 => n2675,
                           A => n926, ZN => n930);
   U964 : OAI22_X1 port map( A1 => n2653, A2 => n117, B1 => n402, B2 => n115, 
                           ZN => n928);
   U965 : AOI221_X1 port map( B1 => n124, B2 => n2676, C1 => n121, C2 => n1648,
                           A => n928, ZN => n929);
   U966 : NAND4_X1 port map( A1 => n932, A2 => n931, A3 => n930, A4 => n929, ZN
                           => n3014);
   U967 : NAND3_X1 port map( A1 => n2342, A2 => n2341, A3 => n67, ZN => n933);
   U968 : NAND2_X1 port map( A1 => n173, A2 => n933, ZN => n944);
   U969 : INV_X1 port map( A => n944, ZN => n1441);
   U970 : OAI211_X1 port map( C1 => n3952, C2 => n125, A => n1927, B => n1926, 
                           ZN => n934);
   U971 : AOI221_X1 port map( B1 => n305, B2 => n1843, C1 => n4030, C2 => n314,
                           A => n934, ZN => n937);
   U972 : NOR2_X1 port map( A1 => n4125, A2 => n128, ZN => n935);
   U973 : NOR4_X1 port map( A1 => n1945, A2 => n1939, A3 => n1920, A4 => n935, 
                           ZN => n936);
   U974 : NAND2_X1 port map( A1 => n937, A2 => n936, ZN => n941);
   U975 : OR2_X1 port map( A1 => n1910, A2 => n944, ZN => n1438);
   U976 : NAND2_X1 port map( A1 => n1911, A2 => n142, ZN => n1436);
   U977 : OAI22_X1 port map( A1 => n134, A2 => n939, B1 => n131, B2 => n938, ZN
                           => n940);
   U978 : AOI221_X1 port map( B1 => n142, B2 => n941, C1 => n137, C2 => n1519, 
                           A => n940, ZN => n949);
   U979 : OR2_X1 port map( A1 => n1914, A2 => n944, ZN => n1443);
   U980 : NAND2_X1 port map( A1 => n1915, A2 => n142, ZN => n1442);
   U981 : OAI22_X1 port map( A1 => n3998, A2 => n149, B1 => n3966, B2 => n146, 
                           ZN => n942);
   U982 : AOI221_X1 port map( B1 => n155, B2 => n1487, C1 => n3957, C2 => n152,
                           A => n942, ZN => n948);
   U983 : NAND2_X1 port map( A1 => n1925, A2 => n142, ZN => n1446);
   U984 : NAND2_X1 port map( A1 => n1918, A2 => n142, ZN => n1445);
   U985 : OAI22_X1 port map( A1 => n3963, A2 => n161, B1 => n3960, B2 => n158, 
                           ZN => n943);
   U986 : AOI221_X1 port map( B1 => n4062, B2 => n167, C1 => n3964, C2 => n164,
                           A => n943, ZN => n947);
   U987 : NAND4_X1 port map( A1 => n67, A2 => n2341, A3 => n173, A4 => n2342, 
                           ZN => n1448);
   U988 : OAI22_X1 port map( A1 => n3943, A2 => n173, B1 => n170, B2 => n371, 
                           ZN => n945);
   U989 : AOI221_X1 port map( B1 => n3965, B2 => n179, C1 => n176, C2 => n1617,
                           A => n945, ZN => n946);
   U990 : NAND4_X1 port map( A1 => n949, A2 => n948, A3 => n947, A4 => n946, ZN
                           => n3046);
   U991 : MUX2_X1 port map( A => n950, B => DATAIN(0), S => n182, Z => n4446);
   U992 : OAI211_X1 port map( C1 => n3929, C2 => n125, A => n1953, B => n1952, 
                           ZN => n951);
   U993 : AOI221_X1 port map( B1 => n305, B2 => n1844, C1 => n4031, C2 => n314,
                           A => n951, ZN => n954);
   U994 : NOR2_X1 port map( A1 => n4124, A2 => n128, ZN => n952);
   U995 : NOR4_X1 port map( A1 => n1959, A2 => n1956, A3 => n1950, A4 => n952, 
                           ZN => n953);
   U996 : NAND2_X1 port map( A1 => n954, A2 => n953, ZN => n958);
   U997 : OAI22_X1 port map( A1 => n134, A2 => n956, B1 => n131, B2 => n955, ZN
                           => n957);
   U998 : AOI221_X1 port map( B1 => n145, B2 => n958, C1 => n137, C2 => n1520, 
                           A => n957, ZN => n965);
   U999 : OAI22_X1 port map( A1 => n3999, A2 => n149, B1 => n3967, B2 => n146, 
                           ZN => n959);
   U1000 : AOI221_X1 port map( B1 => n155, B2 => n1488, C1 => n3934, C2 => n152
                           , A => n959, ZN => n964);
   U1001 : OAI22_X1 port map( A1 => n3940, A2 => n161, B1 => n3937, B2 => n158,
                           ZN => n960);
   U1002 : AOI221_X1 port map( B1 => n4063, B2 => n167, C1 => n3941, C2 => n164
                           , A => n960, ZN => n963);
   U1003 : OAI22_X1 port map( A1 => n3920, A2 => n175, B1 => n170, B2 => n372, 
                           ZN => n961);
   U1004 : AOI221_X1 port map( B1 => n3942, B2 => n179, C1 => n176, C2 => n1618
                           , A => n961, ZN => n962);
   U1005 : NAND4_X1 port map( A1 => n965, A2 => n964, A3 => n963, A4 => n962, 
                           ZN => n3045);
   U1006 : MUX2_X1 port map( A => n966, B => DATAIN(1), S => n182, Z => n4447);
   U1007 : OAI211_X1 port map( C1 => n3906, C2 => n125, A => n1965, B => n1964,
                           ZN => n967);
   U1008 : AOI221_X1 port map( B1 => n305, B2 => n1845, C1 => n4032, C2 => n314
                           , A => n967, ZN => n970);
   U1009 : NOR2_X1 port map( A1 => n4123, A2 => n128, ZN => n968);
   U1010 : NOR4_X1 port map( A1 => n1971, A2 => n1968, A3 => n1962, A4 => n968,
                           ZN => n969);
   U1011 : NAND2_X1 port map( A1 => n970, A2 => n969, ZN => n974);
   U1012 : OAI22_X1 port map( A1 => n134, A2 => n972, B1 => n131, B2 => n971, 
                           ZN => n973);
   U1013 : AOI221_X1 port map( B1 => n145, B2 => n974, C1 => n137, C2 => n1521,
                           A => n973, ZN => n981);
   U1014 : OAI22_X1 port map( A1 => n4000, A2 => n149, B1 => n3968, B2 => n146,
                           ZN => n975);
   U1015 : AOI221_X1 port map( B1 => n155, B2 => n1489, C1 => n3911, C2 => n152
                           , A => n975, ZN => n980);
   U1016 : OAI22_X1 port map( A1 => n3917, A2 => n161, B1 => n3914, B2 => n158,
                           ZN => n976);
   U1017 : AOI221_X1 port map( B1 => n4064, B2 => n167, C1 => n3918, C2 => n164
                           , A => n976, ZN => n979);
   U1018 : OAI22_X1 port map( A1 => n3897, A2 => n175, B1 => n170, B2 => n373, 
                           ZN => n977);
   U1019 : AOI221_X1 port map( B1 => n3919, B2 => n179, C1 => n176, C2 => n1619
                           , A => n977, ZN => n978);
   U1020 : NAND4_X1 port map( A1 => n981, A2 => n980, A3 => n979, A4 => n978, 
                           ZN => n3044);
   U1021 : MUX2_X1 port map( A => n982, B => DATAIN(2), S => n182, Z => n4448);
   U1022 : OAI211_X1 port map( C1 => n3883, C2 => n125, A => n1977, B => n1976,
                           ZN => n983);
   U1023 : AOI221_X1 port map( B1 => n305, B2 => n1846, C1 => n4033, C2 => n314
                           , A => n983, ZN => n986);
   U1024 : NOR2_X1 port map( A1 => n4122, A2 => n128, ZN => n984);
   U1025 : NOR4_X1 port map( A1 => n1983, A2 => n1980, A3 => n1974, A4 => n984,
                           ZN => n985);
   U1026 : NAND2_X1 port map( A1 => n986, A2 => n985, ZN => n990);
   U1027 : OAI22_X1 port map( A1 => n134, A2 => n988, B1 => n131, B2 => n987, 
                           ZN => n989);
   U1028 : AOI221_X1 port map( B1 => n145, B2 => n990, C1 => n137, C2 => n1522,
                           A => n989, ZN => n997);
   U1029 : OAI22_X1 port map( A1 => n4001, A2 => n149, B1 => n3969, B2 => n146,
                           ZN => n991);
   U1030 : AOI221_X1 port map( B1 => n155, B2 => n1490, C1 => n3888, C2 => n152
                           , A => n991, ZN => n996);
   U1031 : OAI22_X1 port map( A1 => n3894, A2 => n161, B1 => n3891, B2 => n158,
                           ZN => n992);
   U1032 : AOI221_X1 port map( B1 => n4065, B2 => n167, C1 => n3895, C2 => n164
                           , A => n992, ZN => n995);
   U1033 : OAI22_X1 port map( A1 => n3874, A2 => n175, B1 => n170, B2 => n374, 
                           ZN => n993);
   U1034 : AOI221_X1 port map( B1 => n3896, B2 => n179, C1 => n176, C2 => n1620
                           , A => n993, ZN => n994);
   U1035 : NAND4_X1 port map( A1 => n997, A2 => n996, A3 => n995, A4 => n994, 
                           ZN => n3043);
   U1036 : MUX2_X1 port map( A => n998, B => DATAIN(3), S => n182, Z => n4449);
   U1037 : OAI211_X1 port map( C1 => n3860, C2 => n125, A => n1989, B => n1988,
                           ZN => n999);
   U1038 : AOI221_X1 port map( B1 => n305, B2 => n1847, C1 => n4034, C2 => n314
                           , A => n999, ZN => n1002);
   U1039 : NOR2_X1 port map( A1 => n4121, A2 => n128, ZN => n1000);
   U1040 : NOR4_X1 port map( A1 => n1995, A2 => n1992, A3 => n1986, A4 => n1000
                           , ZN => n1001);
   U1041 : NAND2_X1 port map( A1 => n1002, A2 => n1001, ZN => n1006);
   U1042 : OAI22_X1 port map( A1 => n134, A2 => n1004, B1 => n131, B2 => n1003,
                           ZN => n1005);
   U1043 : AOI221_X1 port map( B1 => n145, B2 => n1006, C1 => n137, C2 => n1523
                           , A => n1005, ZN => n1013);
   U1044 : OAI22_X1 port map( A1 => n4002, A2 => n149, B1 => n3970, B2 => n146,
                           ZN => n1007);
   U1045 : AOI221_X1 port map( B1 => n155, B2 => n1491, C1 => n3865, C2 => n152
                           , A => n1007, ZN => n1012);
   U1046 : OAI22_X1 port map( A1 => n3871, A2 => n161, B1 => n3868, B2 => n158,
                           ZN => n1008);
   U1047 : AOI221_X1 port map( B1 => n4066, B2 => n167, C1 => n3872, C2 => n164
                           , A => n1008, ZN => n1011);
   U1048 : OAI22_X1 port map( A1 => n3851, A2 => n175, B1 => n170, B2 => n375, 
                           ZN => n1009);
   U1049 : AOI221_X1 port map( B1 => n3873, B2 => n179, C1 => n176, C2 => n1621
                           , A => n1009, ZN => n1010);
   U1050 : NAND4_X1 port map( A1 => n1013, A2 => n1012, A3 => n1011, A4 => 
                           n1010, ZN => n3042);
   U1051 : MUX2_X1 port map( A => n1014, B => DATAIN(4), S => n182, Z => n4450)
                           ;
   U1052 : OAI211_X1 port map( C1 => n3837, C2 => n125, A => n2001, B => n2000,
                           ZN => n1015);
   U1053 : AOI221_X1 port map( B1 => n305, B2 => n1848, C1 => n4035, C2 => n314
                           , A => n1015, ZN => n1018);
   U1054 : NOR2_X1 port map( A1 => n4120, A2 => n128, ZN => n1016);
   U1055 : NOR4_X1 port map( A1 => n2007, A2 => n2004, A3 => n1998, A4 => n1016
                           , ZN => n1017);
   U1056 : NAND2_X1 port map( A1 => n1018, A2 => n1017, ZN => n1022);
   U1057 : OAI22_X1 port map( A1 => n134, A2 => n1020, B1 => n131, B2 => n1019,
                           ZN => n1021);
   U1058 : AOI221_X1 port map( B1 => n144, B2 => n1022, C1 => n137, C2 => n1524
                           , A => n1021, ZN => n1029);
   U1059 : OAI22_X1 port map( A1 => n4003, A2 => n149, B1 => n3971, B2 => n146,
                           ZN => n1023);
   U1060 : AOI221_X1 port map( B1 => n155, B2 => n1492, C1 => n3842, C2 => n152
                           , A => n1023, ZN => n1028);
   U1061 : OAI22_X1 port map( A1 => n3848, A2 => n161, B1 => n3845, B2 => n158,
                           ZN => n1024);
   U1062 : AOI221_X1 port map( B1 => n4067, B2 => n167, C1 => n3849, C2 => n164
                           , A => n1024, ZN => n1027);
   U1063 : OAI22_X1 port map( A1 => n3828, A2 => n175, B1 => n170, B2 => n376, 
                           ZN => n1025);
   U1064 : AOI221_X1 port map( B1 => n3850, B2 => n179, C1 => n176, C2 => n1622
                           , A => n1025, ZN => n1026);
   U1065 : NAND4_X1 port map( A1 => n1029, A2 => n1028, A3 => n1027, A4 => 
                           n1026, ZN => n3041);
   U1066 : MUX2_X1 port map( A => n1030, B => DATAIN(5), S => n182, Z => n4451)
                           ;
   U1067 : OAI211_X1 port map( C1 => n3814, C2 => n125, A => n2013, B => n2012,
                           ZN => n1031);
   U1068 : AOI221_X1 port map( B1 => n305, B2 => n1849, C1 => n4036, C2 => n314
                           , A => n1031, ZN => n1034);
   U1069 : NOR2_X1 port map( A1 => n4119, A2 => n128, ZN => n1032);
   U1070 : NOR4_X1 port map( A1 => n2019, A2 => n2016, A3 => n2010, A4 => n1032
                           , ZN => n1033);
   U1071 : NAND2_X1 port map( A1 => n1034, A2 => n1033, ZN => n1038);
   U1072 : OAI22_X1 port map( A1 => n134, A2 => n1036, B1 => n131, B2 => n1035,
                           ZN => n1037);
   U1073 : AOI221_X1 port map( B1 => n144, B2 => n1038, C1 => n137, C2 => n1525
                           , A => n1037, ZN => n1045);
   U1074 : OAI22_X1 port map( A1 => n4004, A2 => n149, B1 => n3972, B2 => n146,
                           ZN => n1039);
   U1075 : AOI221_X1 port map( B1 => n155, B2 => n1493, C1 => n3819, C2 => n152
                           , A => n1039, ZN => n1044);
   U1076 : OAI22_X1 port map( A1 => n3825, A2 => n161, B1 => n3822, B2 => n158,
                           ZN => n1040);
   U1077 : AOI221_X1 port map( B1 => n4068, B2 => n167, C1 => n3826, C2 => n164
                           , A => n1040, ZN => n1043);
   U1078 : OAI22_X1 port map( A1 => n3805, A2 => n175, B1 => n170, B2 => n377, 
                           ZN => n1041);
   U1079 : AOI221_X1 port map( B1 => n3827, B2 => n179, C1 => n176, C2 => n1623
                           , A => n1041, ZN => n1042);
   U1080 : NAND4_X1 port map( A1 => n1045, A2 => n1044, A3 => n1043, A4 => 
                           n1042, ZN => n3040);
   U1081 : MUX2_X1 port map( A => n1046, B => DATAIN(6), S => n182, Z => n4452)
                           ;
   U1082 : OAI211_X1 port map( C1 => n3791, C2 => n125, A => n2025, B => n2024,
                           ZN => n1047);
   U1083 : AOI221_X1 port map( B1 => n305, B2 => n1850, C1 => n4037, C2 => n314
                           , A => n1047, ZN => n1050);
   U1084 : NOR2_X1 port map( A1 => n4118, A2 => n128, ZN => n1048);
   U1085 : NOR4_X1 port map( A1 => n2031, A2 => n2028, A3 => n2022, A4 => n1048
                           , ZN => n1049);
   U1086 : NAND2_X1 port map( A1 => n1050, A2 => n1049, ZN => n1054);
   U1087 : OAI22_X1 port map( A1 => n134, A2 => n1052, B1 => n131, B2 => n1051,
                           ZN => n1053);
   U1088 : AOI221_X1 port map( B1 => n144, B2 => n1054, C1 => n137, C2 => n1526
                           , A => n1053, ZN => n1061);
   U1089 : OAI22_X1 port map( A1 => n4005, A2 => n149, B1 => n3973, B2 => n146,
                           ZN => n1055);
   U1090 : AOI221_X1 port map( B1 => n155, B2 => n1494, C1 => n3796, C2 => n152
                           , A => n1055, ZN => n1060);
   U1091 : OAI22_X1 port map( A1 => n3802, A2 => n161, B1 => n3799, B2 => n158,
                           ZN => n1056);
   U1092 : AOI221_X1 port map( B1 => n4069, B2 => n167, C1 => n3803, C2 => n164
                           , A => n1056, ZN => n1059);
   U1093 : OAI22_X1 port map( A1 => n3782, A2 => n175, B1 => n170, B2 => n378, 
                           ZN => n1057);
   U1094 : AOI221_X1 port map( B1 => n3804, B2 => n179, C1 => n176, C2 => n1624
                           , A => n1057, ZN => n1058);
   U1095 : NAND4_X1 port map( A1 => n1061, A2 => n1060, A3 => n1059, A4 => 
                           n1058, ZN => n3039);
   U1096 : MUX2_X1 port map( A => n1062, B => DATAIN(7), S => n182, Z => n4453)
                           ;
   U1097 : OAI211_X1 port map( C1 => n3768, C2 => n125, A => n2037, B => n2036,
                           ZN => n1063);
   U1098 : AOI221_X1 port map( B1 => n305, B2 => n1851, C1 => n4038, C2 => n314
                           , A => n1063, ZN => n1066);
   U1099 : NOR2_X1 port map( A1 => n4117, A2 => n128, ZN => n1064);
   U1100 : NOR4_X1 port map( A1 => n2043, A2 => n2040, A3 => n2034, A4 => n1064
                           , ZN => n1065);
   U1101 : NAND2_X1 port map( A1 => n1066, A2 => n1065, ZN => n1070);
   U1102 : OAI22_X1 port map( A1 => n134, A2 => n1068, B1 => n131, B2 => n1067,
                           ZN => n1069);
   U1103 : AOI221_X1 port map( B1 => n144, B2 => n1070, C1 => n137, C2 => n1527
                           , A => n1069, ZN => n1077);
   U1104 : OAI22_X1 port map( A1 => n4006, A2 => n149, B1 => n3974, B2 => n146,
                           ZN => n1071);
   U1105 : AOI221_X1 port map( B1 => n155, B2 => n1495, C1 => n3773, C2 => n152
                           , A => n1071, ZN => n1076);
   U1106 : OAI22_X1 port map( A1 => n3779, A2 => n161, B1 => n3776, B2 => n158,
                           ZN => n1072);
   U1107 : AOI221_X1 port map( B1 => n4070, B2 => n167, C1 => n3780, C2 => n164
                           , A => n1072, ZN => n1075);
   U1108 : OAI22_X1 port map( A1 => n3759, A2 => n175, B1 => n170, B2 => n379, 
                           ZN => n1073);
   U1109 : AOI221_X1 port map( B1 => n3781, B2 => n179, C1 => n176, C2 => n1625
                           , A => n1073, ZN => n1074);
   U1110 : NAND4_X1 port map( A1 => n1077, A2 => n1076, A3 => n1075, A4 => 
                           n1074, ZN => n3038);
   U1111 : MUX2_X1 port map( A => n1078, B => DATAIN(8), S => n182, Z => n4454)
                           ;
   U1112 : OAI211_X1 port map( C1 => n3745, C2 => n125, A => n2049, B => n2048,
                           ZN => n1079);
   U1113 : AOI221_X1 port map( B1 => n305, B2 => n1852, C1 => n4039, C2 => n314
                           , A => n1079, ZN => n1082);
   U1114 : NOR2_X1 port map( A1 => n4116, A2 => n128, ZN => n1080);
   U1115 : NOR4_X1 port map( A1 => n2055, A2 => n2052, A3 => n2046, A4 => n1080
                           , ZN => n1081);
   U1116 : NAND2_X1 port map( A1 => n1082, A2 => n1081, ZN => n1086);
   U1117 : OAI22_X1 port map( A1 => n134, A2 => n1084, B1 => n131, B2 => n1083,
                           ZN => n1085);
   U1118 : AOI221_X1 port map( B1 => n144, B2 => n1086, C1 => n137, C2 => n1528
                           , A => n1085, ZN => n1093);
   U1119 : OAI22_X1 port map( A1 => n4007, A2 => n149, B1 => n3975, B2 => n146,
                           ZN => n1087);
   U1120 : AOI221_X1 port map( B1 => n155, B2 => n1496, C1 => n3750, C2 => n152
                           , A => n1087, ZN => n1092);
   U1121 : OAI22_X1 port map( A1 => n3756, A2 => n161, B1 => n3753, B2 => n158,
                           ZN => n1088);
   U1122 : AOI221_X1 port map( B1 => n4071, B2 => n167, C1 => n3757, C2 => n164
                           , A => n1088, ZN => n1091);
   U1123 : OAI22_X1 port map( A1 => n3736, A2 => n175, B1 => n170, B2 => n380, 
                           ZN => n1089);
   U1124 : AOI221_X1 port map( B1 => n3758, B2 => n179, C1 => n176, C2 => n1626
                           , A => n1089, ZN => n1090);
   U1125 : NAND4_X1 port map( A1 => n1093, A2 => n1092, A3 => n1091, A4 => 
                           n1090, ZN => n3037);
   U1126 : MUX2_X1 port map( A => n1094, B => DATAIN(9), S => n182, Z => n4455)
                           ;
   U1127 : OAI211_X1 port map( C1 => n3722, C2 => n125, A => n2061, B => n2060,
                           ZN => n1095);
   U1128 : AOI221_X1 port map( B1 => n305, B2 => n1853, C1 => n4040, C2 => n314
                           , A => n1095, ZN => n1098);
   U1129 : NOR2_X1 port map( A1 => n4115, A2 => n128, ZN => n1096);
   U1130 : NOR4_X1 port map( A1 => n2067, A2 => n2064, A3 => n2058, A4 => n1096
                           , ZN => n1097);
   U1131 : NAND2_X1 port map( A1 => n1098, A2 => n1097, ZN => n1102);
   U1132 : OAI22_X1 port map( A1 => n134, A2 => n1100, B1 => n131, B2 => n1099,
                           ZN => n1101);
   U1133 : AOI221_X1 port map( B1 => n144, B2 => n1102, C1 => n137, C2 => n1529
                           , A => n1101, ZN => n1109);
   U1134 : OAI22_X1 port map( A1 => n4008, A2 => n149, B1 => n3976, B2 => n146,
                           ZN => n1103);
   U1135 : AOI221_X1 port map( B1 => n155, B2 => n1497, C1 => n3727, C2 => n152
                           , A => n1103, ZN => n1108);
   U1136 : OAI22_X1 port map( A1 => n3733, A2 => n161, B1 => n3730, B2 => n158,
                           ZN => n1104);
   U1137 : AOI221_X1 port map( B1 => n4072, B2 => n167, C1 => n3734, C2 => n164
                           , A => n1104, ZN => n1107);
   U1138 : OAI22_X1 port map( A1 => n3713, A2 => n175, B1 => n170, B2 => n381, 
                           ZN => n1105);
   U1139 : AOI221_X1 port map( B1 => n3735, B2 => n179, C1 => n176, C2 => n1627
                           , A => n1105, ZN => n1106);
   U1140 : NAND4_X1 port map( A1 => n1109, A2 => n1108, A3 => n1107, A4 => 
                           n1106, ZN => n3036);
   U1141 : MUX2_X1 port map( A => n1110, B => DATAIN(10), S => n182, Z => n4456
                           );
   U1142 : OAI211_X1 port map( C1 => n3699, C2 => n125, A => n2073, B => n2072,
                           ZN => n1111);
   U1143 : AOI221_X1 port map( B1 => n305, B2 => n1854, C1 => n4041, C2 => n314
                           , A => n1111, ZN => n1114);
   U1144 : NOR2_X1 port map( A1 => n4114, A2 => n128, ZN => n1112);
   U1145 : NOR4_X1 port map( A1 => n2079, A2 => n2076, A3 => n2070, A4 => n1112
                           , ZN => n1113);
   U1146 : NAND2_X1 port map( A1 => n1114, A2 => n1113, ZN => n1118);
   U1147 : OAI22_X1 port map( A1 => n134, A2 => n1116, B1 => n131, B2 => n1115,
                           ZN => n1117);
   U1148 : AOI221_X1 port map( B1 => n144, B2 => n1118, C1 => n137, C2 => n1530
                           , A => n1117, ZN => n1125);
   U1149 : OAI22_X1 port map( A1 => n4009, A2 => n149, B1 => n3977, B2 => n146,
                           ZN => n1119);
   U1150 : AOI221_X1 port map( B1 => n155, B2 => n1498, C1 => n3704, C2 => n152
                           , A => n1119, ZN => n1124);
   U1151 : OAI22_X1 port map( A1 => n3710, A2 => n161, B1 => n3707, B2 => n158,
                           ZN => n1120);
   U1152 : AOI221_X1 port map( B1 => n4073, B2 => n167, C1 => n3711, C2 => n164
                           , A => n1120, ZN => n1123);
   U1153 : OAI22_X1 port map( A1 => n3690, A2 => n174, B1 => n170, B2 => n382, 
                           ZN => n1121);
   U1154 : AOI221_X1 port map( B1 => n3712, B2 => n179, C1 => n176, C2 => n1628
                           , A => n1121, ZN => n1122);
   U1155 : NAND4_X1 port map( A1 => n1125, A2 => n1124, A3 => n1123, A4 => 
                           n1122, ZN => n3035);
   U1156 : MUX2_X1 port map( A => n1126, B => DATAIN(11), S => n182, Z => n4457
                           );
   U1157 : OAI211_X1 port map( C1 => n3676, C2 => n126, A => n2085, B => n2084,
                           ZN => n1127);
   U1158 : AOI221_X1 port map( B1 => n306, B2 => n1855, C1 => n4042, C2 => n315
                           , A => n1127, ZN => n1130);
   U1159 : NOR2_X1 port map( A1 => n4113, A2 => n129, ZN => n1128);
   U1160 : NOR4_X1 port map( A1 => n2091, A2 => n2088, A3 => n2082, A4 => n1128
                           , ZN => n1129);
   U1161 : NAND2_X1 port map( A1 => n1130, A2 => n1129, ZN => n1134);
   U1162 : OAI22_X1 port map( A1 => n135, A2 => n1132, B1 => n132, B2 => n1131,
                           ZN => n1133);
   U1163 : AOI221_X1 port map( B1 => n144, B2 => n1134, C1 => n138, C2 => n1531
                           , A => n1133, ZN => n1141);
   U1164 : OAI22_X1 port map( A1 => n4010, A2 => n150, B1 => n3978, B2 => n147,
                           ZN => n1135);
   U1165 : AOI221_X1 port map( B1 => n156, B2 => n1499, C1 => n3681, C2 => n153
                           , A => n1135, ZN => n1140);
   U1166 : OAI22_X1 port map( A1 => n3687, A2 => n162, B1 => n3684, B2 => n159,
                           ZN => n1136);
   U1167 : AOI221_X1 port map( B1 => n4074, B2 => n168, C1 => n3688, C2 => n165
                           , A => n1136, ZN => n1139);
   U1168 : OAI22_X1 port map( A1 => n3667, A2 => n174, B1 => n171, B2 => n383, 
                           ZN => n1137);
   U1169 : AOI221_X1 port map( B1 => n3689, B2 => n180, C1 => n177, C2 => n1629
                           , A => n1137, ZN => n1138);
   U1170 : NAND4_X1 port map( A1 => n1141, A2 => n1140, A3 => n1139, A4 => 
                           n1138, ZN => n3034);
   U1171 : MUX2_X1 port map( A => n1142, B => DATAIN(12), S => n183, Z => n4458
                           );
   U1172 : OAI211_X1 port map( C1 => n3653, C2 => n126, A => n2097, B => n2096,
                           ZN => n1143);
   U1173 : AOI221_X1 port map( B1 => n306, B2 => n1856, C1 => n4043, C2 => n315
                           , A => n1143, ZN => n1146);
   U1174 : NOR2_X1 port map( A1 => n4112, A2 => n129, ZN => n1144);
   U1175 : NOR4_X1 port map( A1 => n2103, A2 => n2100, A3 => n2094, A4 => n1144
                           , ZN => n1145);
   U1176 : NAND2_X1 port map( A1 => n1146, A2 => n1145, ZN => n1150);
   U1177 : OAI22_X1 port map( A1 => n135, A2 => n1148, B1 => n132, B2 => n1147,
                           ZN => n1149);
   U1178 : AOI221_X1 port map( B1 => n144, B2 => n1150, C1 => n138, C2 => n1532
                           , A => n1149, ZN => n1157);
   U1179 : OAI22_X1 port map( A1 => n4011, A2 => n150, B1 => n3979, B2 => n147,
                           ZN => n1151);
   U1180 : AOI221_X1 port map( B1 => n156, B2 => n1500, C1 => n3658, C2 => n153
                           , A => n1151, ZN => n1156);
   U1181 : OAI22_X1 port map( A1 => n3664, A2 => n162, B1 => n3661, B2 => n159,
                           ZN => n1152);
   U1182 : AOI221_X1 port map( B1 => n4075, B2 => n168, C1 => n3665, C2 => n165
                           , A => n1152, ZN => n1155);
   U1183 : OAI22_X1 port map( A1 => n3644, A2 => n174, B1 => n171, B2 => n384, 
                           ZN => n1153);
   U1184 : AOI221_X1 port map( B1 => n3666, B2 => n180, C1 => n177, C2 => n1630
                           , A => n1153, ZN => n1154);
   U1185 : NAND4_X1 port map( A1 => n1157, A2 => n1156, A3 => n1155, A4 => 
                           n1154, ZN => n3033);
   U1186 : MUX2_X1 port map( A => n1158, B => DATAIN(13), S => n183, Z => n4459
                           );
   U1187 : OAI211_X1 port map( C1 => n3630, C2 => n126, A => n2109, B => n2108,
                           ZN => n1159);
   U1188 : AOI221_X1 port map( B1 => n306, B2 => n1857, C1 => n4044, C2 => n315
                           , A => n1159, ZN => n1162);
   U1189 : NOR2_X1 port map( A1 => n4111, A2 => n129, ZN => n1160);
   U1190 : NOR4_X1 port map( A1 => n2115, A2 => n2112, A3 => n2106, A4 => n1160
                           , ZN => n1161);
   U1191 : NAND2_X1 port map( A1 => n1162, A2 => n1161, ZN => n1166);
   U1192 : OAI22_X1 port map( A1 => n135, A2 => n1164, B1 => n132, B2 => n1163,
                           ZN => n1165);
   U1193 : AOI221_X1 port map( B1 => n144, B2 => n1166, C1 => n138, C2 => n1533
                           , A => n1165, ZN => n1173);
   U1194 : OAI22_X1 port map( A1 => n4012, A2 => n150, B1 => n3980, B2 => n147,
                           ZN => n1167);
   U1195 : AOI221_X1 port map( B1 => n156, B2 => n1501, C1 => n3635, C2 => n153
                           , A => n1167, ZN => n1172);
   U1196 : OAI22_X1 port map( A1 => n3641, A2 => n162, B1 => n3638, B2 => n159,
                           ZN => n1168);
   U1197 : AOI221_X1 port map( B1 => n4076, B2 => n168, C1 => n3642, C2 => n165
                           , A => n1168, ZN => n1171);
   U1198 : OAI22_X1 port map( A1 => n3621, A2 => n174, B1 => n171, B2 => n385, 
                           ZN => n1169);
   U1199 : AOI221_X1 port map( B1 => n3643, B2 => n180, C1 => n177, C2 => n1631
                           , A => n1169, ZN => n1170);
   U1200 : NAND4_X1 port map( A1 => n1173, A2 => n1172, A3 => n1171, A4 => 
                           n1170, ZN => n3032);
   U1201 : MUX2_X1 port map( A => n1174, B => DATAIN(14), S => n183, Z => n4460
                           );
   U1202 : OAI211_X1 port map( C1 => n3607, C2 => n126, A => n2121, B => n2120,
                           ZN => n1175);
   U1203 : AOI221_X1 port map( B1 => n306, B2 => n1858, C1 => n4045, C2 => n315
                           , A => n1175, ZN => n1178);
   U1204 : NOR2_X1 port map( A1 => n4110, A2 => n129, ZN => n1176);
   U1205 : NOR4_X1 port map( A1 => n2127, A2 => n2124, A3 => n2118, A4 => n1176
                           , ZN => n1177);
   U1206 : NAND2_X1 port map( A1 => n1178, A2 => n1177, ZN => n1182);
   U1207 : OAI22_X1 port map( A1 => n135, A2 => n1180, B1 => n132, B2 => n1179,
                           ZN => n1181);
   U1208 : AOI221_X1 port map( B1 => n144, B2 => n1182, C1 => n138, C2 => n1534
                           , A => n1181, ZN => n1189);
   U1209 : OAI22_X1 port map( A1 => n4013, A2 => n150, B1 => n3981, B2 => n147,
                           ZN => n1183);
   U1210 : AOI221_X1 port map( B1 => n156, B2 => n1502, C1 => n3612, C2 => n153
                           , A => n1183, ZN => n1188);
   U1211 : OAI22_X1 port map( A1 => n3618, A2 => n162, B1 => n3615, B2 => n159,
                           ZN => n1184);
   U1212 : AOI221_X1 port map( B1 => n4077, B2 => n168, C1 => n3619, C2 => n165
                           , A => n1184, ZN => n1187);
   U1213 : OAI22_X1 port map( A1 => n3598, A2 => n174, B1 => n171, B2 => n386, 
                           ZN => n1185);
   U1214 : AOI221_X1 port map( B1 => n3620, B2 => n180, C1 => n177, C2 => n1632
                           , A => n1185, ZN => n1186);
   U1215 : NAND4_X1 port map( A1 => n1189, A2 => n1188, A3 => n1187, A4 => 
                           n1186, ZN => n3031);
   U1216 : MUX2_X1 port map( A => n1190, B => DATAIN(15), S => n183, Z => n4461
                           );
   U1217 : OAI211_X1 port map( C1 => n3584, C2 => n126, A => n2133, B => n2132,
                           ZN => n1191);
   U1218 : AOI221_X1 port map( B1 => n306, B2 => n1859, C1 => n4046, C2 => n315
                           , A => n1191, ZN => n1194);
   U1219 : NOR2_X1 port map( A1 => n4109, A2 => n129, ZN => n1192);
   U1220 : NOR4_X1 port map( A1 => n2139, A2 => n2136, A3 => n2130, A4 => n1192
                           , ZN => n1193);
   U1221 : NAND2_X1 port map( A1 => n1194, A2 => n1193, ZN => n1198);
   U1222 : OAI22_X1 port map( A1 => n135, A2 => n1196, B1 => n132, B2 => n1195,
                           ZN => n1197);
   U1223 : AOI221_X1 port map( B1 => n143, B2 => n1198, C1 => n138, C2 => n1535
                           , A => n1197, ZN => n1205);
   U1224 : OAI22_X1 port map( A1 => n4014, A2 => n150, B1 => n3982, B2 => n147,
                           ZN => n1199);
   U1225 : AOI221_X1 port map( B1 => n156, B2 => n1503, C1 => n3589, C2 => n153
                           , A => n1199, ZN => n1204);
   U1226 : OAI22_X1 port map( A1 => n3595, A2 => n162, B1 => n3592, B2 => n159,
                           ZN => n1200);
   U1227 : AOI221_X1 port map( B1 => n4078, B2 => n168, C1 => n3596, C2 => n165
                           , A => n1200, ZN => n1203);
   U1228 : OAI22_X1 port map( A1 => n3575, A2 => n174, B1 => n171, B2 => n387, 
                           ZN => n1201);
   U1229 : AOI221_X1 port map( B1 => n3597, B2 => n180, C1 => n177, C2 => n1633
                           , A => n1201, ZN => n1202);
   U1230 : NAND4_X1 port map( A1 => n1205, A2 => n1204, A3 => n1203, A4 => 
                           n1202, ZN => n3030);
   U1231 : MUX2_X1 port map( A => n1206, B => DATAIN(16), S => n183, Z => n4462
                           );
   U1232 : OAI211_X1 port map( C1 => n3561, C2 => n126, A => n2145, B => n2144,
                           ZN => n1207);
   U1233 : AOI221_X1 port map( B1 => n306, B2 => n1860, C1 => n4047, C2 => n315
                           , A => n1207, ZN => n1210);
   U1234 : NOR2_X1 port map( A1 => n4108, A2 => n129, ZN => n1208);
   U1235 : NOR4_X1 port map( A1 => n2151, A2 => n2148, A3 => n2142, A4 => n1208
                           , ZN => n1209);
   U1236 : NAND2_X1 port map( A1 => n1210, A2 => n1209, ZN => n1214);
   U1237 : OAI22_X1 port map( A1 => n135, A2 => n1212, B1 => n132, B2 => n1211,
                           ZN => n1213);
   U1238 : AOI221_X1 port map( B1 => n143, B2 => n1214, C1 => n138, C2 => n1536
                           , A => n1213, ZN => n1221);
   U1239 : OAI22_X1 port map( A1 => n4015, A2 => n150, B1 => n3983, B2 => n147,
                           ZN => n1215);
   U1240 : AOI221_X1 port map( B1 => n156, B2 => n1504, C1 => n3566, C2 => n153
                           , A => n1215, ZN => n1220);
   U1241 : OAI22_X1 port map( A1 => n3572, A2 => n162, B1 => n3569, B2 => n159,
                           ZN => n1216);
   U1242 : AOI221_X1 port map( B1 => n4079, B2 => n168, C1 => n3573, C2 => n165
                           , A => n1216, ZN => n1219);
   U1243 : OAI22_X1 port map( A1 => n2976, A2 => n174, B1 => n171, B2 => n388, 
                           ZN => n1217);
   U1244 : AOI221_X1 port map( B1 => n3574, B2 => n180, C1 => n177, C2 => n1634
                           , A => n1217, ZN => n1218);
   U1245 : NAND4_X1 port map( A1 => n1221, A2 => n1220, A3 => n1219, A4 => 
                           n1218, ZN => n3029);
   U1246 : MUX2_X1 port map( A => n1222, B => DATAIN(17), S => n183, Z => n4463
                           );
   U1247 : OAI211_X1 port map( C1 => n2962, C2 => n126, A => n2157, B => n2156,
                           ZN => n1223);
   U1248 : AOI221_X1 port map( B1 => n306, B2 => n1861, C1 => n4048, C2 => n315
                           , A => n1223, ZN => n1226);
   U1249 : NOR2_X1 port map( A1 => n4107, A2 => n129, ZN => n1224);
   U1250 : NOR4_X1 port map( A1 => n2163, A2 => n2160, A3 => n2154, A4 => n1224
                           , ZN => n1225);
   U1251 : NAND2_X1 port map( A1 => n1226, A2 => n1225, ZN => n1230);
   U1252 : OAI22_X1 port map( A1 => n135, A2 => n1228, B1 => n132, B2 => n1227,
                           ZN => n1229);
   U1253 : AOI221_X1 port map( B1 => n143, B2 => n1230, C1 => n138, C2 => n1537
                           , A => n1229, ZN => n1237);
   U1254 : OAI22_X1 port map( A1 => n4016, A2 => n150, B1 => n3984, B2 => n147,
                           ZN => n1231);
   U1255 : AOI221_X1 port map( B1 => n156, B2 => n1505, C1 => n2967, C2 => n153
                           , A => n1231, ZN => n1236);
   U1256 : OAI22_X1 port map( A1 => n2973, A2 => n162, B1 => n2970, B2 => n159,
                           ZN => n1232);
   U1257 : AOI221_X1 port map( B1 => n4080, B2 => n168, C1 => n2974, C2 => n165
                           , A => n1232, ZN => n1235);
   U1258 : OAI22_X1 port map( A1 => n2953, A2 => n174, B1 => n171, B2 => n389, 
                           ZN => n1233);
   U1259 : AOI221_X1 port map( B1 => n2975, B2 => n180, C1 => n177, C2 => n1635
                           , A => n1233, ZN => n1234);
   U1260 : NAND4_X1 port map( A1 => n1237, A2 => n1236, A3 => n1235, A4 => 
                           n1234, ZN => n3028);
   U1261 : MUX2_X1 port map( A => n1238, B => DATAIN(18), S => n183, Z => n4464
                           );
   U1262 : OAI211_X1 port map( C1 => n2939, C2 => n126, A => n2169, B => n2168,
                           ZN => n1239);
   U1263 : AOI221_X1 port map( B1 => n306, B2 => n1862, C1 => n4049, C2 => n315
                           , A => n1239, ZN => n1242);
   U1264 : NOR2_X1 port map( A1 => n4106, A2 => n129, ZN => n1240);
   U1265 : NOR4_X1 port map( A1 => n2175, A2 => n2172, A3 => n2166, A4 => n1240
                           , ZN => n1241);
   U1266 : NAND2_X1 port map( A1 => n1242, A2 => n1241, ZN => n1246);
   U1267 : OAI22_X1 port map( A1 => n135, A2 => n1244, B1 => n132, B2 => n1243,
                           ZN => n1245);
   U1268 : AOI221_X1 port map( B1 => n143, B2 => n1246, C1 => n138, C2 => n1538
                           , A => n1245, ZN => n1253);
   U1269 : OAI22_X1 port map( A1 => n4017, A2 => n150, B1 => n3985, B2 => n147,
                           ZN => n1247);
   U1270 : AOI221_X1 port map( B1 => n156, B2 => n1506, C1 => n2944, C2 => n153
                           , A => n1247, ZN => n1252);
   U1271 : OAI22_X1 port map( A1 => n2950, A2 => n162, B1 => n2947, B2 => n159,
                           ZN => n1248);
   U1272 : AOI221_X1 port map( B1 => n4081, B2 => n168, C1 => n2951, C2 => n165
                           , A => n1248, ZN => n1251);
   U1273 : OAI22_X1 port map( A1 => n2930, A2 => n174, B1 => n171, B2 => n390, 
                           ZN => n1249);
   U1274 : AOI221_X1 port map( B1 => n2952, B2 => n180, C1 => n177, C2 => n1636
                           , A => n1249, ZN => n1250);
   U1275 : NAND4_X1 port map( A1 => n1253, A2 => n1252, A3 => n1251, A4 => 
                           n1250, ZN => n3027);
   U1276 : MUX2_X1 port map( A => n1254, B => DATAIN(19), S => n183, Z => n4465
                           );
   U1277 : OAI211_X1 port map( C1 => n2916, C2 => n126, A => n2181, B => n2180,
                           ZN => n1255);
   U1278 : AOI221_X1 port map( B1 => n306, B2 => n1863, C1 => n4050, C2 => n315
                           , A => n1255, ZN => n1258);
   U1279 : NOR2_X1 port map( A1 => n4105, A2 => n129, ZN => n1256);
   U1280 : NOR4_X1 port map( A1 => n2187, A2 => n2184, A3 => n2178, A4 => n1256
                           , ZN => n1257);
   U1281 : NAND2_X1 port map( A1 => n1258, A2 => n1257, ZN => n1262);
   U1282 : OAI22_X1 port map( A1 => n135, A2 => n1260, B1 => n132, B2 => n1259,
                           ZN => n1261);
   U1283 : AOI221_X1 port map( B1 => n143, B2 => n1262, C1 => n138, C2 => n1539
                           , A => n1261, ZN => n1269);
   U1284 : OAI22_X1 port map( A1 => n4018, A2 => n150, B1 => n3986, B2 => n147,
                           ZN => n1263);
   U1285 : AOI221_X1 port map( B1 => n156, B2 => n1507, C1 => n2921, C2 => n153
                           , A => n1263, ZN => n1268);
   U1286 : OAI22_X1 port map( A1 => n2927, A2 => n162, B1 => n2924, B2 => n159,
                           ZN => n1264);
   U1287 : AOI221_X1 port map( B1 => n4082, B2 => n168, C1 => n2928, C2 => n165
                           , A => n1264, ZN => n1267);
   U1288 : OAI22_X1 port map( A1 => n2907, A2 => n174, B1 => n171, B2 => n391, 
                           ZN => n1265);
   U1289 : AOI221_X1 port map( B1 => n2929, B2 => n180, C1 => n177, C2 => n1637
                           , A => n1265, ZN => n1266);
   U1290 : NAND4_X1 port map( A1 => n1269, A2 => n1268, A3 => n1267, A4 => 
                           n1266, ZN => n3026);
   U1291 : MUX2_X1 port map( A => n1270, B => DATAIN(20), S => n183, Z => n4466
                           );
   U1292 : OAI211_X1 port map( C1 => n2893, C2 => n126, A => n2193, B => n2192,
                           ZN => n1271);
   U1293 : AOI221_X1 port map( B1 => n306, B2 => n1864, C1 => n4051, C2 => n315
                           , A => n1271, ZN => n1274);
   U1294 : NOR2_X1 port map( A1 => n4104, A2 => n129, ZN => n1272);
   U1295 : NOR4_X1 port map( A1 => n2199, A2 => n2196, A3 => n2190, A4 => n1272
                           , ZN => n1273);
   U1296 : NAND2_X1 port map( A1 => n1274, A2 => n1273, ZN => n1278);
   U1297 : OAI22_X1 port map( A1 => n135, A2 => n1276, B1 => n132, B2 => n1275,
                           ZN => n1277);
   U1298 : AOI221_X1 port map( B1 => n143, B2 => n1278, C1 => n138, C2 => n1540
                           , A => n1277, ZN => n1285);
   U1299 : OAI22_X1 port map( A1 => n4019, A2 => n150, B1 => n3987, B2 => n147,
                           ZN => n1279);
   U1300 : AOI221_X1 port map( B1 => n156, B2 => n1508, C1 => n2898, C2 => n153
                           , A => n1279, ZN => n1284);
   U1301 : OAI22_X1 port map( A1 => n2904, A2 => n162, B1 => n2901, B2 => n159,
                           ZN => n1280);
   U1302 : AOI221_X1 port map( B1 => n4083, B2 => n168, C1 => n2905, C2 => n165
                           , A => n1280, ZN => n1283);
   U1303 : OAI22_X1 port map( A1 => n2884, A2 => n174, B1 => n171, B2 => n392, 
                           ZN => n1281);
   U1304 : AOI221_X1 port map( B1 => n2906, B2 => n180, C1 => n177, C2 => n1638
                           , A => n1281, ZN => n1282);
   U1305 : NAND4_X1 port map( A1 => n1285, A2 => n1284, A3 => n1283, A4 => 
                           n1282, ZN => n3025);
   U1306 : MUX2_X1 port map( A => n1286, B => DATAIN(21), S => n183, Z => n4467
                           );
   U1307 : OAI211_X1 port map( C1 => n2870, C2 => n126, A => n2205, B => n2204,
                           ZN => n1287);
   U1308 : AOI221_X1 port map( B1 => n306, B2 => n1865, C1 => n4052, C2 => n315
                           , A => n1287, ZN => n1290);
   U1309 : NOR2_X1 port map( A1 => n4103, A2 => n129, ZN => n1288);
   U1310 : NOR4_X1 port map( A1 => n2211, A2 => n2208, A3 => n2202, A4 => n1288
                           , ZN => n1289);
   U1311 : NAND2_X1 port map( A1 => n1290, A2 => n1289, ZN => n1294);
   U1312 : OAI22_X1 port map( A1 => n135, A2 => n1292, B1 => n132, B2 => n1291,
                           ZN => n1293);
   U1313 : AOI221_X1 port map( B1 => n143, B2 => n1294, C1 => n138, C2 => n1541
                           , A => n1293, ZN => n1301);
   U1314 : OAI22_X1 port map( A1 => n4020, A2 => n150, B1 => n3988, B2 => n147,
                           ZN => n1295);
   U1315 : AOI221_X1 port map( B1 => n156, B2 => n1509, C1 => n2875, C2 => n153
                           , A => n1295, ZN => n1300);
   U1316 : OAI22_X1 port map( A1 => n2881, A2 => n162, B1 => n2878, B2 => n159,
                           ZN => n1296);
   U1317 : AOI221_X1 port map( B1 => n4084, B2 => n168, C1 => n2882, C2 => n165
                           , A => n1296, ZN => n1299);
   U1318 : OAI22_X1 port map( A1 => n2861, A2 => n173, B1 => n171, B2 => n393, 
                           ZN => n1297);
   U1319 : AOI221_X1 port map( B1 => n2883, B2 => n180, C1 => n177, C2 => n1639
                           , A => n1297, ZN => n1298);
   U1320 : NAND4_X1 port map( A1 => n1301, A2 => n1300, A3 => n1299, A4 => 
                           n1298, ZN => n3024);
   U1321 : MUX2_X1 port map( A => n1302, B => DATAIN(22), S => n183, Z => n4468
                           );
   U1322 : OAI211_X1 port map( C1 => n2847, C2 => n126, A => n2217, B => n2216,
                           ZN => n1303);
   U1323 : AOI221_X1 port map( B1 => n306, B2 => n1866, C1 => n4053, C2 => n315
                           , A => n1303, ZN => n1306);
   U1324 : NOR2_X1 port map( A1 => n4102, A2 => n129, ZN => n1304);
   U1325 : NOR4_X1 port map( A1 => n2223, A2 => n2220, A3 => n2214, A4 => n1304
                           , ZN => n1305);
   U1326 : NAND2_X1 port map( A1 => n1306, A2 => n1305, ZN => n1310);
   U1327 : OAI22_X1 port map( A1 => n135, A2 => n1308, B1 => n132, B2 => n1307,
                           ZN => n1309);
   U1328 : AOI221_X1 port map( B1 => n143, B2 => n1310, C1 => n138, C2 => n1542
                           , A => n1309, ZN => n1317);
   U1329 : OAI22_X1 port map( A1 => n4021, A2 => n150, B1 => n3989, B2 => n147,
                           ZN => n1311);
   U1330 : AOI221_X1 port map( B1 => n156, B2 => n1510, C1 => n2852, C2 => n153
                           , A => n1311, ZN => n1316);
   U1331 : OAI22_X1 port map( A1 => n2858, A2 => n162, B1 => n2855, B2 => n159,
                           ZN => n1312);
   U1332 : AOI221_X1 port map( B1 => n4085, B2 => n168, C1 => n2859, C2 => n165
                           , A => n1312, ZN => n1315);
   U1333 : OAI22_X1 port map( A1 => n2838, A2 => n173, B1 => n171, B2 => n394, 
                           ZN => n1313);
   U1334 : AOI221_X1 port map( B1 => n2860, B2 => n180, C1 => n177, C2 => n1640
                           , A => n1313, ZN => n1314);
   U1335 : NAND4_X1 port map( A1 => n1317, A2 => n1316, A3 => n1315, A4 => 
                           n1314, ZN => n3023);
   U1336 : MUX2_X1 port map( A => n1318, B => DATAIN(23), S => n183, Z => n4469
                           );
   U1337 : OAI211_X1 port map( C1 => n2824, C2 => n127, A => n2229, B => n2228,
                           ZN => n1319);
   U1338 : AOI221_X1 port map( B1 => n307, B2 => n1867, C1 => n4054, C2 => n316
                           , A => n1319, ZN => n1322);
   U1339 : NOR2_X1 port map( A1 => n4101, A2 => n130, ZN => n1320);
   U1340 : NOR4_X1 port map( A1 => n2235, A2 => n2232, A3 => n2226, A4 => n1320
                           , ZN => n1321);
   U1341 : NAND2_X1 port map( A1 => n1322, A2 => n1321, ZN => n1326);
   U1342 : OAI22_X1 port map( A1 => n136, A2 => n1324, B1 => n133, B2 => n1323,
                           ZN => n1325);
   U1343 : AOI221_X1 port map( B1 => n143, B2 => n1326, C1 => n139, C2 => n1543
                           , A => n1325, ZN => n1333);
   U1344 : OAI22_X1 port map( A1 => n4022, A2 => n151, B1 => n3990, B2 => n148,
                           ZN => n1327);
   U1345 : AOI221_X1 port map( B1 => n157, B2 => n1511, C1 => n2829, C2 => n154
                           , A => n1327, ZN => n1332);
   U1346 : OAI22_X1 port map( A1 => n2835, A2 => n163, B1 => n2832, B2 => n160,
                           ZN => n1328);
   U1347 : AOI221_X1 port map( B1 => n4086, B2 => n169, C1 => n2836, C2 => n166
                           , A => n1328, ZN => n1331);
   U1348 : OAI22_X1 port map( A1 => n2815, A2 => n173, B1 => n172, B2 => n395, 
                           ZN => n1329);
   U1349 : AOI221_X1 port map( B1 => n2837, B2 => n181, C1 => n178, C2 => n1641
                           , A => n1329, ZN => n1330);
   U1350 : NAND4_X1 port map( A1 => n1333, A2 => n1332, A3 => n1331, A4 => 
                           n1330, ZN => n3022);
   U1351 : MUX2_X1 port map( A => n1334, B => DATAIN(24), S => n184, Z => n4470
                           );
   U1352 : OAI211_X1 port map( C1 => n2801, C2 => n127, A => n2241, B => n2240,
                           ZN => n1335);
   U1353 : AOI221_X1 port map( B1 => n307, B2 => n1868, C1 => n4055, C2 => n316
                           , A => n1335, ZN => n1338);
   U1354 : NOR2_X1 port map( A1 => n4100, A2 => n130, ZN => n1336);
   U1355 : NOR4_X1 port map( A1 => n2247, A2 => n2244, A3 => n2238, A4 => n1336
                           , ZN => n1337);
   U1356 : NAND2_X1 port map( A1 => n1338, A2 => n1337, ZN => n1342);
   U1357 : OAI22_X1 port map( A1 => n136, A2 => n1340, B1 => n133, B2 => n1339,
                           ZN => n1341);
   U1358 : AOI221_X1 port map( B1 => n143, B2 => n1342, C1 => n139, C2 => n1544
                           , A => n1341, ZN => n1349);
   U1359 : OAI22_X1 port map( A1 => n4023, A2 => n151, B1 => n3991, B2 => n148,
                           ZN => n1343);
   U1360 : AOI221_X1 port map( B1 => n157, B2 => n1512, C1 => n2806, C2 => n154
                           , A => n1343, ZN => n1348);
   U1361 : OAI22_X1 port map( A1 => n2812, A2 => n163, B1 => n2809, B2 => n160,
                           ZN => n1344);
   U1362 : AOI221_X1 port map( B1 => n4087, B2 => n169, C1 => n2813, C2 => n166
                           , A => n1344, ZN => n1347);
   U1363 : OAI22_X1 port map( A1 => n2792, A2 => n173, B1 => n172, B2 => n396, 
                           ZN => n1345);
   U1364 : AOI221_X1 port map( B1 => n2814, B2 => n181, C1 => n178, C2 => n1642
                           , A => n1345, ZN => n1346);
   U1365 : NAND4_X1 port map( A1 => n1349, A2 => n1348, A3 => n1347, A4 => 
                           n1346, ZN => n3021);
   U1366 : MUX2_X1 port map( A => n1350, B => DATAIN(25), S => n184, Z => n4471
                           );
   U1367 : OAI211_X1 port map( C1 => n2778, C2 => n127, A => n2253, B => n2252,
                           ZN => n1351);
   U1368 : AOI221_X1 port map( B1 => n307, B2 => n1869, C1 => n4056, C2 => n316
                           , A => n1351, ZN => n1354);
   U1369 : NOR2_X1 port map( A1 => n4099, A2 => n130, ZN => n1352);
   U1370 : NOR4_X1 port map( A1 => n2259, A2 => n2256, A3 => n2250, A4 => n1352
                           , ZN => n1353);
   U1371 : NAND2_X1 port map( A1 => n1354, A2 => n1353, ZN => n1358);
   U1372 : OAI22_X1 port map( A1 => n136, A2 => n1356, B1 => n133, B2 => n1355,
                           ZN => n1357);
   U1373 : AOI221_X1 port map( B1 => n143, B2 => n1358, C1 => n139, C2 => n1545
                           , A => n1357, ZN => n1365);
   U1374 : OAI22_X1 port map( A1 => n4024, A2 => n151, B1 => n3992, B2 => n148,
                           ZN => n1359);
   U1375 : AOI221_X1 port map( B1 => n157, B2 => n1513, C1 => n2783, C2 => n154
                           , A => n1359, ZN => n1364);
   U1376 : OAI22_X1 port map( A1 => n2789, A2 => n163, B1 => n2786, B2 => n160,
                           ZN => n1360);
   U1377 : AOI221_X1 port map( B1 => n4088, B2 => n169, C1 => n2790, C2 => n166
                           , A => n1360, ZN => n1363);
   U1378 : OAI22_X1 port map( A1 => n2769, A2 => n173, B1 => n172, B2 => n397, 
                           ZN => n1361);
   U1379 : AOI221_X1 port map( B1 => n2791, B2 => n181, C1 => n178, C2 => n1643
                           , A => n1361, ZN => n1362);
   U1380 : NAND4_X1 port map( A1 => n1365, A2 => n1364, A3 => n1363, A4 => 
                           n1362, ZN => n3020);
   U1381 : MUX2_X1 port map( A => n1366, B => DATAIN(26), S => n184, Z => n4472
                           );
   U1382 : OAI211_X1 port map( C1 => n2755, C2 => n127, A => n2265, B => n2264,
                           ZN => n1367);
   U1383 : AOI221_X1 port map( B1 => n307, B2 => n1870, C1 => n4057, C2 => n316
                           , A => n1367, ZN => n1370);
   U1384 : NOR2_X1 port map( A1 => n4098, A2 => n130, ZN => n1368);
   U1385 : NOR4_X1 port map( A1 => n2271, A2 => n2268, A3 => n2262, A4 => n1368
                           , ZN => n1369);
   U1386 : NAND2_X1 port map( A1 => n1370, A2 => n1369, ZN => n1374);
   U1387 : OAI22_X1 port map( A1 => n136, A2 => n1372, B1 => n133, B2 => n1371,
                           ZN => n1373);
   U1388 : AOI221_X1 port map( B1 => n143, B2 => n1374, C1 => n139, C2 => n1546
                           , A => n1373, ZN => n1381);
   U1389 : OAI22_X1 port map( A1 => n4025, A2 => n151, B1 => n3993, B2 => n148,
                           ZN => n1375);
   U1390 : AOI221_X1 port map( B1 => n157, B2 => n1514, C1 => n2760, C2 => n154
                           , A => n1375, ZN => n1380);
   U1391 : OAI22_X1 port map( A1 => n2766, A2 => n163, B1 => n2763, B2 => n160,
                           ZN => n1376);
   U1392 : AOI221_X1 port map( B1 => n4089, B2 => n169, C1 => n2767, C2 => n166
                           , A => n1376, ZN => n1379);
   U1393 : OAI22_X1 port map( A1 => n2746, A2 => n173, B1 => n172, B2 => n398, 
                           ZN => n1377);
   U1394 : AOI221_X1 port map( B1 => n2768, B2 => n181, C1 => n178, C2 => n1644
                           , A => n1377, ZN => n1378);
   U1395 : NAND4_X1 port map( A1 => n1381, A2 => n1380, A3 => n1379, A4 => 
                           n1378, ZN => n3019);
   U1396 : MUX2_X1 port map( A => n1382, B => DATAIN(27), S => n184, Z => n4473
                           );
   U1397 : OAI211_X1 port map( C1 => n2732, C2 => n127, A => n2277, B => n2276,
                           ZN => n1383);
   U1398 : AOI221_X1 port map( B1 => n307, B2 => n1871, C1 => n4058, C2 => n316
                           , A => n1383, ZN => n1386);
   U1399 : NOR2_X1 port map( A1 => n4097, A2 => n130, ZN => n1384);
   U1400 : NOR4_X1 port map( A1 => n2283, A2 => n2280, A3 => n2274, A4 => n1384
                           , ZN => n1385);
   U1401 : NAND2_X1 port map( A1 => n1386, A2 => n1385, ZN => n1390);
   U1402 : OAI22_X1 port map( A1 => n136, A2 => n1388, B1 => n133, B2 => n1387,
                           ZN => n1389);
   U1403 : AOI221_X1 port map( B1 => n142, B2 => n1390, C1 => n139, C2 => n1547
                           , A => n1389, ZN => n1397);
   U1404 : OAI22_X1 port map( A1 => n4026, A2 => n151, B1 => n3994, B2 => n148,
                           ZN => n1391);
   U1405 : AOI221_X1 port map( B1 => n157, B2 => n1515, C1 => n2737, C2 => n154
                           , A => n1391, ZN => n1396);
   U1406 : OAI22_X1 port map( A1 => n2743, A2 => n163, B1 => n2740, B2 => n160,
                           ZN => n1392);
   U1407 : AOI221_X1 port map( B1 => n4090, B2 => n169, C1 => n2744, C2 => n166
                           , A => n1392, ZN => n1395);
   U1408 : OAI22_X1 port map( A1 => n2723, A2 => n173, B1 => n172, B2 => n399, 
                           ZN => n1393);
   U1409 : AOI221_X1 port map( B1 => n2745, B2 => n181, C1 => n178, C2 => n1645
                           , A => n1393, ZN => n1394);
   U1410 : NAND4_X1 port map( A1 => n1397, A2 => n1396, A3 => n1395, A4 => 
                           n1394, ZN => n3018);
   U1411 : MUX2_X1 port map( A => n1398, B => DATAIN(28), S => n184, Z => n4474
                           );
   U1412 : OAI211_X1 port map( C1 => n2709, C2 => n127, A => n2289, B => n2288,
                           ZN => n1399);
   U1413 : AOI221_X1 port map( B1 => n307, B2 => n1872, C1 => n4059, C2 => n316
                           , A => n1399, ZN => n1402);
   U1414 : NOR2_X1 port map( A1 => n4096, A2 => n130, ZN => n1400);
   U1415 : NOR4_X1 port map( A1 => n2295, A2 => n2292, A3 => n2286, A4 => n1400
                           , ZN => n1401);
   U1416 : NAND2_X1 port map( A1 => n1402, A2 => n1401, ZN => n1406);
   U1417 : OAI22_X1 port map( A1 => n136, A2 => n1404, B1 => n133, B2 => n1403,
                           ZN => n1405);
   U1418 : AOI221_X1 port map( B1 => n142, B2 => n1406, C1 => n139, C2 => n1548
                           , A => n1405, ZN => n1413);
   U1419 : OAI22_X1 port map( A1 => n4027, A2 => n151, B1 => n3995, B2 => n148,
                           ZN => n1407);
   U1420 : AOI221_X1 port map( B1 => n157, B2 => n1516, C1 => n2714, C2 => n154
                           , A => n1407, ZN => n1412);
   U1421 : OAI22_X1 port map( A1 => n2720, A2 => n163, B1 => n2717, B2 => n160,
                           ZN => n1408);
   U1422 : AOI221_X1 port map( B1 => n4091, B2 => n169, C1 => n2721, C2 => n166
                           , A => n1408, ZN => n1411);
   U1423 : OAI22_X1 port map( A1 => n2700, A2 => n173, B1 => n172, B2 => n400, 
                           ZN => n1409);
   U1424 : AOI221_X1 port map( B1 => n2722, B2 => n181, C1 => n178, C2 => n1646
                           , A => n1409, ZN => n1410);
   U1425 : NAND4_X1 port map( A1 => n1413, A2 => n1412, A3 => n1411, A4 => 
                           n1410, ZN => n3017);
   U1426 : MUX2_X1 port map( A => n1414, B => DATAIN(29), S => n184, Z => n4475
                           );
   U1427 : OAI211_X1 port map( C1 => n2686, C2 => n127, A => n2301, B => n2300,
                           ZN => n1415);
   U1428 : AOI221_X1 port map( B1 => n307, B2 => n1873, C1 => n4060, C2 => n316
                           , A => n1415, ZN => n1418);
   U1429 : NOR2_X1 port map( A1 => n4095, A2 => n130, ZN => n1416);
   U1430 : NOR4_X1 port map( A1 => n2307, A2 => n2304, A3 => n2298, A4 => n1416
                           , ZN => n1417);
   U1431 : NAND2_X1 port map( A1 => n1418, A2 => n1417, ZN => n1422);
   U1432 : OAI22_X1 port map( A1 => n136, A2 => n1420, B1 => n133, B2 => n1419,
                           ZN => n1421);
   U1433 : AOI221_X1 port map( B1 => n142, B2 => n1422, C1 => n139, C2 => n1549
                           , A => n1421, ZN => n1429);
   U1434 : OAI22_X1 port map( A1 => n4028, A2 => n151, B1 => n3996, B2 => n148,
                           ZN => n1423);
   U1435 : AOI221_X1 port map( B1 => n157, B2 => n1517, C1 => n2691, C2 => n154
                           , A => n1423, ZN => n1428);
   U1436 : OAI22_X1 port map( A1 => n2697, A2 => n163, B1 => n2694, B2 => n160,
                           ZN => n1424);
   U1437 : AOI221_X1 port map( B1 => n4092, B2 => n169, C1 => n2698, C2 => n166
                           , A => n1424, ZN => n1427);
   U1438 : OAI22_X1 port map( A1 => n2677, A2 => n173, B1 => n172, B2 => n401, 
                           ZN => n1425);
   U1439 : AOI221_X1 port map( B1 => n2699, B2 => n181, C1 => n178, C2 => n1647
                           , A => n1425, ZN => n1426);
   U1440 : NAND4_X1 port map( A1 => n1429, A2 => n1428, A3 => n1427, A4 => 
                           n1426, ZN => n3016);
   U1441 : MUX2_X1 port map( A => n1430, B => DATAIN(30), S => n184, Z => n4476
                           );
   U1442 : OAI211_X1 port map( C1 => n2663, C2 => n127, A => n2324, B => n2323,
                           ZN => n1431);
   U1443 : AOI221_X1 port map( B1 => n307, B2 => n1874, C1 => n316, C2 => n4061
                           , A => n1431, ZN => n1434);
   U1444 : NOR2_X1 port map( A1 => n4094, A2 => n130, ZN => n1432);
   U1445 : NOR4_X1 port map( A1 => n2336, A2 => n2329, A3 => n2319, A4 => n1432
                           , ZN => n1433);
   U1446 : NAND2_X1 port map( A1 => n1434, A2 => n1433, ZN => n1440);
   U1447 : OAI22_X1 port map( A1 => n136, A2 => n1437, B1 => n133, B2 => n1435,
                           ZN => n1439);
   U1448 : AOI221_X1 port map( B1 => n144, B2 => n1440, C1 => n139, C2 => n1550
                           , A => n1439, ZN => n1453);
   U1449 : OAI22_X1 port map( A1 => n4029, A2 => n151, B1 => n3997, B2 => n148,
                           ZN => n1444);
   U1450 : AOI221_X1 port map( B1 => n157, B2 => n1518, C1 => n2668, C2 => n154
                           , A => n1444, ZN => n1452);
   U1451 : OAI22_X1 port map( A1 => n2674, A2 => n163, B1 => n2671, B2 => n160,
                           ZN => n1447);
   U1452 : AOI221_X1 port map( B1 => n4093, B2 => n169, C1 => n2675, C2 => n166
                           , A => n1447, ZN => n1451);
   U1453 : OAI22_X1 port map( A1 => n2654, A2 => n174, B1 => n172, B2 => n402, 
                           ZN => n1449);
   U1454 : AOI221_X1 port map( B1 => n2676, B2 => n181, C1 => n178, C2 => n1648
                           , A => n1449, ZN => n1450);
   U1455 : NAND4_X1 port map( A1 => n1453, A2 => n1452, A3 => n1451, A4 => 
                           n1450, ZN => n3015);
   U1456 : MUX2_X1 port map( A => n1454, B => DATAIN(31), S => n184, Z => n4477
                           );
   U1457 : MUX2_X1 port map( A => n1455, B => DATAIN(0), S => n185, Z => n4414)
                           ;
   U1458 : MUX2_X1 port map( A => n1456, B => DATAIN(1), S => n185, Z => n4415)
                           ;
   U1459 : MUX2_X1 port map( A => n1457, B => DATAIN(2), S => n185, Z => n4416)
                           ;
   U1460 : MUX2_X1 port map( A => n1458, B => DATAIN(3), S => n185, Z => n4417)
                           ;
   U1461 : MUX2_X1 port map( A => n1459, B => DATAIN(4), S => n185, Z => n4418)
                           ;
   U1462 : MUX2_X1 port map( A => n1460, B => DATAIN(5), S => n185, Z => n4419)
                           ;
   U1463 : MUX2_X1 port map( A => n1461, B => DATAIN(6), S => n185, Z => n4420)
                           ;
   U1464 : MUX2_X1 port map( A => n1462, B => DATAIN(7), S => n185, Z => n4421)
                           ;
   U1465 : MUX2_X1 port map( A => n1463, B => DATAIN(8), S => n185, Z => n4422)
                           ;
   U1466 : MUX2_X1 port map( A => n1464, B => DATAIN(9), S => n185, Z => n4423)
                           ;
   U1467 : MUX2_X1 port map( A => n1465, B => DATAIN(10), S => n185, Z => n4424
                           );
   U1468 : MUX2_X1 port map( A => n1466, B => DATAIN(11), S => n185, Z => n4425
                           );
   U1469 : MUX2_X1 port map( A => n1467, B => DATAIN(12), S => n186, Z => n4426
                           );
   U1470 : MUX2_X1 port map( A => n1468, B => DATAIN(13), S => n186, Z => n4427
                           );
   U1471 : MUX2_X1 port map( A => n1469, B => DATAIN(14), S => n186, Z => n4428
                           );
   U1472 : MUX2_X1 port map( A => n1470, B => DATAIN(15), S => n186, Z => n4429
                           );
   U1473 : MUX2_X1 port map( A => n1471, B => DATAIN(16), S => n186, Z => n4430
                           );
   U1474 : MUX2_X1 port map( A => n1472, B => DATAIN(17), S => n186, Z => n4431
                           );
   U1475 : MUX2_X1 port map( A => n1473, B => DATAIN(18), S => n186, Z => n4432
                           );
   U1476 : MUX2_X1 port map( A => n1474, B => DATAIN(19), S => n186, Z => n4433
                           );
   U1477 : MUX2_X1 port map( A => n1475, B => DATAIN(20), S => n186, Z => n4434
                           );
   U1478 : MUX2_X1 port map( A => n1476, B => DATAIN(21), S => n186, Z => n4435
                           );
   U1479 : MUX2_X1 port map( A => n1477, B => DATAIN(22), S => n186, Z => n4436
                           );
   U1480 : MUX2_X1 port map( A => n1478, B => DATAIN(23), S => n186, Z => n4437
                           );
   U1481 : MUX2_X1 port map( A => n1479, B => DATAIN(24), S => n187, Z => n4438
                           );
   U1482 : MUX2_X1 port map( A => n1480, B => DATAIN(25), S => n187, Z => n4439
                           );
   U1483 : MUX2_X1 port map( A => n1481, B => DATAIN(26), S => n187, Z => n4440
                           );
   U1484 : MUX2_X1 port map( A => n1482, B => DATAIN(27), S => n187, Z => n4441
                           );
   U1485 : MUX2_X1 port map( A => n1483, B => DATAIN(28), S => n187, Z => n4442
                           );
   U1486 : MUX2_X1 port map( A => n1484, B => DATAIN(29), S => n187, Z => n4443
                           );
   U1487 : MUX2_X1 port map( A => n1485, B => DATAIN(30), S => n187, Z => n4444
                           );
   U1488 : MUX2_X1 port map( A => n1486, B => DATAIN(31), S => n187, Z => n4445
                           );
   U1489 : INV_X1 port map( A => ADD_WR(1), ZN => n1552);
   U1490 : MUX2_X1 port map( A => n4030, B => DATAIN(0), S => n188, Z => n3047)
                           ;
   U1491 : MUX2_X1 port map( A => n4031, B => DATAIN(1), S => n188, Z => n3048)
                           ;
   U1492 : MUX2_X1 port map( A => n4032, B => DATAIN(2), S => n188, Z => n3049)
                           ;
   U1493 : MUX2_X1 port map( A => n4033, B => DATAIN(3), S => n188, Z => n3050)
                           ;
   U1494 : MUX2_X1 port map( A => n4034, B => DATAIN(4), S => n188, Z => n3051)
                           ;
   U1495 : MUX2_X1 port map( A => n4035, B => DATAIN(5), S => n188, Z => n3052)
                           ;
   U1496 : MUX2_X1 port map( A => n4036, B => DATAIN(6), S => n188, Z => n3053)
                           ;
   U1497 : MUX2_X1 port map( A => n4037, B => DATAIN(7), S => n188, Z => n3054)
                           ;
   U1498 : MUX2_X1 port map( A => n4038, B => DATAIN(8), S => n188, Z => n3055)
                           ;
   U1499 : MUX2_X1 port map( A => n4039, B => DATAIN(9), S => n188, Z => n3056)
                           ;
   U1500 : MUX2_X1 port map( A => n4040, B => DATAIN(10), S => n188, Z => n3057
                           );
   U1501 : MUX2_X1 port map( A => n4041, B => DATAIN(11), S => n188, Z => n3058
                           );
   U1502 : MUX2_X1 port map( A => n4042, B => DATAIN(12), S => n189, Z => n3059
                           );
   U1503 : MUX2_X1 port map( A => n4043, B => DATAIN(13), S => n189, Z => n3060
                           );
   U1504 : MUX2_X1 port map( A => n4044, B => DATAIN(14), S => n189, Z => n3061
                           );
   U1505 : MUX2_X1 port map( A => n4045, B => DATAIN(15), S => n189, Z => n3062
                           );
   U1506 : MUX2_X1 port map( A => n4046, B => DATAIN(16), S => n189, Z => n3063
                           );
   U1507 : MUX2_X1 port map( A => n4047, B => DATAIN(17), S => n189, Z => n3064
                           );
   U1508 : MUX2_X1 port map( A => n4048, B => DATAIN(18), S => n189, Z => n3065
                           );
   U1509 : MUX2_X1 port map( A => n4049, B => DATAIN(19), S => n189, Z => n3066
                           );
   U1510 : MUX2_X1 port map( A => n4050, B => DATAIN(20), S => n189, Z => n3067
                           );
   U1511 : MUX2_X1 port map( A => n4051, B => DATAIN(21), S => n189, Z => n3068
                           );
   U1512 : MUX2_X1 port map( A => n4052, B => DATAIN(22), S => n189, Z => n3069
                           );
   U1513 : MUX2_X1 port map( A => n4053, B => DATAIN(23), S => n189, Z => n3070
                           );
   U1514 : MUX2_X1 port map( A => n4054, B => DATAIN(24), S => n190, Z => n3071
                           );
   U1515 : MUX2_X1 port map( A => n4055, B => DATAIN(25), S => n190, Z => n3072
                           );
   U1516 : MUX2_X1 port map( A => n4056, B => DATAIN(26), S => n190, Z => n3073
                           );
   U1517 : MUX2_X1 port map( A => n4057, B => DATAIN(27), S => n190, Z => n3074
                           );
   U1518 : MUX2_X1 port map( A => n4058, B => DATAIN(28), S => n190, Z => n3075
                           );
   U1519 : MUX2_X1 port map( A => n4059, B => DATAIN(29), S => n190, Z => n3076
                           );
   U1520 : MUX2_X1 port map( A => n4060, B => DATAIN(30), S => n190, Z => n3077
                           );
   U1521 : MUX2_X1 port map( A => n4061, B => DATAIN(31), S => n190, Z => n3078
                           );
   U1522 : MUX2_X1 port map( A => n4062, B => DATAIN(0), S => n191, Z => n3079)
                           ;
   U1523 : MUX2_X1 port map( A => n4063, B => DATAIN(1), S => n191, Z => n3080)
                           ;
   U1524 : MUX2_X1 port map( A => n4064, B => DATAIN(2), S => n191, Z => n3081)
                           ;
   U1525 : MUX2_X1 port map( A => n4065, B => DATAIN(3), S => n191, Z => n3082)
                           ;
   U1526 : MUX2_X1 port map( A => n4066, B => DATAIN(4), S => n191, Z => n3083)
                           ;
   U1527 : MUX2_X1 port map( A => n4067, B => DATAIN(5), S => n191, Z => n3084)
                           ;
   U1528 : MUX2_X1 port map( A => n4068, B => DATAIN(6), S => n191, Z => n3085)
                           ;
   U1529 : MUX2_X1 port map( A => n4069, B => DATAIN(7), S => n191, Z => n3086)
                           ;
   U1530 : MUX2_X1 port map( A => n4070, B => DATAIN(8), S => n191, Z => n3087)
                           ;
   U1531 : MUX2_X1 port map( A => n4071, B => DATAIN(9), S => n191, Z => n3088)
                           ;
   U1532 : MUX2_X1 port map( A => n4072, B => DATAIN(10), S => n191, Z => n3089
                           );
   U1533 : MUX2_X1 port map( A => n4073, B => DATAIN(11), S => n191, Z => n3090
                           );
   U1534 : MUX2_X1 port map( A => n4074, B => DATAIN(12), S => n192, Z => n3091
                           );
   U1535 : MUX2_X1 port map( A => n4075, B => DATAIN(13), S => n192, Z => n3092
                           );
   U1536 : MUX2_X1 port map( A => n4076, B => DATAIN(14), S => n192, Z => n3093
                           );
   U1537 : MUX2_X1 port map( A => n4077, B => DATAIN(15), S => n192, Z => n3094
                           );
   U1538 : MUX2_X1 port map( A => n4078, B => DATAIN(16), S => n192, Z => n3095
                           );
   U1539 : MUX2_X1 port map( A => n4079, B => DATAIN(17), S => n192, Z => n3096
                           );
   U1540 : MUX2_X1 port map( A => n4080, B => DATAIN(18), S => n192, Z => n3097
                           );
   U1541 : MUX2_X1 port map( A => n4081, B => DATAIN(19), S => n192, Z => n3098
                           );
   U1542 : MUX2_X1 port map( A => n4082, B => DATAIN(20), S => n192, Z => n3099
                           );
   U1543 : MUX2_X1 port map( A => n4083, B => DATAIN(21), S => n192, Z => n3100
                           );
   U1544 : MUX2_X1 port map( A => n4084, B => DATAIN(22), S => n192, Z => n3101
                           );
   U1545 : MUX2_X1 port map( A => n4085, B => DATAIN(23), S => n192, Z => n3102
                           );
   U1546 : MUX2_X1 port map( A => n4086, B => DATAIN(24), S => n193, Z => n3103
                           );
   U1547 : MUX2_X1 port map( A => n4087, B => DATAIN(25), S => n193, Z => n3104
                           );
   U1548 : MUX2_X1 port map( A => n4088, B => DATAIN(26), S => n193, Z => n3105
                           );
   U1549 : MUX2_X1 port map( A => n4089, B => DATAIN(27), S => n193, Z => n3106
                           );
   U1550 : MUX2_X1 port map( A => n4090, B => DATAIN(28), S => n193, Z => n3107
                           );
   U1551 : MUX2_X1 port map( A => n4091, B => DATAIN(29), S => n193, Z => n3108
                           );
   U1552 : MUX2_X1 port map( A => n4092, B => DATAIN(30), S => n193, Z => n3109
                           );
   U1553 : MUX2_X1 port map( A => n4093, B => DATAIN(31), S => n193, Z => n3110
                           );
   U1554 : INV_X1 port map( A => ADD_WR(2), ZN => n1551);
   U1555 : MUX2_X1 port map( A => n1487, B => DATAIN(0), S => n194, Z => n4382)
                           ;
   U1556 : MUX2_X1 port map( A => n1488, B => DATAIN(1), S => n194, Z => n4383)
                           ;
   U1557 : MUX2_X1 port map( A => n1489, B => DATAIN(2), S => n194, Z => n4384)
                           ;
   U1558 : MUX2_X1 port map( A => n1490, B => DATAIN(3), S => n194, Z => n4385)
                           ;
   U1559 : MUX2_X1 port map( A => n1491, B => DATAIN(4), S => n194, Z => n4386)
                           ;
   U1560 : MUX2_X1 port map( A => n1492, B => DATAIN(5), S => n194, Z => n4387)
                           ;
   U1561 : MUX2_X1 port map( A => n1493, B => DATAIN(6), S => n194, Z => n4388)
                           ;
   U1562 : MUX2_X1 port map( A => n1494, B => DATAIN(7), S => n194, Z => n4389)
                           ;
   U1563 : MUX2_X1 port map( A => n1495, B => DATAIN(8), S => n194, Z => n4390)
                           ;
   U1564 : MUX2_X1 port map( A => n1496, B => DATAIN(9), S => n194, Z => n4391)
                           ;
   U1565 : MUX2_X1 port map( A => n1497, B => DATAIN(10), S => n194, Z => n4392
                           );
   U1566 : MUX2_X1 port map( A => n1498, B => DATAIN(11), S => n194, Z => n4393
                           );
   U1567 : MUX2_X1 port map( A => n1499, B => DATAIN(12), S => n195, Z => n4394
                           );
   U1568 : MUX2_X1 port map( A => n1500, B => DATAIN(13), S => n195, Z => n4395
                           );
   U1569 : MUX2_X1 port map( A => n1501, B => DATAIN(14), S => n195, Z => n4396
                           );
   U1570 : MUX2_X1 port map( A => n1502, B => DATAIN(15), S => n195, Z => n4397
                           );
   U1571 : MUX2_X1 port map( A => n1503, B => DATAIN(16), S => n195, Z => n4398
                           );
   U1572 : MUX2_X1 port map( A => n1504, B => DATAIN(17), S => n195, Z => n4399
                           );
   U1573 : MUX2_X1 port map( A => n1505, B => DATAIN(18), S => n195, Z => n4400
                           );
   U1574 : MUX2_X1 port map( A => n1506, B => DATAIN(19), S => n195, Z => n4401
                           );
   U1575 : MUX2_X1 port map( A => n1507, B => DATAIN(20), S => n195, Z => n4402
                           );
   U1576 : MUX2_X1 port map( A => n1508, B => DATAIN(21), S => n195, Z => n4403
                           );
   U1577 : MUX2_X1 port map( A => n1509, B => DATAIN(22), S => n195, Z => n4404
                           );
   U1578 : MUX2_X1 port map( A => n1510, B => DATAIN(23), S => n195, Z => n4405
                           );
   U1579 : MUX2_X1 port map( A => n1511, B => DATAIN(24), S => n196, Z => n4406
                           );
   U1580 : MUX2_X1 port map( A => n1512, B => DATAIN(25), S => n196, Z => n4407
                           );
   U1581 : MUX2_X1 port map( A => n1513, B => DATAIN(26), S => n196, Z => n4408
                           );
   U1582 : MUX2_X1 port map( A => n1514, B => DATAIN(27), S => n196, Z => n4409
                           );
   U1583 : MUX2_X1 port map( A => n1515, B => DATAIN(28), S => n196, Z => n4410
                           );
   U1584 : MUX2_X1 port map( A => n1516, B => DATAIN(29), S => n196, Z => n4411
                           );
   U1585 : MUX2_X1 port map( A => n1517, B => DATAIN(30), S => n196, Z => n4412
                           );
   U1586 : MUX2_X1 port map( A => n1518, B => DATAIN(31), S => n196, Z => n4413
                           );
   U1587 : MUX2_X1 port map( A => n1519, B => DATAIN(0), S => n197, Z => n4351)
                           ;
   U1588 : MUX2_X1 port map( A => n1520, B => DATAIN(1), S => n197, Z => n4352)
                           ;
   U1589 : MUX2_X1 port map( A => n1521, B => DATAIN(2), S => n197, Z => n4353)
                           ;
   U1590 : MUX2_X1 port map( A => n1522, B => DATAIN(3), S => n197, Z => n4354)
                           ;
   U1591 : MUX2_X1 port map( A => n1523, B => DATAIN(4), S => n197, Z => n4355)
                           ;
   U1592 : MUX2_X1 port map( A => n1524, B => DATAIN(5), S => n197, Z => n4356)
                           ;
   U1593 : MUX2_X1 port map( A => n1525, B => DATAIN(6), S => n197, Z => n4357)
                           ;
   U1594 : MUX2_X1 port map( A => n1526, B => DATAIN(7), S => n197, Z => n4358)
                           ;
   U1595 : MUX2_X1 port map( A => n1527, B => DATAIN(8), S => n197, Z => n4359)
                           ;
   U1596 : MUX2_X1 port map( A => n1528, B => DATAIN(9), S => n197, Z => n4360)
                           ;
   U1597 : MUX2_X1 port map( A => n1529, B => DATAIN(10), S => n197, Z => n4361
                           );
   U1598 : MUX2_X1 port map( A => n1530, B => DATAIN(11), S => n197, Z => n4362
                           );
   U1599 : MUX2_X1 port map( A => n1531, B => DATAIN(12), S => n198, Z => n4363
                           );
   U1600 : MUX2_X1 port map( A => n1532, B => DATAIN(13), S => n198, Z => n4364
                           );
   U1601 : MUX2_X1 port map( A => n1533, B => DATAIN(14), S => n198, Z => n4365
                           );
   U1602 : MUX2_X1 port map( A => n1534, B => DATAIN(15), S => n198, Z => n4366
                           );
   U1603 : MUX2_X1 port map( A => n1535, B => DATAIN(16), S => n198, Z => n4367
                           );
   U1604 : MUX2_X1 port map( A => n1536, B => DATAIN(17), S => n198, Z => n4368
                           );
   U1605 : MUX2_X1 port map( A => n1537, B => DATAIN(18), S => n198, Z => n4369
                           );
   U1606 : MUX2_X1 port map( A => n1538, B => DATAIN(19), S => n198, Z => n4370
                           );
   U1607 : MUX2_X1 port map( A => n1539, B => DATAIN(20), S => n198, Z => n4371
                           );
   U1608 : MUX2_X1 port map( A => n1540, B => DATAIN(21), S => n198, Z => n4372
                           );
   U1609 : MUX2_X1 port map( A => n1541, B => DATAIN(22), S => n198, Z => n4373
                           );
   U1610 : MUX2_X1 port map( A => n1542, B => DATAIN(23), S => n198, Z => n4374
                           );
   U1611 : MUX2_X1 port map( A => n1543, B => DATAIN(24), S => n199, Z => n4375
                           );
   U1612 : MUX2_X1 port map( A => n1544, B => DATAIN(25), S => n199, Z => n4376
                           );
   U1613 : MUX2_X1 port map( A => n1545, B => DATAIN(26), S => n199, Z => n4377
                           );
   U1614 : MUX2_X1 port map( A => n1546, B => DATAIN(27), S => n199, Z => n4378
                           );
   U1615 : MUX2_X1 port map( A => n1547, B => DATAIN(28), S => n199, Z => n4379
                           );
   U1616 : MUX2_X1 port map( A => n1548, B => DATAIN(29), S => n199, Z => n4380
                           );
   U1617 : MUX2_X1 port map( A => n1549, B => DATAIN(30), S => n199, Z => n4381
                           );
   U1618 : MUX2_X1 port map( A => n1550, B => DATAIN(31), S => n199, Z => n4350
                           );
   U1619 : MUX2_X1 port map( A => n3957, B => DATAIN(0), S => n200, Z => n3111)
                           ;
   U1620 : MUX2_X1 port map( A => n3934, B => DATAIN(1), S => n200, Z => n3112)
                           ;
   U1621 : MUX2_X1 port map( A => n3911, B => DATAIN(2), S => n200, Z => n3113)
                           ;
   U1622 : MUX2_X1 port map( A => n3888, B => DATAIN(3), S => n200, Z => n3114)
                           ;
   U1623 : MUX2_X1 port map( A => n3865, B => DATAIN(4), S => n200, Z => n3115)
                           ;
   U1624 : MUX2_X1 port map( A => n3842, B => DATAIN(5), S => n200, Z => n3116)
                           ;
   U1625 : MUX2_X1 port map( A => n3819, B => DATAIN(6), S => n200, Z => n3117)
                           ;
   U1626 : MUX2_X1 port map( A => n3796, B => DATAIN(7), S => n200, Z => n3118)
                           ;
   U1627 : MUX2_X1 port map( A => n3773, B => DATAIN(8), S => n200, Z => n3119)
                           ;
   U1628 : MUX2_X1 port map( A => n3750, B => DATAIN(9), S => n200, Z => n3120)
                           ;
   U1629 : MUX2_X1 port map( A => n3727, B => DATAIN(10), S => n200, Z => n3121
                           );
   U1630 : MUX2_X1 port map( A => n3704, B => DATAIN(11), S => n200, Z => n3122
                           );
   U1631 : MUX2_X1 port map( A => n3681, B => DATAIN(12), S => n201, Z => n3123
                           );
   U1632 : MUX2_X1 port map( A => n3658, B => DATAIN(13), S => n201, Z => n3124
                           );
   U1633 : MUX2_X1 port map( A => n3635, B => DATAIN(14), S => n201, Z => n3125
                           );
   U1634 : MUX2_X1 port map( A => n3612, B => DATAIN(15), S => n201, Z => n3126
                           );
   U1635 : MUX2_X1 port map( A => n3589, B => DATAIN(16), S => n201, Z => n3127
                           );
   U1636 : MUX2_X1 port map( A => n3566, B => DATAIN(17), S => n201, Z => n3128
                           );
   U1637 : MUX2_X1 port map( A => n2967, B => DATAIN(18), S => n201, Z => n3129
                           );
   U1638 : MUX2_X1 port map( A => n2944, B => DATAIN(19), S => n201, Z => n3130
                           );
   U1639 : MUX2_X1 port map( A => n2921, B => DATAIN(20), S => n201, Z => n3131
                           );
   U1640 : MUX2_X1 port map( A => n2898, B => DATAIN(21), S => n201, Z => n3132
                           );
   U1641 : MUX2_X1 port map( A => n2875, B => DATAIN(22), S => n201, Z => n3133
                           );
   U1642 : MUX2_X1 port map( A => n2852, B => DATAIN(23), S => n201, Z => n3134
                           );
   U1643 : MUX2_X1 port map( A => n2829, B => DATAIN(24), S => n202, Z => n3135
                           );
   U1644 : MUX2_X1 port map( A => n2806, B => DATAIN(25), S => n202, Z => n3136
                           );
   U1645 : MUX2_X1 port map( A => n2783, B => DATAIN(26), S => n202, Z => n3137
                           );
   U1646 : MUX2_X1 port map( A => n2760, B => DATAIN(27), S => n202, Z => n3138
                           );
   U1647 : MUX2_X1 port map( A => n2737, B => DATAIN(28), S => n202, Z => n3139
                           );
   U1648 : MUX2_X1 port map( A => n2714, B => DATAIN(29), S => n202, Z => n3140
                           );
   U1649 : MUX2_X1 port map( A => n2691, B => DATAIN(30), S => n202, Z => n3141
                           );
   U1650 : MUX2_X1 port map( A => n2668, B => DATAIN(31), S => n202, Z => n3142
                           );
   U1651 : MUX2_X1 port map( A => n3958, B => DATAIN(0), S => n203, Z => n3143)
                           ;
   U1652 : MUX2_X1 port map( A => n3935, B => DATAIN(1), S => n203, Z => n3144)
                           ;
   U1653 : MUX2_X1 port map( A => n3912, B => DATAIN(2), S => n203, Z => n3145)
                           ;
   U1654 : MUX2_X1 port map( A => n3889, B => DATAIN(3), S => n203, Z => n3146)
                           ;
   U1655 : MUX2_X1 port map( A => n3866, B => DATAIN(4), S => n203, Z => n3147)
                           ;
   U1656 : MUX2_X1 port map( A => n3843, B => DATAIN(5), S => n203, Z => n3148)
                           ;
   U1657 : MUX2_X1 port map( A => n3820, B => DATAIN(6), S => n203, Z => n3149)
                           ;
   U1658 : MUX2_X1 port map( A => n3797, B => DATAIN(7), S => n203, Z => n3150)
                           ;
   U1659 : MUX2_X1 port map( A => n3774, B => DATAIN(8), S => n203, Z => n3151)
                           ;
   U1660 : MUX2_X1 port map( A => n3751, B => DATAIN(9), S => n203, Z => n3152)
                           ;
   U1661 : MUX2_X1 port map( A => n3728, B => DATAIN(10), S => n203, Z => n3153
                           );
   U1662 : MUX2_X1 port map( A => n3705, B => DATAIN(11), S => n203, Z => n3154
                           );
   U1663 : MUX2_X1 port map( A => n3682, B => DATAIN(12), S => n204, Z => n3155
                           );
   U1664 : MUX2_X1 port map( A => n3659, B => DATAIN(13), S => n204, Z => n3156
                           );
   U1665 : MUX2_X1 port map( A => n3636, B => DATAIN(14), S => n204, Z => n3157
                           );
   U1666 : MUX2_X1 port map( A => n3613, B => DATAIN(15), S => n204, Z => n3158
                           );
   U1667 : MUX2_X1 port map( A => n3590, B => DATAIN(16), S => n204, Z => n3159
                           );
   U1668 : MUX2_X1 port map( A => n3567, B => DATAIN(17), S => n204, Z => n3160
                           );
   U1669 : MUX2_X1 port map( A => n2968, B => DATAIN(18), S => n204, Z => n3161
                           );
   U1670 : MUX2_X1 port map( A => n2945, B => DATAIN(19), S => n204, Z => n3162
                           );
   U1671 : MUX2_X1 port map( A => n2922, B => DATAIN(20), S => n204, Z => n3163
                           );
   U1672 : MUX2_X1 port map( A => n2899, B => DATAIN(21), S => n204, Z => n3164
                           );
   U1673 : MUX2_X1 port map( A => n2876, B => DATAIN(22), S => n204, Z => n3165
                           );
   U1674 : MUX2_X1 port map( A => n2853, B => DATAIN(23), S => n204, Z => n3166
                           );
   U1675 : MUX2_X1 port map( A => n2830, B => DATAIN(24), S => n205, Z => n3167
                           );
   U1676 : MUX2_X1 port map( A => n2807, B => DATAIN(25), S => n205, Z => n3168
                           );
   U1677 : MUX2_X1 port map( A => n2784, B => DATAIN(26), S => n205, Z => n3169
                           );
   U1678 : MUX2_X1 port map( A => n2761, B => DATAIN(27), S => n205, Z => n3170
                           );
   U1679 : MUX2_X1 port map( A => n2738, B => DATAIN(28), S => n205, Z => n3171
                           );
   U1680 : MUX2_X1 port map( A => n2715, B => DATAIN(29), S => n205, Z => n3172
                           );
   U1681 : MUX2_X1 port map( A => n2692, B => DATAIN(30), S => n205, Z => n3173
                           );
   U1682 : MUX2_X1 port map( A => n2669, B => DATAIN(31), S => n205, Z => n3174
                           );
   U1683 : INV_X1 port map( A => ADD_WR(3), ZN => n1810);
   U1684 : MUX2_X1 port map( A => n3961, B => DATAIN(0), S => n206, Z => n3175)
                           ;
   U1685 : MUX2_X1 port map( A => n3938, B => DATAIN(1), S => n206, Z => n3176)
                           ;
   U1686 : MUX2_X1 port map( A => n3915, B => DATAIN(2), S => n206, Z => n3177)
                           ;
   U1687 : MUX2_X1 port map( A => n3892, B => DATAIN(3), S => n206, Z => n3178)
                           ;
   U1688 : MUX2_X1 port map( A => n3869, B => DATAIN(4), S => n206, Z => n3179)
                           ;
   U1689 : MUX2_X1 port map( A => n3846, B => DATAIN(5), S => n206, Z => n3180)
                           ;
   U1690 : MUX2_X1 port map( A => n3823, B => DATAIN(6), S => n206, Z => n3181)
                           ;
   U1691 : MUX2_X1 port map( A => n3800, B => DATAIN(7), S => n206, Z => n3182)
                           ;
   U1692 : MUX2_X1 port map( A => n3777, B => DATAIN(8), S => n206, Z => n3183)
                           ;
   U1693 : MUX2_X1 port map( A => n3754, B => DATAIN(9), S => n206, Z => n3184)
                           ;
   U1694 : MUX2_X1 port map( A => n3731, B => DATAIN(10), S => n206, Z => n3185
                           );
   U1695 : MUX2_X1 port map( A => n3708, B => DATAIN(11), S => n206, Z => n3186
                           );
   U1696 : MUX2_X1 port map( A => n3685, B => DATAIN(12), S => n207, Z => n3187
                           );
   U1697 : MUX2_X1 port map( A => n3662, B => DATAIN(13), S => n207, Z => n3188
                           );
   U1698 : MUX2_X1 port map( A => n3639, B => DATAIN(14), S => n207, Z => n3189
                           );
   U1699 : MUX2_X1 port map( A => n3616, B => DATAIN(15), S => n207, Z => n3190
                           );
   U1700 : MUX2_X1 port map( A => n3593, B => DATAIN(16), S => n207, Z => n3191
                           );
   U1701 : MUX2_X1 port map( A => n3570, B => DATAIN(17), S => n207, Z => n3192
                           );
   U1702 : MUX2_X1 port map( A => n2971, B => DATAIN(18), S => n207, Z => n3193
                           );
   U1703 : MUX2_X1 port map( A => n2948, B => DATAIN(19), S => n207, Z => n3194
                           );
   U1704 : MUX2_X1 port map( A => n2925, B => DATAIN(20), S => n207, Z => n3195
                           );
   U1705 : MUX2_X1 port map( A => n2902, B => DATAIN(21), S => n207, Z => n3196
                           );
   U1706 : MUX2_X1 port map( A => n2879, B => DATAIN(22), S => n207, Z => n3197
                           );
   U1707 : MUX2_X1 port map( A => n2856, B => DATAIN(23), S => n207, Z => n3198
                           );
   U1708 : MUX2_X1 port map( A => n2833, B => DATAIN(24), S => n208, Z => n3199
                           );
   U1709 : MUX2_X1 port map( A => n2810, B => DATAIN(25), S => n208, Z => n3200
                           );
   U1710 : MUX2_X1 port map( A => n2787, B => DATAIN(26), S => n208, Z => n3201
                           );
   U1711 : MUX2_X1 port map( A => n2764, B => DATAIN(27), S => n208, Z => n3202
                           );
   U1712 : MUX2_X1 port map( A => n2741, B => DATAIN(28), S => n208, Z => n3203
                           );
   U1713 : MUX2_X1 port map( A => n2718, B => DATAIN(29), S => n208, Z => n3204
                           );
   U1714 : MUX2_X1 port map( A => n2695, B => DATAIN(30), S => n208, Z => n3205
                           );
   U1715 : MUX2_X1 port map( A => n2672, B => DATAIN(31), S => n208, Z => n3206
                           );
   U1716 : MUX2_X1 port map( A => n3962, B => DATAIN(0), S => n209, Z => n3207)
                           ;
   U1717 : MUX2_X1 port map( A => n3939, B => DATAIN(1), S => n209, Z => n3208)
                           ;
   U1718 : MUX2_X1 port map( A => n3916, B => DATAIN(2), S => n209, Z => n3209)
                           ;
   U1719 : MUX2_X1 port map( A => n3893, B => DATAIN(3), S => n209, Z => n3210)
                           ;
   U1720 : MUX2_X1 port map( A => n3870, B => DATAIN(4), S => n209, Z => n3211)
                           ;
   U1721 : MUX2_X1 port map( A => n3847, B => DATAIN(5), S => n209, Z => n3212)
                           ;
   U1722 : MUX2_X1 port map( A => n3824, B => DATAIN(6), S => n209, Z => n3213)
                           ;
   U1723 : MUX2_X1 port map( A => n3801, B => DATAIN(7), S => n209, Z => n3214)
                           ;
   U1724 : MUX2_X1 port map( A => n3778, B => DATAIN(8), S => n209, Z => n3215)
                           ;
   U1725 : MUX2_X1 port map( A => n3755, B => DATAIN(9), S => n209, Z => n3216)
                           ;
   U1726 : MUX2_X1 port map( A => n3732, B => DATAIN(10), S => n209, Z => n3217
                           );
   U1727 : MUX2_X1 port map( A => n3709, B => DATAIN(11), S => n209, Z => n3218
                           );
   U1728 : MUX2_X1 port map( A => n3686, B => DATAIN(12), S => n210, Z => n3219
                           );
   U1729 : MUX2_X1 port map( A => n3663, B => DATAIN(13), S => n210, Z => n3220
                           );
   U1730 : MUX2_X1 port map( A => n3640, B => DATAIN(14), S => n210, Z => n3221
                           );
   U1731 : MUX2_X1 port map( A => n3617, B => DATAIN(15), S => n210, Z => n3222
                           );
   U1732 : MUX2_X1 port map( A => n3594, B => DATAIN(16), S => n210, Z => n3223
                           );
   U1733 : MUX2_X1 port map( A => n3571, B => DATAIN(17), S => n210, Z => n3224
                           );
   U1734 : MUX2_X1 port map( A => n2972, B => DATAIN(18), S => n210, Z => n3225
                           );
   U1735 : MUX2_X1 port map( A => n2949, B => DATAIN(19), S => n210, Z => n3226
                           );
   U1736 : MUX2_X1 port map( A => n2926, B => DATAIN(20), S => n210, Z => n3227
                           );
   U1737 : MUX2_X1 port map( A => n2903, B => DATAIN(21), S => n210, Z => n3228
                           );
   U1738 : MUX2_X1 port map( A => n2880, B => DATAIN(22), S => n210, Z => n3229
                           );
   U1739 : MUX2_X1 port map( A => n2857, B => DATAIN(23), S => n210, Z => n3230
                           );
   U1740 : MUX2_X1 port map( A => n2834, B => DATAIN(24), S => n211, Z => n3231
                           );
   U1741 : MUX2_X1 port map( A => n2811, B => DATAIN(25), S => n211, Z => n3232
                           );
   U1742 : MUX2_X1 port map( A => n2788, B => DATAIN(26), S => n211, Z => n3233
                           );
   U1743 : MUX2_X1 port map( A => n2765, B => DATAIN(27), S => n211, Z => n3234
                           );
   U1744 : MUX2_X1 port map( A => n2742, B => DATAIN(28), S => n211, Z => n3235
                           );
   U1745 : MUX2_X1 port map( A => n2719, B => DATAIN(29), S => n211, Z => n3236
                           );
   U1746 : MUX2_X1 port map( A => n2696, B => DATAIN(30), S => n211, Z => n3237
                           );
   U1747 : MUX2_X1 port map( A => n2673, B => DATAIN(31), S => n211, Z => n3238
                           );
   U1748 : MUX2_X1 port map( A => n1553, B => DATAIN(0), S => n212, Z => n4574)
                           ;
   U1749 : MUX2_X1 port map( A => n1554, B => DATAIN(1), S => n212, Z => n4575)
                           ;
   U1750 : MUX2_X1 port map( A => n1555, B => DATAIN(2), S => n212, Z => n4576)
                           ;
   U1751 : MUX2_X1 port map( A => n1556, B => DATAIN(3), S => n212, Z => n4577)
                           ;
   U1752 : MUX2_X1 port map( A => n1557, B => DATAIN(4), S => n212, Z => n4578)
                           ;
   U1753 : MUX2_X1 port map( A => n1558, B => DATAIN(5), S => n212, Z => n4579)
                           ;
   U1754 : MUX2_X1 port map( A => n1559, B => DATAIN(6), S => n212, Z => n4580)
                           ;
   U1755 : MUX2_X1 port map( A => n1560, B => DATAIN(7), S => n212, Z => n4581)
                           ;
   U1756 : MUX2_X1 port map( A => n1561, B => DATAIN(8), S => n212, Z => n4582)
                           ;
   U1757 : MUX2_X1 port map( A => n1562, B => DATAIN(9), S => n212, Z => n4583)
                           ;
   U1758 : MUX2_X1 port map( A => n1563, B => DATAIN(10), S => n212, Z => n4584
                           );
   U1759 : MUX2_X1 port map( A => n1564, B => DATAIN(11), S => n212, Z => n4585
                           );
   U1760 : MUX2_X1 port map( A => n1565, B => DATAIN(12), S => n213, Z => n4586
                           );
   U1761 : MUX2_X1 port map( A => n1566, B => DATAIN(13), S => n213, Z => n4587
                           );
   U1762 : MUX2_X1 port map( A => n1567, B => DATAIN(14), S => n213, Z => n4588
                           );
   U1763 : MUX2_X1 port map( A => n1568, B => DATAIN(15), S => n213, Z => n4589
                           );
   U1764 : MUX2_X1 port map( A => n1569, B => DATAIN(16), S => n213, Z => n4590
                           );
   U1765 : MUX2_X1 port map( A => n1570, B => DATAIN(17), S => n213, Z => n4591
                           );
   U1766 : MUX2_X1 port map( A => n1571, B => DATAIN(18), S => n213, Z => n4592
                           );
   U1767 : MUX2_X1 port map( A => n1572, B => DATAIN(19), S => n213, Z => n4593
                           );
   U1768 : MUX2_X1 port map( A => n1573, B => DATAIN(20), S => n213, Z => n4594
                           );
   U1769 : MUX2_X1 port map( A => n1574, B => DATAIN(21), S => n213, Z => n4595
                           );
   U1770 : MUX2_X1 port map( A => n1575, B => DATAIN(22), S => n213, Z => n4596
                           );
   U1771 : MUX2_X1 port map( A => n1576, B => DATAIN(23), S => n213, Z => n4597
                           );
   U1772 : MUX2_X1 port map( A => n1577, B => DATAIN(24), S => n214, Z => n4598
                           );
   U1773 : MUX2_X1 port map( A => n1578, B => DATAIN(25), S => n214, Z => n4599
                           );
   U1774 : MUX2_X1 port map( A => n1579, B => DATAIN(26), S => n214, Z => n4600
                           );
   U1775 : MUX2_X1 port map( A => n1580, B => DATAIN(27), S => n214, Z => n4601
                           );
   U1776 : MUX2_X1 port map( A => n1581, B => DATAIN(28), S => n214, Z => n4602
                           );
   U1777 : MUX2_X1 port map( A => n1582, B => DATAIN(29), S => n214, Z => n4603
                           );
   U1778 : MUX2_X1 port map( A => n1583, B => DATAIN(30), S => n214, Z => n4604
                           );
   U1779 : MUX2_X1 port map( A => n1584, B => DATAIN(31), S => n214, Z => n4605
                           );
   U1780 : MUX2_X1 port map( A => n1585, B => DATAIN(0), S => n215, Z => n4542)
                           ;
   U1781 : MUX2_X1 port map( A => n1586, B => DATAIN(1), S => n215, Z => n4543)
                           ;
   U1782 : MUX2_X1 port map( A => n1587, B => DATAIN(2), S => n215, Z => n4544)
                           ;
   U1783 : MUX2_X1 port map( A => n1588, B => DATAIN(3), S => n215, Z => n4545)
                           ;
   U1784 : MUX2_X1 port map( A => n1589, B => DATAIN(4), S => n215, Z => n4546)
                           ;
   U1785 : MUX2_X1 port map( A => n1590, B => DATAIN(5), S => n215, Z => n4547)
                           ;
   U1786 : MUX2_X1 port map( A => n1591, B => DATAIN(6), S => n215, Z => n4548)
                           ;
   U1787 : MUX2_X1 port map( A => n1592, B => DATAIN(7), S => n215, Z => n4549)
                           ;
   U1788 : MUX2_X1 port map( A => n1593, B => DATAIN(8), S => n215, Z => n4550)
                           ;
   U1789 : MUX2_X1 port map( A => n1594, B => DATAIN(9), S => n215, Z => n4551)
                           ;
   U1790 : MUX2_X1 port map( A => n1595, B => DATAIN(10), S => n215, Z => n4552
                           );
   U1791 : MUX2_X1 port map( A => n1596, B => DATAIN(11), S => n215, Z => n4553
                           );
   U1792 : MUX2_X1 port map( A => n1597, B => DATAIN(12), S => n216, Z => n4554
                           );
   U1793 : MUX2_X1 port map( A => n1598, B => DATAIN(13), S => n216, Z => n4555
                           );
   U1794 : MUX2_X1 port map( A => n1599, B => DATAIN(14), S => n216, Z => n4556
                           );
   U1795 : MUX2_X1 port map( A => n1600, B => DATAIN(15), S => n216, Z => n4557
                           );
   U1796 : MUX2_X1 port map( A => n1601, B => DATAIN(16), S => n216, Z => n4558
                           );
   U1797 : MUX2_X1 port map( A => n1602, B => DATAIN(17), S => n216, Z => n4559
                           );
   U1798 : MUX2_X1 port map( A => n1603, B => DATAIN(18), S => n216, Z => n4560
                           );
   U1799 : MUX2_X1 port map( A => n1604, B => DATAIN(19), S => n216, Z => n4561
                           );
   U1800 : MUX2_X1 port map( A => n1605, B => DATAIN(20), S => n216, Z => n4562
                           );
   U1801 : MUX2_X1 port map( A => n1606, B => DATAIN(21), S => n216, Z => n4563
                           );
   U1802 : MUX2_X1 port map( A => n1607, B => DATAIN(22), S => n216, Z => n4564
                           );
   U1803 : MUX2_X1 port map( A => n1608, B => DATAIN(23), S => n216, Z => n4565
                           );
   U1804 : MUX2_X1 port map( A => n1609, B => DATAIN(24), S => n217, Z => n4566
                           );
   U1805 : MUX2_X1 port map( A => n1610, B => DATAIN(25), S => n217, Z => n4567
                           );
   U1806 : MUX2_X1 port map( A => n1611, B => DATAIN(26), S => n217, Z => n4568
                           );
   U1807 : MUX2_X1 port map( A => n1612, B => DATAIN(27), S => n217, Z => n4569
                           );
   U1808 : MUX2_X1 port map( A => n1613, B => DATAIN(28), S => n217, Z => n4570
                           );
   U1809 : MUX2_X1 port map( A => n1614, B => DATAIN(29), S => n217, Z => n4571
                           );
   U1810 : MUX2_X1 port map( A => n1615, B => DATAIN(30), S => n217, Z => n4572
                           );
   U1811 : MUX2_X1 port map( A => n1616, B => DATAIN(31), S => n217, Z => n4573
                           );
   U1812 : MUX2_X1 port map( A => n3964, B => DATAIN(0), S => n218, Z => n3239)
                           ;
   U1813 : MUX2_X1 port map( A => n3941, B => DATAIN(1), S => n218, Z => n3240)
                           ;
   U1814 : MUX2_X1 port map( A => n3918, B => DATAIN(2), S => n218, Z => n3241)
                           ;
   U1815 : MUX2_X1 port map( A => n3895, B => DATAIN(3), S => n218, Z => n3242)
                           ;
   U1816 : MUX2_X1 port map( A => n3872, B => DATAIN(4), S => n218, Z => n3243)
                           ;
   U1817 : MUX2_X1 port map( A => n3849, B => DATAIN(5), S => n218, Z => n3244)
                           ;
   U1818 : MUX2_X1 port map( A => n3826, B => DATAIN(6), S => n218, Z => n3245)
                           ;
   U1819 : MUX2_X1 port map( A => n3803, B => DATAIN(7), S => n218, Z => n3246)
                           ;
   U1820 : MUX2_X1 port map( A => n3780, B => DATAIN(8), S => n218, Z => n3247)
                           ;
   U1821 : MUX2_X1 port map( A => n3757, B => DATAIN(9), S => n218, Z => n3248)
                           ;
   U1822 : MUX2_X1 port map( A => n3734, B => DATAIN(10), S => n218, Z => n3249
                           );
   U1823 : MUX2_X1 port map( A => n3711, B => DATAIN(11), S => n218, Z => n3250
                           );
   U1824 : MUX2_X1 port map( A => n3688, B => DATAIN(12), S => n219, Z => n3251
                           );
   U1825 : MUX2_X1 port map( A => n3665, B => DATAIN(13), S => n219, Z => n3252
                           );
   U1826 : MUX2_X1 port map( A => n3642, B => DATAIN(14), S => n219, Z => n3253
                           );
   U1827 : MUX2_X1 port map( A => n3619, B => DATAIN(15), S => n219, Z => n3254
                           );
   U1828 : MUX2_X1 port map( A => n3596, B => DATAIN(16), S => n219, Z => n3255
                           );
   U1829 : MUX2_X1 port map( A => n3573, B => DATAIN(17), S => n219, Z => n3256
                           );
   U1830 : MUX2_X1 port map( A => n2974, B => DATAIN(18), S => n219, Z => n3257
                           );
   U1831 : MUX2_X1 port map( A => n2951, B => DATAIN(19), S => n219, Z => n3258
                           );
   U1832 : MUX2_X1 port map( A => n2928, B => DATAIN(20), S => n219, Z => n3259
                           );
   U1833 : MUX2_X1 port map( A => n2905, B => DATAIN(21), S => n219, Z => n3260
                           );
   U1834 : MUX2_X1 port map( A => n2882, B => DATAIN(22), S => n219, Z => n3261
                           );
   U1835 : MUX2_X1 port map( A => n2859, B => DATAIN(23), S => n219, Z => n3262
                           );
   U1836 : MUX2_X1 port map( A => n2836, B => DATAIN(24), S => n220, Z => n3263
                           );
   U1837 : MUX2_X1 port map( A => n2813, B => DATAIN(25), S => n220, Z => n3264
                           );
   U1838 : MUX2_X1 port map( A => n2790, B => DATAIN(26), S => n220, Z => n3265
                           );
   U1839 : MUX2_X1 port map( A => n2767, B => DATAIN(27), S => n220, Z => n3266
                           );
   U1840 : MUX2_X1 port map( A => n2744, B => DATAIN(28), S => n220, Z => n3267
                           );
   U1841 : MUX2_X1 port map( A => n2721, B => DATAIN(29), S => n220, Z => n3268
                           );
   U1842 : MUX2_X1 port map( A => n2698, B => DATAIN(30), S => n220, Z => n3269
                           );
   U1843 : MUX2_X1 port map( A => n2675, B => DATAIN(31), S => n220, Z => n3270
                           );
   U1844 : MUX2_X1 port map( A => n3965, B => DATAIN(0), S => n221, Z => n3271)
                           ;
   U1845 : MUX2_X1 port map( A => n3942, B => DATAIN(1), S => n221, Z => n3272)
                           ;
   U1846 : MUX2_X1 port map( A => n3919, B => DATAIN(2), S => n221, Z => n3273)
                           ;
   U1847 : MUX2_X1 port map( A => n3896, B => DATAIN(3), S => n221, Z => n3274)
                           ;
   U1848 : MUX2_X1 port map( A => n3873, B => DATAIN(4), S => n221, Z => n3275)
                           ;
   U1849 : MUX2_X1 port map( A => n3850, B => DATAIN(5), S => n221, Z => n3276)
                           ;
   U1850 : MUX2_X1 port map( A => n3827, B => DATAIN(6), S => n221, Z => n3277)
                           ;
   U1851 : MUX2_X1 port map( A => n3804, B => DATAIN(7), S => n221, Z => n3278)
                           ;
   U1852 : MUX2_X1 port map( A => n3781, B => DATAIN(8), S => n221, Z => n3279)
                           ;
   U1853 : MUX2_X1 port map( A => n3758, B => DATAIN(9), S => n221, Z => n3280)
                           ;
   U1854 : MUX2_X1 port map( A => n3735, B => DATAIN(10), S => n221, Z => n3281
                           );
   U1855 : MUX2_X1 port map( A => n3712, B => DATAIN(11), S => n221, Z => n3282
                           );
   U1856 : MUX2_X1 port map( A => n3689, B => DATAIN(12), S => n222, Z => n3283
                           );
   U1857 : MUX2_X1 port map( A => n3666, B => DATAIN(13), S => n222, Z => n3284
                           );
   U1858 : MUX2_X1 port map( A => n3643, B => DATAIN(14), S => n222, Z => n3285
                           );
   U1859 : MUX2_X1 port map( A => n3620, B => DATAIN(15), S => n222, Z => n3286
                           );
   U1860 : MUX2_X1 port map( A => n3597, B => DATAIN(16), S => n222, Z => n3287
                           );
   U1861 : MUX2_X1 port map( A => n3574, B => DATAIN(17), S => n222, Z => n3288
                           );
   U1862 : MUX2_X1 port map( A => n2975, B => DATAIN(18), S => n222, Z => n3289
                           );
   U1863 : MUX2_X1 port map( A => n2952, B => DATAIN(19), S => n222, Z => n3290
                           );
   U1864 : MUX2_X1 port map( A => n2929, B => DATAIN(20), S => n222, Z => n3291
                           );
   U1865 : MUX2_X1 port map( A => n2906, B => DATAIN(21), S => n222, Z => n3292
                           );
   U1866 : MUX2_X1 port map( A => n2883, B => DATAIN(22), S => n222, Z => n3293
                           );
   U1867 : MUX2_X1 port map( A => n2860, B => DATAIN(23), S => n222, Z => n3294
                           );
   U1868 : MUX2_X1 port map( A => n2837, B => DATAIN(24), S => n223, Z => n3295
                           );
   U1869 : MUX2_X1 port map( A => n2814, B => DATAIN(25), S => n223, Z => n3296
                           );
   U1870 : MUX2_X1 port map( A => n2791, B => DATAIN(26), S => n223, Z => n3297
                           );
   U1871 : MUX2_X1 port map( A => n2768, B => DATAIN(27), S => n223, Z => n3298
                           );
   U1872 : MUX2_X1 port map( A => n2745, B => DATAIN(28), S => n223, Z => n3299
                           );
   U1873 : MUX2_X1 port map( A => n2722, B => DATAIN(29), S => n223, Z => n3300
                           );
   U1874 : MUX2_X1 port map( A => n2699, B => DATAIN(30), S => n223, Z => n3301
                           );
   U1875 : MUX2_X1 port map( A => n2676, B => DATAIN(31), S => n223, Z => n3302
                           );
   U1876 : MUX2_X1 port map( A => n1617, B => DATAIN(0), S => n224, Z => n4510)
                           ;
   U1877 : MUX2_X1 port map( A => n1618, B => DATAIN(1), S => n224, Z => n4511)
                           ;
   U1878 : MUX2_X1 port map( A => n1619, B => DATAIN(2), S => n224, Z => n4512)
                           ;
   U1879 : MUX2_X1 port map( A => n1620, B => DATAIN(3), S => n224, Z => n4513)
                           ;
   U1880 : MUX2_X1 port map( A => n1621, B => DATAIN(4), S => n224, Z => n4514)
                           ;
   U1881 : MUX2_X1 port map( A => n1622, B => DATAIN(5), S => n224, Z => n4515)
                           ;
   U1882 : MUX2_X1 port map( A => n1623, B => DATAIN(6), S => n224, Z => n4516)
                           ;
   U1883 : MUX2_X1 port map( A => n1624, B => DATAIN(7), S => n224, Z => n4517)
                           ;
   U1884 : MUX2_X1 port map( A => n1625, B => DATAIN(8), S => n224, Z => n4518)
                           ;
   U1885 : MUX2_X1 port map( A => n1626, B => DATAIN(9), S => n224, Z => n4519)
                           ;
   U1886 : MUX2_X1 port map( A => n1627, B => DATAIN(10), S => n224, Z => n4520
                           );
   U1887 : MUX2_X1 port map( A => n1628, B => DATAIN(11), S => n224, Z => n4521
                           );
   U1888 : MUX2_X1 port map( A => n1629, B => DATAIN(12), S => n225, Z => n4522
                           );
   U1889 : MUX2_X1 port map( A => n1630, B => DATAIN(13), S => n225, Z => n4523
                           );
   U1890 : MUX2_X1 port map( A => n1631, B => DATAIN(14), S => n225, Z => n4524
                           );
   U1891 : MUX2_X1 port map( A => n1632, B => DATAIN(15), S => n225, Z => n4525
                           );
   U1892 : MUX2_X1 port map( A => n1633, B => DATAIN(16), S => n225, Z => n4526
                           );
   U1893 : MUX2_X1 port map( A => n1634, B => DATAIN(17), S => n225, Z => n4527
                           );
   U1894 : MUX2_X1 port map( A => n1635, B => DATAIN(18), S => n225, Z => n4528
                           );
   U1895 : MUX2_X1 port map( A => n1636, B => DATAIN(19), S => n225, Z => n4529
                           );
   U1896 : MUX2_X1 port map( A => n1637, B => DATAIN(20), S => n225, Z => n4530
                           );
   U1897 : MUX2_X1 port map( A => n1638, B => DATAIN(21), S => n225, Z => n4531
                           );
   U1898 : MUX2_X1 port map( A => n1639, B => DATAIN(22), S => n225, Z => n4532
                           );
   U1899 : MUX2_X1 port map( A => n1640, B => DATAIN(23), S => n225, Z => n4533
                           );
   U1900 : MUX2_X1 port map( A => n1641, B => DATAIN(24), S => n226, Z => n4534
                           );
   U1901 : MUX2_X1 port map( A => n1642, B => DATAIN(25), S => n226, Z => n4535
                           );
   U1902 : MUX2_X1 port map( A => n1643, B => DATAIN(26), S => n226, Z => n4536
                           );
   U1903 : MUX2_X1 port map( A => n1644, B => DATAIN(27), S => n226, Z => n4537
                           );
   U1904 : MUX2_X1 port map( A => n1645, B => DATAIN(28), S => n226, Z => n4538
                           );
   U1905 : MUX2_X1 port map( A => n1646, B => DATAIN(29), S => n226, Z => n4539
                           );
   U1906 : MUX2_X1 port map( A => n1647, B => DATAIN(30), S => n226, Z => n4540
                           );
   U1907 : MUX2_X1 port map( A => n1648, B => DATAIN(31), S => n226, Z => n4541
                           );
   U1908 : MUX2_X1 port map( A => n1649, B => DATAIN(0), S => n227, Z => n4478)
                           ;
   U1909 : MUX2_X1 port map( A => n1650, B => DATAIN(1), S => n227, Z => n4479)
                           ;
   U1910 : MUX2_X1 port map( A => n1651, B => DATAIN(2), S => n227, Z => n4480)
                           ;
   U1911 : MUX2_X1 port map( A => n1652, B => DATAIN(3), S => n227, Z => n4481)
                           ;
   U1912 : MUX2_X1 port map( A => n1653, B => DATAIN(4), S => n227, Z => n4482)
                           ;
   U1913 : MUX2_X1 port map( A => n1654, B => DATAIN(5), S => n227, Z => n4483)
                           ;
   U1914 : MUX2_X1 port map( A => n1655, B => DATAIN(6), S => n227, Z => n4484)
                           ;
   U1915 : MUX2_X1 port map( A => n1656, B => DATAIN(7), S => n227, Z => n4485)
                           ;
   U1916 : MUX2_X1 port map( A => n1657, B => DATAIN(8), S => n227, Z => n4486)
                           ;
   U1917 : MUX2_X1 port map( A => n1658, B => DATAIN(9), S => n227, Z => n4487)
                           ;
   U1918 : MUX2_X1 port map( A => n1659, B => DATAIN(10), S => n227, Z => n4488
                           );
   U1919 : MUX2_X1 port map( A => n1660, B => DATAIN(11), S => n227, Z => n4489
                           );
   U1920 : MUX2_X1 port map( A => n1661, B => DATAIN(12), S => n228, Z => n4490
                           );
   U1921 : MUX2_X1 port map( A => n1662, B => DATAIN(13), S => n228, Z => n4491
                           );
   U1922 : MUX2_X1 port map( A => n1663, B => DATAIN(14), S => n228, Z => n4492
                           );
   U1923 : MUX2_X1 port map( A => n1664, B => DATAIN(15), S => n228, Z => n4493
                           );
   U1924 : MUX2_X1 port map( A => n1665, B => DATAIN(16), S => n228, Z => n4494
                           );
   U1925 : MUX2_X1 port map( A => n1666, B => DATAIN(17), S => n228, Z => n4495
                           );
   U1926 : MUX2_X1 port map( A => n1667, B => DATAIN(18), S => n228, Z => n4496
                           );
   U1927 : MUX2_X1 port map( A => n1668, B => DATAIN(19), S => n228, Z => n4497
                           );
   U1928 : MUX2_X1 port map( A => n1669, B => DATAIN(20), S => n228, Z => n4498
                           );
   U1929 : MUX2_X1 port map( A => n1670, B => DATAIN(21), S => n228, Z => n4499
                           );
   U1930 : MUX2_X1 port map( A => n1671, B => DATAIN(22), S => n228, Z => n4500
                           );
   U1931 : MUX2_X1 port map( A => n1672, B => DATAIN(23), S => n228, Z => n4501
                           );
   U1932 : MUX2_X1 port map( A => n1673, B => DATAIN(24), S => n229, Z => n4502
                           );
   U1933 : MUX2_X1 port map( A => n1674, B => DATAIN(25), S => n229, Z => n4503
                           );
   U1934 : MUX2_X1 port map( A => n1675, B => DATAIN(26), S => n229, Z => n4504
                           );
   U1935 : MUX2_X1 port map( A => n1676, B => DATAIN(27), S => n229, Z => n4505
                           );
   U1936 : MUX2_X1 port map( A => n1677, B => DATAIN(28), S => n229, Z => n4506
                           );
   U1937 : MUX2_X1 port map( A => n1678, B => DATAIN(29), S => n229, Z => n4507
                           );
   U1938 : MUX2_X1 port map( A => n1679, B => DATAIN(30), S => n229, Z => n4508
                           );
   U1939 : MUX2_X1 port map( A => n1680, B => DATAIN(31), S => n229, Z => n4509
                           );
   U1940 : INV_X1 port map( A => ADD_WR(4), ZN => n1809);
   U1941 : MUX2_X1 port map( A => n3946, B => DATAIN(0), S => n230, Z => n3303)
                           ;
   U1942 : MUX2_X1 port map( A => n3923, B => DATAIN(1), S => n230, Z => n3304)
                           ;
   U1943 : MUX2_X1 port map( A => n3900, B => DATAIN(2), S => n230, Z => n3305)
                           ;
   U1944 : MUX2_X1 port map( A => n3877, B => DATAIN(3), S => n230, Z => n3306)
                           ;
   U1945 : MUX2_X1 port map( A => n3854, B => DATAIN(4), S => n230, Z => n3307)
                           ;
   U1946 : MUX2_X1 port map( A => n3831, B => DATAIN(5), S => n230, Z => n3308)
                           ;
   U1947 : MUX2_X1 port map( A => n3808, B => DATAIN(6), S => n230, Z => n3309)
                           ;
   U1948 : MUX2_X1 port map( A => n3785, B => DATAIN(7), S => n230, Z => n3310)
                           ;
   U1949 : MUX2_X1 port map( A => n3762, B => DATAIN(8), S => n230, Z => n3311)
                           ;
   U1950 : MUX2_X1 port map( A => n3739, B => DATAIN(9), S => n230, Z => n3312)
                           ;
   U1951 : MUX2_X1 port map( A => n3716, B => DATAIN(10), S => n230, Z => n3313
                           );
   U1952 : MUX2_X1 port map( A => n3693, B => DATAIN(11), S => n230, Z => n3314
                           );
   U1953 : MUX2_X1 port map( A => n3670, B => DATAIN(12), S => n231, Z => n3315
                           );
   U1954 : MUX2_X1 port map( A => n3647, B => DATAIN(13), S => n231, Z => n3316
                           );
   U1955 : MUX2_X1 port map( A => n3624, B => DATAIN(14), S => n231, Z => n3317
                           );
   U1956 : MUX2_X1 port map( A => n3601, B => DATAIN(15), S => n231, Z => n3318
                           );
   U1957 : MUX2_X1 port map( A => n3578, B => DATAIN(16), S => n231, Z => n3319
                           );
   U1958 : MUX2_X1 port map( A => n2979, B => DATAIN(17), S => n231, Z => n3320
                           );
   U1959 : MUX2_X1 port map( A => n2956, B => DATAIN(18), S => n231, Z => n3321
                           );
   U1960 : MUX2_X1 port map( A => n2933, B => DATAIN(19), S => n231, Z => n3322
                           );
   U1961 : MUX2_X1 port map( A => n2910, B => DATAIN(20), S => n231, Z => n3323
                           );
   U1962 : MUX2_X1 port map( A => n2887, B => DATAIN(21), S => n231, Z => n3324
                           );
   U1963 : MUX2_X1 port map( A => n2864, B => DATAIN(22), S => n231, Z => n3325
                           );
   U1964 : MUX2_X1 port map( A => n2841, B => DATAIN(23), S => n231, Z => n3326
                           );
   U1965 : MUX2_X1 port map( A => n2818, B => DATAIN(24), S => n232, Z => n3327
                           );
   U1966 : MUX2_X1 port map( A => n2795, B => DATAIN(25), S => n232, Z => n3328
                           );
   U1967 : MUX2_X1 port map( A => n2772, B => DATAIN(26), S => n232, Z => n3329
                           );
   U1968 : MUX2_X1 port map( A => n2749, B => DATAIN(27), S => n232, Z => n3330
                           );
   U1969 : MUX2_X1 port map( A => n2726, B => DATAIN(28), S => n232, Z => n3331
                           );
   U1970 : MUX2_X1 port map( A => n2703, B => DATAIN(29), S => n232, Z => n3332
                           );
   U1971 : MUX2_X1 port map( A => n2680, B => DATAIN(30), S => n232, Z => n3333
                           );
   U1972 : MUX2_X1 port map( A => n2657, B => DATAIN(31), S => n232, Z => n3334
                           );
   U1973 : MUX2_X1 port map( A => n3947, B => DATAIN(0), S => n233, Z => n3335)
                           ;
   U1974 : MUX2_X1 port map( A => n3924, B => DATAIN(1), S => n233, Z => n3336)
                           ;
   U1975 : MUX2_X1 port map( A => n3901, B => DATAIN(2), S => n233, Z => n3337)
                           ;
   U1976 : MUX2_X1 port map( A => n3878, B => DATAIN(3), S => n233, Z => n3338)
                           ;
   U1977 : MUX2_X1 port map( A => n3855, B => DATAIN(4), S => n233, Z => n3339)
                           ;
   U1978 : MUX2_X1 port map( A => n3832, B => DATAIN(5), S => n233, Z => n3340)
                           ;
   U1979 : MUX2_X1 port map( A => n3809, B => DATAIN(6), S => n233, Z => n3341)
                           ;
   U1980 : MUX2_X1 port map( A => n3786, B => DATAIN(7), S => n233, Z => n3342)
                           ;
   U1981 : MUX2_X1 port map( A => n3763, B => DATAIN(8), S => n233, Z => n3343)
                           ;
   U1982 : MUX2_X1 port map( A => n3740, B => DATAIN(9), S => n233, Z => n3344)
                           ;
   U1983 : MUX2_X1 port map( A => n3717, B => DATAIN(10), S => n233, Z => n3345
                           );
   U1984 : MUX2_X1 port map( A => n3694, B => DATAIN(11), S => n233, Z => n3346
                           );
   U1985 : MUX2_X1 port map( A => n3671, B => DATAIN(12), S => n234, Z => n3347
                           );
   U1986 : MUX2_X1 port map( A => n3648, B => DATAIN(13), S => n234, Z => n3348
                           );
   U1987 : MUX2_X1 port map( A => n3625, B => DATAIN(14), S => n234, Z => n3349
                           );
   U1988 : MUX2_X1 port map( A => n3602, B => DATAIN(15), S => n234, Z => n3350
                           );
   U1989 : MUX2_X1 port map( A => n3579, B => DATAIN(16), S => n234, Z => n3351
                           );
   U1990 : MUX2_X1 port map( A => n2980, B => DATAIN(17), S => n234, Z => n3352
                           );
   U1991 : MUX2_X1 port map( A => n2957, B => DATAIN(18), S => n234, Z => n3353
                           );
   U1992 : MUX2_X1 port map( A => n2934, B => DATAIN(19), S => n234, Z => n3354
                           );
   U1993 : MUX2_X1 port map( A => n2911, B => DATAIN(20), S => n234, Z => n3355
                           );
   U1994 : MUX2_X1 port map( A => n2888, B => DATAIN(21), S => n234, Z => n3356
                           );
   U1995 : MUX2_X1 port map( A => n2865, B => DATAIN(22), S => n234, Z => n3357
                           );
   U1996 : MUX2_X1 port map( A => n2842, B => DATAIN(23), S => n234, Z => n3358
                           );
   U1997 : MUX2_X1 port map( A => n2819, B => DATAIN(24), S => n235, Z => n3359
                           );
   U1998 : MUX2_X1 port map( A => n2796, B => DATAIN(25), S => n235, Z => n3360
                           );
   U1999 : MUX2_X1 port map( A => n2773, B => DATAIN(26), S => n235, Z => n3361
                           );
   U2000 : MUX2_X1 port map( A => n2750, B => DATAIN(27), S => n235, Z => n3362
                           );
   U2001 : MUX2_X1 port map( A => n2727, B => DATAIN(28), S => n235, Z => n3363
                           );
   U2002 : MUX2_X1 port map( A => n2704, B => DATAIN(29), S => n235, Z => n3364
                           );
   U2003 : MUX2_X1 port map( A => n2681, B => DATAIN(30), S => n235, Z => n3365
                           );
   U2004 : MUX2_X1 port map( A => n2658, B => DATAIN(31), S => n235, Z => n3366
                           );
   U2005 : MUX2_X1 port map( A => n1681, B => DATAIN(0), S => n236, Z => n4222)
                           ;
   U2006 : MUX2_X1 port map( A => n1682, B => DATAIN(1), S => n236, Z => n4223)
                           ;
   U2007 : MUX2_X1 port map( A => n1683, B => DATAIN(2), S => n236, Z => n4224)
                           ;
   U2008 : MUX2_X1 port map( A => n1684, B => DATAIN(3), S => n236, Z => n4225)
                           ;
   U2009 : MUX2_X1 port map( A => n1685, B => DATAIN(4), S => n236, Z => n4226)
                           ;
   U2010 : MUX2_X1 port map( A => n1686, B => DATAIN(5), S => n236, Z => n4227)
                           ;
   U2011 : MUX2_X1 port map( A => n1687, B => DATAIN(6), S => n236, Z => n4228)
                           ;
   U2012 : MUX2_X1 port map( A => n1688, B => DATAIN(7), S => n236, Z => n4229)
                           ;
   U2013 : MUX2_X1 port map( A => n1689, B => DATAIN(8), S => n236, Z => n4230)
                           ;
   U2014 : MUX2_X1 port map( A => n1690, B => DATAIN(9), S => n236, Z => n4231)
                           ;
   U2015 : MUX2_X1 port map( A => n1691, B => DATAIN(10), S => n236, Z => n4232
                           );
   U2016 : MUX2_X1 port map( A => n1692, B => DATAIN(11), S => n236, Z => n4233
                           );
   U2017 : MUX2_X1 port map( A => n1693, B => DATAIN(12), S => n237, Z => n4234
                           );
   U2018 : MUX2_X1 port map( A => n1694, B => DATAIN(13), S => n237, Z => n4235
                           );
   U2019 : MUX2_X1 port map( A => n1695, B => DATAIN(14), S => n237, Z => n4236
                           );
   U2020 : MUX2_X1 port map( A => n1696, B => DATAIN(15), S => n237, Z => n4237
                           );
   U2021 : MUX2_X1 port map( A => n1697, B => DATAIN(16), S => n237, Z => n4238
                           );
   U2022 : MUX2_X1 port map( A => n1698, B => DATAIN(17), S => n237, Z => n4239
                           );
   U2023 : MUX2_X1 port map( A => n1699, B => DATAIN(18), S => n237, Z => n4240
                           );
   U2024 : MUX2_X1 port map( A => n1700, B => DATAIN(19), S => n237, Z => n4241
                           );
   U2025 : MUX2_X1 port map( A => n1701, B => DATAIN(20), S => n237, Z => n4242
                           );
   U2026 : MUX2_X1 port map( A => n1702, B => DATAIN(21), S => n237, Z => n4243
                           );
   U2027 : MUX2_X1 port map( A => n1703, B => DATAIN(22), S => n237, Z => n4244
                           );
   U2028 : MUX2_X1 port map( A => n1704, B => DATAIN(23), S => n237, Z => n4245
                           );
   U2029 : MUX2_X1 port map( A => n1705, B => DATAIN(24), S => n238, Z => n4246
                           );
   U2030 : MUX2_X1 port map( A => n1706, B => DATAIN(25), S => n238, Z => n4247
                           );
   U2031 : MUX2_X1 port map( A => n1707, B => DATAIN(26), S => n238, Z => n4248
                           );
   U2032 : MUX2_X1 port map( A => n1708, B => DATAIN(27), S => n238, Z => n4249
                           );
   U2033 : MUX2_X1 port map( A => n1709, B => DATAIN(28), S => n238, Z => n4250
                           );
   U2034 : MUX2_X1 port map( A => n1710, B => DATAIN(29), S => n238, Z => n4251
                           );
   U2035 : MUX2_X1 port map( A => n1711, B => DATAIN(30), S => n238, Z => n4252
                           );
   U2036 : MUX2_X1 port map( A => n1712, B => DATAIN(31), S => n238, Z => n4253
                           );
   U2037 : MUX2_X1 port map( A => n1713, B => DATAIN(0), S => n239, Z => n4190)
                           ;
   U2038 : MUX2_X1 port map( A => n1714, B => DATAIN(1), S => n239, Z => n4191)
                           ;
   U2039 : MUX2_X1 port map( A => n1715, B => DATAIN(2), S => n239, Z => n4192)
                           ;
   U2040 : MUX2_X1 port map( A => n1716, B => DATAIN(3), S => n239, Z => n4193)
                           ;
   U2041 : MUX2_X1 port map( A => n1717, B => DATAIN(4), S => n239, Z => n4194)
                           ;
   U2042 : MUX2_X1 port map( A => n1718, B => DATAIN(5), S => n239, Z => n4195)
                           ;
   U2043 : MUX2_X1 port map( A => n1719, B => DATAIN(6), S => n239, Z => n4196)
                           ;
   U2044 : MUX2_X1 port map( A => n1720, B => DATAIN(7), S => n239, Z => n4197)
                           ;
   U2045 : MUX2_X1 port map( A => n1721, B => DATAIN(8), S => n239, Z => n4198)
                           ;
   U2046 : MUX2_X1 port map( A => n1722, B => DATAIN(9), S => n239, Z => n4199)
                           ;
   U2047 : MUX2_X1 port map( A => n1723, B => DATAIN(10), S => n239, Z => n4200
                           );
   U2048 : MUX2_X1 port map( A => n1724, B => DATAIN(11), S => n239, Z => n4201
                           );
   U2049 : MUX2_X1 port map( A => n1725, B => DATAIN(12), S => n240, Z => n4202
                           );
   U2050 : MUX2_X1 port map( A => n1726, B => DATAIN(13), S => n240, Z => n4203
                           );
   U2051 : MUX2_X1 port map( A => n1727, B => DATAIN(14), S => n240, Z => n4204
                           );
   U2052 : MUX2_X1 port map( A => n1728, B => DATAIN(15), S => n240, Z => n4205
                           );
   U2053 : MUX2_X1 port map( A => n1729, B => DATAIN(16), S => n240, Z => n4206
                           );
   U2054 : MUX2_X1 port map( A => n1730, B => DATAIN(17), S => n240, Z => n4207
                           );
   U2055 : MUX2_X1 port map( A => n1731, B => DATAIN(18), S => n240, Z => n4208
                           );
   U2056 : MUX2_X1 port map( A => n1732, B => DATAIN(19), S => n240, Z => n4209
                           );
   U2057 : MUX2_X1 port map( A => n1733, B => DATAIN(20), S => n240, Z => n4210
                           );
   U2058 : MUX2_X1 port map( A => n1734, B => DATAIN(21), S => n240, Z => n4211
                           );
   U2059 : MUX2_X1 port map( A => n1735, B => DATAIN(22), S => n240, Z => n4212
                           );
   U2060 : MUX2_X1 port map( A => n1736, B => DATAIN(23), S => n240, Z => n4213
                           );
   U2061 : MUX2_X1 port map( A => n1737, B => DATAIN(24), S => n241, Z => n4214
                           );
   U2062 : MUX2_X1 port map( A => n1738, B => DATAIN(25), S => n241, Z => n4215
                           );
   U2063 : MUX2_X1 port map( A => n1739, B => DATAIN(26), S => n241, Z => n4216
                           );
   U2064 : MUX2_X1 port map( A => n1740, B => DATAIN(27), S => n241, Z => n4217
                           );
   U2065 : MUX2_X1 port map( A => n1741, B => DATAIN(28), S => n241, Z => n4218
                           );
   U2066 : MUX2_X1 port map( A => n1742, B => DATAIN(29), S => n241, Z => n4219
                           );
   U2067 : MUX2_X1 port map( A => n1743, B => DATAIN(30), S => n241, Z => n4220
                           );
   U2068 : MUX2_X1 port map( A => n1744, B => DATAIN(31), S => n241, Z => n4221
                           );
   U2069 : MUX2_X1 port map( A => n3950, B => DATAIN(0), S => n242, Z => n3367)
                           ;
   U2070 : MUX2_X1 port map( A => n3927, B => DATAIN(1), S => n242, Z => n3368)
                           ;
   U2071 : MUX2_X1 port map( A => n3904, B => DATAIN(2), S => n242, Z => n3369)
                           ;
   U2072 : MUX2_X1 port map( A => n3881, B => DATAIN(3), S => n242, Z => n3370)
                           ;
   U2073 : MUX2_X1 port map( A => n3858, B => DATAIN(4), S => n242, Z => n3371)
                           ;
   U2074 : MUX2_X1 port map( A => n3835, B => DATAIN(5), S => n242, Z => n3372)
                           ;
   U2075 : MUX2_X1 port map( A => n3812, B => DATAIN(6), S => n242, Z => n3373)
                           ;
   U2076 : MUX2_X1 port map( A => n3789, B => DATAIN(7), S => n242, Z => n3374)
                           ;
   U2077 : MUX2_X1 port map( A => n3766, B => DATAIN(8), S => n242, Z => n3375)
                           ;
   U2078 : MUX2_X1 port map( A => n3743, B => DATAIN(9), S => n242, Z => n3376)
                           ;
   U2079 : MUX2_X1 port map( A => n3720, B => DATAIN(10), S => n242, Z => n3377
                           );
   U2080 : MUX2_X1 port map( A => n3697, B => DATAIN(11), S => n242, Z => n3378
                           );
   U2081 : MUX2_X1 port map( A => n3674, B => DATAIN(12), S => n243, Z => n3379
                           );
   U2082 : MUX2_X1 port map( A => n3651, B => DATAIN(13), S => n243, Z => n3380
                           );
   U2083 : MUX2_X1 port map( A => n3628, B => DATAIN(14), S => n243, Z => n3381
                           );
   U2084 : MUX2_X1 port map( A => n3605, B => DATAIN(15), S => n243, Z => n3382
                           );
   U2085 : MUX2_X1 port map( A => n3582, B => DATAIN(16), S => n243, Z => n3383
                           );
   U2086 : MUX2_X1 port map( A => n3559, B => DATAIN(17), S => n243, Z => n3384
                           );
   U2087 : MUX2_X1 port map( A => n2960, B => DATAIN(18), S => n243, Z => n3385
                           );
   U2088 : MUX2_X1 port map( A => n2937, B => DATAIN(19), S => n243, Z => n3386
                           );
   U2089 : MUX2_X1 port map( A => n2914, B => DATAIN(20), S => n243, Z => n3387
                           );
   U2090 : MUX2_X1 port map( A => n2891, B => DATAIN(21), S => n243, Z => n3388
                           );
   U2091 : MUX2_X1 port map( A => n2868, B => DATAIN(22), S => n243, Z => n3389
                           );
   U2092 : MUX2_X1 port map( A => n2845, B => DATAIN(23), S => n243, Z => n3390
                           );
   U2093 : MUX2_X1 port map( A => n2822, B => DATAIN(24), S => n244, Z => n3391
                           );
   U2094 : MUX2_X1 port map( A => n2799, B => DATAIN(25), S => n244, Z => n3392
                           );
   U2095 : MUX2_X1 port map( A => n2776, B => DATAIN(26), S => n244, Z => n3393
                           );
   U2096 : MUX2_X1 port map( A => n2753, B => DATAIN(27), S => n244, Z => n3394
                           );
   U2097 : MUX2_X1 port map( A => n2730, B => DATAIN(28), S => n244, Z => n3395
                           );
   U2098 : MUX2_X1 port map( A => n2707, B => DATAIN(29), S => n244, Z => n3396
                           );
   U2099 : MUX2_X1 port map( A => n2684, B => DATAIN(30), S => n244, Z => n3397
                           );
   U2100 : MUX2_X1 port map( A => n2661, B => DATAIN(31), S => n244, Z => n3398
                           );
   U2101 : MUX2_X1 port map( A => n3951, B => DATAIN(0), S => n245, Z => n3399)
                           ;
   U2102 : MUX2_X1 port map( A => n3928, B => DATAIN(1), S => n245, Z => n3400)
                           ;
   U2103 : MUX2_X1 port map( A => n3905, B => DATAIN(2), S => n245, Z => n3401)
                           ;
   U2104 : MUX2_X1 port map( A => n3882, B => DATAIN(3), S => n245, Z => n3402)
                           ;
   U2105 : MUX2_X1 port map( A => n3859, B => DATAIN(4), S => n245, Z => n3403)
                           ;
   U2106 : MUX2_X1 port map( A => n3836, B => DATAIN(5), S => n245, Z => n3404)
                           ;
   U2107 : MUX2_X1 port map( A => n3813, B => DATAIN(6), S => n245, Z => n3405)
                           ;
   U2108 : MUX2_X1 port map( A => n3790, B => DATAIN(7), S => n245, Z => n3406)
                           ;
   U2109 : MUX2_X1 port map( A => n3767, B => DATAIN(8), S => n245, Z => n3407)
                           ;
   U2110 : MUX2_X1 port map( A => n3744, B => DATAIN(9), S => n245, Z => n3408)
                           ;
   U2111 : MUX2_X1 port map( A => n3721, B => DATAIN(10), S => n245, Z => n3409
                           );
   U2112 : MUX2_X1 port map( A => n3698, B => DATAIN(11), S => n245, Z => n3410
                           );
   U2113 : MUX2_X1 port map( A => n3675, B => DATAIN(12), S => n246, Z => n3411
                           );
   U2114 : MUX2_X1 port map( A => n3652, B => DATAIN(13), S => n246, Z => n3412
                           );
   U2115 : MUX2_X1 port map( A => n3629, B => DATAIN(14), S => n246, Z => n3413
                           );
   U2116 : MUX2_X1 port map( A => n3606, B => DATAIN(15), S => n246, Z => n3414
                           );
   U2117 : MUX2_X1 port map( A => n3583, B => DATAIN(16), S => n246, Z => n3415
                           );
   U2118 : MUX2_X1 port map( A => n3560, B => DATAIN(17), S => n246, Z => n3416
                           );
   U2119 : MUX2_X1 port map( A => n2961, B => DATAIN(18), S => n246, Z => n3417
                           );
   U2120 : MUX2_X1 port map( A => n2938, B => DATAIN(19), S => n246, Z => n3418
                           );
   U2121 : MUX2_X1 port map( A => n2915, B => DATAIN(20), S => n246, Z => n3419
                           );
   U2122 : MUX2_X1 port map( A => n2892, B => DATAIN(21), S => n246, Z => n3420
                           );
   U2123 : MUX2_X1 port map( A => n2869, B => DATAIN(22), S => n246, Z => n3421
                           );
   U2124 : MUX2_X1 port map( A => n2846, B => DATAIN(23), S => n246, Z => n3422
                           );
   U2125 : MUX2_X1 port map( A => n2823, B => DATAIN(24), S => n247, Z => n3423
                           );
   U2126 : MUX2_X1 port map( A => n2800, B => DATAIN(25), S => n247, Z => n3424
                           );
   U2127 : MUX2_X1 port map( A => n2777, B => DATAIN(26), S => n247, Z => n3425
                           );
   U2128 : MUX2_X1 port map( A => n2754, B => DATAIN(27), S => n247, Z => n3426
                           );
   U2129 : MUX2_X1 port map( A => n2731, B => DATAIN(28), S => n247, Z => n3427
                           );
   U2130 : MUX2_X1 port map( A => n2708, B => DATAIN(29), S => n247, Z => n3428
                           );
   U2131 : MUX2_X1 port map( A => n2685, B => DATAIN(30), S => n247, Z => n3429
                           );
   U2132 : MUX2_X1 port map( A => n2662, B => DATAIN(31), S => n247, Z => n3430
                           );
   U2133 : MUX2_X1 port map( A => n1745, B => DATAIN(0), S => n248, Z => n4158)
                           ;
   U2134 : MUX2_X1 port map( A => n1746, B => DATAIN(1), S => n248, Z => n4159)
                           ;
   U2135 : MUX2_X1 port map( A => n1747, B => DATAIN(2), S => n248, Z => n4160)
                           ;
   U2136 : MUX2_X1 port map( A => n1748, B => DATAIN(3), S => n248, Z => n4161)
                           ;
   U2137 : MUX2_X1 port map( A => n1749, B => DATAIN(4), S => n248, Z => n4162)
                           ;
   U2138 : MUX2_X1 port map( A => n1750, B => DATAIN(5), S => n248, Z => n4163)
                           ;
   U2139 : MUX2_X1 port map( A => n1751, B => DATAIN(6), S => n248, Z => n4164)
                           ;
   U2140 : MUX2_X1 port map( A => n1752, B => DATAIN(7), S => n248, Z => n4165)
                           ;
   U2141 : MUX2_X1 port map( A => n1753, B => DATAIN(8), S => n248, Z => n4166)
                           ;
   U2142 : MUX2_X1 port map( A => n1754, B => DATAIN(9), S => n248, Z => n4167)
                           ;
   U2143 : MUX2_X1 port map( A => n1755, B => DATAIN(10), S => n248, Z => n4168
                           );
   U2144 : MUX2_X1 port map( A => n1756, B => DATAIN(11), S => n248, Z => n4169
                           );
   U2145 : MUX2_X1 port map( A => n1757, B => DATAIN(12), S => n249, Z => n4170
                           );
   U2146 : MUX2_X1 port map( A => n1758, B => DATAIN(13), S => n249, Z => n4171
                           );
   U2147 : MUX2_X1 port map( A => n1759, B => DATAIN(14), S => n249, Z => n4172
                           );
   U2148 : MUX2_X1 port map( A => n1760, B => DATAIN(15), S => n249, Z => n4173
                           );
   U2149 : MUX2_X1 port map( A => n1761, B => DATAIN(16), S => n249, Z => n4174
                           );
   U2150 : MUX2_X1 port map( A => n1762, B => DATAIN(17), S => n249, Z => n4175
                           );
   U2151 : MUX2_X1 port map( A => n1763, B => DATAIN(18), S => n249, Z => n4176
                           );
   U2152 : MUX2_X1 port map( A => n1764, B => DATAIN(19), S => n249, Z => n4177
                           );
   U2153 : MUX2_X1 port map( A => n1765, B => DATAIN(20), S => n249, Z => n4178
                           );
   U2154 : MUX2_X1 port map( A => n1766, B => DATAIN(21), S => n249, Z => n4179
                           );
   U2155 : MUX2_X1 port map( A => n1767, B => DATAIN(22), S => n249, Z => n4180
                           );
   U2156 : MUX2_X1 port map( A => n1768, B => DATAIN(23), S => n249, Z => n4181
                           );
   U2157 : MUX2_X1 port map( A => n1769, B => DATAIN(24), S => n250, Z => n4182
                           );
   U2158 : MUX2_X1 port map( A => n1770, B => DATAIN(25), S => n250, Z => n4183
                           );
   U2159 : MUX2_X1 port map( A => n1771, B => DATAIN(26), S => n250, Z => n4184
                           );
   U2160 : MUX2_X1 port map( A => n1772, B => DATAIN(27), S => n250, Z => n4185
                           );
   U2161 : MUX2_X1 port map( A => n1773, B => DATAIN(28), S => n250, Z => n4186
                           );
   U2162 : MUX2_X1 port map( A => n1774, B => DATAIN(29), S => n250, Z => n4187
                           );
   U2163 : MUX2_X1 port map( A => n1775, B => DATAIN(30), S => n250, Z => n4188
                           );
   U2164 : MUX2_X1 port map( A => n1776, B => DATAIN(31), S => n250, Z => n4189
                           );
   U2165 : MUX2_X1 port map( A => n1777, B => DATAIN(0), S => n251, Z => n4126)
                           ;
   U2166 : MUX2_X1 port map( A => n1778, B => DATAIN(1), S => n251, Z => n4127)
                           ;
   U2167 : MUX2_X1 port map( A => n1779, B => DATAIN(2), S => n251, Z => n4128)
                           ;
   U2168 : MUX2_X1 port map( A => n1780, B => DATAIN(3), S => n251, Z => n4129)
                           ;
   U2169 : MUX2_X1 port map( A => n1781, B => DATAIN(4), S => n251, Z => n4130)
                           ;
   U2170 : MUX2_X1 port map( A => n1782, B => DATAIN(5), S => n251, Z => n4131)
                           ;
   U2171 : MUX2_X1 port map( A => n1783, B => DATAIN(6), S => n251, Z => n4132)
                           ;
   U2172 : MUX2_X1 port map( A => n1784, B => DATAIN(7), S => n251, Z => n4133)
                           ;
   U2173 : MUX2_X1 port map( A => n1785, B => DATAIN(8), S => n251, Z => n4134)
                           ;
   U2174 : MUX2_X1 port map( A => n1786, B => DATAIN(9), S => n251, Z => n4135)
                           ;
   U2175 : MUX2_X1 port map( A => n1787, B => DATAIN(10), S => n251, Z => n4136
                           );
   U2176 : MUX2_X1 port map( A => n1788, B => DATAIN(11), S => n251, Z => n4137
                           );
   U2177 : MUX2_X1 port map( A => n1789, B => DATAIN(12), S => n252, Z => n4138
                           );
   U2178 : MUX2_X1 port map( A => n1790, B => DATAIN(13), S => n252, Z => n4139
                           );
   U2179 : MUX2_X1 port map( A => n1791, B => DATAIN(14), S => n252, Z => n4140
                           );
   U2180 : MUX2_X1 port map( A => n1792, B => DATAIN(15), S => n252, Z => n4141
                           );
   U2181 : MUX2_X1 port map( A => n1793, B => DATAIN(16), S => n252, Z => n4142
                           );
   U2182 : MUX2_X1 port map( A => n1794, B => DATAIN(17), S => n252, Z => n4143
                           );
   U2183 : MUX2_X1 port map( A => n1795, B => DATAIN(18), S => n252, Z => n4144
                           );
   U2184 : MUX2_X1 port map( A => n1796, B => DATAIN(19), S => n252, Z => n4145
                           );
   U2185 : MUX2_X1 port map( A => n1797, B => DATAIN(20), S => n252, Z => n4146
                           );
   U2186 : MUX2_X1 port map( A => n1798, B => DATAIN(21), S => n252, Z => n4147
                           );
   U2187 : MUX2_X1 port map( A => n1799, B => DATAIN(22), S => n252, Z => n4148
                           );
   U2188 : MUX2_X1 port map( A => n1800, B => DATAIN(23), S => n252, Z => n4149
                           );
   U2189 : MUX2_X1 port map( A => n1801, B => DATAIN(24), S => n253, Z => n4150
                           );
   U2190 : MUX2_X1 port map( A => n1802, B => DATAIN(25), S => n253, Z => n4151
                           );
   U2191 : MUX2_X1 port map( A => n1803, B => DATAIN(26), S => n253, Z => n4152
                           );
   U2192 : MUX2_X1 port map( A => n1804, B => DATAIN(27), S => n253, Z => n4153
                           );
   U2193 : MUX2_X1 port map( A => n1805, B => DATAIN(28), S => n253, Z => n4154
                           );
   U2194 : MUX2_X1 port map( A => n1806, B => DATAIN(29), S => n253, Z => n4155
                           );
   U2195 : MUX2_X1 port map( A => n1807, B => DATAIN(30), S => n253, Z => n4156
                           );
   U2196 : MUX2_X1 port map( A => n1808, B => DATAIN(31), S => n253, Z => n4157
                           );
   U2197 : MUX2_X1 port map( A => n3953, B => DATAIN(0), S => n254, Z => n3431)
                           ;
   U2198 : MUX2_X1 port map( A => n3930, B => DATAIN(1), S => n254, Z => n3432)
                           ;
   U2199 : MUX2_X1 port map( A => n3907, B => DATAIN(2), S => n254, Z => n3433)
                           ;
   U2200 : MUX2_X1 port map( A => n3884, B => DATAIN(3), S => n254, Z => n3434)
                           ;
   U2201 : MUX2_X1 port map( A => n3861, B => DATAIN(4), S => n254, Z => n3435)
                           ;
   U2202 : MUX2_X1 port map( A => n3838, B => DATAIN(5), S => n254, Z => n3436)
                           ;
   U2203 : MUX2_X1 port map( A => n3815, B => DATAIN(6), S => n254, Z => n3437)
                           ;
   U2204 : MUX2_X1 port map( A => n3792, B => DATAIN(7), S => n254, Z => n3438)
                           ;
   U2205 : MUX2_X1 port map( A => n3769, B => DATAIN(8), S => n254, Z => n3439)
                           ;
   U2206 : MUX2_X1 port map( A => n3746, B => DATAIN(9), S => n254, Z => n3440)
                           ;
   U2207 : MUX2_X1 port map( A => n3723, B => DATAIN(10), S => n254, Z => n3441
                           );
   U2208 : MUX2_X1 port map( A => n3700, B => DATAIN(11), S => n254, Z => n3442
                           );
   U2209 : MUX2_X1 port map( A => n3677, B => DATAIN(12), S => n255, Z => n3443
                           );
   U2210 : MUX2_X1 port map( A => n3654, B => DATAIN(13), S => n255, Z => n3444
                           );
   U2211 : MUX2_X1 port map( A => n3631, B => DATAIN(14), S => n255, Z => n3445
                           );
   U2212 : MUX2_X1 port map( A => n3608, B => DATAIN(15), S => n255, Z => n3446
                           );
   U2213 : MUX2_X1 port map( A => n3585, B => DATAIN(16), S => n255, Z => n3447
                           );
   U2214 : MUX2_X1 port map( A => n3562, B => DATAIN(17), S => n255, Z => n3448
                           );
   U2215 : MUX2_X1 port map( A => n2963, B => DATAIN(18), S => n255, Z => n3449
                           );
   U2216 : MUX2_X1 port map( A => n2940, B => DATAIN(19), S => n255, Z => n3450
                           );
   U2217 : MUX2_X1 port map( A => n2917, B => DATAIN(20), S => n255, Z => n3451
                           );
   U2218 : MUX2_X1 port map( A => n2894, B => DATAIN(21), S => n255, Z => n3452
                           );
   U2219 : MUX2_X1 port map( A => n2871, B => DATAIN(22), S => n255, Z => n3453
                           );
   U2220 : MUX2_X1 port map( A => n2848, B => DATAIN(23), S => n255, Z => n3454
                           );
   U2221 : MUX2_X1 port map( A => n2825, B => DATAIN(24), S => n256, Z => n3455
                           );
   U2222 : MUX2_X1 port map( A => n2802, B => DATAIN(25), S => n256, Z => n3456
                           );
   U2223 : MUX2_X1 port map( A => n2779, B => DATAIN(26), S => n256, Z => n3457
                           );
   U2224 : MUX2_X1 port map( A => n2756, B => DATAIN(27), S => n256, Z => n3458
                           );
   U2225 : MUX2_X1 port map( A => n2733, B => DATAIN(28), S => n256, Z => n3459
                           );
   U2226 : MUX2_X1 port map( A => n2710, B => DATAIN(29), S => n256, Z => n3460
                           );
   U2227 : MUX2_X1 port map( A => n2687, B => DATAIN(30), S => n256, Z => n3461
                           );
   U2228 : MUX2_X1 port map( A => n2664, B => DATAIN(31), S => n256, Z => n3462
                           );
   U2229 : MUX2_X1 port map( A => n3954, B => DATAIN(0), S => n257, Z => n3463)
                           ;
   U2230 : MUX2_X1 port map( A => n3931, B => DATAIN(1), S => n257, Z => n3464)
                           ;
   U2231 : MUX2_X1 port map( A => n3908, B => DATAIN(2), S => n257, Z => n3465)
                           ;
   U2232 : MUX2_X1 port map( A => n3885, B => DATAIN(3), S => n257, Z => n3466)
                           ;
   U2233 : MUX2_X1 port map( A => n3862, B => DATAIN(4), S => n257, Z => n3467)
                           ;
   U2234 : MUX2_X1 port map( A => n3839, B => DATAIN(5), S => n257, Z => n3468)
                           ;
   U2235 : MUX2_X1 port map( A => n3816, B => DATAIN(6), S => n257, Z => n3469)
                           ;
   U2236 : MUX2_X1 port map( A => n3793, B => DATAIN(7), S => n257, Z => n3470)
                           ;
   U2237 : MUX2_X1 port map( A => n3770, B => DATAIN(8), S => n257, Z => n3471)
                           ;
   U2238 : MUX2_X1 port map( A => n3747, B => DATAIN(9), S => n257, Z => n3472)
                           ;
   U2239 : MUX2_X1 port map( A => n3724, B => DATAIN(10), S => n257, Z => n3473
                           );
   U2240 : MUX2_X1 port map( A => n3701, B => DATAIN(11), S => n257, Z => n3474
                           );
   U2241 : MUX2_X1 port map( A => n3678, B => DATAIN(12), S => n258, Z => n3475
                           );
   U2242 : MUX2_X1 port map( A => n3655, B => DATAIN(13), S => n258, Z => n3476
                           );
   U2243 : MUX2_X1 port map( A => n3632, B => DATAIN(14), S => n258, Z => n3477
                           );
   U2244 : MUX2_X1 port map( A => n3609, B => DATAIN(15), S => n258, Z => n3478
                           );
   U2245 : MUX2_X1 port map( A => n3586, B => DATAIN(16), S => n258, Z => n3479
                           );
   U2246 : MUX2_X1 port map( A => n3563, B => DATAIN(17), S => n258, Z => n3480
                           );
   U2247 : MUX2_X1 port map( A => n2964, B => DATAIN(18), S => n258, Z => n3481
                           );
   U2248 : MUX2_X1 port map( A => n2941, B => DATAIN(19), S => n258, Z => n3482
                           );
   U2249 : MUX2_X1 port map( A => n2918, B => DATAIN(20), S => n258, Z => n3483
                           );
   U2250 : MUX2_X1 port map( A => n2895, B => DATAIN(21), S => n258, Z => n3484
                           );
   U2251 : MUX2_X1 port map( A => n2872, B => DATAIN(22), S => n258, Z => n3485
                           );
   U2252 : MUX2_X1 port map( A => n2849, B => DATAIN(23), S => n258, Z => n3486
                           );
   U2253 : MUX2_X1 port map( A => n2826, B => DATAIN(24), S => n259, Z => n3487
                           );
   U2254 : MUX2_X1 port map( A => n2803, B => DATAIN(25), S => n259, Z => n3488
                           );
   U2255 : MUX2_X1 port map( A => n2780, B => DATAIN(26), S => n259, Z => n3489
                           );
   U2256 : MUX2_X1 port map( A => n2757, B => DATAIN(27), S => n259, Z => n3490
                           );
   U2257 : MUX2_X1 port map( A => n2734, B => DATAIN(28), S => n259, Z => n3491
                           );
   U2258 : MUX2_X1 port map( A => n2711, B => DATAIN(29), S => n259, Z => n3492
                           );
   U2259 : MUX2_X1 port map( A => n2688, B => DATAIN(30), S => n259, Z => n3493
                           );
   U2260 : MUX2_X1 port map( A => n2665, B => DATAIN(31), S => n259, Z => n3494
                           );
   U2261 : MUX2_X1 port map( A => n1811, B => DATAIN(0), S => n260, Z => n4318)
                           ;
   U2262 : MUX2_X1 port map( A => n1812, B => DATAIN(1), S => n260, Z => n4319)
                           ;
   U2263 : MUX2_X1 port map( A => n1813, B => DATAIN(2), S => n260, Z => n4320)
                           ;
   U2264 : MUX2_X1 port map( A => n1814, B => DATAIN(3), S => n260, Z => n4321)
                           ;
   U2265 : MUX2_X1 port map( A => n1815, B => DATAIN(4), S => n260, Z => n4322)
                           ;
   U2266 : MUX2_X1 port map( A => n1816, B => DATAIN(5), S => n260, Z => n4323)
                           ;
   U2267 : MUX2_X1 port map( A => n1817, B => DATAIN(6), S => n260, Z => n4324)
                           ;
   U2268 : MUX2_X1 port map( A => n1818, B => DATAIN(7), S => n260, Z => n4325)
                           ;
   U2269 : MUX2_X1 port map( A => n1819, B => DATAIN(8), S => n260, Z => n4326)
                           ;
   U2270 : MUX2_X1 port map( A => n1820, B => DATAIN(9), S => n260, Z => n4327)
                           ;
   U2271 : MUX2_X1 port map( A => n1821, B => DATAIN(10), S => n260, Z => n4328
                           );
   U2272 : MUX2_X1 port map( A => n1822, B => DATAIN(11), S => n260, Z => n4329
                           );
   U2273 : MUX2_X1 port map( A => n1823, B => DATAIN(12), S => n261, Z => n4330
                           );
   U2274 : MUX2_X1 port map( A => n1824, B => DATAIN(13), S => n261, Z => n4331
                           );
   U2275 : MUX2_X1 port map( A => n1825, B => DATAIN(14), S => n261, Z => n4332
                           );
   U2276 : MUX2_X1 port map( A => n1826, B => DATAIN(15), S => n261, Z => n4333
                           );
   U2277 : MUX2_X1 port map( A => n1827, B => DATAIN(16), S => n261, Z => n4334
                           );
   U2278 : MUX2_X1 port map( A => n1828, B => DATAIN(17), S => n261, Z => n4335
                           );
   U2279 : MUX2_X1 port map( A => n1829, B => DATAIN(18), S => n261, Z => n4336
                           );
   U2280 : MUX2_X1 port map( A => n1830, B => DATAIN(19), S => n261, Z => n4337
                           );
   U2281 : MUX2_X1 port map( A => n1831, B => DATAIN(20), S => n261, Z => n4338
                           );
   U2282 : MUX2_X1 port map( A => n1832, B => DATAIN(21), S => n261, Z => n4339
                           );
   U2283 : MUX2_X1 port map( A => n1833, B => DATAIN(22), S => n261, Z => n4340
                           );
   U2284 : MUX2_X1 port map( A => n1834, B => DATAIN(23), S => n261, Z => n4341
                           );
   U2285 : MUX2_X1 port map( A => n1835, B => DATAIN(24), S => n262, Z => n4342
                           );
   U2286 : MUX2_X1 port map( A => n1836, B => DATAIN(25), S => n262, Z => n4343
                           );
   U2287 : MUX2_X1 port map( A => n1837, B => DATAIN(26), S => n262, Z => n4344
                           );
   U2288 : MUX2_X1 port map( A => n1838, B => DATAIN(27), S => n262, Z => n4345
                           );
   U2289 : MUX2_X1 port map( A => n1839, B => DATAIN(28), S => n262, Z => n4346
                           );
   U2290 : MUX2_X1 port map( A => n1840, B => DATAIN(29), S => n262, Z => n4347
                           );
   U2291 : MUX2_X1 port map( A => n1841, B => DATAIN(30), S => n262, Z => n4348
                           );
   U2292 : MUX2_X1 port map( A => n1842, B => DATAIN(31), S => n262, Z => n4349
                           );
   U2293 : MUX2_X1 port map( A => n1843, B => DATAIN(0), S => n263, Z => n4286)
                           ;
   U2294 : MUX2_X1 port map( A => n1844, B => DATAIN(1), S => n263, Z => n4287)
                           ;
   U2295 : MUX2_X1 port map( A => n1845, B => DATAIN(2), S => n263, Z => n4288)
                           ;
   U2296 : MUX2_X1 port map( A => n1846, B => DATAIN(3), S => n263, Z => n4289)
                           ;
   U2297 : MUX2_X1 port map( A => n1847, B => DATAIN(4), S => n263, Z => n4290)
                           ;
   U2298 : MUX2_X1 port map( A => n1848, B => DATAIN(5), S => n263, Z => n4291)
                           ;
   U2299 : MUX2_X1 port map( A => n1849, B => DATAIN(6), S => n263, Z => n4292)
                           ;
   U2300 : MUX2_X1 port map( A => n1850, B => DATAIN(7), S => n263, Z => n4293)
                           ;
   U2301 : MUX2_X1 port map( A => n1851, B => DATAIN(8), S => n263, Z => n4294)
                           ;
   U2302 : MUX2_X1 port map( A => n1852, B => DATAIN(9), S => n263, Z => n4295)
                           ;
   U2303 : MUX2_X1 port map( A => n1853, B => DATAIN(10), S => n263, Z => n4296
                           );
   U2304 : MUX2_X1 port map( A => n1854, B => DATAIN(11), S => n263, Z => n4297
                           );
   U2305 : MUX2_X1 port map( A => n1855, B => DATAIN(12), S => n264, Z => n4298
                           );
   U2306 : MUX2_X1 port map( A => n1856, B => DATAIN(13), S => n264, Z => n4299
                           );
   U2307 : MUX2_X1 port map( A => n1857, B => DATAIN(14), S => n264, Z => n4300
                           );
   U2308 : MUX2_X1 port map( A => n1858, B => DATAIN(15), S => n264, Z => n4301
                           );
   U2309 : MUX2_X1 port map( A => n1859, B => DATAIN(16), S => n264, Z => n4302
                           );
   U2310 : MUX2_X1 port map( A => n1860, B => DATAIN(17), S => n264, Z => n4303
                           );
   U2311 : MUX2_X1 port map( A => n1861, B => DATAIN(18), S => n264, Z => n4304
                           );
   U2312 : MUX2_X1 port map( A => n1862, B => DATAIN(19), S => n264, Z => n4305
                           );
   U2313 : MUX2_X1 port map( A => n1863, B => DATAIN(20), S => n264, Z => n4306
                           );
   U2314 : MUX2_X1 port map( A => n1864, B => DATAIN(21), S => n264, Z => n4307
                           );
   U2315 : MUX2_X1 port map( A => n1865, B => DATAIN(22), S => n264, Z => n4308
                           );
   U2316 : MUX2_X1 port map( A => n1866, B => DATAIN(23), S => n264, Z => n4309
                           );
   U2317 : MUX2_X1 port map( A => n1867, B => DATAIN(24), S => n265, Z => n4310
                           );
   U2318 : MUX2_X1 port map( A => n1868, B => DATAIN(25), S => n265, Z => n4311
                           );
   U2319 : MUX2_X1 port map( A => n1869, B => DATAIN(26), S => n265, Z => n4312
                           );
   U2320 : MUX2_X1 port map( A => n1870, B => DATAIN(27), S => n265, Z => n4313
                           );
   U2321 : MUX2_X1 port map( A => n1871, B => DATAIN(28), S => n265, Z => n4314
                           );
   U2322 : MUX2_X1 port map( A => n1872, B => DATAIN(29), S => n265, Z => n4315
                           );
   U2323 : MUX2_X1 port map( A => n1873, B => DATAIN(30), S => n265, Z => n4316
                           );
   U2324 : MUX2_X1 port map( A => n1874, B => DATAIN(31), S => n265, Z => n4317
                           );
   U2325 : MUX2_X1 port map( A => n3955, B => DATAIN(0), S => n266, Z => n3495)
                           ;
   U2326 : MUX2_X1 port map( A => n3932, B => DATAIN(1), S => n266, Z => n3496)
                           ;
   U2327 : MUX2_X1 port map( A => n3909, B => DATAIN(2), S => n266, Z => n3497)
                           ;
   U2328 : MUX2_X1 port map( A => n3886, B => DATAIN(3), S => n266, Z => n3498)
                           ;
   U2329 : MUX2_X1 port map( A => n3863, B => DATAIN(4), S => n266, Z => n3499)
                           ;
   U2330 : MUX2_X1 port map( A => n3840, B => DATAIN(5), S => n266, Z => n3500)
                           ;
   U2331 : MUX2_X1 port map( A => n3817, B => DATAIN(6), S => n266, Z => n3501)
                           ;
   U2332 : MUX2_X1 port map( A => n3794, B => DATAIN(7), S => n266, Z => n3502)
                           ;
   U2333 : MUX2_X1 port map( A => n3771, B => DATAIN(8), S => n266, Z => n3503)
                           ;
   U2334 : MUX2_X1 port map( A => n3748, B => DATAIN(9), S => n266, Z => n3504)
                           ;
   U2335 : MUX2_X1 port map( A => n3725, B => DATAIN(10), S => n266, Z => n3505
                           );
   U2336 : MUX2_X1 port map( A => n3702, B => DATAIN(11), S => n266, Z => n3506
                           );
   U2337 : MUX2_X1 port map( A => n3679, B => DATAIN(12), S => n267, Z => n3507
                           );
   U2338 : MUX2_X1 port map( A => n3656, B => DATAIN(13), S => n267, Z => n3508
                           );
   U2339 : MUX2_X1 port map( A => n3633, B => DATAIN(14), S => n267, Z => n3509
                           );
   U2340 : MUX2_X1 port map( A => n3610, B => DATAIN(15), S => n267, Z => n3510
                           );
   U2341 : MUX2_X1 port map( A => n3587, B => DATAIN(16), S => n267, Z => n3511
                           );
   U2342 : MUX2_X1 port map( A => n3564, B => DATAIN(17), S => n267, Z => n3512
                           );
   U2343 : MUX2_X1 port map( A => n2965, B => DATAIN(18), S => n267, Z => n3513
                           );
   U2344 : MUX2_X1 port map( A => n2942, B => DATAIN(19), S => n267, Z => n3514
                           );
   U2345 : MUX2_X1 port map( A => n2919, B => DATAIN(20), S => n267, Z => n3515
                           );
   U2346 : MUX2_X1 port map( A => n2896, B => DATAIN(21), S => n267, Z => n3516
                           );
   U2347 : MUX2_X1 port map( A => n2873, B => DATAIN(22), S => n267, Z => n3517
                           );
   U2348 : MUX2_X1 port map( A => n2850, B => DATAIN(23), S => n267, Z => n3518
                           );
   U2349 : MUX2_X1 port map( A => n2827, B => DATAIN(24), S => n268, Z => n3519
                           );
   U2350 : MUX2_X1 port map( A => n2804, B => DATAIN(25), S => n268, Z => n3520
                           );
   U2351 : MUX2_X1 port map( A => n2781, B => DATAIN(26), S => n268, Z => n3521
                           );
   U2352 : MUX2_X1 port map( A => n2758, B => DATAIN(27), S => n268, Z => n3522
                           );
   U2353 : MUX2_X1 port map( A => n2735, B => DATAIN(28), S => n268, Z => n3523
                           );
   U2354 : MUX2_X1 port map( A => n2712, B => DATAIN(29), S => n268, Z => n3524
                           );
   U2355 : MUX2_X1 port map( A => n2689, B => DATAIN(30), S => n268, Z => n3525
                           );
   U2356 : MUX2_X1 port map( A => n2666, B => DATAIN(31), S => n268, Z => n3526
                           );
   U2357 : MUX2_X1 port map( A => n3956, B => DATAIN(0), S => n269, Z => n3527)
                           ;
   U2358 : MUX2_X1 port map( A => n3933, B => DATAIN(1), S => n269, Z => n3528)
                           ;
   U2359 : MUX2_X1 port map( A => n3910, B => DATAIN(2), S => n269, Z => n3529)
                           ;
   U2360 : MUX2_X1 port map( A => n3887, B => DATAIN(3), S => n269, Z => n3530)
                           ;
   U2361 : MUX2_X1 port map( A => n3864, B => DATAIN(4), S => n269, Z => n3531)
                           ;
   U2362 : MUX2_X1 port map( A => n3841, B => DATAIN(5), S => n269, Z => n3532)
                           ;
   U2363 : MUX2_X1 port map( A => n3818, B => DATAIN(6), S => n269, Z => n3533)
                           ;
   U2364 : MUX2_X1 port map( A => n3795, B => DATAIN(7), S => n269, Z => n3534)
                           ;
   U2365 : MUX2_X1 port map( A => n3772, B => DATAIN(8), S => n269, Z => n3535)
                           ;
   U2366 : MUX2_X1 port map( A => n3749, B => DATAIN(9), S => n269, Z => n3536)
                           ;
   U2367 : MUX2_X1 port map( A => n3726, B => DATAIN(10), S => n269, Z => n3537
                           );
   U2368 : MUX2_X1 port map( A => n3703, B => DATAIN(11), S => n269, Z => n3538
                           );
   U2369 : MUX2_X1 port map( A => n3680, B => DATAIN(12), S => n270, Z => n3539
                           );
   U2370 : MUX2_X1 port map( A => n3657, B => DATAIN(13), S => n270, Z => n3540
                           );
   U2371 : MUX2_X1 port map( A => n3634, B => DATAIN(14), S => n270, Z => n3541
                           );
   U2372 : MUX2_X1 port map( A => n3611, B => DATAIN(15), S => n270, Z => n3542
                           );
   U2373 : MUX2_X1 port map( A => n3588, B => DATAIN(16), S => n270, Z => n3543
                           );
   U2374 : MUX2_X1 port map( A => n3565, B => DATAIN(17), S => n270, Z => n3544
                           );
   U2375 : MUX2_X1 port map( A => n2966, B => DATAIN(18), S => n270, Z => n3545
                           );
   U2376 : MUX2_X1 port map( A => n2943, B => DATAIN(19), S => n270, Z => n3546
                           );
   U2377 : MUX2_X1 port map( A => n2920, B => DATAIN(20), S => n270, Z => n3547
                           );
   U2378 : MUX2_X1 port map( A => n2897, B => DATAIN(21), S => n270, Z => n3548
                           );
   U2379 : MUX2_X1 port map( A => n2874, B => DATAIN(22), S => n270, Z => n3549
                           );
   U2380 : MUX2_X1 port map( A => n2851, B => DATAIN(23), S => n270, Z => n3550
                           );
   U2381 : MUX2_X1 port map( A => n2828, B => DATAIN(24), S => n271, Z => n3551
                           );
   U2382 : MUX2_X1 port map( A => n2805, B => DATAIN(25), S => n271, Z => n3552
                           );
   U2383 : MUX2_X1 port map( A => n2782, B => DATAIN(26), S => n271, Z => n3553
                           );
   U2384 : MUX2_X1 port map( A => n2759, B => DATAIN(27), S => n271, Z => n3554
                           );
   U2385 : MUX2_X1 port map( A => n2736, B => DATAIN(28), S => n271, Z => n3555
                           );
   U2386 : MUX2_X1 port map( A => n2713, B => DATAIN(29), S => n271, Z => n3556
                           );
   U2387 : MUX2_X1 port map( A => n2690, B => DATAIN(30), S => n271, Z => n3557
                           );
   U2388 : MUX2_X1 port map( A => n2667, B => DATAIN(31), S => n271, Z => n3558
                           );
   U2389 : MUX2_X1 port map( A => n1875, B => DATAIN(0), S => n272, Z => n4254)
                           ;
   U2390 : MUX2_X1 port map( A => n1876, B => DATAIN(1), S => n272, Z => n4255)
                           ;
   U2391 : MUX2_X1 port map( A => n1877, B => DATAIN(2), S => n272, Z => n4256)
                           ;
   U2392 : MUX2_X1 port map( A => n1878, B => DATAIN(3), S => n272, Z => n4257)
                           ;
   U2393 : MUX2_X1 port map( A => n1879, B => DATAIN(4), S => n272, Z => n4258)
                           ;
   U2394 : MUX2_X1 port map( A => n1880, B => DATAIN(5), S => n272, Z => n4259)
                           ;
   U2395 : MUX2_X1 port map( A => n1881, B => DATAIN(6), S => n272, Z => n4260)
                           ;
   U2396 : MUX2_X1 port map( A => n1882, B => DATAIN(7), S => n272, Z => n4261)
                           ;
   U2397 : MUX2_X1 port map( A => n1883, B => DATAIN(8), S => n272, Z => n4262)
                           ;
   U2398 : MUX2_X1 port map( A => n1884, B => DATAIN(9), S => n272, Z => n4263)
                           ;
   U2399 : MUX2_X1 port map( A => n1885, B => DATAIN(10), S => n272, Z => n4264
                           );
   U2400 : MUX2_X1 port map( A => n1886, B => DATAIN(11), S => n272, Z => n4265
                           );
   U2401 : MUX2_X1 port map( A => n1887, B => DATAIN(12), S => n273, Z => n4266
                           );
   U2402 : MUX2_X1 port map( A => n1888, B => DATAIN(13), S => n273, Z => n4267
                           );
   U2403 : MUX2_X1 port map( A => n1889, B => DATAIN(14), S => n273, Z => n4268
                           );
   U2404 : MUX2_X1 port map( A => n1890, B => DATAIN(15), S => n273, Z => n4269
                           );
   U2405 : MUX2_X1 port map( A => n1891, B => DATAIN(16), S => n273, Z => n4270
                           );
   U2406 : MUX2_X1 port map( A => n1892, B => DATAIN(17), S => n273, Z => n4271
                           );
   U2407 : MUX2_X1 port map( A => n1893, B => DATAIN(18), S => n273, Z => n4272
                           );
   U2408 : MUX2_X1 port map( A => n1894, B => DATAIN(19), S => n273, Z => n4273
                           );
   U2409 : MUX2_X1 port map( A => n1895, B => DATAIN(20), S => n273, Z => n4274
                           );
   U2410 : MUX2_X1 port map( A => n1896, B => DATAIN(21), S => n273, Z => n4275
                           );
   U2411 : MUX2_X1 port map( A => n1897, B => DATAIN(22), S => n273, Z => n4276
                           );
   U2412 : MUX2_X1 port map( A => n1898, B => DATAIN(23), S => n273, Z => n4277
                           );
   U2413 : MUX2_X1 port map( A => n1899, B => DATAIN(24), S => n274, Z => n4278
                           );
   U2414 : MUX2_X1 port map( A => n1900, B => DATAIN(25), S => n274, Z => n4279
                           );
   U2415 : MUX2_X1 port map( A => n1901, B => DATAIN(26), S => n274, Z => n4280
                           );
   U2416 : MUX2_X1 port map( A => n1902, B => DATAIN(27), S => n274, Z => n4281
                           );
   U2417 : MUX2_X1 port map( A => n1903, B => DATAIN(28), S => n274, Z => n4282
                           );
   U2418 : MUX2_X1 port map( A => n1904, B => DATAIN(29), S => n274, Z => n4283
                           );
   U2419 : MUX2_X1 port map( A => n1905, B => DATAIN(30), S => n274, Z => n4284
                           );
   U2420 : MUX2_X1 port map( A => n1906, B => DATAIN(31), S => n274, Z => n4285
                           );
   U2421 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n1908);
   U2422 : OAI22_X1 port map( A1 => n3959, A2 => n277, B1 => n1922, B2 => n280,
                           ZN => n1920);
   U2423 : AOI221_X1 port map( B1 => n283, B2 => n3946, C1 => n286, C2 => n3947
                           , A => n1930, ZN => n1927);
   U2424 : OAI22_X1 port map( A1 => n3945, A2 => n289, B1 => n3944, B2 => n292,
                           ZN => n1930);
   U2425 : AOI221_X1 port map( B1 => n295, B2 => n3950, C1 => n298, C2 => n3951
                           , A => n1935, ZN => n1926);
   U2426 : OAI22_X1 port map( A1 => n3949, A2 => n301, B1 => n3948, B2 => n304,
                           ZN => n1935);
   U2427 : OAI22_X1 port map( A1 => n1940, A2 => n310, B1 => n1942, B2 => n313,
                           ZN => n1939);
   U2428 : OAI22_X1 port map( A1 => n1946, A2 => n319, B1 => n1948, B2 => n322,
                           ZN => n1945);
   U2429 : OAI22_X1 port map( A1 => n3936, A2 => n277, B1 => n1951, B2 => n280,
                           ZN => n1950);
   U2430 : AOI221_X1 port map( B1 => n283, B2 => n3923, C1 => n286, C2 => n3924
                           , A => n1954, ZN => n1953);
   U2431 : OAI22_X1 port map( A1 => n3922, A2 => n289, B1 => n3921, B2 => n292,
                           ZN => n1954);
   U2432 : AOI221_X1 port map( B1 => n295, B2 => n3927, C1 => n298, C2 => n3928
                           , A => n1955, ZN => n1952);
   U2433 : OAI22_X1 port map( A1 => n3926, A2 => n301, B1 => n3925, B2 => n304,
                           ZN => n1955);
   U2434 : OAI22_X1 port map( A1 => n1957, A2 => n310, B1 => n1958, B2 => n313,
                           ZN => n1956);
   U2435 : OAI22_X1 port map( A1 => n1960, A2 => n319, B1 => n1961, B2 => n322,
                           ZN => n1959);
   U2436 : OAI22_X1 port map( A1 => n3913, A2 => n277, B1 => n1963, B2 => n280,
                           ZN => n1962);
   U2437 : AOI221_X1 port map( B1 => n283, B2 => n3900, C1 => n286, C2 => n3901
                           , A => n1966, ZN => n1965);
   U2438 : OAI22_X1 port map( A1 => n3899, A2 => n289, B1 => n3898, B2 => n292,
                           ZN => n1966);
   U2439 : AOI221_X1 port map( B1 => n295, B2 => n3904, C1 => n298, C2 => n3905
                           , A => n1967, ZN => n1964);
   U2440 : OAI22_X1 port map( A1 => n3903, A2 => n301, B1 => n3902, B2 => n304,
                           ZN => n1967);
   U2441 : OAI22_X1 port map( A1 => n1969, A2 => n310, B1 => n1970, B2 => n313,
                           ZN => n1968);
   U2442 : OAI22_X1 port map( A1 => n1972, A2 => n319, B1 => n1973, B2 => n322,
                           ZN => n1971);
   U2443 : OAI22_X1 port map( A1 => n3890, A2 => n277, B1 => n1975, B2 => n280,
                           ZN => n1974);
   U2444 : AOI221_X1 port map( B1 => n283, B2 => n3877, C1 => n286, C2 => n3878
                           , A => n1978, ZN => n1977);
   U2445 : OAI22_X1 port map( A1 => n3876, A2 => n289, B1 => n3875, B2 => n292,
                           ZN => n1978);
   U2446 : AOI221_X1 port map( B1 => n295, B2 => n3881, C1 => n298, C2 => n3882
                           , A => n1979, ZN => n1976);
   U2447 : OAI22_X1 port map( A1 => n3880, A2 => n301, B1 => n3879, B2 => n304,
                           ZN => n1979);
   U2448 : OAI22_X1 port map( A1 => n1981, A2 => n310, B1 => n1982, B2 => n313,
                           ZN => n1980);
   U2449 : OAI22_X1 port map( A1 => n1984, A2 => n319, B1 => n1985, B2 => n322,
                           ZN => n1983);
   U2450 : OAI22_X1 port map( A1 => n3867, A2 => n277, B1 => n1987, B2 => n280,
                           ZN => n1986);
   U2451 : AOI221_X1 port map( B1 => n283, B2 => n3854, C1 => n286, C2 => n3855
                           , A => n1990, ZN => n1989);
   U2452 : OAI22_X1 port map( A1 => n3853, A2 => n289, B1 => n3852, B2 => n292,
                           ZN => n1990);
   U2453 : AOI221_X1 port map( B1 => n295, B2 => n3858, C1 => n298, C2 => n3859
                           , A => n1991, ZN => n1988);
   U2454 : OAI22_X1 port map( A1 => n3857, A2 => n301, B1 => n3856, B2 => n304,
                           ZN => n1991);
   U2455 : OAI22_X1 port map( A1 => n1993, A2 => n310, B1 => n1994, B2 => n313,
                           ZN => n1992);
   U2456 : OAI22_X1 port map( A1 => n1996, A2 => n319, B1 => n1997, B2 => n322,
                           ZN => n1995);
   U2457 : OAI22_X1 port map( A1 => n3844, A2 => n277, B1 => n1999, B2 => n280,
                           ZN => n1998);
   U2458 : AOI221_X1 port map( B1 => n283, B2 => n3831, C1 => n286, C2 => n3832
                           , A => n2002, ZN => n2001);
   U2459 : OAI22_X1 port map( A1 => n3830, A2 => n289, B1 => n3829, B2 => n292,
                           ZN => n2002);
   U2460 : AOI221_X1 port map( B1 => n295, B2 => n3835, C1 => n298, C2 => n3836
                           , A => n2003, ZN => n2000);
   U2461 : OAI22_X1 port map( A1 => n3834, A2 => n301, B1 => n3833, B2 => n304,
                           ZN => n2003);
   U2462 : OAI22_X1 port map( A1 => n2005, A2 => n310, B1 => n2006, B2 => n313,
                           ZN => n2004);
   U2463 : OAI22_X1 port map( A1 => n2008, A2 => n319, B1 => n2009, B2 => n322,
                           ZN => n2007);
   U2464 : OAI22_X1 port map( A1 => n3821, A2 => n277, B1 => n2011, B2 => n280,
                           ZN => n2010);
   U2465 : AOI221_X1 port map( B1 => n283, B2 => n3808, C1 => n286, C2 => n3809
                           , A => n2014, ZN => n2013);
   U2466 : OAI22_X1 port map( A1 => n3807, A2 => n289, B1 => n3806, B2 => n292,
                           ZN => n2014);
   U2467 : AOI221_X1 port map( B1 => n295, B2 => n3812, C1 => n298, C2 => n3813
                           , A => n2015, ZN => n2012);
   U2468 : OAI22_X1 port map( A1 => n3811, A2 => n301, B1 => n3810, B2 => n304,
                           ZN => n2015);
   U2469 : OAI22_X1 port map( A1 => n2017, A2 => n310, B1 => n2018, B2 => n313,
                           ZN => n2016);
   U2470 : OAI22_X1 port map( A1 => n2020, A2 => n319, B1 => n2021, B2 => n322,
                           ZN => n2019);
   U2471 : OAI22_X1 port map( A1 => n3798, A2 => n277, B1 => n2023, B2 => n280,
                           ZN => n2022);
   U2472 : AOI221_X1 port map( B1 => n283, B2 => n3785, C1 => n286, C2 => n3786
                           , A => n2026, ZN => n2025);
   U2473 : OAI22_X1 port map( A1 => n3784, A2 => n289, B1 => n3783, B2 => n292,
                           ZN => n2026);
   U2474 : AOI221_X1 port map( B1 => n295, B2 => n3789, C1 => n298, C2 => n3790
                           , A => n2027, ZN => n2024);
   U2475 : OAI22_X1 port map( A1 => n3788, A2 => n301, B1 => n3787, B2 => n304,
                           ZN => n2027);
   U2476 : OAI22_X1 port map( A1 => n2029, A2 => n310, B1 => n2030, B2 => n313,
                           ZN => n2028);
   U2477 : OAI22_X1 port map( A1 => n2032, A2 => n319, B1 => n2033, B2 => n322,
                           ZN => n2031);
   U2478 : OAI22_X1 port map( A1 => n3775, A2 => n276, B1 => n2035, B2 => n279,
                           ZN => n2034);
   U2479 : AOI221_X1 port map( B1 => n282, B2 => n3762, C1 => n285, C2 => n3763
                           , A => n2038, ZN => n2037);
   U2480 : OAI22_X1 port map( A1 => n3761, A2 => n288, B1 => n3760, B2 => n291,
                           ZN => n2038);
   U2481 : AOI221_X1 port map( B1 => n294, B2 => n3766, C1 => n297, C2 => n3767
                           , A => n2039, ZN => n2036);
   U2482 : OAI22_X1 port map( A1 => n3765, A2 => n300, B1 => n3764, B2 => n303,
                           ZN => n2039);
   U2483 : OAI22_X1 port map( A1 => n2041, A2 => n309, B1 => n2042, B2 => n312,
                           ZN => n2040);
   U2484 : OAI22_X1 port map( A1 => n2044, A2 => n318, B1 => n2045, B2 => n321,
                           ZN => n2043);
   U2485 : OAI22_X1 port map( A1 => n3752, A2 => n276, B1 => n2047, B2 => n279,
                           ZN => n2046);
   U2486 : AOI221_X1 port map( B1 => n282, B2 => n3739, C1 => n285, C2 => n3740
                           , A => n2050, ZN => n2049);
   U2487 : OAI22_X1 port map( A1 => n3738, A2 => n288, B1 => n3737, B2 => n291,
                           ZN => n2050);
   U2488 : AOI221_X1 port map( B1 => n294, B2 => n3743, C1 => n297, C2 => n3744
                           , A => n2051, ZN => n2048);
   U2489 : OAI22_X1 port map( A1 => n3742, A2 => n300, B1 => n3741, B2 => n303,
                           ZN => n2051);
   U2490 : OAI22_X1 port map( A1 => n2053, A2 => n309, B1 => n2054, B2 => n312,
                           ZN => n2052);
   U2491 : OAI22_X1 port map( A1 => n2056, A2 => n318, B1 => n2057, B2 => n321,
                           ZN => n2055);
   U2492 : OAI22_X1 port map( A1 => n3729, A2 => n276, B1 => n2059, B2 => n279,
                           ZN => n2058);
   U2493 : AOI221_X1 port map( B1 => n282, B2 => n3716, C1 => n285, C2 => n3717
                           , A => n2062, ZN => n2061);
   U2494 : OAI22_X1 port map( A1 => n3715, A2 => n288, B1 => n3714, B2 => n291,
                           ZN => n2062);
   U2495 : AOI221_X1 port map( B1 => n294, B2 => n3720, C1 => n297, C2 => n3721
                           , A => n2063, ZN => n2060);
   U2496 : OAI22_X1 port map( A1 => n3719, A2 => n300, B1 => n3718, B2 => n303,
                           ZN => n2063);
   U2497 : OAI22_X1 port map( A1 => n2065, A2 => n309, B1 => n2066, B2 => n312,
                           ZN => n2064);
   U2498 : OAI22_X1 port map( A1 => n2068, A2 => n318, B1 => n2069, B2 => n321,
                           ZN => n2067);
   U2499 : OAI22_X1 port map( A1 => n3706, A2 => n276, B1 => n2071, B2 => n279,
                           ZN => n2070);
   U2500 : AOI221_X1 port map( B1 => n282, B2 => n3693, C1 => n285, C2 => n3694
                           , A => n2074, ZN => n2073);
   U2501 : OAI22_X1 port map( A1 => n3692, A2 => n288, B1 => n3691, B2 => n291,
                           ZN => n2074);
   U2502 : AOI221_X1 port map( B1 => n294, B2 => n3697, C1 => n297, C2 => n3698
                           , A => n2075, ZN => n2072);
   U2503 : OAI22_X1 port map( A1 => n3696, A2 => n300, B1 => n3695, B2 => n303,
                           ZN => n2075);
   U2504 : OAI22_X1 port map( A1 => n2077, A2 => n309, B1 => n2078, B2 => n312,
                           ZN => n2076);
   U2505 : OAI22_X1 port map( A1 => n2080, A2 => n318, B1 => n2081, B2 => n321,
                           ZN => n2079);
   U2506 : OAI22_X1 port map( A1 => n3683, A2 => n276, B1 => n2083, B2 => n279,
                           ZN => n2082);
   U2507 : AOI221_X1 port map( B1 => n282, B2 => n3670, C1 => n285, C2 => n3671
                           , A => n2086, ZN => n2085);
   U2508 : OAI22_X1 port map( A1 => n3669, A2 => n288, B1 => n3668, B2 => n291,
                           ZN => n2086);
   U2509 : AOI221_X1 port map( B1 => n294, B2 => n3674, C1 => n297, C2 => n3675
                           , A => n2087, ZN => n2084);
   U2510 : OAI22_X1 port map( A1 => n3673, A2 => n300, B1 => n3672, B2 => n303,
                           ZN => n2087);
   U2511 : OAI22_X1 port map( A1 => n2089, A2 => n309, B1 => n2090, B2 => n312,
                           ZN => n2088);
   U2512 : OAI22_X1 port map( A1 => n2092, A2 => n318, B1 => n2093, B2 => n321,
                           ZN => n2091);
   U2513 : OAI22_X1 port map( A1 => n3660, A2 => n276, B1 => n2095, B2 => n279,
                           ZN => n2094);
   U2514 : AOI221_X1 port map( B1 => n282, B2 => n3647, C1 => n285, C2 => n3648
                           , A => n2098, ZN => n2097);
   U2515 : OAI22_X1 port map( A1 => n3646, A2 => n288, B1 => n3645, B2 => n291,
                           ZN => n2098);
   U2516 : AOI221_X1 port map( B1 => n294, B2 => n3651, C1 => n297, C2 => n3652
                           , A => n2099, ZN => n2096);
   U2517 : OAI22_X1 port map( A1 => n3650, A2 => n300, B1 => n3649, B2 => n303,
                           ZN => n2099);
   U2518 : OAI22_X1 port map( A1 => n2101, A2 => n309, B1 => n2102, B2 => n312,
                           ZN => n2100);
   U2519 : OAI22_X1 port map( A1 => n2104, A2 => n318, B1 => n2105, B2 => n321,
                           ZN => n2103);
   U2520 : OAI22_X1 port map( A1 => n3637, A2 => n276, B1 => n2107, B2 => n279,
                           ZN => n2106);
   U2521 : AOI221_X1 port map( B1 => n282, B2 => n3624, C1 => n285, C2 => n3625
                           , A => n2110, ZN => n2109);
   U2522 : OAI22_X1 port map( A1 => n3623, A2 => n288, B1 => n3622, B2 => n291,
                           ZN => n2110);
   U2523 : AOI221_X1 port map( B1 => n294, B2 => n3628, C1 => n297, C2 => n3629
                           , A => n2111, ZN => n2108);
   U2524 : OAI22_X1 port map( A1 => n3627, A2 => n300, B1 => n3626, B2 => n303,
                           ZN => n2111);
   U2525 : OAI22_X1 port map( A1 => n2113, A2 => n309, B1 => n2114, B2 => n312,
                           ZN => n2112);
   U2526 : OAI22_X1 port map( A1 => n2116, A2 => n318, B1 => n2117, B2 => n321,
                           ZN => n2115);
   U2527 : OAI22_X1 port map( A1 => n3614, A2 => n276, B1 => n2119, B2 => n279,
                           ZN => n2118);
   U2528 : AOI221_X1 port map( B1 => n282, B2 => n3601, C1 => n285, C2 => n3602
                           , A => n2122, ZN => n2121);
   U2529 : OAI22_X1 port map( A1 => n3600, A2 => n288, B1 => n3599, B2 => n291,
                           ZN => n2122);
   U2530 : AOI221_X1 port map( B1 => n294, B2 => n3605, C1 => n297, C2 => n3606
                           , A => n2123, ZN => n2120);
   U2531 : OAI22_X1 port map( A1 => n3604, A2 => n300, B1 => n3603, B2 => n303,
                           ZN => n2123);
   U2532 : OAI22_X1 port map( A1 => n2125, A2 => n309, B1 => n2126, B2 => n312,
                           ZN => n2124);
   U2533 : OAI22_X1 port map( A1 => n2128, A2 => n318, B1 => n2129, B2 => n321,
                           ZN => n2127);
   U2534 : OAI22_X1 port map( A1 => n3591, A2 => n276, B1 => n2131, B2 => n279,
                           ZN => n2130);
   U2535 : AOI221_X1 port map( B1 => n282, B2 => n3578, C1 => n285, C2 => n3579
                           , A => n2134, ZN => n2133);
   U2536 : OAI22_X1 port map( A1 => n3577, A2 => n288, B1 => n3576, B2 => n291,
                           ZN => n2134);
   U2537 : AOI221_X1 port map( B1 => n294, B2 => n3582, C1 => n297, C2 => n3583
                           , A => n2135, ZN => n2132);
   U2538 : OAI22_X1 port map( A1 => n3581, A2 => n300, B1 => n3580, B2 => n303,
                           ZN => n2135);
   U2539 : OAI22_X1 port map( A1 => n2137, A2 => n309, B1 => n2138, B2 => n312,
                           ZN => n2136);
   U2540 : OAI22_X1 port map( A1 => n2140, A2 => n318, B1 => n2141, B2 => n321,
                           ZN => n2139);
   U2541 : OAI22_X1 port map( A1 => n3568, A2 => n276, B1 => n2143, B2 => n279,
                           ZN => n2142);
   U2542 : AOI221_X1 port map( B1 => n282, B2 => n2979, C1 => n285, C2 => n2980
                           , A => n2146, ZN => n2145);
   U2543 : OAI22_X1 port map( A1 => n2978, A2 => n288, B1 => n2977, B2 => n291,
                           ZN => n2146);
   U2544 : AOI221_X1 port map( B1 => n294, B2 => n3559, C1 => n297, C2 => n3560
                           , A => n2147, ZN => n2144);
   U2545 : OAI22_X1 port map( A1 => n2982, A2 => n300, B1 => n2981, B2 => n303,
                           ZN => n2147);
   U2546 : OAI22_X1 port map( A1 => n2149, A2 => n309, B1 => n2150, B2 => n312,
                           ZN => n2148);
   U2547 : OAI22_X1 port map( A1 => n2152, A2 => n318, B1 => n2153, B2 => n321,
                           ZN => n2151);
   U2548 : OAI22_X1 port map( A1 => n2969, A2 => n276, B1 => n2155, B2 => n279,
                           ZN => n2154);
   U2549 : AOI221_X1 port map( B1 => n282, B2 => n2956, C1 => n285, C2 => n2957
                           , A => n2158, ZN => n2157);
   U2550 : OAI22_X1 port map( A1 => n2955, A2 => n288, B1 => n2954, B2 => n291,
                           ZN => n2158);
   U2551 : AOI221_X1 port map( B1 => n294, B2 => n2960, C1 => n297, C2 => n2961
                           , A => n2159, ZN => n2156);
   U2552 : OAI22_X1 port map( A1 => n2959, A2 => n300, B1 => n2958, B2 => n303,
                           ZN => n2159);
   U2553 : OAI22_X1 port map( A1 => n2161, A2 => n309, B1 => n2162, B2 => n312,
                           ZN => n2160);
   U2554 : OAI22_X1 port map( A1 => n2164, A2 => n318, B1 => n2165, B2 => n321,
                           ZN => n2163);
   U2555 : OAI22_X1 port map( A1 => n2946, A2 => n276, B1 => n2167, B2 => n279,
                           ZN => n2166);
   U2556 : AOI221_X1 port map( B1 => n282, B2 => n2933, C1 => n285, C2 => n2934
                           , A => n2170, ZN => n2169);
   U2557 : OAI22_X1 port map( A1 => n2932, A2 => n288, B1 => n2931, B2 => n291,
                           ZN => n2170);
   U2558 : AOI221_X1 port map( B1 => n294, B2 => n2937, C1 => n297, C2 => n2938
                           , A => n2171, ZN => n2168);
   U2559 : OAI22_X1 port map( A1 => n2936, A2 => n300, B1 => n2935, B2 => n303,
                           ZN => n2171);
   U2560 : OAI22_X1 port map( A1 => n2173, A2 => n309, B1 => n2174, B2 => n312,
                           ZN => n2172);
   U2561 : OAI22_X1 port map( A1 => n2176, A2 => n318, B1 => n2177, B2 => n321,
                           ZN => n2175);
   U2562 : OAI22_X1 port map( A1 => n2923, A2 => n275, B1 => n2179, B2 => n278,
                           ZN => n2178);
   U2563 : AOI221_X1 port map( B1 => n281, B2 => n2910, C1 => n284, C2 => n2911
                           , A => n2182, ZN => n2181);
   U2564 : OAI22_X1 port map( A1 => n2909, A2 => n287, B1 => n2908, B2 => n290,
                           ZN => n2182);
   U2565 : AOI221_X1 port map( B1 => n293, B2 => n2914, C1 => n296, C2 => n2915
                           , A => n2183, ZN => n2180);
   U2566 : OAI22_X1 port map( A1 => n2913, A2 => n299, B1 => n2912, B2 => n302,
                           ZN => n2183);
   U2567 : OAI22_X1 port map( A1 => n2185, A2 => n308, B1 => n2186, B2 => n311,
                           ZN => n2184);
   U2568 : OAI22_X1 port map( A1 => n2188, A2 => n317, B1 => n2189, B2 => n320,
                           ZN => n2187);
   U2569 : OAI22_X1 port map( A1 => n2900, A2 => n275, B1 => n2191, B2 => n278,
                           ZN => n2190);
   U2570 : AOI221_X1 port map( B1 => n281, B2 => n2887, C1 => n284, C2 => n2888
                           , A => n2194, ZN => n2193);
   U2571 : OAI22_X1 port map( A1 => n2886, A2 => n287, B1 => n2885, B2 => n290,
                           ZN => n2194);
   U2572 : AOI221_X1 port map( B1 => n293, B2 => n2891, C1 => n296, C2 => n2892
                           , A => n2195, ZN => n2192);
   U2573 : OAI22_X1 port map( A1 => n2890, A2 => n299, B1 => n2889, B2 => n302,
                           ZN => n2195);
   U2574 : OAI22_X1 port map( A1 => n2197, A2 => n308, B1 => n2198, B2 => n311,
                           ZN => n2196);
   U2575 : OAI22_X1 port map( A1 => n2200, A2 => n317, B1 => n2201, B2 => n320,
                           ZN => n2199);
   U2576 : OAI22_X1 port map( A1 => n2877, A2 => n275, B1 => n2203, B2 => n278,
                           ZN => n2202);
   U2577 : AOI221_X1 port map( B1 => n281, B2 => n2864, C1 => n284, C2 => n2865
                           , A => n2206, ZN => n2205);
   U2578 : OAI22_X1 port map( A1 => n2863, A2 => n287, B1 => n2862, B2 => n290,
                           ZN => n2206);
   U2579 : AOI221_X1 port map( B1 => n293, B2 => n2868, C1 => n296, C2 => n2869
                           , A => n2207, ZN => n2204);
   U2580 : OAI22_X1 port map( A1 => n2867, A2 => n299, B1 => n2866, B2 => n302,
                           ZN => n2207);
   U2581 : OAI22_X1 port map( A1 => n2209, A2 => n308, B1 => n2210, B2 => n311,
                           ZN => n2208);
   U2582 : OAI22_X1 port map( A1 => n2212, A2 => n317, B1 => n2213, B2 => n320,
                           ZN => n2211);
   U2583 : OAI22_X1 port map( A1 => n2854, A2 => n275, B1 => n2215, B2 => n278,
                           ZN => n2214);
   U2584 : AOI221_X1 port map( B1 => n281, B2 => n2841, C1 => n284, C2 => n2842
                           , A => n2218, ZN => n2217);
   U2585 : OAI22_X1 port map( A1 => n2840, A2 => n287, B1 => n2839, B2 => n290,
                           ZN => n2218);
   U2586 : AOI221_X1 port map( B1 => n293, B2 => n2845, C1 => n296, C2 => n2846
                           , A => n2219, ZN => n2216);
   U2587 : OAI22_X1 port map( A1 => n2844, A2 => n299, B1 => n2843, B2 => n302,
                           ZN => n2219);
   U2588 : OAI22_X1 port map( A1 => n2221, A2 => n308, B1 => n2222, B2 => n311,
                           ZN => n2220);
   U2589 : OAI22_X1 port map( A1 => n2224, A2 => n317, B1 => n2225, B2 => n320,
                           ZN => n2223);
   U2590 : OAI22_X1 port map( A1 => n2831, A2 => n275, B1 => n2227, B2 => n278,
                           ZN => n2226);
   U2591 : AOI221_X1 port map( B1 => n281, B2 => n2818, C1 => n284, C2 => n2819
                           , A => n2230, ZN => n2229);
   U2592 : OAI22_X1 port map( A1 => n2817, A2 => n287, B1 => n2816, B2 => n290,
                           ZN => n2230);
   U2593 : AOI221_X1 port map( B1 => n293, B2 => n2822, C1 => n296, C2 => n2823
                           , A => n2231, ZN => n2228);
   U2594 : OAI22_X1 port map( A1 => n2821, A2 => n299, B1 => n2820, B2 => n302,
                           ZN => n2231);
   U2595 : OAI22_X1 port map( A1 => n2233, A2 => n308, B1 => n2234, B2 => n311,
                           ZN => n2232);
   U2596 : OAI22_X1 port map( A1 => n2236, A2 => n317, B1 => n2237, B2 => n320,
                           ZN => n2235);
   U2597 : OAI22_X1 port map( A1 => n2808, A2 => n275, B1 => n2239, B2 => n278,
                           ZN => n2238);
   U2598 : AOI221_X1 port map( B1 => n281, B2 => n2795, C1 => n284, C2 => n2796
                           , A => n2242, ZN => n2241);
   U2599 : OAI22_X1 port map( A1 => n2794, A2 => n287, B1 => n2793, B2 => n290,
                           ZN => n2242);
   U2600 : AOI221_X1 port map( B1 => n293, B2 => n2799, C1 => n296, C2 => n2800
                           , A => n2243, ZN => n2240);
   U2601 : OAI22_X1 port map( A1 => n2798, A2 => n299, B1 => n2797, B2 => n302,
                           ZN => n2243);
   U2602 : OAI22_X1 port map( A1 => n2245, A2 => n308, B1 => n2246, B2 => n311,
                           ZN => n2244);
   U2603 : OAI22_X1 port map( A1 => n2248, A2 => n317, B1 => n2249, B2 => n320,
                           ZN => n2247);
   U2604 : OAI22_X1 port map( A1 => n2785, A2 => n275, B1 => n2251, B2 => n278,
                           ZN => n2250);
   U2605 : AOI221_X1 port map( B1 => n281, B2 => n2772, C1 => n284, C2 => n2773
                           , A => n2254, ZN => n2253);
   U2606 : OAI22_X1 port map( A1 => n2771, A2 => n287, B1 => n2770, B2 => n290,
                           ZN => n2254);
   U2607 : AOI221_X1 port map( B1 => n293, B2 => n2776, C1 => n296, C2 => n2777
                           , A => n2255, ZN => n2252);
   U2608 : OAI22_X1 port map( A1 => n2775, A2 => n299, B1 => n2774, B2 => n302,
                           ZN => n2255);
   U2609 : OAI22_X1 port map( A1 => n2257, A2 => n308, B1 => n2258, B2 => n311,
                           ZN => n2256);
   U2610 : OAI22_X1 port map( A1 => n2260, A2 => n317, B1 => n2261, B2 => n320,
                           ZN => n2259);
   U2611 : OAI22_X1 port map( A1 => n2762, A2 => n275, B1 => n2263, B2 => n278,
                           ZN => n2262);
   U2612 : AOI221_X1 port map( B1 => n281, B2 => n2749, C1 => n284, C2 => n2750
                           , A => n2266, ZN => n2265);
   U2613 : OAI22_X1 port map( A1 => n2748, A2 => n287, B1 => n2747, B2 => n290,
                           ZN => n2266);
   U2614 : AOI221_X1 port map( B1 => n293, B2 => n2753, C1 => n296, C2 => n2754
                           , A => n2267, ZN => n2264);
   U2615 : OAI22_X1 port map( A1 => n2752, A2 => n299, B1 => n2751, B2 => n302,
                           ZN => n2267);
   U2616 : OAI22_X1 port map( A1 => n2269, A2 => n308, B1 => n2270, B2 => n311,
                           ZN => n2268);
   U2617 : OAI22_X1 port map( A1 => n2272, A2 => n317, B1 => n2273, B2 => n320,
                           ZN => n2271);
   U2618 : OAI22_X1 port map( A1 => n2739, A2 => n275, B1 => n2275, B2 => n278,
                           ZN => n2274);
   U2619 : AOI221_X1 port map( B1 => n281, B2 => n2726, C1 => n284, C2 => n2727
                           , A => n2278, ZN => n2277);
   U2620 : OAI22_X1 port map( A1 => n2725, A2 => n287, B1 => n2724, B2 => n290,
                           ZN => n2278);
   U2621 : AOI221_X1 port map( B1 => n293, B2 => n2730, C1 => n296, C2 => n2731
                           , A => n2279, ZN => n2276);
   U2622 : OAI22_X1 port map( A1 => n2729, A2 => n299, B1 => n2728, B2 => n302,
                           ZN => n2279);
   U2623 : OAI22_X1 port map( A1 => n2281, A2 => n308, B1 => n2282, B2 => n311,
                           ZN => n2280);
   U2624 : OAI22_X1 port map( A1 => n2284, A2 => n317, B1 => n2285, B2 => n320,
                           ZN => n2283);
   U2625 : OAI22_X1 port map( A1 => n2716, A2 => n275, B1 => n2287, B2 => n278,
                           ZN => n2286);
   U2626 : AOI221_X1 port map( B1 => n281, B2 => n2703, C1 => n284, C2 => n2704
                           , A => n2290, ZN => n2289);
   U2627 : OAI22_X1 port map( A1 => n2702, A2 => n287, B1 => n2701, B2 => n290,
                           ZN => n2290);
   U2628 : AOI221_X1 port map( B1 => n293, B2 => n2707, C1 => n296, C2 => n2708
                           , A => n2291, ZN => n2288);
   U2629 : OAI22_X1 port map( A1 => n2706, A2 => n299, B1 => n2705, B2 => n302,
                           ZN => n2291);
   U2630 : OAI22_X1 port map( A1 => n2293, A2 => n308, B1 => n2294, B2 => n311,
                           ZN => n2292);
   U2631 : OAI22_X1 port map( A1 => n2296, A2 => n317, B1 => n2297, B2 => n320,
                           ZN => n2295);
   U2632 : OAI22_X1 port map( A1 => n2693, A2 => n275, B1 => n2299, B2 => n278,
                           ZN => n2298);
   U2633 : AOI221_X1 port map( B1 => n281, B2 => n2680, C1 => n284, C2 => n2681
                           , A => n2302, ZN => n2301);
   U2634 : OAI22_X1 port map( A1 => n2679, A2 => n287, B1 => n2678, B2 => n290,
                           ZN => n2302);
   U2635 : AOI221_X1 port map( B1 => n293, B2 => n2684, C1 => n296, C2 => n2685
                           , A => n2303, ZN => n2300);
   U2636 : OAI22_X1 port map( A1 => n2683, A2 => n299, B1 => n2682, B2 => n302,
                           ZN => n2303);
   U2637 : OAI22_X1 port map( A1 => n2305, A2 => n308, B1 => n2306, B2 => n311,
                           ZN => n2304);
   U2638 : OAI22_X1 port map( A1 => n2308, A2 => n317, B1 => n2309, B2 => n320,
                           ZN => n2307);
   U2639 : AND2_X1 port map( A1 => n2310, A2 => n2311, ZN => n1912);
   U2640 : AND2_X1 port map( A1 => n2310, A2 => n2312, ZN => n1911);
   U2641 : NAND2_X1 port map( A1 => n2313, A2 => n2314, ZN => n1910);
   U2642 : NAND2_X1 port map( A1 => n2315, A2 => n2311, ZN => n1909);
   U2643 : AND2_X1 port map( A1 => n2315, A2 => n2312, ZN => n1916);
   U2644 : AND2_X1 port map( A1 => n2315, A2 => n2314, ZN => n1915);
   U2645 : NAND2_X1 port map( A1 => n2310, A2 => n2314, ZN => n1914);
   U2646 : NAND2_X1 port map( A1 => n2310, A2 => n2316, ZN => n1913);
   U2647 : NOR3_X1 port map( A1 => n2317, A2 => ADD_RS2(0), A3 => n2318, ZN => 
                           n2310);
   U2648 : OAI22_X1 port map( A1 => n2670, A2 => n275, B1 => n2320, B2 => n278,
                           ZN => n2319);
   U2649 : NAND2_X1 port map( A1 => n2321, A2 => n2314, ZN => n1923);
   U2650 : NAND2_X1 port map( A1 => n2321, A2 => n2316, ZN => n1921);
   U2651 : AND2_X1 port map( A1 => n2313, A2 => n2311, ZN => n1919);
   U2652 : AND2_X1 port map( A1 => n2313, A2 => n2316, ZN => n1918);
   U2653 : AND2_X1 port map( A1 => n2321, A2 => n2312, ZN => n1925);
   U2654 : AND2_X1 port map( A1 => n2321, A2 => n2311, ZN => n1924);
   U2655 : NOR3_X1 port map( A1 => ADD_RS2(0), A2 => ADD_RS2(3), A3 => n2317, 
                           ZN => n2321);
   U2656 : NAND2_X1 port map( A1 => n2313, A2 => n2312, ZN => n1917);
   U2657 : NOR3_X1 port map( A1 => n2322, A2 => ADD_RS2(3), A3 => n2317, ZN => 
                           n2313);
   U2658 : AOI221_X1 port map( B1 => n281, B2 => n2657, C1 => n284, C2 => n2658
                           , A => n2325, ZN => n2324);
   U2659 : OAI22_X1 port map( A1 => n2656, A2 => n287, B1 => n2655, B2 => n290,
                           ZN => n2325);
   U2660 : NAND2_X1 port map( A1 => n2316, A2 => n2326, ZN => n1932);
   U2661 : NAND2_X1 port map( A1 => n2316, A2 => n2327, ZN => n1931);
   U2662 : AND2_X1 port map( A1 => n2326, A2 => n2314, ZN => n1929);
   U2663 : AND2_X1 port map( A1 => n2314, A2 => n2327, ZN => n1928);
   U2664 : AOI221_X1 port map( B1 => n293, B2 => n2661, C1 => n296, C2 => n2662
                           , A => n2328, ZN => n2323);
   U2665 : OAI22_X1 port map( A1 => n2660, A2 => n299, B1 => n2659, B2 => n302,
                           ZN => n2328);
   U2666 : NAND2_X1 port map( A1 => n2312, A2 => n2326, ZN => n1937);
   U2667 : NAND2_X1 port map( A1 => n2312, A2 => n2327, ZN => n1936);
   U2668 : AND2_X1 port map( A1 => n2311, A2 => n2326, ZN => n1934);
   U2669 : NOR3_X1 port map( A1 => ADD_RS2(0), A2 => ADD_RS2(4), A3 => n2318, 
                           ZN => n2326);
   U2670 : AND2_X1 port map( A1 => n2311, A2 => n2327, ZN => n1933);
   U2671 : NOR3_X1 port map( A1 => n2322, A2 => ADD_RS2(4), A3 => n2318, ZN => 
                           n2327);
   U2672 : OAI22_X1 port map( A1 => n2330, A2 => n308, B1 => n2331, B2 => n311,
                           ZN => n2329);
   U2673 : NAND2_X1 port map( A1 => n2332, A2 => n2314, ZN => n1943);
   U2674 : NAND2_X1 port map( A1 => n2333, A2 => n2314, ZN => n1941);
   U2675 : NOR2_X1 port map( A1 => n2334, A2 => n2335, ZN => n2314);
   U2676 : AND2_X1 port map( A1 => n2333, A2 => n2316, ZN => n1938);
   U2677 : OAI22_X1 port map( A1 => n2337, A2 => n317, B1 => n2338, B2 => n320,
                           ZN => n2336);
   U2678 : NAND2_X1 port map( A1 => n2332, A2 => n2311, ZN => n1949);
   U2679 : NAND2_X1 port map( A1 => n2333, A2 => n2311, ZN => n1947);
   U2680 : NOR2_X1 port map( A1 => n2335, A2 => ADD_RS2(2), ZN => n2311);
   U2681 : NOR3_X1 port map( A1 => ADD_RS2(3), A2 => ADD_RS2(4), A3 => 
                           ADD_RS2(0), ZN => n2333);
   U2682 : AND2_X1 port map( A1 => n2315, A2 => n2316, ZN => n1944);
   U2683 : NOR2_X1 port map( A1 => n2334, A2 => ADD_RS2(1), ZN => n2316);
   U2684 : INV_X1 port map( A => ADD_RS2(2), ZN => n2334);
   U2685 : NOR3_X1 port map( A1 => n2317, A2 => n2322, A3 => n2318, ZN => n2315
                           );
   U2686 : INV_X1 port map( A => ADD_RS2(3), ZN => n2318);
   U2687 : INV_X1 port map( A => ADD_RS2(4), ZN => n2317);
   U2688 : NOR2_X1 port map( A1 => ADD_RS2(1), A2 => ADD_RS2(2), ZN => n2312);
   U2689 : NOR3_X1 port map( A1 => ADD_RS2(3), A2 => ADD_RS2(4), A3 => n2322, 
                           ZN => n2332);
   U2690 : INV_X1 port map( A => ADD_RS2(0), ZN => n2322);
   U2691 : NOR3_X1 port map( A1 => n2343, A2 => n2344, A3 => n2345, ZN => n2342
                           );
   U2692 : XNOR2_X1 port map( A => ADD_WR(1), B => n2335, ZN => n2345);
   U2693 : INV_X1 port map( A => ADD_RS2(1), ZN => n2335);
   U2694 : XNOR2_X1 port map( A => n1907, B => ADD_RS2(0), ZN => n2343);
   U2695 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS2(3), ZN => n2341);
   U2696 : XNOR2_X1 port map( A => ADD_WR(4), B => ADD_RS2(4), ZN => n2340);
   U2697 : XNOR2_X1 port map( A => ADD_RS2(2), B => ADD_WR(2), ZN => n2339);
   U2698 : OAI22_X1 port map( A1 => n2670, A2 => n325, B1 => n2320, B2 => n328,
                           ZN => n2357);
   U2699 : AOI221_X1 port map( B1 => n331, B2 => n2657, C1 => n334, C2 => n2658
                           , A => n2366, ZN => n2363);
   U2700 : OAI22_X1 port map( A1 => n2656, A2 => n337, B1 => n2655, B2 => n340,
                           ZN => n2366);
   U2701 : AOI221_X1 port map( B1 => n343, B2 => n2661, C1 => n346, C2 => n2662
                           , A => n2371, ZN => n2362);
   U2702 : OAI22_X1 port map( A1 => n2660, A2 => n349, B1 => n2659, B2 => n352,
                           ZN => n2371);
   U2703 : OAI22_X1 port map( A1 => n2330, A2 => n358, B1 => n2331, B2 => n361,
                           ZN => n2375);
   U2704 : OAI22_X1 port map( A1 => n2337, A2 => n367, B1 => n2338, B2 => n370,
                           ZN => n2379);
   U2705 : OAI22_X1 port map( A1 => n2693, A2 => n325, B1 => n2299, B2 => n328,
                           ZN => n2382);
   U2706 : AOI221_X1 port map( B1 => n331, B2 => n2680, C1 => n334, C2 => n2681
                           , A => n2385, ZN => n2384);
   U2707 : OAI22_X1 port map( A1 => n2679, A2 => n337, B1 => n2678, B2 => n340,
                           ZN => n2385);
   U2708 : AOI221_X1 port map( B1 => n343, B2 => n2684, C1 => n346, C2 => n2685
                           , A => n2386, ZN => n2383);
   U2709 : OAI22_X1 port map( A1 => n2683, A2 => n349, B1 => n2682, B2 => n352,
                           ZN => n2386);
   U2710 : OAI22_X1 port map( A1 => n2305, A2 => n358, B1 => n2306, B2 => n361,
                           ZN => n2387);
   U2711 : OAI22_X1 port map( A1 => n2308, A2 => n367, B1 => n2309, B2 => n370,
                           ZN => n2388);
   U2712 : OAI22_X1 port map( A1 => n2716, A2 => n325, B1 => n2287, B2 => n328,
                           ZN => n2389);
   U2713 : AOI221_X1 port map( B1 => n331, B2 => n2703, C1 => n334, C2 => n2704
                           , A => n2392, ZN => n2391);
   U2714 : OAI22_X1 port map( A1 => n2702, A2 => n337, B1 => n2701, B2 => n340,
                           ZN => n2392);
   U2715 : AOI221_X1 port map( B1 => n343, B2 => n2707, C1 => n346, C2 => n2708
                           , A => n2393, ZN => n2390);
   U2716 : OAI22_X1 port map( A1 => n2706, A2 => n349, B1 => n2705, B2 => n352,
                           ZN => n2393);
   U2717 : OAI22_X1 port map( A1 => n2293, A2 => n358, B1 => n2294, B2 => n361,
                           ZN => n2394);
   U2718 : OAI22_X1 port map( A1 => n2296, A2 => n367, B1 => n2297, B2 => n370,
                           ZN => n2395);
   U2719 : OAI22_X1 port map( A1 => n2739, A2 => n325, B1 => n2275, B2 => n328,
                           ZN => n2396);
   U2720 : AOI221_X1 port map( B1 => n331, B2 => n2726, C1 => n334, C2 => n2727
                           , A => n2399, ZN => n2398);
   U2721 : OAI22_X1 port map( A1 => n2725, A2 => n337, B1 => n2724, B2 => n340,
                           ZN => n2399);
   U2722 : AOI221_X1 port map( B1 => n343, B2 => n2730, C1 => n346, C2 => n2731
                           , A => n2400, ZN => n2397);
   U2723 : OAI22_X1 port map( A1 => n2729, A2 => n349, B1 => n2728, B2 => n352,
                           ZN => n2400);
   U2724 : OAI22_X1 port map( A1 => n2281, A2 => n358, B1 => n2282, B2 => n361,
                           ZN => n2401);
   U2725 : OAI22_X1 port map( A1 => n2284, A2 => n367, B1 => n2285, B2 => n370,
                           ZN => n2402);
   U2726 : OAI22_X1 port map( A1 => n2762, A2 => n325, B1 => n2263, B2 => n328,
                           ZN => n2403);
   U2727 : AOI221_X1 port map( B1 => n331, B2 => n2749, C1 => n334, C2 => n2750
                           , A => n2406, ZN => n2405);
   U2728 : OAI22_X1 port map( A1 => n2748, A2 => n337, B1 => n2747, B2 => n340,
                           ZN => n2406);
   U2729 : AOI221_X1 port map( B1 => n343, B2 => n2753, C1 => n346, C2 => n2754
                           , A => n2407, ZN => n2404);
   U2730 : OAI22_X1 port map( A1 => n2752, A2 => n349, B1 => n2751, B2 => n352,
                           ZN => n2407);
   U2731 : OAI22_X1 port map( A1 => n2269, A2 => n358, B1 => n2270, B2 => n361,
                           ZN => n2408);
   U2732 : OAI22_X1 port map( A1 => n2272, A2 => n367, B1 => n2273, B2 => n370,
                           ZN => n2409);
   U2733 : OAI22_X1 port map( A1 => n2785, A2 => n325, B1 => n2251, B2 => n328,
                           ZN => n2410);
   U2734 : AOI221_X1 port map( B1 => n331, B2 => n2772, C1 => n334, C2 => n2773
                           , A => n2413, ZN => n2412);
   U2735 : OAI22_X1 port map( A1 => n2771, A2 => n337, B1 => n2770, B2 => n340,
                           ZN => n2413);
   U2736 : AOI221_X1 port map( B1 => n343, B2 => n2776, C1 => n346, C2 => n2777
                           , A => n2414, ZN => n2411);
   U2737 : OAI22_X1 port map( A1 => n2775, A2 => n349, B1 => n2774, B2 => n352,
                           ZN => n2414);
   U2738 : OAI22_X1 port map( A1 => n2257, A2 => n358, B1 => n2258, B2 => n361,
                           ZN => n2415);
   U2739 : OAI22_X1 port map( A1 => n2260, A2 => n367, B1 => n2261, B2 => n370,
                           ZN => n2416);
   U2740 : OAI22_X1 port map( A1 => n2808, A2 => n325, B1 => n2239, B2 => n328,
                           ZN => n2417);
   U2741 : AOI221_X1 port map( B1 => n331, B2 => n2795, C1 => n334, C2 => n2796
                           , A => n2420, ZN => n2419);
   U2742 : OAI22_X1 port map( A1 => n2794, A2 => n337, B1 => n2793, B2 => n340,
                           ZN => n2420);
   U2743 : AOI221_X1 port map( B1 => n343, B2 => n2799, C1 => n346, C2 => n2800
                           , A => n2421, ZN => n2418);
   U2744 : OAI22_X1 port map( A1 => n2798, A2 => n349, B1 => n2797, B2 => n352,
                           ZN => n2421);
   U2745 : OAI22_X1 port map( A1 => n2245, A2 => n358, B1 => n2246, B2 => n361,
                           ZN => n2422);
   U2746 : OAI22_X1 port map( A1 => n2248, A2 => n367, B1 => n2249, B2 => n370,
                           ZN => n2423);
   U2747 : OAI22_X1 port map( A1 => n2831, A2 => n325, B1 => n2227, B2 => n328,
                           ZN => n2424);
   U2748 : AOI221_X1 port map( B1 => n331, B2 => n2818, C1 => n334, C2 => n2819
                           , A => n2427, ZN => n2426);
   U2749 : OAI22_X1 port map( A1 => n2817, A2 => n337, B1 => n2816, B2 => n340,
                           ZN => n2427);
   U2750 : AOI221_X1 port map( B1 => n343, B2 => n2822, C1 => n346, C2 => n2823
                           , A => n2428, ZN => n2425);
   U2751 : OAI22_X1 port map( A1 => n2821, A2 => n349, B1 => n2820, B2 => n352,
                           ZN => n2428);
   U2752 : OAI22_X1 port map( A1 => n2233, A2 => n358, B1 => n2234, B2 => n361,
                           ZN => n2429);
   U2753 : OAI22_X1 port map( A1 => n2236, A2 => n367, B1 => n2237, B2 => n370,
                           ZN => n2430);
   U2754 : OAI22_X1 port map( A1 => n2854, A2 => n324, B1 => n2215, B2 => n327,
                           ZN => n2431);
   U2755 : AOI221_X1 port map( B1 => n330, B2 => n2841, C1 => n333, C2 => n2842
                           , A => n2434, ZN => n2433);
   U2756 : OAI22_X1 port map( A1 => n2840, A2 => n336, B1 => n2839, B2 => n339,
                           ZN => n2434);
   U2757 : AOI221_X1 port map( B1 => n342, B2 => n2845, C1 => n345, C2 => n2846
                           , A => n2435, ZN => n2432);
   U2758 : OAI22_X1 port map( A1 => n2844, A2 => n348, B1 => n2843, B2 => n351,
                           ZN => n2435);
   U2759 : OAI22_X1 port map( A1 => n2221, A2 => n357, B1 => n2222, B2 => n360,
                           ZN => n2436);
   U2760 : OAI22_X1 port map( A1 => n2224, A2 => n366, B1 => n2225, B2 => n369,
                           ZN => n2437);
   U2761 : OAI22_X1 port map( A1 => n2877, A2 => n324, B1 => n2203, B2 => n327,
                           ZN => n2438);
   U2762 : AOI221_X1 port map( B1 => n330, B2 => n2864, C1 => n333, C2 => n2865
                           , A => n2441, ZN => n2440);
   U2763 : OAI22_X1 port map( A1 => n2863, A2 => n336, B1 => n2862, B2 => n339,
                           ZN => n2441);
   U2764 : AOI221_X1 port map( B1 => n342, B2 => n2868, C1 => n345, C2 => n2869
                           , A => n2442, ZN => n2439);
   U2765 : OAI22_X1 port map( A1 => n2867, A2 => n348, B1 => n2866, B2 => n351,
                           ZN => n2442);
   U2766 : OAI22_X1 port map( A1 => n2209, A2 => n357, B1 => n2210, B2 => n360,
                           ZN => n2443);
   U2767 : OAI22_X1 port map( A1 => n2212, A2 => n366, B1 => n2213, B2 => n369,
                           ZN => n2444);
   U2768 : OAI22_X1 port map( A1 => n2900, A2 => n324, B1 => n2191, B2 => n327,
                           ZN => n2445);
   U2769 : AOI221_X1 port map( B1 => n330, B2 => n2887, C1 => n333, C2 => n2888
                           , A => n2448, ZN => n2447);
   U2770 : OAI22_X1 port map( A1 => n2886, A2 => n336, B1 => n2885, B2 => n339,
                           ZN => n2448);
   U2771 : AOI221_X1 port map( B1 => n342, B2 => n2891, C1 => n345, C2 => n2892
                           , A => n2449, ZN => n2446);
   U2772 : OAI22_X1 port map( A1 => n2890, A2 => n348, B1 => n2889, B2 => n351,
                           ZN => n2449);
   U2773 : OAI22_X1 port map( A1 => n2197, A2 => n357, B1 => n2198, B2 => n360,
                           ZN => n2450);
   U2774 : OAI22_X1 port map( A1 => n2200, A2 => n366, B1 => n2201, B2 => n369,
                           ZN => n2451);
   U2775 : OAI22_X1 port map( A1 => n2923, A2 => n324, B1 => n2179, B2 => n327,
                           ZN => n2452);
   U2776 : AOI221_X1 port map( B1 => n330, B2 => n2910, C1 => n333, C2 => n2911
                           , A => n2455, ZN => n2454);
   U2777 : OAI22_X1 port map( A1 => n2909, A2 => n336, B1 => n2908, B2 => n339,
                           ZN => n2455);
   U2778 : AOI221_X1 port map( B1 => n342, B2 => n2914, C1 => n345, C2 => n2915
                           , A => n2456, ZN => n2453);
   U2779 : OAI22_X1 port map( A1 => n2913, A2 => n348, B1 => n2912, B2 => n351,
                           ZN => n2456);
   U2780 : OAI22_X1 port map( A1 => n2185, A2 => n357, B1 => n2186, B2 => n360,
                           ZN => n2457);
   U2781 : OAI22_X1 port map( A1 => n2188, A2 => n366, B1 => n2189, B2 => n369,
                           ZN => n2458);
   U2782 : OAI22_X1 port map( A1 => n2946, A2 => n324, B1 => n2167, B2 => n327,
                           ZN => n2459);
   U2783 : AOI221_X1 port map( B1 => n330, B2 => n2933, C1 => n333, C2 => n2934
                           , A => n2462, ZN => n2461);
   U2784 : OAI22_X1 port map( A1 => n2932, A2 => n336, B1 => n2931, B2 => n339,
                           ZN => n2462);
   U2785 : AOI221_X1 port map( B1 => n342, B2 => n2937, C1 => n345, C2 => n2938
                           , A => n2463, ZN => n2460);
   U2786 : OAI22_X1 port map( A1 => n2936, A2 => n348, B1 => n2935, B2 => n351,
                           ZN => n2463);
   U2787 : OAI22_X1 port map( A1 => n2173, A2 => n357, B1 => n2174, B2 => n360,
                           ZN => n2464);
   U2788 : OAI22_X1 port map( A1 => n2176, A2 => n366, B1 => n2177, B2 => n369,
                           ZN => n2465);
   U2789 : OAI22_X1 port map( A1 => n2969, A2 => n324, B1 => n2155, B2 => n327,
                           ZN => n2466);
   U2790 : AOI221_X1 port map( B1 => n330, B2 => n2956, C1 => n333, C2 => n2957
                           , A => n2469, ZN => n2468);
   U2791 : OAI22_X1 port map( A1 => n2955, A2 => n336, B1 => n2954, B2 => n339,
                           ZN => n2469);
   U2792 : AOI221_X1 port map( B1 => n342, B2 => n2960, C1 => n345, C2 => n2961
                           , A => n2470, ZN => n2467);
   U2793 : OAI22_X1 port map( A1 => n2959, A2 => n348, B1 => n2958, B2 => n351,
                           ZN => n2470);
   U2794 : OAI22_X1 port map( A1 => n2161, A2 => n357, B1 => n2162, B2 => n360,
                           ZN => n2471);
   U2795 : OAI22_X1 port map( A1 => n2164, A2 => n366, B1 => n2165, B2 => n369,
                           ZN => n2472);
   U2796 : OAI22_X1 port map( A1 => n3568, A2 => n324, B1 => n2143, B2 => n327,
                           ZN => n2473);
   U2797 : AOI221_X1 port map( B1 => n330, B2 => n2979, C1 => n333, C2 => n2980
                           , A => n2476, ZN => n2475);
   U2798 : OAI22_X1 port map( A1 => n2978, A2 => n336, B1 => n2977, B2 => n339,
                           ZN => n2476);
   U2799 : AOI221_X1 port map( B1 => n342, B2 => n3559, C1 => n345, C2 => n3560
                           , A => n2477, ZN => n2474);
   U2800 : OAI22_X1 port map( A1 => n2982, A2 => n348, B1 => n2981, B2 => n351,
                           ZN => n2477);
   U2801 : OAI22_X1 port map( A1 => n2149, A2 => n357, B1 => n2150, B2 => n360,
                           ZN => n2478);
   U2802 : OAI22_X1 port map( A1 => n2152, A2 => n366, B1 => n2153, B2 => n369,
                           ZN => n2479);
   U2803 : OAI22_X1 port map( A1 => n3591, A2 => n324, B1 => n2131, B2 => n327,
                           ZN => n2480);
   U2804 : AOI221_X1 port map( B1 => n330, B2 => n3578, C1 => n333, C2 => n3579
                           , A => n2483, ZN => n2482);
   U2805 : OAI22_X1 port map( A1 => n3577, A2 => n336, B1 => n3576, B2 => n339,
                           ZN => n2483);
   U2806 : AOI221_X1 port map( B1 => n342, B2 => n3582, C1 => n345, C2 => n3583
                           , A => n2484, ZN => n2481);
   U2807 : OAI22_X1 port map( A1 => n3581, A2 => n348, B1 => n3580, B2 => n351,
                           ZN => n2484);
   U2808 : OAI22_X1 port map( A1 => n2137, A2 => n357, B1 => n2138, B2 => n360,
                           ZN => n2485);
   U2809 : OAI22_X1 port map( A1 => n2140, A2 => n366, B1 => n2141, B2 => n369,
                           ZN => n2486);
   U2810 : OAI22_X1 port map( A1 => n3614, A2 => n324, B1 => n2119, B2 => n327,
                           ZN => n2487);
   U2811 : AOI221_X1 port map( B1 => n330, B2 => n3601, C1 => n333, C2 => n3602
                           , A => n2490, ZN => n2489);
   U2812 : OAI22_X1 port map( A1 => n3600, A2 => n336, B1 => n3599, B2 => n339,
                           ZN => n2490);
   U2813 : AOI221_X1 port map( B1 => n342, B2 => n3605, C1 => n345, C2 => n3606
                           , A => n2491, ZN => n2488);
   U2814 : OAI22_X1 port map( A1 => n3604, A2 => n348, B1 => n3603, B2 => n351,
                           ZN => n2491);
   U2815 : OAI22_X1 port map( A1 => n2125, A2 => n357, B1 => n2126, B2 => n360,
                           ZN => n2492);
   U2816 : OAI22_X1 port map( A1 => n2128, A2 => n366, B1 => n2129, B2 => n369,
                           ZN => n2493);
   U2817 : OAI22_X1 port map( A1 => n3637, A2 => n324, B1 => n2107, B2 => n327,
                           ZN => n2494);
   U2818 : AOI221_X1 port map( B1 => n330, B2 => n3624, C1 => n333, C2 => n3625
                           , A => n2497, ZN => n2496);
   U2819 : OAI22_X1 port map( A1 => n3623, A2 => n336, B1 => n3622, B2 => n339,
                           ZN => n2497);
   U2820 : AOI221_X1 port map( B1 => n342, B2 => n3628, C1 => n345, C2 => n3629
                           , A => n2498, ZN => n2495);
   U2821 : OAI22_X1 port map( A1 => n3627, A2 => n348, B1 => n3626, B2 => n351,
                           ZN => n2498);
   U2822 : OAI22_X1 port map( A1 => n2113, A2 => n357, B1 => n2114, B2 => n360,
                           ZN => n2499);
   U2823 : OAI22_X1 port map( A1 => n2116, A2 => n366, B1 => n2117, B2 => n369,
                           ZN => n2500);
   U2824 : OAI22_X1 port map( A1 => n3660, A2 => n324, B1 => n2095, B2 => n327,
                           ZN => n2501);
   U2825 : AOI221_X1 port map( B1 => n330, B2 => n3647, C1 => n333, C2 => n3648
                           , A => n2504, ZN => n2503);
   U2826 : OAI22_X1 port map( A1 => n3646, A2 => n336, B1 => n3645, B2 => n339,
                           ZN => n2504);
   U2827 : AOI221_X1 port map( B1 => n342, B2 => n3651, C1 => n345, C2 => n3652
                           , A => n2505, ZN => n2502);
   U2828 : OAI22_X1 port map( A1 => n3650, A2 => n348, B1 => n3649, B2 => n351,
                           ZN => n2505);
   U2829 : OAI22_X1 port map( A1 => n2101, A2 => n357, B1 => n2102, B2 => n360,
                           ZN => n2506);
   U2830 : OAI22_X1 port map( A1 => n2104, A2 => n366, B1 => n2105, B2 => n369,
                           ZN => n2507);
   U2831 : OAI22_X1 port map( A1 => n3683, A2 => n324, B1 => n2083, B2 => n327,
                           ZN => n2508);
   U2832 : AOI221_X1 port map( B1 => n330, B2 => n3670, C1 => n333, C2 => n3671
                           , A => n2511, ZN => n2510);
   U2833 : OAI22_X1 port map( A1 => n3669, A2 => n336, B1 => n3668, B2 => n339,
                           ZN => n2511);
   U2834 : AOI221_X1 port map( B1 => n342, B2 => n3674, C1 => n345, C2 => n3675
                           , A => n2512, ZN => n2509);
   U2835 : OAI22_X1 port map( A1 => n3673, A2 => n348, B1 => n3672, B2 => n351,
                           ZN => n2512);
   U2836 : OAI22_X1 port map( A1 => n2089, A2 => n357, B1 => n2090, B2 => n360,
                           ZN => n2513);
   U2837 : OAI22_X1 port map( A1 => n2092, A2 => n366, B1 => n2093, B2 => n369,
                           ZN => n2514);
   U2838 : OAI22_X1 port map( A1 => n3706, A2 => n323, B1 => n2071, B2 => n326,
                           ZN => n2515);
   U2839 : AOI221_X1 port map( B1 => n329, B2 => n3693, C1 => n332, C2 => n3694
                           , A => n2518, ZN => n2517);
   U2840 : OAI22_X1 port map( A1 => n3692, A2 => n335, B1 => n3691, B2 => n338,
                           ZN => n2518);
   U2841 : AOI221_X1 port map( B1 => n341, B2 => n3697, C1 => n344, C2 => n3698
                           , A => n2519, ZN => n2516);
   U2842 : OAI22_X1 port map( A1 => n3696, A2 => n347, B1 => n3695, B2 => n350,
                           ZN => n2519);
   U2843 : OAI22_X1 port map( A1 => n2077, A2 => n356, B1 => n2078, B2 => n359,
                           ZN => n2520);
   U2844 : OAI22_X1 port map( A1 => n2080, A2 => n365, B1 => n2081, B2 => n368,
                           ZN => n2521);
   U2845 : OAI22_X1 port map( A1 => n3729, A2 => n323, B1 => n2059, B2 => n326,
                           ZN => n2522);
   U2846 : AOI221_X1 port map( B1 => n329, B2 => n3716, C1 => n332, C2 => n3717
                           , A => n2525, ZN => n2524);
   U2847 : OAI22_X1 port map( A1 => n3715, A2 => n335, B1 => n3714, B2 => n338,
                           ZN => n2525);
   U2848 : AOI221_X1 port map( B1 => n341, B2 => n3720, C1 => n344, C2 => n3721
                           , A => n2526, ZN => n2523);
   U2849 : OAI22_X1 port map( A1 => n3719, A2 => n347, B1 => n3718, B2 => n350,
                           ZN => n2526);
   U2850 : OAI22_X1 port map( A1 => n2065, A2 => n356, B1 => n2066, B2 => n359,
                           ZN => n2527);
   U2851 : OAI22_X1 port map( A1 => n2068, A2 => n365, B1 => n2069, B2 => n368,
                           ZN => n2528);
   U2852 : OAI22_X1 port map( A1 => n3752, A2 => n323, B1 => n2047, B2 => n326,
                           ZN => n2529);
   U2853 : AOI221_X1 port map( B1 => n329, B2 => n3739, C1 => n332, C2 => n3740
                           , A => n2532, ZN => n2531);
   U2854 : OAI22_X1 port map( A1 => n3738, A2 => n335, B1 => n3737, B2 => n338,
                           ZN => n2532);
   U2855 : AOI221_X1 port map( B1 => n341, B2 => n3743, C1 => n344, C2 => n3744
                           , A => n2533, ZN => n2530);
   U2856 : OAI22_X1 port map( A1 => n3742, A2 => n347, B1 => n3741, B2 => n350,
                           ZN => n2533);
   U2857 : OAI22_X1 port map( A1 => n2053, A2 => n356, B1 => n2054, B2 => n359,
                           ZN => n2534);
   U2858 : OAI22_X1 port map( A1 => n2056, A2 => n365, B1 => n2057, B2 => n368,
                           ZN => n2535);
   U2859 : OAI22_X1 port map( A1 => n3775, A2 => n323, B1 => n2035, B2 => n326,
                           ZN => n2536);
   U2860 : AOI221_X1 port map( B1 => n329, B2 => n3762, C1 => n332, C2 => n3763
                           , A => n2539, ZN => n2538);
   U2861 : OAI22_X1 port map( A1 => n3761, A2 => n335, B1 => n3760, B2 => n338,
                           ZN => n2539);
   U2862 : AOI221_X1 port map( B1 => n341, B2 => n3766, C1 => n344, C2 => n3767
                           , A => n2540, ZN => n2537);
   U2863 : OAI22_X1 port map( A1 => n3765, A2 => n347, B1 => n3764, B2 => n350,
                           ZN => n2540);
   U2864 : OAI22_X1 port map( A1 => n2041, A2 => n356, B1 => n2042, B2 => n359,
                           ZN => n2541);
   U2865 : OAI22_X1 port map( A1 => n2044, A2 => n365, B1 => n2045, B2 => n368,
                           ZN => n2542);
   U2866 : OAI22_X1 port map( A1 => n3798, A2 => n323, B1 => n2023, B2 => n326,
                           ZN => n2543);
   U2867 : AOI221_X1 port map( B1 => n329, B2 => n3785, C1 => n332, C2 => n3786
                           , A => n2546, ZN => n2545);
   U2868 : OAI22_X1 port map( A1 => n3784, A2 => n335, B1 => n3783, B2 => n338,
                           ZN => n2546);
   U2869 : AOI221_X1 port map( B1 => n341, B2 => n3789, C1 => n344, C2 => n3790
                           , A => n2547, ZN => n2544);
   U2870 : OAI22_X1 port map( A1 => n3788, A2 => n347, B1 => n3787, B2 => n350,
                           ZN => n2547);
   U2871 : OAI22_X1 port map( A1 => n2029, A2 => n356, B1 => n2030, B2 => n359,
                           ZN => n2548);
   U2872 : OAI22_X1 port map( A1 => n2032, A2 => n365, B1 => n2033, B2 => n368,
                           ZN => n2549);
   U2873 : OAI22_X1 port map( A1 => n3821, A2 => n323, B1 => n2011, B2 => n326,
                           ZN => n2550);
   U2874 : AOI221_X1 port map( B1 => n329, B2 => n3808, C1 => n332, C2 => n3809
                           , A => n2553, ZN => n2552);
   U2875 : OAI22_X1 port map( A1 => n3807, A2 => n335, B1 => n3806, B2 => n338,
                           ZN => n2553);
   U2876 : AOI221_X1 port map( B1 => n341, B2 => n3812, C1 => n344, C2 => n3813
                           , A => n2554, ZN => n2551);
   U2877 : OAI22_X1 port map( A1 => n3811, A2 => n347, B1 => n3810, B2 => n350,
                           ZN => n2554);
   U2878 : OAI22_X1 port map( A1 => n2017, A2 => n356, B1 => n2018, B2 => n359,
                           ZN => n2555);
   U2879 : OAI22_X1 port map( A1 => n2020, A2 => n365, B1 => n2021, B2 => n368,
                           ZN => n2556);
   U2880 : OAI22_X1 port map( A1 => n3844, A2 => n323, B1 => n1999, B2 => n326,
                           ZN => n2557);
   U2881 : AOI221_X1 port map( B1 => n329, B2 => n3831, C1 => n332, C2 => n3832
                           , A => n2560, ZN => n2559);
   U2882 : OAI22_X1 port map( A1 => n3830, A2 => n335, B1 => n3829, B2 => n338,
                           ZN => n2560);
   U2883 : AOI221_X1 port map( B1 => n341, B2 => n3835, C1 => n344, C2 => n3836
                           , A => n2561, ZN => n2558);
   U2884 : OAI22_X1 port map( A1 => n3834, A2 => n347, B1 => n3833, B2 => n350,
                           ZN => n2561);
   U2885 : OAI22_X1 port map( A1 => n2005, A2 => n356, B1 => n2006, B2 => n359,
                           ZN => n2562);
   U2886 : OAI22_X1 port map( A1 => n2008, A2 => n365, B1 => n2009, B2 => n368,
                           ZN => n2563);
   U2887 : OAI22_X1 port map( A1 => n3867, A2 => n323, B1 => n1987, B2 => n326,
                           ZN => n2564);
   U2888 : AOI221_X1 port map( B1 => n329, B2 => n3854, C1 => n332, C2 => n3855
                           , A => n2567, ZN => n2566);
   U2889 : OAI22_X1 port map( A1 => n3853, A2 => n335, B1 => n3852, B2 => n338,
                           ZN => n2567);
   U2890 : AOI221_X1 port map( B1 => n341, B2 => n3858, C1 => n344, C2 => n3859
                           , A => n2568, ZN => n2565);
   U2891 : OAI22_X1 port map( A1 => n3857, A2 => n347, B1 => n3856, B2 => n350,
                           ZN => n2568);
   U2892 : OAI22_X1 port map( A1 => n1993, A2 => n356, B1 => n1994, B2 => n359,
                           ZN => n2569);
   U2893 : OAI22_X1 port map( A1 => n1996, A2 => n365, B1 => n1997, B2 => n368,
                           ZN => n2570);
   U2894 : OAI22_X1 port map( A1 => n3890, A2 => n323, B1 => n1975, B2 => n326,
                           ZN => n2571);
   U2895 : AOI221_X1 port map( B1 => n329, B2 => n3877, C1 => n332, C2 => n3878
                           , A => n2574, ZN => n2573);
   U2896 : OAI22_X1 port map( A1 => n3876, A2 => n335, B1 => n3875, B2 => n338,
                           ZN => n2574);
   U2897 : AOI221_X1 port map( B1 => n341, B2 => n3881, C1 => n344, C2 => n3882
                           , A => n2575, ZN => n2572);
   U2898 : OAI22_X1 port map( A1 => n3880, A2 => n347, B1 => n3879, B2 => n350,
                           ZN => n2575);
   U2899 : OAI22_X1 port map( A1 => n1981, A2 => n356, B1 => n1982, B2 => n359,
                           ZN => n2576);
   U2900 : OAI22_X1 port map( A1 => n1984, A2 => n365, B1 => n1985, B2 => n368,
                           ZN => n2577);
   U2901 : OAI22_X1 port map( A1 => n3913, A2 => n323, B1 => n1963, B2 => n326,
                           ZN => n2578);
   U2902 : AOI221_X1 port map( B1 => n329, B2 => n3900, C1 => n332, C2 => n3901
                           , A => n2581, ZN => n2580);
   U2903 : OAI22_X1 port map( A1 => n3899, A2 => n335, B1 => n3898, B2 => n338,
                           ZN => n2581);
   U2904 : AOI221_X1 port map( B1 => n341, B2 => n3904, C1 => n344, C2 => n3905
                           , A => n2582, ZN => n2579);
   U2905 : OAI22_X1 port map( A1 => n3903, A2 => n347, B1 => n3902, B2 => n350,
                           ZN => n2582);
   U2906 : OAI22_X1 port map( A1 => n1969, A2 => n356, B1 => n1970, B2 => n359,
                           ZN => n2583);
   U2907 : OAI22_X1 port map( A1 => n1972, A2 => n365, B1 => n1973, B2 => n368,
                           ZN => n2584);
   U2908 : OAI22_X1 port map( A1 => n3936, A2 => n323, B1 => n1951, B2 => n326,
                           ZN => n2585);
   U2909 : AOI221_X1 port map( B1 => n329, B2 => n3923, C1 => n332, C2 => n3924
                           , A => n2588, ZN => n2587);
   U2910 : OAI22_X1 port map( A1 => n3922, A2 => n335, B1 => n3921, B2 => n338,
                           ZN => n2588);
   U2911 : AOI221_X1 port map( B1 => n341, B2 => n3927, C1 => n344, C2 => n3928
                           , A => n2589, ZN => n2586);
   U2912 : OAI22_X1 port map( A1 => n3926, A2 => n347, B1 => n3925, B2 => n350,
                           ZN => n2589);
   U2913 : OAI22_X1 port map( A1 => n1957, A2 => n356, B1 => n1958, B2 => n359,
                           ZN => n2590);
   U2914 : OAI22_X1 port map( A1 => n1960, A2 => n365, B1 => n1961, B2 => n368,
                           ZN => n2591);
   U2915 : AND2_X1 port map( A1 => n2592, A2 => n2593, ZN => n2349);
   U2916 : AND2_X1 port map( A1 => n2592, A2 => n2594, ZN => n2348);
   U2917 : NAND2_X1 port map( A1 => n2595, A2 => n2596, ZN => n2347);
   U2918 : NAND2_X1 port map( A1 => n2597, A2 => n2593, ZN => n2346);
   U2919 : AND2_X1 port map( A1 => n2597, A2 => n2594, ZN => n2353);
   U2920 : AND2_X1 port map( A1 => n2597, A2 => n2596, ZN => n2352);
   U2921 : NAND2_X1 port map( A1 => n2592, A2 => n2596, ZN => n2351);
   U2922 : NAND2_X1 port map( A1 => n2592, A2 => n2598, ZN => n2350);
   U2923 : NOR3_X1 port map( A1 => n2599, A2 => ADD_RS1(0), A3 => n2600, ZN => 
                           n2592);
   U2924 : OAI22_X1 port map( A1 => n3959, A2 => n323, B1 => n1922, B2 => n326,
                           ZN => n2601);
   U2925 : NAND2_X1 port map( A1 => n2602, A2 => n2596, ZN => n2359);
   U2926 : NAND2_X1 port map( A1 => n2602, A2 => n2598, ZN => n2358);
   U2927 : AND2_X1 port map( A1 => n2595, A2 => n2593, ZN => n2356);
   U2928 : AND2_X1 port map( A1 => n2595, A2 => n2598, ZN => n2355);
   U2929 : AND2_X1 port map( A1 => n2602, A2 => n2594, ZN => n2361);
   U2930 : AND2_X1 port map( A1 => n2602, A2 => n2593, ZN => n2360);
   U2931 : NOR3_X1 port map( A1 => ADD_RS1(0), A2 => ADD_RS1(3), A3 => n2599, 
                           ZN => n2602);
   U2932 : NAND2_X1 port map( A1 => n2595, A2 => n2594, ZN => n2354);
   U2933 : NOR3_X1 port map( A1 => n2603, A2 => ADD_RS1(3), A3 => n2599, ZN => 
                           n2595);
   U2934 : AOI221_X1 port map( B1 => n329, B2 => n3946, C1 => n332, C2 => n3947
                           , A => n2606, ZN => n2605);
   U2935 : OAI22_X1 port map( A1 => n3945, A2 => n335, B1 => n3944, B2 => n338,
                           ZN => n2606);
   U2936 : NAND2_X1 port map( A1 => n2598, A2 => n2607, ZN => n2368);
   U2937 : NAND2_X1 port map( A1 => n2598, A2 => n2608, ZN => n2367);
   U2938 : AND2_X1 port map( A1 => n2607, A2 => n2596, ZN => n2365);
   U2939 : AND2_X1 port map( A1 => n2596, A2 => n2608, ZN => n2364);
   U2940 : AOI221_X1 port map( B1 => n341, B2 => n3950, C1 => n344, C2 => n3951
                           , A => n2609, ZN => n2604);
   U2941 : OAI22_X1 port map( A1 => n3949, A2 => n347, B1 => n3948, B2 => n350,
                           ZN => n2609);
   U2942 : NAND2_X1 port map( A1 => n2594, A2 => n2607, ZN => n2373);
   U2943 : NAND2_X1 port map( A1 => n2594, A2 => n2608, ZN => n2372);
   U2944 : AND2_X1 port map( A1 => n2593, A2 => n2607, ZN => n2370);
   U2945 : NOR3_X1 port map( A1 => ADD_RS1(0), A2 => ADD_RS1(4), A3 => n2600, 
                           ZN => n2607);
   U2946 : AND2_X1 port map( A1 => n2593, A2 => n2608, ZN => n2369);
   U2947 : NOR3_X1 port map( A1 => n2603, A2 => ADD_RS1(4), A3 => n2600, ZN => 
                           n2608);
   U2948 : OAI22_X1 port map( A1 => n1940, A2 => n356, B1 => n1942, B2 => n359,
                           ZN => n2610);
   U2949 : NAND2_X1 port map( A1 => n2611, A2 => n2596, ZN => n2377);
   U2950 : NAND2_X1 port map( A1 => n2612, A2 => n2596, ZN => n2376);
   U2951 : NOR2_X1 port map( A1 => n2613, A2 => n2614, ZN => n2596);
   U2952 : AND2_X1 port map( A1 => n2612, A2 => n2598, ZN => n2374);
   U2953 : OAI22_X1 port map( A1 => n1946, A2 => n365, B1 => n1948, B2 => n368,
                           ZN => n2615);
   U2954 : NAND2_X1 port map( A1 => n2611, A2 => n2593, ZN => n2381);
   U2955 : NAND2_X1 port map( A1 => n2612, A2 => n2593, ZN => n2380);
   U2956 : NOR2_X1 port map( A1 => n2614, A2 => ADD_RS1(2), ZN => n2593);
   U2957 : NOR3_X1 port map( A1 => ADD_RS1(3), A2 => ADD_RS1(4), A3 => 
                           ADD_RS1(0), ZN => n2612);
   U2958 : AND2_X1 port map( A1 => n2597, A2 => n2598, ZN => n2378);
   U2959 : NOR2_X1 port map( A1 => n2613, A2 => ADD_RS1(1), ZN => n2598);
   U2960 : INV_X1 port map( A => ADD_RS1(2), ZN => n2613);
   U2961 : NOR3_X1 port map( A1 => n2599, A2 => n2603, A3 => n2600, ZN => n2597
                           );
   U2962 : INV_X1 port map( A => ADD_RS1(3), ZN => n2600);
   U2963 : INV_X1 port map( A => ADD_RS1(4), ZN => n2599);
   U2964 : NOR2_X1 port map( A1 => ADD_RS1(1), A2 => ADD_RS1(2), ZN => n2594);
   U2965 : NOR3_X1 port map( A1 => ADD_RS1(3), A2 => ADD_RS1(4), A3 => n2603, 
                           ZN => n2611);
   U2966 : INV_X1 port map( A => ADD_RS1(0), ZN => n2603);
   U2967 : NOR3_X1 port map( A1 => n2620, A2 => n2344, A3 => n2621, ZN => n2619
                           );
   U2968 : XNOR2_X1 port map( A => ADD_WR(1), B => n2614, ZN => n2621);
   U2969 : INV_X1 port map( A => ADD_RS1(1), ZN => n2614);
   U2970 : INV_X1 port map( A => WR, ZN => n2344);
   U2971 : XNOR2_X1 port map( A => n1907, B => ADD_RS1(0), ZN => n2620);
   U2972 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS1(3), ZN => n2618);
   U2973 : XNOR2_X1 port map( A => ADD_WR(4), B => ADD_RS1(4), ZN => n2617);
   U2974 : XNOR2_X1 port map( A => ADD_RS1(2), B => ADD_WR(2), ZN => n2616);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_0 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_0;

architecture SYN_bhv of regn_N5_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n11, n12, n13, n14, n15, DOUT_0_port, DOUT_1_port, DOUT_2_port, 
      DOUT_3_port, DOUT_4_port, n_1819, n_1820, n_1821, n_1822, n_1823 : 
      std_logic;

begin
   DOUT <= ( DOUT_4_port, DOUT_3_port, DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n15, CK => CLK, RN => RST, Q => 
                           DOUT_4_port, QN => n_1819);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n14, CK => CLK, RN => RST, Q => 
                           DOUT_3_port, QN => n_1820);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n13, CK => CLK, RN => RST, Q => 
                           DOUT_2_port, QN => n_1821);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n12, CK => CLK, RN => RST, Q => 
                           DOUT_1_port, QN => n_1822);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n11, CK => CLK, RN => RST, Q => 
                           DOUT_0_port, QN => n_1823);
   U2 : MUX2_X1 port map( A => DOUT_0_port, B => DIN(0), S => EN, Z => n11);
   U3 : MUX2_X1 port map( A => DOUT_1_port, B => DIN(1), S => EN, Z => n12);
   U4 : MUX2_X1 port map( A => DOUT_2_port, B => DIN(2), S => EN, Z => n13);
   U5 : MUX2_X1 port map( A => DOUT_3_port, B => DIN(3), S => EN, Z => n14);
   U6 : MUX2_X1 port map( A => DOUT_4_port, B => DIN(4), S => EN, Z => n15);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity instruction_decomposition is

   port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype : in
         std_logic;  ADD_RS1, ADD_RS2, ADD_WR : out std_logic_vector (4 downto 
         0);  IMM : out std_logic_vector (31 downto 0));

end instruction_decomposition;

architecture SYN_bhv of instruction_decomposition is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal IMM_24_port, IMM_23_port, IMM_22_port, IMM_21_port, IMM_20_port, 
      IMM_19_port, IMM_18_port, IMM_17_port, IMM_16_port, IMM_15_port, 
      IMM_14_port, IMM_13_port, IMM_12_port, IMM_11_port, IMM_10_port, 
      IMM_9_port, IMM_8_port, IMM_7_port, IMM_6_port, IMM_5_port, IMM_4_port, 
      IMM_3_port, IMM_2_port, IMM_1_port, IMM_0_port, n21, n22, n23, n24, n25, 
      n26, n27, n28, n29, n30, n31, n32, n1, n2, IMM_31_port, n4, n5, n6, n7, 
      n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20 : std_logic
      ;

begin
   IMM <= ( IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, 
      IMM_31_port, IMM_31_port, IMM_24_port, IMM_23_port, IMM_22_port, 
      IMM_21_port, IMM_20_port, IMM_19_port, IMM_18_port, IMM_17_port, 
      IMM_16_port, IMM_15_port, IMM_14_port, IMM_13_port, IMM_12_port, 
      IMM_11_port, IMM_10_port, IMM_9_port, IMM_8_port, IMM_7_port, IMM_6_port,
      IMM_5_port, IMM_4_port, IMM_3_port, IMM_2_port, IMM_1_port, IMM_0_port );
   
   U72 : NAND3_X1 port map( A1 => INST_IN(29), A2 => INST_IN(27), A3 => 
                           INST_IN(31), ZN => n31);
   U73 : NAND3_X1 port map( A1 => INST_IN(26), A2 => Itype, A3 => n32, ZN => 
                           n30);
   U2 : INV_X1 port map( A => Rtype, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n28, A2 => Jtype, ZN => n24);
   U4 : INV_X1 port map( A => n27, ZN => n2);
   U5 : OAI21_X1 port map( B1 => Itype, B2 => Jtype, A => n4, ZN => n27);
   U6 : NOR2_X1 port map( A1 => Rtype, A2 => Itype, ZN => n28);
   U7 : NOR2_X1 port map( A1 => n28, A2 => n7, ZN => ADD_RS1(3));
   U8 : NOR2_X1 port map( A1 => n1, A2 => n12, ZN => ADD_RS2(3));
   U9 : NOR2_X1 port map( A1 => n28, A2 => n10, ZN => ADD_RS1(0));
   U10 : NOR2_X1 port map( A1 => n1, A2 => n15, ZN => ADD_RS2(0));
   U11 : NOR2_X1 port map( A1 => n1, A2 => n11, ZN => ADD_RS2(4));
   U12 : OR2_X1 port map( A1 => n26, A2 => n16, ZN => n25);
   U13 : NOR2_X1 port map( A1 => n28, A2 => n8, ZN => ADD_RS1(2));
   U14 : NOR2_X1 port map( A1 => n1, A2 => n13, ZN => ADD_RS2(2));
   U15 : NOR2_X1 port map( A1 => n28, A2 => n9, ZN => ADD_RS1(1));
   U16 : NOR2_X1 port map( A1 => n1, A2 => n14, ZN => ADD_RS2(1));
   U17 : NAND2_X1 port map( A1 => Itype, A2 => n4, ZN => n26);
   U18 : INV_X1 port map( A => Itype, ZN => n5);
   U19 : AND2_X1 port map( A1 => INST_IN(0), A2 => n2, ZN => IMM_0_port);
   U20 : AND2_X1 port map( A1 => INST_IN(1), A2 => n2, ZN => IMM_1_port);
   U21 : AND2_X1 port map( A1 => INST_IN(2), A2 => n2, ZN => IMM_2_port);
   U22 : AND2_X1 port map( A1 => INST_IN(3), A2 => n2, ZN => IMM_3_port);
   U23 : AND2_X1 port map( A1 => INST_IN(4), A2 => n2, ZN => IMM_4_port);
   U24 : AND2_X1 port map( A1 => INST_IN(5), A2 => n2, ZN => IMM_5_port);
   U25 : AND2_X1 port map( A1 => INST_IN(6), A2 => n2, ZN => IMM_6_port);
   U26 : AND2_X1 port map( A1 => INST_IN(7), A2 => n2, ZN => IMM_7_port);
   U27 : AND2_X1 port map( A1 => INST_IN(8), A2 => n2, ZN => IMM_8_port);
   U28 : AND2_X1 port map( A1 => INST_IN(9), A2 => n2, ZN => IMM_9_port);
   U29 : AND2_X1 port map( A1 => INST_IN(10), A2 => n2, ZN => IMM_10_port);
   U30 : NOR2_X1 port map( A1 => n27, A2 => n20, ZN => IMM_11_port);
   U31 : NOR2_X1 port map( A1 => n27, A2 => n19, ZN => IMM_12_port);
   U32 : NOR2_X1 port map( A1 => n27, A2 => n18, ZN => IMM_13_port);
   U33 : NOR2_X1 port map( A1 => n27, A2 => n17, ZN => IMM_14_port);
   U34 : NOR2_X1 port map( A1 => n27, A2 => n16, ZN => IMM_15_port);
   U35 : OAI21_X1 port map( B1 => n24, B2 => n15, A => n25, ZN => IMM_16_port);
   U36 : OAI21_X1 port map( B1 => n24, B2 => n14, A => n25, ZN => IMM_17_port);
   U37 : OAI21_X1 port map( B1 => n24, B2 => n13, A => n25, ZN => IMM_18_port);
   U38 : OAI21_X1 port map( B1 => n24, B2 => n12, A => n25, ZN => IMM_19_port);
   U39 : OAI21_X1 port map( B1 => n24, B2 => n11, A => n25, ZN => IMM_20_port);
   U40 : OAI21_X1 port map( B1 => n24, B2 => n10, A => n25, ZN => IMM_21_port);
   U41 : OAI21_X1 port map( B1 => n24, B2 => n9, A => n25, ZN => IMM_22_port);
   U42 : OAI21_X1 port map( B1 => n24, B2 => n8, A => n25, ZN => IMM_23_port);
   U43 : OAI21_X1 port map( B1 => n24, B2 => n7, A => n25, ZN => IMM_24_port);
   U44 : OAI221_X1 port map( B1 => n26, B2 => n15, C1 => n20, C2 => n4, A => 
                           n24, ZN => ADD_WR(0));
   U45 : OAI221_X1 port map( B1 => n26, B2 => n14, C1 => n19, C2 => n4, A => 
                           n24, ZN => ADD_WR(1));
   U46 : OAI221_X1 port map( B1 => n26, B2 => n13, C1 => n18, C2 => n4, A => 
                           n24, ZN => ADD_WR(2));
   U47 : OAI221_X1 port map( B1 => n26, B2 => n12, C1 => n17, C2 => n4, A => 
                           n24, ZN => ADD_WR(3));
   U48 : OAI221_X1 port map( B1 => n26, B2 => n11, C1 => n16, C2 => n4, A => 
                           n24, ZN => ADD_WR(4));
   U49 : NOR2_X1 port map( A1 => n28, A2 => n6, ZN => ADD_RS1(4));
   U50 : INV_X1 port map( A => INST_IN(25), ZN => n6);
   U51 : INV_X1 port map( A => n29, ZN => n1);
   U52 : OAI21_X1 port map( B1 => n30, B2 => n31, A => n4, ZN => n29);
   U53 : INV_X1 port map( A => INST_IN(15), ZN => n16);
   U54 : INV_X1 port map( A => INST_IN(16), ZN => n15);
   U55 : INV_X1 port map( A => INST_IN(17), ZN => n14);
   U56 : INV_X1 port map( A => INST_IN(19), ZN => n12);
   U57 : INV_X1 port map( A => INST_IN(18), ZN => n13);
   U58 : INV_X1 port map( A => INST_IN(20), ZN => n11);
   U59 : NOR2_X1 port map( A1 => INST_IN(30), A2 => INST_IN(28), ZN => n32);
   U60 : INV_X1 port map( A => n21, ZN => IMM_31_port);
   U61 : OAI21_X1 port map( B1 => n22, B2 => n23, A => n4, ZN => n21);
   U62 : AND3_X1 port map( A1 => Jtype, A2 => n5, A3 => INST_IN(25), ZN => n22)
                           ;
   U63 : NOR2_X1 port map( A1 => n16, A2 => n5, ZN => n23);
   U64 : INV_X1 port map( A => INST_IN(21), ZN => n10);
   U65 : INV_X1 port map( A => INST_IN(24), ZN => n7);
   U66 : INV_X1 port map( A => INST_IN(22), ZN => n9);
   U67 : INV_X1 port map( A => INST_IN(23), ZN => n8);
   U68 : INV_X1 port map( A => INST_IN(11), ZN => n20);
   U69 : INV_X1 port map( A => INST_IN(12), ZN => n19);
   U70 : INV_X1 port map( A => INST_IN(13), ZN => n18);
   U71 : INV_X1 port map( A => INST_IN(14), ZN => n17);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity instruction_type is

   port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype : 
         out std_logic);

end instruction_type;

architecture SYN_bhv of instruction_type is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n1, n2, n3, n4, n5, 
      n6, n7, n8 : std_logic;

begin
   
   U21 : OAI33_X1 port map( A1 => n5, A2 => INST_IN(29), A3 => n2, B1 => n4, B2
                           => INST_IN(30), B3 => INST_IN(26), ZN => n17);
   U1 : NOR2_X1 port map( A1 => n9, A2 => n10, ZN => Rtype);
   U2 : OAI22_X1 port map( A1 => n10, A2 => n5, B1 => n7, B2 => n4, ZN => n16);
   U3 : NOR2_X1 port map( A1 => n9, A2 => n6, ZN => Jtype);
   U4 : NAND4_X1 port map( A1 => n5, A2 => n4, A3 => n3, A4 => n1, ZN => n9);
   U5 : NAND2_X1 port map( A1 => n6, A2 => n8, ZN => n10);
   U6 : INV_X1 port map( A => n14, ZN => n7);
   U7 : INV_X1 port map( A => n18, ZN => n2);
   U8 : OAI221_X1 port map( B1 => n7, B2 => INST_IN(30), C1 => n3, C2 => 
                           INST_IN(26), A => n10, ZN => n18);
   U9 : OAI211_X1 port map( C1 => INST_IN(31), C2 => n11, A => n12, B => n13, 
                           ZN => Itype);
   U10 : NAND4_X1 port map( A1 => INST_IN(29), A2 => INST_IN(28), A3 => n14, A4
                           => n1, ZN => n13);
   U11 : NAND4_X1 port map( A1 => INST_IN(31), A2 => INST_IN(27), A3 => n15, A4
                           => INST_IN(26), ZN => n12);
   U12 : AOI21_X1 port map( B1 => INST_IN(30), B2 => n16, A => n17, ZN => n11);
   U13 : NOR2_X1 port map( A1 => n8, A2 => INST_IN(27), ZN => n14);
   U14 : NOR2_X1 port map( A1 => INST_IN(30), A2 => INST_IN(28), ZN => n15);
   U15 : INV_X1 port map( A => INST_IN(30), ZN => n3);
   U16 : INV_X1 port map( A => INST_IN(28), ZN => n5);
   U17 : INV_X1 port map( A => INST_IN(29), ZN => n4);
   U18 : INV_X1 port map( A => INST_IN(26), ZN => n8);
   U19 : INV_X1 port map( A => INST_IN(31), ZN => n1);
   U20 : INV_X1 port map( A => INST_IN(27), ZN => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_0 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_0;

architecture SYN_bhv of regn_N32_0 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, DOUT_27_port,
      DOUT_26_port, DOUT_25_port, n117, DOUT_23_port, DOUT_22_port, 
      DOUT_21_port, DOUT_20_port, DOUT_19_port, DOUT_18_port, DOUT_17_port, 
      n118, DOUT_15_port, n119, n120, DOUT_11_port, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, DOUT_1_port, DOUT_0_port, n33, n34, n35, 
      n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50
      , n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, 
      n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79
      , n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, 
      n94, n95, n96, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, DOUT_2_port, DOUT_3_port, 
      DOUT_4_port, DOUT_5_port, DOUT_6_port, DOUT_7_port, DOUT_8_port, 
      DOUT_9_port, DOUT_10_port, n31, DOUT_12_port, DOUT_13_port, DOUT_14_port,
      n99, DOUT_16_port, n101, n102, n103, n104, n105, n106, n107, n108, 
      DOUT_24_port, n110, n111, n112, n113, n114, n115, n116, n_1824 : 
      std_logic;

begin
   DOUT <= ( DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, 
      DOUT_27_port, DOUT_26_port, DOUT_25_port, DOUT_24_port, DOUT_23_port, 
      DOUT_22_port, DOUT_21_port, DOUT_20_port, DOUT_19_port, DOUT_18_port, 
      DOUT_17_port, DOUT_16_port, DOUT_15_port, DOUT_14_port, DOUT_13_port, 
      DOUT_12_port, DOUT_11_port, DOUT_10_port, DOUT_9_port, DOUT_8_port, 
      DOUT_7_port, DOUT_6_port, DOUT_5_port, DOUT_4_port, DOUT_3_port, 
      DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n96, CK => CLK, RN => n19, Q => 
                           DOUT_31_port, QN => n64);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n95, CK => CLK, RN => n19, Q => 
                           DOUT_30_port, QN => n63);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n93, CK => CLK, RN => n19, Q => 
                           DOUT_28_port, QN => n61);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n91, CK => CLK, RN => n19, Q => 
                           DOUT_26_port, QN => n59);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n90, CK => CLK, RN => n19, Q => 
                           DOUT_25_port, QN => n58);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n89, CK => CLK, RN => n19, Q => 
                           n117, QN => n57);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n88, CK => CLK, RN => n18, Q => 
                           DOUT_23_port, QN => n56);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n87, CK => CLK, RN => n18, Q => 
                           DOUT_22_port, QN => n55);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n86, CK => CLK, RN => n18, Q => 
                           DOUT_21_port, QN => n54);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n85, CK => CLK, RN => n18, Q => 
                           DOUT_20_port, QN => n53);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n84, CK => CLK, RN => n18, Q => 
                           DOUT_19_port, QN => n52);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n83, CK => CLK, RN => n18, Q => 
                           DOUT_18_port, QN => n51);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n82, CK => CLK, RN => n18, Q => 
                           DOUT_17_port, QN => n50);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n81, CK => CLK, RN => n18, Q => 
                           n118, QN => n49);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n80, CK => CLK, RN => n18, Q => 
                           DOUT_15_port, QN => n48);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n79, CK => CLK, RN => n18, Q => 
                           n_1824, QN => n47);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n78, CK => CLK, RN => n18, Q => 
                           n119, QN => n46);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n77, CK => CLK, RN => n18, Q => 
                           n120, QN => n45);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n76, CK => CLK, RN => n17, Q => 
                           DOUT_11_port, QN => n44);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n75, CK => CLK, RN => n17, Q => 
                           n121, QN => n43);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n74, CK => CLK, RN => n17, Q => 
                           n122, QN => n42);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n73, CK => CLK, RN => n17, Q => 
                           n123, QN => n41);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n72, CK => CLK, RN => n17, Q => 
                           n124, QN => n40);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n71, CK => CLK, RN => n17, Q => 
                           n125, QN => n39);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n70, CK => CLK, RN => n17, Q => 
                           n126, QN => n38);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n69, CK => CLK, RN => n17, Q => 
                           n127, QN => n37);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n68, CK => CLK, RN => n17, Q => 
                           n128, QN => n36);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n67, CK => CLK, RN => n17, Q => 
                           n129, QN => n35);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n66, CK => CLK, RN => n17, Q => 
                           DOUT_1_port, QN => n34);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n65, CK => CLK, RN => n17, Q => 
                           DOUT_0_port, QN => n33);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n92, CK => CLK, RN => n19, Q => 
                           DOUT_27_port, QN => n60);
   DOUT_reg_29_inst : DFFR_X2 port map( D => n94, CK => CLK, RN => n19, Q => 
                           DOUT_29_port, QN => n62);
   U2 : INV_X1 port map( A => EN, ZN => n5);
   U3 : INV_X1 port map( A => EN, ZN => n4);
   U4 : INV_X1 port map( A => EN, ZN => n6);
   U5 : INV_X1 port map( A => EN, ZN => n7);
   U6 : INV_X1 port map( A => EN, ZN => n3);
   U7 : INV_X1 port map( A => EN, ZN => n2);
   U8 : INV_X1 port map( A => EN, ZN => n1);
   U9 : MUX2_X1 port map( A => DIN(0), B => n20, S => n1, Z => n65);
   U10 : MUX2_X1 port map( A => DIN(4), B => n127, S => n2, Z => n69);
   U11 : MUX2_X1 port map( A => DIN(3), B => n128, S => n3, Z => n68);
   U12 : MUX2_X1 port map( A => DIN(5), B => n126, S => n4, Z => n70);
   U13 : MUX2_X1 port map( A => DIN(1), B => n21, S => n5, Z => n66);
   U14 : MUX2_X1 port map( A => DIN(6), B => n125, S => n5, Z => n71);
   U15 : MUX2_X1 port map( A => DIN(10), B => n121, S => n6, Z => n75);
   U16 : MUX2_X1 port map( A => DIN(16), B => n118, S => n7, Z => n81);
   U17 : INV_X1 port map( A => n49, ZN => DOUT_16_port);
   U18 : MUX2_X1 port map( A => DIN(24), B => n117, S => n3, Z => n89);
   U19 : MUX2_X1 port map( A => DIN(8), B => n123, S => n2, Z => n73);
   U20 : MUX2_X1 port map( A => DIN(12), B => n120, S => n1, Z => n77);
   U21 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n8);
   U22 : NAND2_X1 port map( A1 => n124, A2 => n108, ZN => n9);
   U23 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => n72);
   U24 : OR2_X1 port map( A1 => n58, A2 => EN, ZN => n10);
   U25 : NAND2_X1 port map( A1 => n110, A2 => n10, ZN => n90);
   U26 : OR2_X2 port map( A1 => n62, A2 => EN, ZN => n11);
   U27 : NAND2_X1 port map( A1 => n114, A2 => n11, ZN => n94);
   U28 : OR2_X1 port map( A1 => n61, A2 => EN, ZN => n12);
   U29 : NAND2_X1 port map( A1 => n113, A2 => n12, ZN => n93);
   U30 : OR2_X1 port map( A1 => n63, A2 => EN, ZN => n13);
   U31 : NAND2_X1 port map( A1 => n115, A2 => n13, ZN => n95);
   U32 : OR2_X2 port map( A1 => n50, A2 => EN, ZN => n14);
   U33 : NAND2_X1 port map( A1 => n101, A2 => n14, ZN => n82);
   U34 : OR2_X2 port map( A1 => n44, A2 => EN, ZN => n15);
   U35 : NAND2_X1 port map( A1 => n31, A2 => n15, ZN => n76);
   U36 : OR2_X2 port map( A1 => n59, A2 => EN, ZN => n16);
   U37 : NAND2_X1 port map( A1 => n111, A2 => n16, ZN => n91);
   U38 : BUF_X1 port map( A => RST, Z => n17);
   U39 : BUF_X1 port map( A => RST, Z => n18);
   U40 : BUF_X1 port map( A => RST, Z => n19);
   U41 : INV_X1 port map( A => EN, ZN => n108);
   U42 : OAI22_X1 port map( A1 => n107, A2 => n108, B1 => n56, B2 => EN, ZN => 
                           n88);
   U43 : INV_X1 port map( A => DIN(23), ZN => n107);
   U44 : INV_X1 port map( A => n33, ZN => n20);
   U45 : INV_X1 port map( A => n34, ZN => n21);
   U46 : INV_X1 port map( A => n35, ZN => DOUT_2_port);
   U47 : MUX2_X1 port map( A => n129, B => DIN(2), S => EN, Z => n67);
   U48 : INV_X1 port map( A => n36, ZN => DOUT_3_port);
   U49 : INV_X1 port map( A => n37, ZN => DOUT_4_port);
   U50 : INV_X1 port map( A => n38, ZN => DOUT_5_port);
   U51 : INV_X1 port map( A => n39, ZN => DOUT_6_port);
   U52 : INV_X1 port map( A => n40, ZN => DOUT_7_port);
   U53 : INV_X1 port map( A => n41, ZN => DOUT_8_port);
   U54 : INV_X1 port map( A => n42, ZN => DOUT_9_port);
   U55 : MUX2_X1 port map( A => n122, B => DIN(9), S => EN, Z => n74);
   U56 : INV_X1 port map( A => n43, ZN => DOUT_10_port);
   U57 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n31);
   U58 : INV_X1 port map( A => n45, ZN => DOUT_12_port);
   U59 : INV_X1 port map( A => n46, ZN => DOUT_13_port);
   U60 : MUX2_X1 port map( A => n119, B => DIN(13), S => EN, Z => n78);
   U61 : INV_X1 port map( A => n47, ZN => DOUT_14_port);
   U62 : MUX2_X1 port map( A => DOUT_14_port, B => DIN(14), S => EN, Z => n79);
   U63 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n99);
   U64 : OAI21_X1 port map( B1 => n48, B2 => EN, A => n99, ZN => n80);
   U65 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n102);
   U67 : OAI21_X1 port map( B1 => n51, B2 => EN, A => n102, ZN => n83);
   U68 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n103);
   U69 : OAI21_X1 port map( B1 => n52, B2 => EN, A => n103, ZN => n84);
   U70 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n104);
   U71 : OAI21_X1 port map( B1 => n53, B2 => EN, A => n104, ZN => n85);
   U72 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n105);
   U73 : OAI21_X1 port map( B1 => n54, B2 => EN, A => n105, ZN => n86);
   U74 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n106);
   U75 : OAI21_X1 port map( B1 => n55, B2 => EN, A => n106, ZN => n87);
   U76 : INV_X1 port map( A => n57, ZN => DOUT_24_port);
   U77 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n110);
   U78 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n111);
   U79 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n112);
   U80 : OAI21_X1 port map( B1 => n60, B2 => EN, A => n112, ZN => n92);
   U81 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n113);
   U82 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n114);
   U83 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n115);
   U84 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n116);
   U85 : OAI21_X1 port map( B1 => n64, B2 => EN, A => n116, ZN => n96);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_0;

architecture SYN_bhv of mux21_NBIT32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => B(29), B => A(29), S => n1, Z => Z(29));
   U2 : INV_X32 port map( A => n12, ZN => n1);
   U3 : NAND2_X1 port map( A1 => B(26), A2 => n12, ZN => n9);
   U4 : INV_X1 port map( A => n13, ZN => n11);
   U5 : INV_X1 port map( A => n13, ZN => n12);
   U6 : MUX2_X1 port map( A => A(19), B => B(19), S => S, Z => Z(19));
   U7 : MUX2_X1 port map( A => A(15), B => B(15), S => S, Z => Z(15));
   U8 : NAND2_X1 port map( A1 => A(17), A2 => n14, ZN => n2);
   U9 : NAND2_X1 port map( A1 => B(17), A2 => n11, ZN => n3);
   U10 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Z(17));
   U11 : NAND2_X1 port map( A1 => A(28), A2 => n14, ZN => n4);
   U12 : NAND2_X1 port map( A1 => B(28), A2 => n11, ZN => n5);
   U13 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Z(28));
   U14 : NAND2_X1 port map( A1 => A(30), A2 => n13, ZN => n6);
   U15 : NAND2_X1 port map( A1 => B(30), A2 => n11, ZN => n7);
   U16 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Z(30));
   U17 : NAND2_X1 port map( A1 => A(26), A2 => n14, ZN => n8);
   U18 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => Z(26));
   U19 : INV_X1 port map( A => n14, ZN => n10);
   U20 : INV_X1 port map( A => S, ZN => n13);
   U21 : INV_X1 port map( A => S, ZN => n14);
   U22 : MUX2_X1 port map( A => A(0), B => B(0), S => n10, Z => Z(0));
   U23 : MUX2_X1 port map( A => A(1), B => B(1), S => n10, Z => Z(1));
   U24 : MUX2_X1 port map( A => A(2), B => B(2), S => n10, Z => Z(2));
   U25 : MUX2_X1 port map( A => A(3), B => B(3), S => n10, Z => Z(3));
   U26 : MUX2_X1 port map( A => A(4), B => B(4), S => n10, Z => Z(4));
   U27 : MUX2_X1 port map( A => A(5), B => B(5), S => n10, Z => Z(5));
   U28 : MUX2_X1 port map( A => A(6), B => B(6), S => n10, Z => Z(6));
   U29 : MUX2_X1 port map( A => A(7), B => B(7), S => n10, Z => Z(7));
   U30 : MUX2_X1 port map( A => A(8), B => B(8), S => n10, Z => Z(8));
   U31 : MUX2_X1 port map( A => A(9), B => B(9), S => n10, Z => Z(9));
   U32 : MUX2_X1 port map( A => A(10), B => B(10), S => n10, Z => Z(10));
   U33 : MUX2_X1 port map( A => A(11), B => B(11), S => n10, Z => Z(11));
   U34 : MUX2_X1 port map( A => A(12), B => B(12), S => n11, Z => Z(12));
   U35 : MUX2_X1 port map( A => A(13), B => B(13), S => n11, Z => Z(13));
   U36 : MUX2_X1 port map( A => A(14), B => B(14), S => n11, Z => Z(14));
   U37 : MUX2_X1 port map( A => A(16), B => B(16), S => n11, Z => Z(16));
   U38 : MUX2_X1 port map( A => A(18), B => B(18), S => n11, Z => Z(18));
   U39 : MUX2_X1 port map( A => A(20), B => B(20), S => n11, Z => Z(20));
   U40 : MUX2_X1 port map( A => A(21), B => B(21), S => n11, Z => Z(21));
   U41 : MUX2_X1 port map( A => A(22), B => B(22), S => n11, Z => Z(22));
   U42 : AOI22_X1 port map( A1 => B(23), A2 => n12, B1 => A(23), B2 => n14, ZN 
                           => n15);
   U43 : INV_X1 port map( A => n15, ZN => Z(23));
   U44 : MUX2_X1 port map( A => A(24), B => B(24), S => n11, Z => Z(24));
   U45 : MUX2_X1 port map( A => A(25), B => B(25), S => n12, Z => Z(25));
   U46 : AOI22_X1 port map( A1 => A(27), A2 => n13, B1 => B(27), B2 => n12, ZN 
                           => n16);
   U47 : INV_X1 port map( A => n16, ZN => Z(27));
   U48 : AOI22_X1 port map( A1 => A(31), A2 => n13, B1 => B(31), B2 => n12, ZN 
                           => n17);
   U49 : INV_X1 port map( A => n17, ZN => Z(31));

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HazardDetection is

   port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : in std_logic_vector (4
         downto 0);  DRAM_R : in std_logic;  INS_IN, PC_IN : in 
         std_logic_vector (31 downto 0);  Bubble : out std_logic;  HDU_INS_OUT,
         HDU_PC_OUT, HDU_NPC_OUT : out std_logic_vector (31 downto 0));

end HazardDetection;

architecture SYN_arch of HazardDetection is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component HazardDetection_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n7, n8, n11, n1, n2, n3, n4, n5, n6, n9, n10, n12, n13, n14, n15, n16
      , n_1825 : std_logic;

begin
   HDU_INS_OUT <= ( INS_IN(31), INS_IN(30), INS_IN(29), INS_IN(28), INS_IN(27),
      INS_IN(26), INS_IN(25), INS_IN(24), INS_IN(23), INS_IN(22), INS_IN(21), 
      INS_IN(20), INS_IN(19), INS_IN(18), INS_IN(17), INS_IN(16), INS_IN(15), 
      INS_IN(14), INS_IN(13), INS_IN(12), INS_IN(11), INS_IN(10), INS_IN(9), 
      INS_IN(8), INS_IN(7), INS_IN(6), INS_IN(5), INS_IN(4), INS_IN(3), 
      INS_IN(2), INS_IN(1), INS_IN(0) );
   HDU_NPC_OUT <= ( PC_IN(31), PC_IN(30), PC_IN(29), PC_IN(28), PC_IN(27), 
      PC_IN(26), PC_IN(25), PC_IN(24), PC_IN(23), PC_IN(22), PC_IN(21), 
      PC_IN(20), PC_IN(19), PC_IN(18), PC_IN(17), PC_IN(16), PC_IN(15), 
      PC_IN(14), PC_IN(13), PC_IN(12), PC_IN(11), PC_IN(10), PC_IN(9), PC_IN(8)
      , PC_IN(7), PC_IN(6), PC_IN(5), PC_IN(4), PC_IN(3), PC_IN(2), PC_IN(1), 
      PC_IN(0) );
   
   n7 <= '0';
   n8 <= '1';
   n11 <= '0';
   sub_25 : HazardDetection_DW01_sub_0 port map( A(31) => PC_IN(31), A(30) => 
                           PC_IN(30), A(29) => PC_IN(29), A(28) => PC_IN(28), 
                           A(27) => PC_IN(27), A(26) => PC_IN(26), A(25) => 
                           PC_IN(25), A(24) => PC_IN(24), A(23) => PC_IN(23), 
                           A(22) => PC_IN(22), A(21) => PC_IN(21), A(20) => 
                           PC_IN(20), A(19) => PC_IN(19), A(18) => PC_IN(18), 
                           A(17) => PC_IN(17), A(16) => PC_IN(16), A(15) => 
                           PC_IN(15), A(14) => PC_IN(14), A(13) => PC_IN(13), 
                           A(12) => PC_IN(12), A(11) => PC_IN(11), A(10) => 
                           PC_IN(10), A(9) => PC_IN(9), A(8) => PC_IN(8), A(7) 
                           => PC_IN(7), A(6) => PC_IN(6), A(5) => PC_IN(5), 
                           A(4) => PC_IN(4), A(3) => PC_IN(3), A(2) => PC_IN(2)
                           , A(1) => PC_IN(1), A(0) => PC_IN(0), B(31) => n7, 
                           B(30) => n7, B(29) => n7, B(28) => n7, B(27) => n7, 
                           B(26) => n7, B(25) => n7, B(24) => n7, B(23) => n7, 
                           B(22) => n7, B(21) => n7, B(20) => n7, B(19) => n7, 
                           B(18) => n7, B(17) => n7, B(16) => n7, B(15) => n7, 
                           B(14) => n7, B(13) => n7, B(12) => n7, B(11) => n7, 
                           B(10) => n7, B(9) => n7, B(8) => n7, B(7) => n7, 
                           B(6) => n7, B(5) => n7, B(4) => n7, B(3) => n7, B(2)
                           => n8, B(1) => n7, B(0) => n7, CI => n11, DIFF(31) 
                           => HDU_PC_OUT(31), DIFF(30) => HDU_PC_OUT(30), 
                           DIFF(29) => HDU_PC_OUT(29), DIFF(28) => 
                           HDU_PC_OUT(28), DIFF(27) => HDU_PC_OUT(27), DIFF(26)
                           => HDU_PC_OUT(26), DIFF(25) => HDU_PC_OUT(25), 
                           DIFF(24) => HDU_PC_OUT(24), DIFF(23) => 
                           HDU_PC_OUT(23), DIFF(22) => HDU_PC_OUT(22), DIFF(21)
                           => HDU_PC_OUT(21), DIFF(20) => HDU_PC_OUT(20), 
                           DIFF(19) => HDU_PC_OUT(19), DIFF(18) => 
                           HDU_PC_OUT(18), DIFF(17) => HDU_PC_OUT(17), DIFF(16)
                           => HDU_PC_OUT(16), DIFF(15) => HDU_PC_OUT(15), 
                           DIFF(14) => HDU_PC_OUT(14), DIFF(13) => 
                           HDU_PC_OUT(13), DIFF(12) => HDU_PC_OUT(12), DIFF(11)
                           => HDU_PC_OUT(11), DIFF(10) => HDU_PC_OUT(10), 
                           DIFF(9) => HDU_PC_OUT(9), DIFF(8) => HDU_PC_OUT(8), 
                           DIFF(7) => HDU_PC_OUT(7), DIFF(6) => HDU_PC_OUT(6), 
                           DIFF(5) => HDU_PC_OUT(5), DIFF(4) => HDU_PC_OUT(4), 
                           DIFF(3) => HDU_PC_OUT(3), DIFF(2) => HDU_PC_OUT(2), 
                           DIFF(1) => HDU_PC_OUT(1), DIFF(0) => HDU_PC_OUT(0), 
                           CO => n_1825);
   U4 : AND3_X1 port map( A1 => DRAM_R, A2 => n1, A3 => RST, ZN => Bubble);
   U5 : OAI33_X1 port map( A1 => n2, A2 => n3, A3 => n4, B1 => n5, B2 => n6, B3
                           => n9, ZN => n1);
   U6 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RS2(4), Z => n9);
   U8 : XOR2_X1 port map( A => ADD_WR(2), B => ADD_RS2(2), Z => n6);
   U9 : NAND3_X1 port map( A1 => n10, A2 => n12, A3 => n13, ZN => n5);
   U11 : XNOR2_X1 port map( A => ADD_WR(0), B => ADD_RS2(0), ZN => n13);
   U12 : XNOR2_X1 port map( A => ADD_WR(1), B => ADD_RS2(1), ZN => n12);
   U13 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS2(3), ZN => n10);
   U14 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RS1(4), Z => n4);
   U15 : XOR2_X1 port map( A => ADD_WR(2), B => ADD_RS1(2), Z => n3);
   U16 : NAND3_X1 port map( A1 => n14, A2 => n15, A3 => n16, ZN => n2);
   U17 : XNOR2_X1 port map( A => ADD_WR(0), B => ADD_RS1(0), ZN => n16);
   U18 : XNOR2_X1 port map( A => ADD_WR(1), B => ADD_RS1(1), ZN => n15);
   U19 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS1(3), ZN => n14);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Writeback is

   port( WB_MUX_SEL : in std_logic;  DATA_IN, ALU_RES_IN : in std_logic_vector 
         (31 downto 0);  ADD_WR_IN : in std_logic_vector (4 downto 0);  
         DATA_OUT : out std_logic_vector (31 downto 0);  ADD_WR_OUT : out 
         std_logic_vector (4 downto 0));

end Writeback;

architecture SYN_struct of Writeback is

   component mux21_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;

begin
   ADD_WR_OUT <= ( ADD_WR_IN(4), ADD_WR_IN(3), ADD_WR_IN(2), ADD_WR_IN(1), 
      ADD_WR_IN(0) );
   
   WBmux : mux21_NBIT32_2 port map( A(31) => DATA_IN(31), A(30) => DATA_IN(30),
                           A(29) => DATA_IN(29), A(28) => DATA_IN(28), A(27) =>
                           DATA_IN(27), A(26) => DATA_IN(26), A(25) => 
                           DATA_IN(25), A(24) => DATA_IN(24), A(23) => 
                           DATA_IN(23), A(22) => DATA_IN(22), A(21) => 
                           DATA_IN(21), A(20) => DATA_IN(20), A(19) => 
                           DATA_IN(19), A(18) => DATA_IN(18), A(17) => 
                           DATA_IN(17), A(16) => DATA_IN(16), A(15) => 
                           DATA_IN(15), A(14) => DATA_IN(14), A(13) => 
                           DATA_IN(13), A(12) => DATA_IN(12), A(11) => 
                           DATA_IN(11), A(10) => DATA_IN(10), A(9) => 
                           DATA_IN(9), A(8) => DATA_IN(8), A(7) => DATA_IN(7), 
                           A(6) => DATA_IN(6), A(5) => DATA_IN(5), A(4) => 
                           DATA_IN(4), A(3) => DATA_IN(3), A(2) => DATA_IN(2), 
                           A(1) => DATA_IN(1), A(0) => DATA_IN(0), B(31) => 
                           ALU_RES_IN(31), B(30) => ALU_RES_IN(30), B(29) => 
                           ALU_RES_IN(29), B(28) => ALU_RES_IN(28), B(27) => 
                           ALU_RES_IN(27), B(26) => ALU_RES_IN(26), B(25) => 
                           ALU_RES_IN(25), B(24) => ALU_RES_IN(24), B(23) => 
                           ALU_RES_IN(23), B(22) => ALU_RES_IN(22), B(21) => 
                           ALU_RES_IN(21), B(20) => ALU_RES_IN(20), B(19) => 
                           ALU_RES_IN(19), B(18) => ALU_RES_IN(18), B(17) => 
                           ALU_RES_IN(17), B(16) => ALU_RES_IN(16), B(15) => 
                           ALU_RES_IN(15), B(14) => ALU_RES_IN(14), B(13) => 
                           ALU_RES_IN(13), B(12) => ALU_RES_IN(12), B(11) => 
                           ALU_RES_IN(11), B(10) => ALU_RES_IN(10), B(9) => 
                           ALU_RES_IN(9), B(8) => ALU_RES_IN(8), B(7) => 
                           ALU_RES_IN(7), B(6) => ALU_RES_IN(6), B(5) => 
                           ALU_RES_IN(5), B(4) => ALU_RES_IN(4), B(3) => 
                           ALU_RES_IN(3), B(2) => ALU_RES_IN(2), B(1) => 
                           ALU_RES_IN(1), B(0) => ALU_RES_IN(0), S => 
                           WB_MUX_SEL, Z(31) => DATA_OUT(31), Z(30) => 
                           DATA_OUT(30), Z(29) => DATA_OUT(29), Z(28) => 
                           DATA_OUT(28), Z(27) => DATA_OUT(27), Z(26) => 
                           DATA_OUT(26), Z(25) => DATA_OUT(25), Z(24) => 
                           DATA_OUT(24), Z(23) => DATA_OUT(23), Z(22) => 
                           DATA_OUT(22), Z(21) => DATA_OUT(21), Z(20) => 
                           DATA_OUT(20), Z(19) => DATA_OUT(19), Z(18) => 
                           DATA_OUT(18), Z(17) => DATA_OUT(17), Z(16) => 
                           DATA_OUT(16), Z(15) => DATA_OUT(15), Z(14) => 
                           DATA_OUT(14), Z(13) => DATA_OUT(13), Z(12) => 
                           DATA_OUT(12), Z(11) => DATA_OUT(11), Z(10) => 
                           DATA_OUT(10), Z(9) => DATA_OUT(9), Z(8) => 
                           DATA_OUT(8), Z(7) => DATA_OUT(7), Z(6) => 
                           DATA_OUT(6), Z(5) => DATA_OUT(5), Z(4) => 
                           DATA_OUT(4), Z(3) => DATA_OUT(3), Z(2) => 
                           DATA_OUT(2), Z(1) => DATA_OUT(1), Z(0) => 
                           DATA_OUT(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Memory is

   port( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, DRAM_EN_IN : in std_logic; 
         PC_SEL : in std_logic_vector (1 downto 0);  NPC_IN, NPC_ABS, NPC_REL, 
         ALU_RES_IN, B_IN : in std_logic_vector (31 downto 0);  ADD_WR_IN : in 
         std_logic_vector (4 downto 0);  DRAM_DATA_IN : in std_logic_vector (31
         downto 0);  PC_OUT : out std_logic_vector (31 downto 0);  DRAM_EN_OUT,
         DRAM_R_OUT, DRAM_W_OUT : out std_logic;  DRAM_ADDR_OUT, DRAM_DATA_OUT,
         DATA_OUT, ALU_RES_OUT, OP_MEM : out std_logic_vector (31 downto 0);  
         ADD_WR_MEM, ADD_WR_OUT : out std_logic_vector (4 downto 0));

end Memory;

architecture SYN_struct of Memory is

   component mux41_NBIT32_2
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component regn_N32_1
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N5_1
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N32_2
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port : std_logic;

begin
   DRAM_EN_OUT <= DRAM_EN_IN;
   DRAM_R_OUT <= DRAM_R_IN;
   DRAM_W_OUT <= DRAM_W_IN;
   DRAM_ADDR_OUT <= ( ALU_RES_IN(31), ALU_RES_IN(30), ALU_RES_IN(29), 
      ALU_RES_IN(28), ALU_RES_IN(27), ALU_RES_IN(26), ALU_RES_IN(25), 
      ALU_RES_IN(24), ALU_RES_IN(23), ALU_RES_IN(22), ALU_RES_IN(21), 
      ALU_RES_IN(20), ALU_RES_IN(19), ALU_RES_IN(18), ALU_RES_IN(17), 
      ALU_RES_IN(16), ALU_RES_IN(15), ALU_RES_IN(14), ALU_RES_IN(13), 
      ALU_RES_IN(12), ALU_RES_IN(11), ALU_RES_IN(10), ALU_RES_IN(9), 
      ALU_RES_IN(8), ALU_RES_IN(7), ALU_RES_IN(6), ALU_RES_IN(5), ALU_RES_IN(4)
      , ALU_RES_IN(3), ALU_RES_IN(2), ALU_RES_IN(1), ALU_RES_IN(0) );
   DRAM_DATA_OUT <= ( B_IN(31), B_IN(30), B_IN(29), B_IN(28), B_IN(27), 
      B_IN(26), B_IN(25), B_IN(24), B_IN(23), B_IN(22), B_IN(21), B_IN(20), 
      B_IN(19), B_IN(18), B_IN(17), B_IN(16), B_IN(15), B_IN(14), B_IN(13), 
      B_IN(12), B_IN(11), B_IN(10), B_IN(9), B_IN(8), B_IN(7), B_IN(6), B_IN(5)
      , B_IN(4), B_IN(3), B_IN(2), B_IN(1), B_IN(0) );
   OP_MEM <= ( ALU_RES_IN(31), ALU_RES_IN(30), ALU_RES_IN(29), ALU_RES_IN(28), 
      ALU_RES_IN(27), ALU_RES_IN(26), ALU_RES_IN(25), ALU_RES_IN(24), 
      ALU_RES_IN(23), ALU_RES_IN(22), ALU_RES_IN(21), ALU_RES_IN(20), 
      ALU_RES_IN(19), ALU_RES_IN(18), ALU_RES_IN(17), ALU_RES_IN(16), 
      ALU_RES_IN(15), ALU_RES_IN(14), ALU_RES_IN(13), ALU_RES_IN(12), 
      ALU_RES_IN(11), ALU_RES_IN(10), ALU_RES_IN(9), ALU_RES_IN(8), 
      ALU_RES_IN(7), ALU_RES_IN(6), ALU_RES_IN(5), ALU_RES_IN(4), ALU_RES_IN(3)
      , ALU_RES_IN(2), ALU_RES_IN(1), ALU_RES_IN(0) );
   ADD_WR_MEM <= ( ADD_WR_IN(4), ADD_WR_IN(3), ADD_WR_IN(2), ADD_WR_IN(1), 
      ADD_WR_IN(0) );
   
   X_Logic0_port <= '0';
   LMD : regn_N32_2 port map( DIN(31) => DRAM_DATA_IN(31), DIN(30) => 
                           DRAM_DATA_IN(30), DIN(29) => DRAM_DATA_IN(29), 
                           DIN(28) => DRAM_DATA_IN(28), DIN(27) => 
                           DRAM_DATA_IN(27), DIN(26) => DRAM_DATA_IN(26), 
                           DIN(25) => DRAM_DATA_IN(25), DIN(24) => 
                           DRAM_DATA_IN(24), DIN(23) => DRAM_DATA_IN(23), 
                           DIN(22) => DRAM_DATA_IN(22), DIN(21) => 
                           DRAM_DATA_IN(21), DIN(20) => DRAM_DATA_IN(20), 
                           DIN(19) => DRAM_DATA_IN(19), DIN(18) => 
                           DRAM_DATA_IN(18), DIN(17) => DRAM_DATA_IN(17), 
                           DIN(16) => DRAM_DATA_IN(16), DIN(15) => 
                           DRAM_DATA_IN(15), DIN(14) => DRAM_DATA_IN(14), 
                           DIN(13) => DRAM_DATA_IN(13), DIN(12) => 
                           DRAM_DATA_IN(12), DIN(11) => DRAM_DATA_IN(11), 
                           DIN(10) => DRAM_DATA_IN(10), DIN(9) => 
                           DRAM_DATA_IN(9), DIN(8) => DRAM_DATA_IN(8), DIN(7) 
                           => DRAM_DATA_IN(7), DIN(6) => DRAM_DATA_IN(6), 
                           DIN(5) => DRAM_DATA_IN(5), DIN(4) => DRAM_DATA_IN(4)
                           , DIN(3) => DRAM_DATA_IN(3), DIN(2) => 
                           DRAM_DATA_IN(2), DIN(1) => DRAM_DATA_IN(1), DIN(0) 
                           => DRAM_DATA_IN(0), CLK => CLK, EN => MEM_EN_IN, RST
                           => RST, DOUT(31) => DATA_OUT(31), DOUT(30) => 
                           DATA_OUT(30), DOUT(29) => DATA_OUT(29), DOUT(28) => 
                           DATA_OUT(28), DOUT(27) => DATA_OUT(27), DOUT(26) => 
                           DATA_OUT(26), DOUT(25) => DATA_OUT(25), DOUT(24) => 
                           DATA_OUT(24), DOUT(23) => DATA_OUT(23), DOUT(22) => 
                           DATA_OUT(22), DOUT(21) => DATA_OUT(21), DOUT(20) => 
                           DATA_OUT(20), DOUT(19) => DATA_OUT(19), DOUT(18) => 
                           DATA_OUT(18), DOUT(17) => DATA_OUT(17), DOUT(16) => 
                           DATA_OUT(16), DOUT(15) => DATA_OUT(15), DOUT(14) => 
                           DATA_OUT(14), DOUT(13) => DATA_OUT(13), DOUT(12) => 
                           DATA_OUT(12), DOUT(11) => DATA_OUT(11), DOUT(10) => 
                           DATA_OUT(10), DOUT(9) => DATA_OUT(9), DOUT(8) => 
                           DATA_OUT(8), DOUT(7) => DATA_OUT(7), DOUT(6) => 
                           DATA_OUT(6), DOUT(5) => DATA_OUT(5), DOUT(4) => 
                           DATA_OUT(4), DOUT(3) => DATA_OUT(3), DOUT(2) => 
                           DATA_OUT(2), DOUT(1) => DATA_OUT(1), DOUT(0) => 
                           DATA_OUT(0));
   reg0 : regn_N5_1 port map( DIN(4) => ADD_WR_IN(4), DIN(3) => ADD_WR_IN(3), 
                           DIN(2) => ADD_WR_IN(2), DIN(1) => ADD_WR_IN(1), 
                           DIN(0) => ADD_WR_IN(0), CLK => CLK, EN => MEM_EN_IN,
                           RST => RST, DOUT(4) => ADD_WR_OUT(4), DOUT(3) => 
                           ADD_WR_OUT(3), DOUT(2) => ADD_WR_OUT(2), DOUT(1) => 
                           ADD_WR_OUT(1), DOUT(0) => ADD_WR_OUT(0));
   reg1 : regn_N32_1 port map( DIN(31) => ALU_RES_IN(31), DIN(30) => 
                           ALU_RES_IN(30), DIN(29) => ALU_RES_IN(29), DIN(28) 
                           => ALU_RES_IN(28), DIN(27) => ALU_RES_IN(27), 
                           DIN(26) => ALU_RES_IN(26), DIN(25) => ALU_RES_IN(25)
                           , DIN(24) => ALU_RES_IN(24), DIN(23) => 
                           ALU_RES_IN(23), DIN(22) => ALU_RES_IN(22), DIN(21) 
                           => ALU_RES_IN(21), DIN(20) => ALU_RES_IN(20), 
                           DIN(19) => ALU_RES_IN(19), DIN(18) => ALU_RES_IN(18)
                           , DIN(17) => ALU_RES_IN(17), DIN(16) => 
                           ALU_RES_IN(16), DIN(15) => ALU_RES_IN(15), DIN(14) 
                           => ALU_RES_IN(14), DIN(13) => ALU_RES_IN(13), 
                           DIN(12) => ALU_RES_IN(12), DIN(11) => ALU_RES_IN(11)
                           , DIN(10) => ALU_RES_IN(10), DIN(9) => ALU_RES_IN(9)
                           , DIN(8) => ALU_RES_IN(8), DIN(7) => ALU_RES_IN(7), 
                           DIN(6) => ALU_RES_IN(6), DIN(5) => ALU_RES_IN(5), 
                           DIN(4) => ALU_RES_IN(4), DIN(3) => ALU_RES_IN(3), 
                           DIN(2) => ALU_RES_IN(2), DIN(1) => ALU_RES_IN(1), 
                           DIN(0) => ALU_RES_IN(0), CLK => CLK, EN => MEM_EN_IN
                           , RST => RST, DOUT(31) => ALU_RES_OUT(31), DOUT(30) 
                           => ALU_RES_OUT(30), DOUT(29) => ALU_RES_OUT(29), 
                           DOUT(28) => ALU_RES_OUT(28), DOUT(27) => 
                           ALU_RES_OUT(27), DOUT(26) => ALU_RES_OUT(26), 
                           DOUT(25) => ALU_RES_OUT(25), DOUT(24) => 
                           ALU_RES_OUT(24), DOUT(23) => ALU_RES_OUT(23), 
                           DOUT(22) => ALU_RES_OUT(22), DOUT(21) => 
                           ALU_RES_OUT(21), DOUT(20) => ALU_RES_OUT(20), 
                           DOUT(19) => ALU_RES_OUT(19), DOUT(18) => 
                           ALU_RES_OUT(18), DOUT(17) => ALU_RES_OUT(17), 
                           DOUT(16) => ALU_RES_OUT(16), DOUT(15) => 
                           ALU_RES_OUT(15), DOUT(14) => ALU_RES_OUT(14), 
                           DOUT(13) => ALU_RES_OUT(13), DOUT(12) => 
                           ALU_RES_OUT(12), DOUT(11) => ALU_RES_OUT(11), 
                           DOUT(10) => ALU_RES_OUT(10), DOUT(9) => 
                           ALU_RES_OUT(9), DOUT(8) => ALU_RES_OUT(8), DOUT(7) 
                           => ALU_RES_OUT(7), DOUT(6) => ALU_RES_OUT(6), 
                           DOUT(5) => ALU_RES_OUT(5), DOUT(4) => ALU_RES_OUT(4)
                           , DOUT(3) => ALU_RES_OUT(3), DOUT(2) => 
                           ALU_RES_OUT(2), DOUT(1) => ALU_RES_OUT(1), DOUT(0) 
                           => ALU_RES_OUT(0));
   PCsel : mux41_NBIT32_2 port map( A(31) => NPC_IN(31), A(30) => NPC_IN(30), 
                           A(29) => NPC_IN(29), A(28) => NPC_IN(28), A(27) => 
                           NPC_IN(27), A(26) => NPC_IN(26), A(25) => NPC_IN(25)
                           , A(24) => NPC_IN(24), A(23) => NPC_IN(23), A(22) =>
                           NPC_IN(22), A(21) => NPC_IN(21), A(20) => NPC_IN(20)
                           , A(19) => NPC_IN(19), A(18) => NPC_IN(18), A(17) =>
                           NPC_IN(17), A(16) => NPC_IN(16), A(15) => NPC_IN(15)
                           , A(14) => NPC_IN(14), A(13) => NPC_IN(13), A(12) =>
                           NPC_IN(12), A(11) => NPC_IN(11), A(10) => NPC_IN(10)
                           , A(9) => NPC_IN(9), A(8) => NPC_IN(8), A(7) => 
                           NPC_IN(7), A(6) => NPC_IN(6), A(5) => NPC_IN(5), 
                           A(4) => NPC_IN(4), A(3) => NPC_IN(3), A(2) => 
                           NPC_IN(2), A(1) => NPC_IN(1), A(0) => NPC_IN(0), 
                           B(31) => NPC_REL(31), B(30) => NPC_REL(30), B(29) =>
                           NPC_REL(29), B(28) => NPC_REL(28), B(27) => 
                           NPC_REL(27), B(26) => NPC_REL(26), B(25) => 
                           NPC_REL(25), B(24) => NPC_REL(24), B(23) => 
                           NPC_REL(23), B(22) => NPC_REL(22), B(21) => 
                           NPC_REL(21), B(20) => NPC_REL(20), B(19) => 
                           NPC_REL(19), B(18) => NPC_REL(18), B(17) => 
                           NPC_REL(17), B(16) => NPC_REL(16), B(15) => 
                           NPC_REL(15), B(14) => NPC_REL(14), B(13) => 
                           NPC_REL(13), B(12) => NPC_REL(12), B(11) => 
                           NPC_REL(11), B(10) => NPC_REL(10), B(9) => 
                           NPC_REL(9), B(8) => NPC_REL(8), B(7) => NPC_REL(7), 
                           B(6) => NPC_REL(6), B(5) => NPC_REL(5), B(4) => 
                           NPC_REL(4), B(3) => NPC_REL(3), B(2) => NPC_REL(2), 
                           B(1) => NPC_REL(1), B(0) => NPC_REL(0), C(31) => 
                           NPC_ABS(31), C(30) => NPC_ABS(30), C(29) => 
                           NPC_ABS(29), C(28) => NPC_ABS(28), C(27) => 
                           NPC_ABS(27), C(26) => NPC_ABS(26), C(25) => 
                           NPC_ABS(25), C(24) => NPC_ABS(24), C(23) => 
                           NPC_ABS(23), C(22) => NPC_ABS(22), C(21) => 
                           NPC_ABS(21), C(20) => NPC_ABS(20), C(19) => 
                           NPC_ABS(19), C(18) => NPC_ABS(18), C(17) => 
                           NPC_ABS(17), C(16) => NPC_ABS(16), C(15) => 
                           NPC_ABS(15), C(14) => NPC_ABS(14), C(13) => 
                           NPC_ABS(13), C(12) => NPC_ABS(12), C(11) => 
                           NPC_ABS(11), C(10) => NPC_ABS(10), C(9) => 
                           NPC_ABS(9), C(8) => NPC_ABS(8), C(7) => NPC_ABS(7), 
                           C(6) => NPC_ABS(6), C(5) => NPC_ABS(5), C(4) => 
                           NPC_ABS(4), C(3) => NPC_ABS(3), C(2) => NPC_ABS(2), 
                           C(1) => NPC_ABS(1), C(0) => NPC_ABS(0), D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => X_Logic0_port, D(25) => 
                           X_Logic0_port, D(24) => X_Logic0_port, D(23) => 
                           X_Logic0_port, D(22) => X_Logic0_port, D(21) => 
                           X_Logic0_port, D(20) => X_Logic0_port, D(19) => 
                           X_Logic0_port, D(18) => X_Logic0_port, D(17) => 
                           X_Logic0_port, D(16) => X_Logic0_port, D(15) => 
                           X_Logic0_port, D(14) => X_Logic0_port, D(13) => 
                           X_Logic0_port, D(12) => X_Logic0_port, D(11) => 
                           X_Logic0_port, D(10) => X_Logic0_port, D(9) => 
                           X_Logic0_port, D(8) => X_Logic0_port, D(7) => 
                           X_Logic0_port, D(6) => X_Logic0_port, D(5) => 
                           X_Logic0_port, D(4) => X_Logic0_port, D(3) => 
                           X_Logic0_port, D(2) => X_Logic0_port, D(1) => 
                           X_Logic0_port, D(0) => X_Logic0_port, S(1) => 
                           PC_SEL(1), S(0) => PC_SEL(0), Z(31) => PC_OUT(31), 
                           Z(30) => PC_OUT(30), Z(29) => PC_OUT(29), Z(28) => 
                           PC_OUT(28), Z(27) => PC_OUT(27), Z(26) => PC_OUT(26)
                           , Z(25) => PC_OUT(25), Z(24) => PC_OUT(24), Z(23) =>
                           PC_OUT(23), Z(22) => PC_OUT(22), Z(21) => PC_OUT(21)
                           , Z(20) => PC_OUT(20), Z(19) => PC_OUT(19), Z(18) =>
                           PC_OUT(18), Z(17) => PC_OUT(17), Z(16) => PC_OUT(16)
                           , Z(15) => PC_OUT(15), Z(14) => PC_OUT(14), Z(13) =>
                           PC_OUT(13), Z(12) => PC_OUT(12), Z(11) => PC_OUT(11)
                           , Z(10) => PC_OUT(10), Z(9) => PC_OUT(9), Z(8) => 
                           PC_OUT(8), Z(7) => PC_OUT(7), Z(6) => PC_OUT(6), 
                           Z(5) => PC_OUT(5), Z(4) => PC_OUT(4), Z(3) => 
                           PC_OUT(3), Z(2) => PC_OUT(2), Z(1) => PC_OUT(1), 
                           Z(0) => PC_OUT(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ff_0 is

   port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);

end ff_0;

architecture SYN_bhv of ff_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n3, CK => CLK, RN => RST, Q => Q, QN => n2);
   U2 : OAI21_X1 port map( B1 => n2, B2 => EN, A => n1, ZN => n3);
   U3 : NAND2_X1 port map( A1 => EN, A2 => D, ZN => n1);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute is

   port( CLK, RST, MUX_A_SEL : in std_logic;  MUX_B_SEL : in std_logic_vector 
         (1 downto 0);  ALU_OPC : in std_logic_vector (0 to 3);  ALU_OUTREG_EN 
         : in std_logic;  JUMP_TYPE : in std_logic_vector (1 downto 0);  PC_IN,
         A_IN, B_IN, IMM_IN : in std_logic_vector (31 downto 0);  ADD_WR_IN, 
         ADD_RS1_IN, ADD_RS2_IN, ADD_WR_MEM, ADD_WR_WB : in std_logic_vector (4
         downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;  OP_MEM, OP_WB : in 
         std_logic_vector (31 downto 0);  PC_SEL : out std_logic_vector (1 
         downto 0);  ZERO_FLAG : out std_logic;  NPC_ABS, NPC_REL, ALU_RES, 
         B_OUT : out std_logic_vector (31 downto 0);  ADD_WR_OUT : out 
         std_logic_vector (4 downto 0));

end Execute;

architecture SYN_struct of Execute is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component Execute_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component Execute_DW01_add_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component regn_N32_3
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_4
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N5_2
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N32_5
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_6
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component ALU_NBIT32
      port( OP1, OP2 : in std_logic_vector (31 downto 0);  ALU_OPC : in 
            std_logic_vector (0 to 3);  ALU_RES : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux41_NBIT32_3
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux21_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux41_NBIT32_4
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux41_NBIT32_0
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component FWD_Unit
      port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB : in 
            std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;
            FWDA, FWDB : out std_logic_vector (1 downto 0));
   end component;
   
   component regn_N2
      port( DIN : in std_logic_vector (1 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (1 downto 0));
   end component;
   
   component ff_1
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Branch_Cond_Unit_NBIT32
      port( RST : in std_logic;  A : in std_logic_vector (31 downto 0);  
            ALU_OPC : in std_logic_vector (0 to 3);  JUMP_TYPE : in 
            std_logic_vector (1 downto 0);  PC_SEL : out std_logic_vector (1 
            downto 0);  ZERO : out std_logic);
   end component;
   
   signal ZERO_FLAG_port, sig_RST, sig_NPC_ABS_31_port, sig_NPC_ABS_30_port, 
      sig_NPC_ABS_29_port, sig_NPC_ABS_28_port, sig_NPC_ABS_27_port, 
      sig_NPC_ABS_26_port, sig_NPC_ABS_25_port, sig_NPC_ABS_24_port, 
      sig_NPC_ABS_23_port, sig_NPC_ABS_22_port, sig_NPC_ABS_21_port, 
      sig_NPC_ABS_20_port, sig_NPC_ABS_19_port, sig_NPC_ABS_18_port, 
      sig_NPC_ABS_17_port, sig_NPC_ABS_16_port, sig_NPC_ABS_15_port, 
      sig_NPC_ABS_14_port, sig_NPC_ABS_13_port, sig_NPC_ABS_12_port, 
      sig_NPC_ABS_11_port, sig_NPC_ABS_10_port, sig_NPC_ABS_9_port, 
      sig_NPC_ABS_8_port, sig_NPC_ABS_7_port, sig_NPC_ABS_6_port, 
      sig_NPC_ABS_5_port, sig_NPC_ABS_4_port, sig_NPC_ABS_3_port, 
      sig_NPC_ABS_2_port, sig_NPC_ABS_1_port, sig_NPC_ABS_0_port, 
      sig_NPC_REL_31_port, sig_NPC_REL_30_port, sig_NPC_REL_29_port, 
      sig_NPC_REL_28_port, sig_NPC_REL_27_port, sig_NPC_REL_26_port, 
      sig_NPC_REL_25_port, sig_NPC_REL_24_port, sig_NPC_REL_23_port, 
      sig_NPC_REL_22_port, sig_NPC_REL_21_port, sig_NPC_REL_20_port, 
      sig_NPC_REL_19_port, sig_NPC_REL_18_port, sig_NPC_REL_17_port, 
      sig_NPC_REL_16_port, sig_NPC_REL_15_port, sig_NPC_REL_14_port, 
      sig_NPC_REL_13_port, sig_NPC_REL_12_port, sig_NPC_REL_11_port, 
      sig_NPC_REL_10_port, sig_NPC_REL_9_port, sig_NPC_REL_8_port, 
      sig_NPC_REL_7_port, sig_NPC_REL_6_port, sig_NPC_REL_5_port, 
      sig_NPC_REL_4_port, sig_NPC_REL_3_port, sig_NPC_REL_2_port, 
      sig_NPC_REL_1_port, sig_NPC_REL_0_port, sig_PC_SEL_1_port, 
      sig_PC_SEL_0_port, sig_ZERO_FLAG, FWDA_1_port, FWDA_0_port, FWDB_1_port, 
      FWDB_0_port, OP2_FW_31_port, OP2_FW_30_port, OP2_FW_29_port, 
      OP2_FW_28_port, OP2_FW_27_port, OP2_FW_26_port, OP2_FW_25_port, 
      OP2_FW_24_port, OP2_FW_23_port, OP2_FW_22_port, OP2_FW_21_port, 
      OP2_FW_20_port, OP2_FW_19_port, OP2_FW_18_port, OP2_FW_17_port, 
      OP2_FW_16_port, OP2_FW_15_port, OP2_FW_14_port, OP2_FW_13_port, 
      OP2_FW_12_port, OP2_FW_11_port, OP2_FW_10_port, OP2_FW_9_port, 
      OP2_FW_8_port, OP2_FW_7_port, OP2_FW_6_port, OP2_FW_5_port, OP2_FW_4_port
      , OP2_FW_3_port, OP2_FW_2_port, OP2_FW_1_port, OP2_FW_0_port, 
      sig_OP1_31_port, sig_OP1_30_port, sig_OP1_29_port, sig_OP1_28_port, 
      sig_OP1_27_port, sig_OP1_26_port, sig_OP1_25_port, sig_OP1_24_port, 
      sig_OP1_23_port, sig_OP1_22_port, sig_OP1_21_port, sig_OP1_20_port, 
      sig_OP1_19_port, sig_OP1_18_port, sig_OP1_17_port, sig_OP1_16_port, 
      sig_OP1_15_port, sig_OP1_14_port, sig_OP1_13_port, sig_OP1_12_port, 
      sig_OP1_11_port, sig_OP1_10_port, sig_OP1_9_port, sig_OP1_8_port, 
      sig_OP1_7_port, sig_OP1_6_port, sig_OP1_5_port, sig_OP1_4_port, 
      sig_OP1_3_port, sig_OP1_2_port, sig_OP1_1_port, sig_OP1_0_port, 
      sig_OP2_31_port, sig_OP2_30_port, sig_OP2_29_port, sig_OP2_28_port, 
      sig_OP2_27_port, sig_OP2_26_port, sig_OP2_25_port, sig_OP2_24_port, 
      sig_OP2_23_port, sig_OP2_22_port, sig_OP2_21_port, sig_OP2_20_port, 
      sig_OP2_19_port, sig_OP2_18_port, sig_OP2_17_port, sig_OP2_16_port, 
      sig_OP2_15_port, sig_OP2_14_port, sig_OP2_13_port, sig_OP2_12_port, 
      sig_OP2_11_port, sig_OP2_10_port, sig_OP2_9_port, sig_OP2_8_port, 
      sig_OP2_7_port, sig_OP2_6_port, sig_OP2_5_port, sig_OP2_4_port, 
      sig_OP2_3_port, sig_OP2_2_port, sig_OP2_1_port, sig_OP2_0_port, 
      sig_ALU_RES_31_port, sig_ALU_RES_30_port, sig_ALU_RES_29_port, 
      sig_ALU_RES_28_port, sig_ALU_RES_27_port, sig_ALU_RES_26_port, 
      sig_ALU_RES_25_port, sig_ALU_RES_24_port, sig_ALU_RES_23_port, 
      sig_ALU_RES_22_port, sig_ALU_RES_21_port, sig_ALU_RES_20_port, 
      sig_ALU_RES_19_port, sig_ALU_RES_18_port, sig_ALU_RES_17_port, 
      sig_ALU_RES_16_port, sig_ALU_RES_15_port, sig_ALU_RES_14_port, 
      sig_ALU_RES_13_port, sig_ALU_RES_12_port, sig_ALU_RES_11_port, 
      sig_ALU_RES_10_port, sig_ALU_RES_9_port, sig_ALU_RES_8_port, 
      sig_ALU_RES_7_port, sig_ALU_RES_6_port, sig_ALU_RES_5_port, 
      sig_ALU_RES_4_port, sig_ALU_RES_3_port, sig_ALU_RES_2_port, 
      sig_ALU_RES_1_port, sig_ALU_RES_0_port, N9, N8, N7, N6, N5, N4, N31, N30,
      N3, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N2, N19, N18, N17, 
      N16, N15, N14, N13, N12, N11, N10, N1, N0, n1_port, n2_port, n3_port, 
      n4_port, n5_port, n6_port, n7_port, n_1826, n_1827 : std_logic;

begin
   ZERO_FLAG <= ZERO_FLAG_port;
   
   n7_port <= '1';
   n6_port <= '0';
   Branch_Cond : Branch_Cond_Unit_NBIT32 port map( RST => sig_RST, A(31) => 
                           sig_NPC_ABS_31_port, A(30) => sig_NPC_ABS_30_port, 
                           A(29) => sig_NPC_ABS_29_port, A(28) => 
                           sig_NPC_ABS_28_port, A(27) => sig_NPC_ABS_27_port, 
                           A(26) => sig_NPC_ABS_26_port, A(25) => 
                           sig_NPC_ABS_25_port, A(24) => sig_NPC_ABS_24_port, 
                           A(23) => sig_NPC_ABS_23_port, A(22) => 
                           sig_NPC_ABS_22_port, A(21) => sig_NPC_ABS_21_port, 
                           A(20) => sig_NPC_ABS_20_port, A(19) => 
                           sig_NPC_ABS_19_port, A(18) => sig_NPC_ABS_18_port, 
                           A(17) => sig_NPC_ABS_17_port, A(16) => 
                           sig_NPC_ABS_16_port, A(15) => sig_NPC_ABS_15_port, 
                           A(14) => sig_NPC_ABS_14_port, A(13) => 
                           sig_NPC_ABS_13_port, A(12) => sig_NPC_ABS_12_port, 
                           A(11) => sig_NPC_ABS_11_port, A(10) => 
                           sig_NPC_ABS_10_port, A(9) => sig_NPC_ABS_9_port, 
                           A(8) => sig_NPC_ABS_8_port, A(7) => 
                           sig_NPC_ABS_7_port, A(6) => sig_NPC_ABS_6_port, A(5)
                           => sig_NPC_ABS_5_port, A(4) => sig_NPC_ABS_4_port, 
                           A(3) => sig_NPC_ABS_3_port, A(2) => 
                           sig_NPC_ABS_2_port, A(1) => sig_NPC_ABS_1_port, A(0)
                           => sig_NPC_ABS_0_port, ALU_OPC(0) => ALU_OPC(0), 
                           ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => ALU_OPC(2), 
                           ALU_OPC(3) => ALU_OPC(3), JUMP_TYPE(1) => 
                           JUMP_TYPE(1), JUMP_TYPE(0) => JUMP_TYPE(0), 
                           PC_SEL(1) => sig_PC_SEL_1_port, PC_SEL(0) => 
                           sig_PC_SEL_0_port, ZERO => sig_ZERO_FLAG);
   ff0 : ff_1 port map( D => sig_ZERO_FLAG, CLK => CLK, EN => n7_port, RST => 
                           RST, Q => ZERO_FLAG_port);
   reg0 : regn_N2 port map( DIN(1) => sig_PC_SEL_1_port, DIN(0) => 
                           sig_PC_SEL_0_port, CLK => CLK, EN => n7_port, RST =>
                           RST, DOUT(1) => PC_SEL(1), DOUT(0) => PC_SEL(0));
   FWD : FWD_Unit port map( RST => sig_RST, ADD_RS1(4) => ADD_RS1_IN(4), 
                           ADD_RS1(3) => ADD_RS1_IN(3), ADD_RS1(2) => 
                           ADD_RS1_IN(2), ADD_RS1(1) => ADD_RS1_IN(1), 
                           ADD_RS1(0) => ADD_RS1_IN(0), ADD_RS2(4) => 
                           ADD_RS2_IN(4), ADD_RS2(3) => ADD_RS2_IN(3), 
                           ADD_RS2(2) => ADD_RS2_IN(2), ADD_RS2(1) => 
                           ADD_RS2_IN(1), ADD_RS2(0) => ADD_RS2_IN(0), 
                           ADD_WR_MEM(4) => ADD_WR_MEM(4), ADD_WR_MEM(3) => 
                           ADD_WR_MEM(3), ADD_WR_MEM(2) => ADD_WR_MEM(2), 
                           ADD_WR_MEM(1) => ADD_WR_MEM(1), ADD_WR_MEM(0) => 
                           ADD_WR_MEM(0), ADD_WR_WB(4) => ADD_WR_WB(4), 
                           ADD_WR_WB(3) => ADD_WR_WB(3), ADD_WR_WB(2) => 
                           ADD_WR_WB(2), ADD_WR_WB(1) => ADD_WR_WB(1), 
                           ADD_WR_WB(0) => ADD_WR_WB(0), RF_WE_MEM => RF_WE_MEM
                           , RF_WE_WB => RF_WE_WB, FWDA(1) => FWDA_1_port, 
                           FWDA(0) => FWDA_0_port, FWDB(1) => FWDB_1_port, 
                           FWDB(0) => FWDB_0_port);
   FW1 : mux41_NBIT32_0 port map( A(31) => A_IN(31), A(30) => A_IN(30), A(29) 
                           => A_IN(29), A(28) => A_IN(28), A(27) => A_IN(27), 
                           A(26) => A_IN(26), A(25) => A_IN(25), A(24) => 
                           A_IN(24), A(23) => A_IN(23), A(22) => A_IN(22), 
                           A(21) => A_IN(21), A(20) => A_IN(20), A(19) => 
                           A_IN(19), A(18) => A_IN(18), A(17) => A_IN(17), 
                           A(16) => A_IN(16), A(15) => A_IN(15), A(14) => 
                           A_IN(14), A(13) => A_IN(13), A(12) => A_IN(12), 
                           A(11) => A_IN(11), A(10) => A_IN(10), A(9) => 
                           A_IN(9), A(8) => A_IN(8), A(7) => A_IN(7), A(6) => 
                           A_IN(6), A(5) => A_IN(5), A(4) => A_IN(4), A(3) => 
                           A_IN(3), A(2) => A_IN(2), A(1) => A_IN(1), A(0) => 
                           A_IN(0), B(31) => OP_WB(31), B(30) => OP_WB(30), 
                           B(29) => OP_WB(29), B(28) => OP_WB(28), B(27) => 
                           OP_WB(27), B(26) => OP_WB(26), B(25) => OP_WB(25), 
                           B(24) => OP_WB(24), B(23) => OP_WB(23), B(22) => 
                           OP_WB(22), B(21) => OP_WB(21), B(20) => OP_WB(20), 
                           B(19) => OP_WB(19), B(18) => OP_WB(18), B(17) => 
                           OP_WB(17), B(16) => OP_WB(16), B(15) => OP_WB(15), 
                           B(14) => OP_WB(14), B(13) => OP_WB(13), B(12) => 
                           OP_WB(12), B(11) => OP_WB(11), B(10) => OP_WB(10), 
                           B(9) => OP_WB(9), B(8) => OP_WB(8), B(7) => OP_WB(7)
                           , B(6) => OP_WB(6), B(5) => OP_WB(5), B(4) => 
                           OP_WB(4), B(3) => OP_WB(3), B(2) => OP_WB(2), B(1) 
                           => OP_WB(1), B(0) => OP_WB(0), C(31) => OP_MEM(31), 
                           C(30) => OP_MEM(30), C(29) => OP_MEM(29), C(28) => 
                           OP_MEM(28), C(27) => OP_MEM(27), C(26) => OP_MEM(26)
                           , C(25) => OP_MEM(25), C(24) => OP_MEM(24), C(23) =>
                           OP_MEM(23), C(22) => OP_MEM(22), C(21) => OP_MEM(21)
                           , C(20) => OP_MEM(20), C(19) => OP_MEM(19), C(18) =>
                           OP_MEM(18), C(17) => OP_MEM(17), C(16) => OP_MEM(16)
                           , C(15) => OP_MEM(15), C(14) => OP_MEM(14), C(13) =>
                           OP_MEM(13), C(12) => OP_MEM(12), C(11) => OP_MEM(11)
                           , C(10) => OP_MEM(10), C(9) => OP_MEM(9), C(8) => 
                           OP_MEM(8), C(7) => OP_MEM(7), C(6) => OP_MEM(6), 
                           C(5) => OP_MEM(5), C(4) => OP_MEM(4), C(3) => 
                           OP_MEM(3), C(2) => OP_MEM(2), C(1) => OP_MEM(1), 
                           C(0) => OP_MEM(0), D(31) => n6_port, D(30) => 
                           n6_port, D(29) => n6_port, D(28) => n6_port, D(27) 
                           => n6_port, D(26) => n6_port, D(25) => n6_port, 
                           D(24) => n6_port, D(23) => n6_port, D(22) => n6_port
                           , D(21) => n6_port, D(20) => n6_port, D(19) => 
                           n6_port, D(18) => n6_port, D(17) => n6_port, D(16) 
                           => n6_port, D(15) => n6_port, D(14) => n6_port, 
                           D(13) => n6_port, D(12) => n6_port, D(11) => n6_port
                           , D(10) => n6_port, D(9) => n6_port, D(8) => n6_port
                           , D(7) => n6_port, D(6) => n6_port, D(5) => n6_port,
                           D(4) => n6_port, D(3) => n6_port, D(2) => n6_port, 
                           D(1) => n6_port, D(0) => n6_port, S(1) => 
                           FWDA_1_port, S(0) => FWDA_0_port, Z(31) => 
                           sig_NPC_ABS_31_port, Z(30) => sig_NPC_ABS_30_port, 
                           Z(29) => sig_NPC_ABS_29_port, Z(28) => 
                           sig_NPC_ABS_28_port, Z(27) => sig_NPC_ABS_27_port, 
                           Z(26) => sig_NPC_ABS_26_port, Z(25) => 
                           sig_NPC_ABS_25_port, Z(24) => sig_NPC_ABS_24_port, 
                           Z(23) => sig_NPC_ABS_23_port, Z(22) => 
                           sig_NPC_ABS_22_port, Z(21) => sig_NPC_ABS_21_port, 
                           Z(20) => sig_NPC_ABS_20_port, Z(19) => 
                           sig_NPC_ABS_19_port, Z(18) => sig_NPC_ABS_18_port, 
                           Z(17) => sig_NPC_ABS_17_port, Z(16) => 
                           sig_NPC_ABS_16_port, Z(15) => sig_NPC_ABS_15_port, 
                           Z(14) => sig_NPC_ABS_14_port, Z(13) => 
                           sig_NPC_ABS_13_port, Z(12) => sig_NPC_ABS_12_port, 
                           Z(11) => sig_NPC_ABS_11_port, Z(10) => 
                           sig_NPC_ABS_10_port, Z(9) => sig_NPC_ABS_9_port, 
                           Z(8) => sig_NPC_ABS_8_port, Z(7) => 
                           sig_NPC_ABS_7_port, Z(6) => sig_NPC_ABS_6_port, Z(5)
                           => sig_NPC_ABS_5_port, Z(4) => sig_NPC_ABS_4_port, 
                           Z(3) => sig_NPC_ABS_3_port, Z(2) => 
                           sig_NPC_ABS_2_port, Z(1) => sig_NPC_ABS_1_port, Z(0)
                           => sig_NPC_ABS_0_port);
   FW2 : mux41_NBIT32_4 port map( A(31) => B_IN(31), A(30) => B_IN(30), A(29) 
                           => B_IN(29), A(28) => B_IN(28), A(27) => B_IN(27), 
                           A(26) => B_IN(26), A(25) => B_IN(25), A(24) => 
                           B_IN(24), A(23) => B_IN(23), A(22) => B_IN(22), 
                           A(21) => B_IN(21), A(20) => B_IN(20), A(19) => 
                           B_IN(19), A(18) => B_IN(18), A(17) => B_IN(17), 
                           A(16) => B_IN(16), A(15) => B_IN(15), A(14) => 
                           B_IN(14), A(13) => B_IN(13), A(12) => B_IN(12), 
                           A(11) => B_IN(11), A(10) => B_IN(10), A(9) => 
                           B_IN(9), A(8) => B_IN(8), A(7) => B_IN(7), A(6) => 
                           B_IN(6), A(5) => B_IN(5), A(4) => B_IN(4), A(3) => 
                           B_IN(3), A(2) => B_IN(2), A(1) => B_IN(1), A(0) => 
                           B_IN(0), B(31) => OP_WB(31), B(30) => OP_WB(30), 
                           B(29) => OP_WB(29), B(28) => OP_WB(28), B(27) => 
                           OP_WB(27), B(26) => OP_WB(26), B(25) => OP_WB(25), 
                           B(24) => OP_WB(24), B(23) => OP_WB(23), B(22) => 
                           OP_WB(22), B(21) => OP_WB(21), B(20) => OP_WB(20), 
                           B(19) => OP_WB(19), B(18) => OP_WB(18), B(17) => 
                           OP_WB(17), B(16) => OP_WB(16), B(15) => OP_WB(15), 
                           B(14) => OP_WB(14), B(13) => OP_WB(13), B(12) => 
                           OP_WB(12), B(11) => OP_WB(11), B(10) => OP_WB(10), 
                           B(9) => OP_WB(9), B(8) => OP_WB(8), B(7) => OP_WB(7)
                           , B(6) => OP_WB(6), B(5) => OP_WB(5), B(4) => 
                           OP_WB(4), B(3) => OP_WB(3), B(2) => OP_WB(2), B(1) 
                           => OP_WB(1), B(0) => OP_WB(0), C(31) => OP_MEM(31), 
                           C(30) => OP_MEM(30), C(29) => OP_MEM(29), C(28) => 
                           OP_MEM(28), C(27) => OP_MEM(27), C(26) => OP_MEM(26)
                           , C(25) => OP_MEM(25), C(24) => OP_MEM(24), C(23) =>
                           OP_MEM(23), C(22) => OP_MEM(22), C(21) => OP_MEM(21)
                           , C(20) => OP_MEM(20), C(19) => OP_MEM(19), C(18) =>
                           OP_MEM(18), C(17) => OP_MEM(17), C(16) => OP_MEM(16)
                           , C(15) => OP_MEM(15), C(14) => OP_MEM(14), C(13) =>
                           OP_MEM(13), C(12) => OP_MEM(12), C(11) => OP_MEM(11)
                           , C(10) => OP_MEM(10), C(9) => OP_MEM(9), C(8) => 
                           OP_MEM(8), C(7) => OP_MEM(7), C(6) => OP_MEM(6), 
                           C(5) => OP_MEM(5), C(4) => OP_MEM(4), C(3) => 
                           OP_MEM(3), C(2) => OP_MEM(2), C(1) => OP_MEM(1), 
                           C(0) => OP_MEM(0), D(31) => n6_port, D(30) => 
                           n6_port, D(29) => n6_port, D(28) => n6_port, D(27) 
                           => n6_port, D(26) => n6_port, D(25) => n6_port, 
                           D(24) => n6_port, D(23) => n6_port, D(22) => n6_port
                           , D(21) => n6_port, D(20) => n6_port, D(19) => 
                           n6_port, D(18) => n6_port, D(17) => n6_port, D(16) 
                           => n6_port, D(15) => n6_port, D(14) => n6_port, 
                           D(13) => n6_port, D(12) => n6_port, D(11) => n6_port
                           , D(10) => n6_port, D(9) => n6_port, D(8) => n6_port
                           , D(7) => n6_port, D(6) => n6_port, D(5) => n6_port,
                           D(4) => n6_port, D(3) => n6_port, D(2) => n6_port, 
                           D(1) => n6_port, D(0) => n6_port, S(1) => 
                           FWDB_1_port, S(0) => FWDB_0_port, Z(31) => 
                           OP2_FW_31_port, Z(30) => OP2_FW_30_port, Z(29) => 
                           OP2_FW_29_port, Z(28) => OP2_FW_28_port, Z(27) => 
                           OP2_FW_27_port, Z(26) => OP2_FW_26_port, Z(25) => 
                           OP2_FW_25_port, Z(24) => OP2_FW_24_port, Z(23) => 
                           OP2_FW_23_port, Z(22) => OP2_FW_22_port, Z(21) => 
                           OP2_FW_21_port, Z(20) => OP2_FW_20_port, Z(19) => 
                           OP2_FW_19_port, Z(18) => OP2_FW_18_port, Z(17) => 
                           OP2_FW_17_port, Z(16) => OP2_FW_16_port, Z(15) => 
                           OP2_FW_15_port, Z(14) => OP2_FW_14_port, Z(13) => 
                           OP2_FW_13_port, Z(12) => OP2_FW_12_port, Z(11) => 
                           OP2_FW_11_port, Z(10) => OP2_FW_10_port, Z(9) => 
                           OP2_FW_9_port, Z(8) => OP2_FW_8_port, Z(7) => 
                           OP2_FW_7_port, Z(6) => OP2_FW_6_port, Z(5) => 
                           OP2_FW_5_port, Z(4) => OP2_FW_4_port, Z(3) => 
                           OP2_FW_3_port, Z(2) => OP2_FW_2_port, Z(1) => 
                           OP2_FW_1_port, Z(0) => OP2_FW_0_port);
   muxA : mux21_NBIT32_3 port map( A(31) => sig_NPC_ABS_31_port, A(30) => 
                           sig_NPC_ABS_30_port, A(29) => sig_NPC_ABS_29_port, 
                           A(28) => sig_NPC_ABS_28_port, A(27) => 
                           sig_NPC_ABS_27_port, A(26) => sig_NPC_ABS_26_port, 
                           A(25) => sig_NPC_ABS_25_port, A(24) => 
                           sig_NPC_ABS_24_port, A(23) => sig_NPC_ABS_23_port, 
                           A(22) => sig_NPC_ABS_22_port, A(21) => 
                           sig_NPC_ABS_21_port, A(20) => sig_NPC_ABS_20_port, 
                           A(19) => sig_NPC_ABS_19_port, A(18) => 
                           sig_NPC_ABS_18_port, A(17) => sig_NPC_ABS_17_port, 
                           A(16) => sig_NPC_ABS_16_port, A(15) => 
                           sig_NPC_ABS_15_port, A(14) => sig_NPC_ABS_14_port, 
                           A(13) => sig_NPC_ABS_13_port, A(12) => 
                           sig_NPC_ABS_12_port, A(11) => sig_NPC_ABS_11_port, 
                           A(10) => sig_NPC_ABS_10_port, A(9) => 
                           sig_NPC_ABS_9_port, A(8) => sig_NPC_ABS_8_port, A(7)
                           => sig_NPC_ABS_7_port, A(6) => sig_NPC_ABS_6_port, 
                           A(5) => sig_NPC_ABS_5_port, A(4) => 
                           sig_NPC_ABS_4_port, A(3) => sig_NPC_ABS_3_port, A(2)
                           => sig_NPC_ABS_2_port, A(1) => sig_NPC_ABS_1_port, 
                           A(0) => sig_NPC_ABS_0_port, B(31) => PC_IN(31), 
                           B(30) => PC_IN(30), B(29) => PC_IN(29), B(28) => 
                           PC_IN(28), B(27) => PC_IN(27), B(26) => PC_IN(26), 
                           B(25) => PC_IN(25), B(24) => PC_IN(24), B(23) => 
                           PC_IN(23), B(22) => PC_IN(22), B(21) => PC_IN(21), 
                           B(20) => PC_IN(20), B(19) => PC_IN(19), B(18) => 
                           PC_IN(18), B(17) => PC_IN(17), B(16) => PC_IN(16), 
                           B(15) => PC_IN(15), B(14) => PC_IN(14), B(13) => 
                           PC_IN(13), B(12) => PC_IN(12), B(11) => PC_IN(11), 
                           B(10) => PC_IN(10), B(9) => PC_IN(9), B(8) => 
                           PC_IN(8), B(7) => PC_IN(7), B(6) => PC_IN(6), B(5) 
                           => PC_IN(5), B(4) => PC_IN(4), B(3) => PC_IN(3), 
                           B(2) => PC_IN(2), B(1) => PC_IN(1), B(0) => PC_IN(0)
                           , S => MUX_A_SEL, Z(31) => sig_OP1_31_port, Z(30) =>
                           sig_OP1_30_port, Z(29) => sig_OP1_29_port, Z(28) => 
                           sig_OP1_28_port, Z(27) => sig_OP1_27_port, Z(26) => 
                           sig_OP1_26_port, Z(25) => sig_OP1_25_port, Z(24) => 
                           sig_OP1_24_port, Z(23) => sig_OP1_23_port, Z(22) => 
                           sig_OP1_22_port, Z(21) => sig_OP1_21_port, Z(20) => 
                           sig_OP1_20_port, Z(19) => sig_OP1_19_port, Z(18) => 
                           sig_OP1_18_port, Z(17) => sig_OP1_17_port, Z(16) => 
                           sig_OP1_16_port, Z(15) => sig_OP1_15_port, Z(14) => 
                           sig_OP1_14_port, Z(13) => sig_OP1_13_port, Z(12) => 
                           sig_OP1_12_port, Z(11) => sig_OP1_11_port, Z(10) => 
                           sig_OP1_10_port, Z(9) => sig_OP1_9_port, Z(8) => 
                           sig_OP1_8_port, Z(7) => sig_OP1_7_port, Z(6) => 
                           sig_OP1_6_port, Z(5) => sig_OP1_5_port, Z(4) => 
                           sig_OP1_4_port, Z(3) => sig_OP1_3_port, Z(2) => 
                           sig_OP1_2_port, Z(1) => sig_OP1_1_port, Z(0) => 
                           sig_OP1_0_port);
   muxB : mux41_NBIT32_3 port map( A(31) => OP2_FW_31_port, A(30) => 
                           OP2_FW_30_port, A(29) => OP2_FW_29_port, A(28) => 
                           OP2_FW_28_port, A(27) => OP2_FW_27_port, A(26) => 
                           OP2_FW_26_port, A(25) => OP2_FW_25_port, A(24) => 
                           OP2_FW_24_port, A(23) => OP2_FW_23_port, A(22) => 
                           OP2_FW_22_port, A(21) => OP2_FW_21_port, A(20) => 
                           OP2_FW_20_port, A(19) => OP2_FW_19_port, A(18) => 
                           OP2_FW_18_port, A(17) => OP2_FW_17_port, A(16) => 
                           OP2_FW_16_port, A(15) => OP2_FW_15_port, A(14) => 
                           OP2_FW_14_port, A(13) => OP2_FW_13_port, A(12) => 
                           OP2_FW_12_port, A(11) => OP2_FW_11_port, A(10) => 
                           OP2_FW_10_port, A(9) => OP2_FW_9_port, A(8) => 
                           OP2_FW_8_port, A(7) => OP2_FW_7_port, A(6) => 
                           OP2_FW_6_port, A(5) => OP2_FW_5_port, A(4) => 
                           OP2_FW_4_port, A(3) => OP2_FW_3_port, A(2) => 
                           OP2_FW_2_port, A(1) => OP2_FW_1_port, A(0) => 
                           OP2_FW_0_port, B(31) => IMM_IN(31), B(30) => 
                           IMM_IN(30), B(29) => IMM_IN(29), B(28) => IMM_IN(28)
                           , B(27) => IMM_IN(27), B(26) => IMM_IN(26), B(25) =>
                           IMM_IN(25), B(24) => IMM_IN(24), B(23) => IMM_IN(23)
                           , B(22) => IMM_IN(22), B(21) => IMM_IN(21), B(20) =>
                           IMM_IN(20), B(19) => IMM_IN(19), B(18) => IMM_IN(18)
                           , B(17) => IMM_IN(17), B(16) => IMM_IN(16), B(15) =>
                           IMM_IN(15), B(14) => IMM_IN(14), B(13) => IMM_IN(13)
                           , B(12) => IMM_IN(12), B(11) => IMM_IN(11), B(10) =>
                           IMM_IN(10), B(9) => IMM_IN(9), B(8) => IMM_IN(8), 
                           B(7) => IMM_IN(7), B(6) => IMM_IN(6), B(5) => 
                           IMM_IN(5), B(4) => IMM_IN(4), B(3) => IMM_IN(3), 
                           B(2) => IMM_IN(2), B(1) => IMM_IN(1), B(0) => 
                           IMM_IN(0), C(31) => n6_port, C(30) => n6_port, C(29)
                           => n6_port, C(28) => n6_port, C(27) => n6_port, 
                           C(26) => n6_port, C(25) => n6_port, C(24) => n6_port
                           , C(23) => n6_port, C(22) => n6_port, C(21) => 
                           n6_port, C(20) => n6_port, C(19) => n6_port, C(18) 
                           => n6_port, C(17) => n6_port, C(16) => n6_port, 
                           C(15) => n6_port, C(14) => n6_port, C(13) => n6_port
                           , C(12) => n6_port, C(11) => n6_port, C(10) => 
                           n6_port, C(9) => n6_port, C(8) => n6_port, C(7) => 
                           n6_port, C(6) => n6_port, C(5) => n6_port, C(4) => 
                           n6_port, C(3) => n6_port, C(2) => n7_port, C(1) => 
                           n6_port, C(0) => n6_port, D(31) => n6_port, D(30) =>
                           n6_port, D(29) => n6_port, D(28) => n6_port, D(27) 
                           => n6_port, D(26) => n6_port, D(25) => n6_port, 
                           D(24) => n6_port, D(23) => n6_port, D(22) => n6_port
                           , D(21) => n6_port, D(20) => n6_port, D(19) => 
                           n6_port, D(18) => n6_port, D(17) => n6_port, D(16) 
                           => n6_port, D(15) => n6_port, D(14) => n6_port, 
                           D(13) => n6_port, D(12) => n6_port, D(11) => n6_port
                           , D(10) => n6_port, D(9) => n6_port, D(8) => n6_port
                           , D(7) => n6_port, D(6) => n6_port, D(5) => n6_port,
                           D(4) => n6_port, D(3) => n6_port, D(2) => n6_port, 
                           D(1) => n6_port, D(0) => n6_port, S(1) => 
                           MUX_B_SEL(1), S(0) => MUX_B_SEL(0), Z(31) => 
                           sig_OP2_31_port, Z(30) => sig_OP2_30_port, Z(29) => 
                           sig_OP2_29_port, Z(28) => sig_OP2_28_port, Z(27) => 
                           sig_OP2_27_port, Z(26) => sig_OP2_26_port, Z(25) => 
                           sig_OP2_25_port, Z(24) => sig_OP2_24_port, Z(23) => 
                           sig_OP2_23_port, Z(22) => sig_OP2_22_port, Z(21) => 
                           sig_OP2_21_port, Z(20) => sig_OP2_20_port, Z(19) => 
                           sig_OP2_19_port, Z(18) => sig_OP2_18_port, Z(17) => 
                           sig_OP2_17_port, Z(16) => sig_OP2_16_port, Z(15) => 
                           sig_OP2_15_port, Z(14) => sig_OP2_14_port, Z(13) => 
                           sig_OP2_13_port, Z(12) => sig_OP2_12_port, Z(11) => 
                           sig_OP2_11_port, Z(10) => sig_OP2_10_port, Z(9) => 
                           sig_OP2_9_port, Z(8) => sig_OP2_8_port, Z(7) => 
                           sig_OP2_7_port, Z(6) => sig_OP2_6_port, Z(5) => 
                           sig_OP2_5_port, Z(4) => sig_OP2_4_port, Z(3) => 
                           sig_OP2_3_port, Z(2) => sig_OP2_2_port, Z(1) => 
                           sig_OP2_1_port, Z(0) => sig_OP2_0_port);
   alu0 : ALU_NBIT32 port map( OP1(31) => sig_OP1_31_port, OP1(30) => 
                           sig_OP1_30_port, OP1(29) => sig_OP1_29_port, OP1(28)
                           => sig_OP1_28_port, OP1(27) => sig_OP1_27_port, 
                           OP1(26) => sig_OP1_26_port, OP1(25) => 
                           sig_OP1_25_port, OP1(24) => sig_OP1_24_port, OP1(23)
                           => sig_OP1_23_port, OP1(22) => sig_OP1_22_port, 
                           OP1(21) => sig_OP1_21_port, OP1(20) => 
                           sig_OP1_20_port, OP1(19) => sig_OP1_19_port, OP1(18)
                           => sig_OP1_18_port, OP1(17) => sig_OP1_17_port, 
                           OP1(16) => sig_OP1_16_port, OP1(15) => 
                           sig_OP1_15_port, OP1(14) => sig_OP1_14_port, OP1(13)
                           => sig_OP1_13_port, OP1(12) => sig_OP1_12_port, 
                           OP1(11) => sig_OP1_11_port, OP1(10) => 
                           sig_OP1_10_port, OP1(9) => sig_OP1_9_port, OP1(8) =>
                           sig_OP1_8_port, OP1(7) => sig_OP1_7_port, OP1(6) => 
                           sig_OP1_6_port, OP1(5) => sig_OP1_5_port, OP1(4) => 
                           sig_OP1_4_port, OP1(3) => sig_OP1_3_port, OP1(2) => 
                           sig_OP1_2_port, OP1(1) => sig_OP1_1_port, OP1(0) => 
                           sig_OP1_0_port, OP2(31) => sig_OP2_31_port, OP2(30) 
                           => sig_OP2_30_port, OP2(29) => sig_OP2_29_port, 
                           OP2(28) => sig_OP2_28_port, OP2(27) => 
                           sig_OP2_27_port, OP2(26) => sig_OP2_26_port, OP2(25)
                           => sig_OP2_25_port, OP2(24) => sig_OP2_24_port, 
                           OP2(23) => sig_OP2_23_port, OP2(22) => 
                           sig_OP2_22_port, OP2(21) => sig_OP2_21_port, OP2(20)
                           => sig_OP2_20_port, OP2(19) => sig_OP2_19_port, 
                           OP2(18) => sig_OP2_18_port, OP2(17) => 
                           sig_OP2_17_port, OP2(16) => sig_OP2_16_port, OP2(15)
                           => sig_OP2_15_port, OP2(14) => sig_OP2_14_port, 
                           OP2(13) => sig_OP2_13_port, OP2(12) => 
                           sig_OP2_12_port, OP2(11) => sig_OP2_11_port, OP2(10)
                           => sig_OP2_10_port, OP2(9) => sig_OP2_9_port, OP2(8)
                           => sig_OP2_8_port, OP2(7) => sig_OP2_7_port, OP2(6) 
                           => sig_OP2_6_port, OP2(5) => sig_OP2_5_port, OP2(4) 
                           => sig_OP2_4_port, OP2(3) => sig_OP2_3_port, OP2(2) 
                           => sig_OP2_2_port, OP2(1) => sig_OP2_1_port, OP2(0) 
                           => sig_OP2_0_port, ALU_OPC(0) => ALU_OPC(0), 
                           ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => ALU_OPC(2), 
                           ALU_OPC(3) => ALU_OPC(3), ALU_RES(31) => 
                           sig_ALU_RES_31_port, ALU_RES(30) => 
                           sig_ALU_RES_30_port, ALU_RES(29) => 
                           sig_ALU_RES_29_port, ALU_RES(28) => 
                           sig_ALU_RES_28_port, ALU_RES(27) => 
                           sig_ALU_RES_27_port, ALU_RES(26) => 
                           sig_ALU_RES_26_port, ALU_RES(25) => 
                           sig_ALU_RES_25_port, ALU_RES(24) => 
                           sig_ALU_RES_24_port, ALU_RES(23) => 
                           sig_ALU_RES_23_port, ALU_RES(22) => 
                           sig_ALU_RES_22_port, ALU_RES(21) => 
                           sig_ALU_RES_21_port, ALU_RES(20) => 
                           sig_ALU_RES_20_port, ALU_RES(19) => 
                           sig_ALU_RES_19_port, ALU_RES(18) => 
                           sig_ALU_RES_18_port, ALU_RES(17) => 
                           sig_ALU_RES_17_port, ALU_RES(16) => 
                           sig_ALU_RES_16_port, ALU_RES(15) => 
                           sig_ALU_RES_15_port, ALU_RES(14) => 
                           sig_ALU_RES_14_port, ALU_RES(13) => 
                           sig_ALU_RES_13_port, ALU_RES(12) => 
                           sig_ALU_RES_12_port, ALU_RES(11) => 
                           sig_ALU_RES_11_port, ALU_RES(10) => 
                           sig_ALU_RES_10_port, ALU_RES(9) => 
                           sig_ALU_RES_9_port, ALU_RES(8) => sig_ALU_RES_8_port
                           , ALU_RES(7) => sig_ALU_RES_7_port, ALU_RES(6) => 
                           sig_ALU_RES_6_port, ALU_RES(5) => sig_ALU_RES_5_port
                           , ALU_RES(4) => sig_ALU_RES_4_port, ALU_RES(3) => 
                           sig_ALU_RES_3_port, ALU_RES(2) => sig_ALU_RES_2_port
                           , ALU_RES(1) => sig_ALU_RES_1_port, ALU_RES(0) => 
                           sig_ALU_RES_0_port);
   alureg : regn_N32_6 port map( DIN(31) => sig_ALU_RES_31_port, DIN(30) => 
                           sig_ALU_RES_30_port, DIN(29) => sig_ALU_RES_29_port,
                           DIN(28) => sig_ALU_RES_28_port, DIN(27) => 
                           sig_ALU_RES_27_port, DIN(26) => sig_ALU_RES_26_port,
                           DIN(25) => sig_ALU_RES_25_port, DIN(24) => 
                           sig_ALU_RES_24_port, DIN(23) => sig_ALU_RES_23_port,
                           DIN(22) => sig_ALU_RES_22_port, DIN(21) => 
                           sig_ALU_RES_21_port, DIN(20) => sig_ALU_RES_20_port,
                           DIN(19) => sig_ALU_RES_19_port, DIN(18) => 
                           sig_ALU_RES_18_port, DIN(17) => sig_ALU_RES_17_port,
                           DIN(16) => sig_ALU_RES_16_port, DIN(15) => 
                           sig_ALU_RES_15_port, DIN(14) => sig_ALU_RES_14_port,
                           DIN(13) => sig_ALU_RES_13_port, DIN(12) => 
                           sig_ALU_RES_12_port, DIN(11) => sig_ALU_RES_11_port,
                           DIN(10) => sig_ALU_RES_10_port, DIN(9) => 
                           sig_ALU_RES_9_port, DIN(8) => sig_ALU_RES_8_port, 
                           DIN(7) => sig_ALU_RES_7_port, DIN(6) => 
                           sig_ALU_RES_6_port, DIN(5) => sig_ALU_RES_5_port, 
                           DIN(4) => sig_ALU_RES_4_port, DIN(3) => 
                           sig_ALU_RES_3_port, DIN(2) => sig_ALU_RES_2_port, 
                           DIN(1) => sig_ALU_RES_1_port, DIN(0) => 
                           sig_ALU_RES_0_port, CLK => CLK, EN => ALU_OUTREG_EN,
                           RST => RST, DOUT(31) => ALU_RES(31), DOUT(30) => 
                           ALU_RES(30), DOUT(29) => ALU_RES(29), DOUT(28) => 
                           ALU_RES(28), DOUT(27) => ALU_RES(27), DOUT(26) => 
                           ALU_RES(26), DOUT(25) => ALU_RES(25), DOUT(24) => 
                           ALU_RES(24), DOUT(23) => ALU_RES(23), DOUT(22) => 
                           ALU_RES(22), DOUT(21) => ALU_RES(21), DOUT(20) => 
                           ALU_RES(20), DOUT(19) => ALU_RES(19), DOUT(18) => 
                           ALU_RES(18), DOUT(17) => ALU_RES(17), DOUT(16) => 
                           ALU_RES(16), DOUT(15) => ALU_RES(15), DOUT(14) => 
                           ALU_RES(14), DOUT(13) => ALU_RES(13), DOUT(12) => 
                           ALU_RES(12), DOUT(11) => ALU_RES(11), DOUT(10) => 
                           ALU_RES(10), DOUT(9) => ALU_RES(9), DOUT(8) => 
                           ALU_RES(8), DOUT(7) => ALU_RES(7), DOUT(6) => 
                           ALU_RES(6), DOUT(5) => ALU_RES(5), DOUT(4) => 
                           ALU_RES(4), DOUT(3) => ALU_RES(3), DOUT(2) => 
                           ALU_RES(2), DOUT(1) => ALU_RES(1), DOUT(0) => 
                           ALU_RES(0));
   B_reg : regn_N32_5 port map( DIN(31) => OP2_FW_31_port, DIN(30) => 
                           OP2_FW_30_port, DIN(29) => OP2_FW_29_port, DIN(28) 
                           => OP2_FW_28_port, DIN(27) => OP2_FW_27_port, 
                           DIN(26) => OP2_FW_26_port, DIN(25) => OP2_FW_25_port
                           , DIN(24) => OP2_FW_24_port, DIN(23) => 
                           OP2_FW_23_port, DIN(22) => OP2_FW_22_port, DIN(21) 
                           => OP2_FW_21_port, DIN(20) => OP2_FW_20_port, 
                           DIN(19) => OP2_FW_19_port, DIN(18) => OP2_FW_18_port
                           , DIN(17) => OP2_FW_17_port, DIN(16) => 
                           OP2_FW_16_port, DIN(15) => OP2_FW_15_port, DIN(14) 
                           => OP2_FW_14_port, DIN(13) => OP2_FW_13_port, 
                           DIN(12) => OP2_FW_12_port, DIN(11) => OP2_FW_11_port
                           , DIN(10) => OP2_FW_10_port, DIN(9) => OP2_FW_9_port
                           , DIN(8) => OP2_FW_8_port, DIN(7) => OP2_FW_7_port, 
                           DIN(6) => OP2_FW_6_port, DIN(5) => OP2_FW_5_port, 
                           DIN(4) => OP2_FW_4_port, DIN(3) => OP2_FW_3_port, 
                           DIN(2) => OP2_FW_2_port, DIN(1) => OP2_FW_1_port, 
                           DIN(0) => OP2_FW_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => B_OUT(31), 
                           DOUT(30) => B_OUT(30), DOUT(29) => B_OUT(29), 
                           DOUT(28) => B_OUT(28), DOUT(27) => B_OUT(27), 
                           DOUT(26) => B_OUT(26), DOUT(25) => B_OUT(25), 
                           DOUT(24) => B_OUT(24), DOUT(23) => B_OUT(23), 
                           DOUT(22) => B_OUT(22), DOUT(21) => B_OUT(21), 
                           DOUT(20) => B_OUT(20), DOUT(19) => B_OUT(19), 
                           DOUT(18) => B_OUT(18), DOUT(17) => B_OUT(17), 
                           DOUT(16) => B_OUT(16), DOUT(15) => B_OUT(15), 
                           DOUT(14) => B_OUT(14), DOUT(13) => B_OUT(13), 
                           DOUT(12) => B_OUT(12), DOUT(11) => B_OUT(11), 
                           DOUT(10) => B_OUT(10), DOUT(9) => B_OUT(9), DOUT(8) 
                           => B_OUT(8), DOUT(7) => B_OUT(7), DOUT(6) => 
                           B_OUT(6), DOUT(5) => B_OUT(5), DOUT(4) => B_OUT(4), 
                           DOUT(3) => B_OUT(3), DOUT(2) => B_OUT(2), DOUT(1) =>
                           B_OUT(1), DOUT(0) => B_OUT(0));
   ADD_WR_reg : regn_N5_2 port map( DIN(4) => ADD_WR_IN(4), DIN(3) => 
                           ADD_WR_IN(3), DIN(2) => ADD_WR_IN(2), DIN(1) => 
                           ADD_WR_IN(1), DIN(0) => ADD_WR_IN(0), CLK => CLK, EN
                           => ALU_OUTREG_EN, RST => RST, DOUT(4) => 
                           ADD_WR_OUT(4), DOUT(3) => ADD_WR_OUT(3), DOUT(2) => 
                           ADD_WR_OUT(2), DOUT(1) => ADD_WR_OUT(1), DOUT(0) => 
                           ADD_WR_OUT(0));
   NPC_ABS_reg : regn_N32_4 port map( DIN(31) => sig_NPC_ABS_31_port, DIN(30) 
                           => sig_NPC_ABS_30_port, DIN(29) => 
                           sig_NPC_ABS_29_port, DIN(28) => sig_NPC_ABS_28_port,
                           DIN(27) => sig_NPC_ABS_27_port, DIN(26) => 
                           sig_NPC_ABS_26_port, DIN(25) => sig_NPC_ABS_25_port,
                           DIN(24) => sig_NPC_ABS_24_port, DIN(23) => 
                           sig_NPC_ABS_23_port, DIN(22) => sig_NPC_ABS_22_port,
                           DIN(21) => sig_NPC_ABS_21_port, DIN(20) => 
                           sig_NPC_ABS_20_port, DIN(19) => sig_NPC_ABS_19_port,
                           DIN(18) => sig_NPC_ABS_18_port, DIN(17) => 
                           sig_NPC_ABS_17_port, DIN(16) => sig_NPC_ABS_16_port,
                           DIN(15) => sig_NPC_ABS_15_port, DIN(14) => 
                           sig_NPC_ABS_14_port, DIN(13) => sig_NPC_ABS_13_port,
                           DIN(12) => sig_NPC_ABS_12_port, DIN(11) => 
                           sig_NPC_ABS_11_port, DIN(10) => sig_NPC_ABS_10_port,
                           DIN(9) => sig_NPC_ABS_9_port, DIN(8) => 
                           sig_NPC_ABS_8_port, DIN(7) => sig_NPC_ABS_7_port, 
                           DIN(6) => sig_NPC_ABS_6_port, DIN(5) => 
                           sig_NPC_ABS_5_port, DIN(4) => sig_NPC_ABS_4_port, 
                           DIN(3) => sig_NPC_ABS_3_port, DIN(2) => 
                           sig_NPC_ABS_2_port, DIN(1) => sig_NPC_ABS_1_port, 
                           DIN(0) => sig_NPC_ABS_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => NPC_ABS(31), 
                           DOUT(30) => NPC_ABS(30), DOUT(29) => NPC_ABS(29), 
                           DOUT(28) => NPC_ABS(28), DOUT(27) => NPC_ABS(27), 
                           DOUT(26) => NPC_ABS(26), DOUT(25) => NPC_ABS(25), 
                           DOUT(24) => NPC_ABS(24), DOUT(23) => NPC_ABS(23), 
                           DOUT(22) => NPC_ABS(22), DOUT(21) => NPC_ABS(21), 
                           DOUT(20) => NPC_ABS(20), DOUT(19) => NPC_ABS(19), 
                           DOUT(18) => NPC_ABS(18), DOUT(17) => NPC_ABS(17), 
                           DOUT(16) => NPC_ABS(16), DOUT(15) => NPC_ABS(15), 
                           DOUT(14) => NPC_ABS(14), DOUT(13) => NPC_ABS(13), 
                           DOUT(12) => NPC_ABS(12), DOUT(11) => NPC_ABS(11), 
                           DOUT(10) => NPC_ABS(10), DOUT(9) => NPC_ABS(9), 
                           DOUT(8) => NPC_ABS(8), DOUT(7) => NPC_ABS(7), 
                           DOUT(6) => NPC_ABS(6), DOUT(5) => NPC_ABS(5), 
                           DOUT(4) => NPC_ABS(4), DOUT(3) => NPC_ABS(3), 
                           DOUT(2) => NPC_ABS(2), DOUT(1) => NPC_ABS(1), 
                           DOUT(0) => NPC_ABS(0));
   NPC_REL_reg : regn_N32_3 port map( DIN(31) => sig_NPC_REL_31_port, DIN(30) 
                           => sig_NPC_REL_30_port, DIN(29) => 
                           sig_NPC_REL_29_port, DIN(28) => sig_NPC_REL_28_port,
                           DIN(27) => sig_NPC_REL_27_port, DIN(26) => 
                           sig_NPC_REL_26_port, DIN(25) => sig_NPC_REL_25_port,
                           DIN(24) => sig_NPC_REL_24_port, DIN(23) => 
                           sig_NPC_REL_23_port, DIN(22) => sig_NPC_REL_22_port,
                           DIN(21) => sig_NPC_REL_21_port, DIN(20) => 
                           sig_NPC_REL_20_port, DIN(19) => sig_NPC_REL_19_port,
                           DIN(18) => sig_NPC_REL_18_port, DIN(17) => 
                           sig_NPC_REL_17_port, DIN(16) => sig_NPC_REL_16_port,
                           DIN(15) => sig_NPC_REL_15_port, DIN(14) => 
                           sig_NPC_REL_14_port, DIN(13) => sig_NPC_REL_13_port,
                           DIN(12) => sig_NPC_REL_12_port, DIN(11) => 
                           sig_NPC_REL_11_port, DIN(10) => sig_NPC_REL_10_port,
                           DIN(9) => sig_NPC_REL_9_port, DIN(8) => 
                           sig_NPC_REL_8_port, DIN(7) => sig_NPC_REL_7_port, 
                           DIN(6) => sig_NPC_REL_6_port, DIN(5) => 
                           sig_NPC_REL_5_port, DIN(4) => sig_NPC_REL_4_port, 
                           DIN(3) => sig_NPC_REL_3_port, DIN(2) => 
                           sig_NPC_REL_2_port, DIN(1) => sig_NPC_REL_1_port, 
                           DIN(0) => sig_NPC_REL_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => NPC_REL(31), 
                           DOUT(30) => NPC_REL(30), DOUT(29) => NPC_REL(29), 
                           DOUT(28) => NPC_REL(28), DOUT(27) => NPC_REL(27), 
                           DOUT(26) => NPC_REL(26), DOUT(25) => NPC_REL(25), 
                           DOUT(24) => NPC_REL(24), DOUT(23) => NPC_REL(23), 
                           DOUT(22) => NPC_REL(22), DOUT(21) => NPC_REL(21), 
                           DOUT(20) => NPC_REL(20), DOUT(19) => NPC_REL(19), 
                           DOUT(18) => NPC_REL(18), DOUT(17) => NPC_REL(17), 
                           DOUT(16) => NPC_REL(16), DOUT(15) => NPC_REL(15), 
                           DOUT(14) => NPC_REL(14), DOUT(13) => NPC_REL(13), 
                           DOUT(12) => NPC_REL(12), DOUT(11) => NPC_REL(11), 
                           DOUT(10) => NPC_REL(10), DOUT(9) => NPC_REL(9), 
                           DOUT(8) => NPC_REL(8), DOUT(7) => NPC_REL(7), 
                           DOUT(6) => NPC_REL(6), DOUT(5) => NPC_REL(5), 
                           DOUT(4) => NPC_REL(4), DOUT(3) => NPC_REL(3), 
                           DOUT(2) => NPC_REL(2), DOUT(1) => NPC_REL(1), 
                           DOUT(0) => NPC_REL(0));
   add_1_root_add_0_root_add_118_2 : Execute_DW01_add_1 port map( A(31) => 
                           n2_port, A(30) => n2_port, A(29) => n2_port, A(28) 
                           => n2_port, A(27) => n2_port, A(26) => n2_port, 
                           A(25) => n2_port, A(24) => n2_port, A(23) => n2_port
                           , A(22) => n2_port, A(21) => n2_port, A(20) => 
                           n2_port, A(19) => n2_port, A(18) => n2_port, A(17) 
                           => n2_port, A(16) => n2_port, A(15) => n2_port, 
                           A(14) => n2_port, A(13) => n2_port, A(12) => n2_port
                           , A(11) => n2_port, A(10) => n2_port, A(9) => 
                           n2_port, A(8) => n2_port, A(7) => n2_port, A(6) => 
                           n2_port, A(5) => n2_port, A(4) => n2_port, A(3) => 
                           n2_port, A(2) => n3_port, A(1) => n2_port, A(0) => 
                           n2_port, B(31) => IMM_IN(31), B(30) => IMM_IN(30), 
                           B(29) => IMM_IN(29), B(28) => IMM_IN(28), B(27) => 
                           IMM_IN(27), B(26) => IMM_IN(26), B(25) => IMM_IN(25)
                           , B(24) => IMM_IN(24), B(23) => IMM_IN(23), B(22) =>
                           IMM_IN(22), B(21) => IMM_IN(21), B(20) => IMM_IN(20)
                           , B(19) => IMM_IN(19), B(18) => IMM_IN(18), B(17) =>
                           IMM_IN(17), B(16) => IMM_IN(16), B(15) => IMM_IN(15)
                           , B(14) => IMM_IN(14), B(13) => IMM_IN(13), B(12) =>
                           IMM_IN(12), B(11) => IMM_IN(11), B(10) => IMM_IN(10)
                           , B(9) => IMM_IN(9), B(8) => IMM_IN(8), B(7) => 
                           IMM_IN(7), B(6) => IMM_IN(6), B(5) => IMM_IN(5), 
                           B(4) => IMM_IN(4), B(3) => IMM_IN(3), B(2) => 
                           IMM_IN(2), B(1) => IMM_IN(1), B(0) => IMM_IN(0), CI 
                           => n4_port, SUM(31) => N31, SUM(30) => N30, SUM(29) 
                           => N29, SUM(28) => N28, SUM(27) => N27, SUM(26) => 
                           N26, SUM(25) => N25, SUM(24) => N24, SUM(23) => N23,
                           SUM(22) => N22, SUM(21) => N21, SUM(20) => N20, 
                           SUM(19) => N19, SUM(18) => N18, SUM(17) => N17, 
                           SUM(16) => N16, SUM(15) => N15, SUM(14) => N14, 
                           SUM(13) => N13, SUM(12) => N12, SUM(11) => N11, 
                           SUM(10) => N10, SUM(9) => N9, SUM(8) => N8, SUM(7) 
                           => N7, SUM(6) => N6, SUM(5) => N5, SUM(4) => N4, 
                           SUM(3) => N3, SUM(2) => N2, SUM(1) => N1, SUM(0) => 
                           N0, CO => n_1826);
   add_0_root_add_0_root_add_118_2 : Execute_DW01_add_0 port map( A(31) => 
                           PC_IN(31), A(30) => PC_IN(30), A(29) => PC_IN(29), 
                           A(28) => PC_IN(28), A(27) => PC_IN(27), A(26) => 
                           PC_IN(26), A(25) => PC_IN(25), A(24) => PC_IN(24), 
                           A(23) => PC_IN(23), A(22) => PC_IN(22), A(21) => 
                           PC_IN(21), A(20) => PC_IN(20), A(19) => PC_IN(19), 
                           A(18) => PC_IN(18), A(17) => PC_IN(17), A(16) => 
                           PC_IN(16), A(15) => PC_IN(15), A(14) => PC_IN(14), 
                           A(13) => PC_IN(13), A(12) => PC_IN(12), A(11) => 
                           PC_IN(11), A(10) => PC_IN(10), A(9) => PC_IN(9), 
                           A(8) => PC_IN(8), A(7) => PC_IN(7), A(6) => PC_IN(6)
                           , A(5) => PC_IN(5), A(4) => PC_IN(4), A(3) => 
                           PC_IN(3), A(2) => PC_IN(2), A(1) => PC_IN(1), A(0) 
                           => PC_IN(0), B(31) => N31, B(30) => N30, B(29) => 
                           N29, B(28) => N28, B(27) => N27, B(26) => N26, B(25)
                           => N25, B(24) => N24, B(23) => N23, B(22) => N22, 
                           B(21) => N21, B(20) => N20, B(19) => N19, B(18) => 
                           N18, B(17) => N17, B(16) => N16, B(15) => N15, B(14)
                           => N14, B(13) => N13, B(12) => N12, B(11) => N11, 
                           B(10) => N10, B(9) => N9, B(8) => N8, B(7) => N7, 
                           B(6) => N6, B(5) => N5, B(4) => N4, B(3) => N3, B(2)
                           => N2, B(1) => N1, B(0) => N0, CI => n5_port, 
                           SUM(31) => sig_NPC_REL_31_port, SUM(30) => 
                           sig_NPC_REL_30_port, SUM(29) => sig_NPC_REL_29_port,
                           SUM(28) => sig_NPC_REL_28_port, SUM(27) => 
                           sig_NPC_REL_27_port, SUM(26) => sig_NPC_REL_26_port,
                           SUM(25) => sig_NPC_REL_25_port, SUM(24) => 
                           sig_NPC_REL_24_port, SUM(23) => sig_NPC_REL_23_port,
                           SUM(22) => sig_NPC_REL_22_port, SUM(21) => 
                           sig_NPC_REL_21_port, SUM(20) => sig_NPC_REL_20_port,
                           SUM(19) => sig_NPC_REL_19_port, SUM(18) => 
                           sig_NPC_REL_18_port, SUM(17) => sig_NPC_REL_17_port,
                           SUM(16) => sig_NPC_REL_16_port, SUM(15) => 
                           sig_NPC_REL_15_port, SUM(14) => sig_NPC_REL_14_port,
                           SUM(13) => sig_NPC_REL_13_port, SUM(12) => 
                           sig_NPC_REL_12_port, SUM(11) => sig_NPC_REL_11_port,
                           SUM(10) => sig_NPC_REL_10_port, SUM(9) => 
                           sig_NPC_REL_9_port, SUM(8) => sig_NPC_REL_8_port, 
                           SUM(7) => sig_NPC_REL_7_port, SUM(6) => 
                           sig_NPC_REL_6_port, SUM(5) => sig_NPC_REL_5_port, 
                           SUM(4) => sig_NPC_REL_4_port, SUM(3) => 
                           sig_NPC_REL_3_port, SUM(2) => sig_NPC_REL_2_port, 
                           SUM(1) => sig_NPC_REL_1_port, SUM(0) => 
                           sig_NPC_REL_0_port, CO => n_1827);
   U3 : NOR2_X1 port map( A1 => ZERO_FLAG_port, A2 => n1_port, ZN => sig_RST);
   U4 : INV_X1 port map( A => RST, ZN => n1_port);
   n2_port <= '0';
   n3_port <= '1';
   n4_port <= '0';
   n5_port <= '0';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Decode is

   port( CLK, RST, REG_LATCH_EN, RD1, RD2, RF_WE, ZERO_FLAG : in std_logic;  
         PC_IN, INS_IN : in std_logic_vector (31 downto 0);  ADD_WR : in 
         std_logic_vector (4 downto 0);  DATA_WR_IN : in std_logic_vector (31 
         downto 0);  PC_OUT, A_OUT, B_OUT, IMM_OUT : out std_logic_vector (31 
         downto 0);  ADD_RS1_HDU, ADD_RS2_HDU, ADD_WR_OUT, ADD_RS1_OUT, 
         ADD_RS2_OUT : out std_logic_vector (4 downto 0));

end Decode;

architecture SYN_struct of Decode is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component register_file_NBIT_ADD5_NBIT_DATA32
      port( CLK, RST, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RS1, 
            ADD_RS2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component regn_N5_3
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N5_4
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N5_0
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N32_7
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_8
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component instruction_decomposition
      port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype :
            in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : out std_logic_vector (4 
            downto 0);  IMM : out std_logic_vector (31 downto 0));
   end component;
   
   component instruction_type
      port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype :
            out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic1_port, ADD_RS1_HDU_4_port, ADD_RS1_HDU_3_port, 
      ADD_RS1_HDU_2_port, ADD_RS1_HDU_1_port, ADD_RS1_HDU_0_port, 
      ADD_RS2_HDU_4_port, ADD_RS2_HDU_3_port, ADD_RS2_HDU_2_port, 
      ADD_RS2_HDU_1_port, ADD_RS2_HDU_0_port, sig_RST, sig_Rtype, sig_Itype, 
      sig_Jtype, sig_ADD_WR_4_port, sig_ADD_WR_3_port, sig_ADD_WR_2_port, 
      sig_ADD_WR_1_port, sig_ADD_WR_0_port, sig_IMM_31_port, sig_IMM_30_port, 
      sig_IMM_29_port, sig_IMM_28_port, sig_IMM_27_port, sig_IMM_26_port, 
      sig_IMM_25_port, sig_IMM_24_port, sig_IMM_23_port, sig_IMM_22_port, 
      sig_IMM_21_port, sig_IMM_20_port, sig_IMM_19_port, sig_IMM_18_port, 
      sig_IMM_17_port, sig_IMM_16_port, sig_IMM_15_port, sig_IMM_14_port, 
      sig_IMM_13_port, sig_IMM_12_port, sig_IMM_11_port, sig_IMM_10_port, 
      sig_IMM_9_port, sig_IMM_8_port, sig_IMM_7_port, sig_IMM_6_port, 
      sig_IMM_5_port, sig_IMM_4_port, sig_IMM_3_port, sig_IMM_2_port, 
      sig_IMM_1_port, sig_IMM_0_port, n1 : std_logic;

begin
   ADD_RS1_HDU <= ( ADD_RS1_HDU_4_port, ADD_RS1_HDU_3_port, ADD_RS1_HDU_2_port,
      ADD_RS1_HDU_1_port, ADD_RS1_HDU_0_port );
   ADD_RS2_HDU <= ( ADD_RS2_HDU_4_port, ADD_RS2_HDU_3_port, ADD_RS2_HDU_2_port,
      ADD_RS2_HDU_1_port, ADD_RS2_HDU_0_port );
   
   X_Logic1_port <= '1';
   U2 : NOR2_X2 port map( A1 => ZERO_FLAG, A2 => n1, ZN => sig_RST);
   ins_type : instruction_type port map( INST_IN(31) => INS_IN(31), INST_IN(30)
                           => INS_IN(30), INST_IN(29) => INS_IN(29), 
                           INST_IN(28) => INS_IN(28), INST_IN(27) => INS_IN(27)
                           , INST_IN(26) => INS_IN(26), INST_IN(25) => 
                           INS_IN(25), INST_IN(24) => INS_IN(24), INST_IN(23) 
                           => INS_IN(23), INST_IN(22) => INS_IN(22), 
                           INST_IN(21) => INS_IN(21), INST_IN(20) => INS_IN(20)
                           , INST_IN(19) => INS_IN(19), INST_IN(18) => 
                           INS_IN(18), INST_IN(17) => INS_IN(17), INST_IN(16) 
                           => INS_IN(16), INST_IN(15) => INS_IN(15), 
                           INST_IN(14) => INS_IN(14), INST_IN(13) => INS_IN(13)
                           , INST_IN(12) => INS_IN(12), INST_IN(11) => 
                           INS_IN(11), INST_IN(10) => INS_IN(10), INST_IN(9) =>
                           INS_IN(9), INST_IN(8) => INS_IN(8), INST_IN(7) => 
                           INS_IN(7), INST_IN(6) => INS_IN(6), INST_IN(5) => 
                           INS_IN(5), INST_IN(4) => INS_IN(4), INST_IN(3) => 
                           INS_IN(3), INST_IN(2) => INS_IN(2), INST_IN(1) => 
                           INS_IN(1), INST_IN(0) => INS_IN(0), Rtype => 
                           sig_Rtype, Itype => sig_Itype, Jtype => sig_Jtype);
   ins_dec : instruction_decomposition port map( INST_IN(31) => INS_IN(31), 
                           INST_IN(30) => INS_IN(30), INST_IN(29) => INS_IN(29)
                           , INST_IN(28) => INS_IN(28), INST_IN(27) => 
                           INS_IN(27), INST_IN(26) => INS_IN(26), INST_IN(25) 
                           => INS_IN(25), INST_IN(24) => INS_IN(24), 
                           INST_IN(23) => INS_IN(23), INST_IN(22) => INS_IN(22)
                           , INST_IN(21) => INS_IN(21), INST_IN(20) => 
                           INS_IN(20), INST_IN(19) => INS_IN(19), INST_IN(18) 
                           => INS_IN(18), INST_IN(17) => INS_IN(17), 
                           INST_IN(16) => INS_IN(16), INST_IN(15) => INS_IN(15)
                           , INST_IN(14) => INS_IN(14), INST_IN(13) => 
                           INS_IN(13), INST_IN(12) => INS_IN(12), INST_IN(11) 
                           => INS_IN(11), INST_IN(10) => INS_IN(10), INST_IN(9)
                           => INS_IN(9), INST_IN(8) => INS_IN(8), INST_IN(7) =>
                           INS_IN(7), INST_IN(6) => INS_IN(6), INST_IN(5) => 
                           INS_IN(5), INST_IN(4) => INS_IN(4), INST_IN(3) => 
                           INS_IN(3), INST_IN(2) => INS_IN(2), INST_IN(1) => 
                           INS_IN(1), INST_IN(0) => INS_IN(0), Rtype => 
                           sig_Rtype, Itype => sig_Itype, Jtype => sig_Jtype, 
                           ADD_RS1(4) => ADD_RS1_HDU_4_port, ADD_RS1(3) => 
                           ADD_RS1_HDU_3_port, ADD_RS1(2) => ADD_RS1_HDU_2_port
                           , ADD_RS1(1) => ADD_RS1_HDU_1_port, ADD_RS1(0) => 
                           ADD_RS1_HDU_0_port, ADD_RS2(4) => ADD_RS2_HDU_4_port
                           , ADD_RS2(3) => ADD_RS2_HDU_3_port, ADD_RS2(2) => 
                           ADD_RS2_HDU_2_port, ADD_RS2(1) => ADD_RS2_HDU_1_port
                           , ADD_RS2(0) => ADD_RS2_HDU_0_port, ADD_WR(4) => 
                           sig_ADD_WR_4_port, ADD_WR(3) => sig_ADD_WR_3_port, 
                           ADD_WR(2) => sig_ADD_WR_2_port, ADD_WR(1) => 
                           sig_ADD_WR_1_port, ADD_WR(0) => sig_ADD_WR_0_port, 
                           IMM(31) => sig_IMM_31_port, IMM(30) => 
                           sig_IMM_30_port, IMM(29) => sig_IMM_29_port, IMM(28)
                           => sig_IMM_28_port, IMM(27) => sig_IMM_27_port, 
                           IMM(26) => sig_IMM_26_port, IMM(25) => 
                           sig_IMM_25_port, IMM(24) => sig_IMM_24_port, IMM(23)
                           => sig_IMM_23_port, IMM(22) => sig_IMM_22_port, 
                           IMM(21) => sig_IMM_21_port, IMM(20) => 
                           sig_IMM_20_port, IMM(19) => sig_IMM_19_port, IMM(18)
                           => sig_IMM_18_port, IMM(17) => sig_IMM_17_port, 
                           IMM(16) => sig_IMM_16_port, IMM(15) => 
                           sig_IMM_15_port, IMM(14) => sig_IMM_14_port, IMM(13)
                           => sig_IMM_13_port, IMM(12) => sig_IMM_12_port, 
                           IMM(11) => sig_IMM_11_port, IMM(10) => 
                           sig_IMM_10_port, IMM(9) => sig_IMM_9_port, IMM(8) =>
                           sig_IMM_8_port, IMM(7) => sig_IMM_7_port, IMM(6) => 
                           sig_IMM_6_port, IMM(5) => sig_IMM_5_port, IMM(4) => 
                           sig_IMM_4_port, IMM(3) => sig_IMM_3_port, IMM(2) => 
                           sig_IMM_2_port, IMM(1) => sig_IMM_1_port, IMM(0) => 
                           sig_IMM_0_port);
   regPC : regn_N32_8 port map( DIN(31) => PC_IN(31), DIN(30) => PC_IN(30), 
                           DIN(29) => PC_IN(29), DIN(28) => PC_IN(28), DIN(27) 
                           => PC_IN(27), DIN(26) => PC_IN(26), DIN(25) => 
                           PC_IN(25), DIN(24) => PC_IN(24), DIN(23) => 
                           PC_IN(23), DIN(22) => PC_IN(22), DIN(21) => 
                           PC_IN(21), DIN(20) => PC_IN(20), DIN(19) => 
                           PC_IN(19), DIN(18) => PC_IN(18), DIN(17) => 
                           PC_IN(17), DIN(16) => PC_IN(16), DIN(15) => 
                           PC_IN(15), DIN(14) => PC_IN(14), DIN(13) => 
                           PC_IN(13), DIN(12) => PC_IN(12), DIN(11) => 
                           PC_IN(11), DIN(10) => PC_IN(10), DIN(9) => PC_IN(9),
                           DIN(8) => PC_IN(8), DIN(7) => PC_IN(7), DIN(6) => 
                           PC_IN(6), DIN(5) => PC_IN(5), DIN(4) => PC_IN(4), 
                           DIN(3) => PC_IN(3), DIN(2) => PC_IN(2), DIN(1) => 
                           PC_IN(1), DIN(0) => PC_IN(0), CLK => CLK, EN => 
                           X_Logic1_port, RST => sig_RST, DOUT(31) => 
                           PC_OUT(31), DOUT(30) => PC_OUT(30), DOUT(29) => 
                           PC_OUT(29), DOUT(28) => PC_OUT(28), DOUT(27) => 
                           PC_OUT(27), DOUT(26) => PC_OUT(26), DOUT(25) => 
                           PC_OUT(25), DOUT(24) => PC_OUT(24), DOUT(23) => 
                           PC_OUT(23), DOUT(22) => PC_OUT(22), DOUT(21) => 
                           PC_OUT(21), DOUT(20) => PC_OUT(20), DOUT(19) => 
                           PC_OUT(19), DOUT(18) => PC_OUT(18), DOUT(17) => 
                           PC_OUT(17), DOUT(16) => PC_OUT(16), DOUT(15) => 
                           PC_OUT(15), DOUT(14) => PC_OUT(14), DOUT(13) => 
                           PC_OUT(13), DOUT(12) => PC_OUT(12), DOUT(11) => 
                           PC_OUT(11), DOUT(10) => PC_OUT(10), DOUT(9) => 
                           PC_OUT(9), DOUT(8) => PC_OUT(8), DOUT(7) => 
                           PC_OUT(7), DOUT(6) => PC_OUT(6), DOUT(5) => 
                           PC_OUT(5), DOUT(4) => PC_OUT(4), DOUT(3) => 
                           PC_OUT(3), DOUT(2) => PC_OUT(2), DOUT(1) => 
                           PC_OUT(1), DOUT(0) => PC_OUT(0));
   regIMM : regn_N32_7 port map( DIN(31) => sig_IMM_31_port, DIN(30) => 
                           sig_IMM_30_port, DIN(29) => sig_IMM_29_port, DIN(28)
                           => sig_IMM_28_port, DIN(27) => sig_IMM_27_port, 
                           DIN(26) => sig_IMM_26_port, DIN(25) => 
                           sig_IMM_25_port, DIN(24) => sig_IMM_24_port, DIN(23)
                           => sig_IMM_23_port, DIN(22) => sig_IMM_22_port, 
                           DIN(21) => sig_IMM_21_port, DIN(20) => 
                           sig_IMM_20_port, DIN(19) => sig_IMM_19_port, DIN(18)
                           => sig_IMM_18_port, DIN(17) => sig_IMM_17_port, 
                           DIN(16) => sig_IMM_16_port, DIN(15) => 
                           sig_IMM_15_port, DIN(14) => sig_IMM_14_port, DIN(13)
                           => sig_IMM_13_port, DIN(12) => sig_IMM_12_port, 
                           DIN(11) => sig_IMM_11_port, DIN(10) => 
                           sig_IMM_10_port, DIN(9) => sig_IMM_9_port, DIN(8) =>
                           sig_IMM_8_port, DIN(7) => sig_IMM_7_port, DIN(6) => 
                           sig_IMM_6_port, DIN(5) => sig_IMM_5_port, DIN(4) => 
                           sig_IMM_4_port, DIN(3) => sig_IMM_3_port, DIN(2) => 
                           sig_IMM_2_port, DIN(1) => sig_IMM_1_port, DIN(0) => 
                           sig_IMM_0_port, CLK => CLK, EN => REG_LATCH_EN, RST 
                           => sig_RST, DOUT(31) => IMM_OUT(31), DOUT(30) => 
                           IMM_OUT(30), DOUT(29) => IMM_OUT(29), DOUT(28) => 
                           IMM_OUT(28), DOUT(27) => IMM_OUT(27), DOUT(26) => 
                           IMM_OUT(26), DOUT(25) => IMM_OUT(25), DOUT(24) => 
                           IMM_OUT(24), DOUT(23) => IMM_OUT(23), DOUT(22) => 
                           IMM_OUT(22), DOUT(21) => IMM_OUT(21), DOUT(20) => 
                           IMM_OUT(20), DOUT(19) => IMM_OUT(19), DOUT(18) => 
                           IMM_OUT(18), DOUT(17) => IMM_OUT(17), DOUT(16) => 
                           IMM_OUT(16), DOUT(15) => IMM_OUT(15), DOUT(14) => 
                           IMM_OUT(14), DOUT(13) => IMM_OUT(13), DOUT(12) => 
                           IMM_OUT(12), DOUT(11) => IMM_OUT(11), DOUT(10) => 
                           IMM_OUT(10), DOUT(9) => IMM_OUT(9), DOUT(8) => 
                           IMM_OUT(8), DOUT(7) => IMM_OUT(7), DOUT(6) => 
                           IMM_OUT(6), DOUT(5) => IMM_OUT(5), DOUT(4) => 
                           IMM_OUT(4), DOUT(3) => IMM_OUT(3), DOUT(2) => 
                           IMM_OUT(2), DOUT(1) => IMM_OUT(1), DOUT(0) => 
                           IMM_OUT(0));
   regWR : regn_N5_0 port map( DIN(4) => sig_ADD_WR_4_port, DIN(3) => 
                           sig_ADD_WR_3_port, DIN(2) => sig_ADD_WR_2_port, 
                           DIN(1) => sig_ADD_WR_1_port, DIN(0) => 
                           sig_ADD_WR_0_port, CLK => CLK, EN => REG_LATCH_EN, 
                           RST => sig_RST, DOUT(4) => ADD_WR_OUT(4), DOUT(3) =>
                           ADD_WR_OUT(3), DOUT(2) => ADD_WR_OUT(2), DOUT(1) => 
                           ADD_WR_OUT(1), DOUT(0) => ADD_WR_OUT(0));
   regRS1 : regn_N5_4 port map( DIN(4) => ADD_RS1_HDU_4_port, DIN(3) => 
                           ADD_RS1_HDU_3_port, DIN(2) => ADD_RS1_HDU_2_port, 
                           DIN(1) => ADD_RS1_HDU_1_port, DIN(0) => 
                           ADD_RS1_HDU_0_port, CLK => CLK, EN => REG_LATCH_EN, 
                           RST => sig_RST, DOUT(4) => ADD_RS1_OUT(4), DOUT(3) 
                           => ADD_RS1_OUT(3), DOUT(2) => ADD_RS1_OUT(2), 
                           DOUT(1) => ADD_RS1_OUT(1), DOUT(0) => ADD_RS1_OUT(0)
                           );
   regRS2 : regn_N5_3 port map( DIN(4) => ADD_RS2_HDU_4_port, DIN(3) => 
                           ADD_RS2_HDU_3_port, DIN(2) => ADD_RS2_HDU_2_port, 
                           DIN(1) => ADD_RS2_HDU_1_port, DIN(0) => 
                           ADD_RS2_HDU_0_port, CLK => CLK, EN => REG_LATCH_EN, 
                           RST => sig_RST, DOUT(4) => ADD_RS2_OUT(4), DOUT(3) 
                           => ADD_RS2_OUT(3), DOUT(2) => ADD_RS2_OUT(2), 
                           DOUT(1) => ADD_RS2_OUT(1), DOUT(0) => ADD_RS2_OUT(0)
                           );
   rf : register_file_NBIT_ADD5_NBIT_DATA32 port map( CLK => CLK, RST => RST, 
                           ENABLE => REG_LATCH_EN, RD1 => RD1, RD2 => RD2, WR 
                           => RF_WE, ADD_WR(4) => ADD_WR(4), ADD_WR(3) => 
                           ADD_WR(3), ADD_WR(2) => ADD_WR(2), ADD_WR(1) => 
                           ADD_WR(1), ADD_WR(0) => ADD_WR(0), ADD_RS1(4) => 
                           ADD_RS1_HDU_4_port, ADD_RS1(3) => ADD_RS1_HDU_3_port
                           , ADD_RS1(2) => ADD_RS1_HDU_2_port, ADD_RS1(1) => 
                           ADD_RS1_HDU_1_port, ADD_RS1(0) => ADD_RS1_HDU_0_port
                           , ADD_RS2(4) => ADD_RS2_HDU_4_port, ADD_RS2(3) => 
                           ADD_RS2_HDU_3_port, ADD_RS2(2) => ADD_RS2_HDU_2_port
                           , ADD_RS2(1) => ADD_RS2_HDU_1_port, ADD_RS2(0) => 
                           ADD_RS2_HDU_0_port, DATAIN(31) => DATA_WR_IN(31), 
                           DATAIN(30) => DATA_WR_IN(30), DATAIN(29) => 
                           DATA_WR_IN(29), DATAIN(28) => DATA_WR_IN(28), 
                           DATAIN(27) => DATA_WR_IN(27), DATAIN(26) => 
                           DATA_WR_IN(26), DATAIN(25) => DATA_WR_IN(25), 
                           DATAIN(24) => DATA_WR_IN(24), DATAIN(23) => 
                           DATA_WR_IN(23), DATAIN(22) => DATA_WR_IN(22), 
                           DATAIN(21) => DATA_WR_IN(21), DATAIN(20) => 
                           DATA_WR_IN(20), DATAIN(19) => DATA_WR_IN(19), 
                           DATAIN(18) => DATA_WR_IN(18), DATAIN(17) => 
                           DATA_WR_IN(17), DATAIN(16) => DATA_WR_IN(16), 
                           DATAIN(15) => DATA_WR_IN(15), DATAIN(14) => 
                           DATA_WR_IN(14), DATAIN(13) => DATA_WR_IN(13), 
                           DATAIN(12) => DATA_WR_IN(12), DATAIN(11) => 
                           DATA_WR_IN(11), DATAIN(10) => DATA_WR_IN(10), 
                           DATAIN(9) => DATA_WR_IN(9), DATAIN(8) => 
                           DATA_WR_IN(8), DATAIN(7) => DATA_WR_IN(7), DATAIN(6)
                           => DATA_WR_IN(6), DATAIN(5) => DATA_WR_IN(5), 
                           DATAIN(4) => DATA_WR_IN(4), DATAIN(3) => 
                           DATA_WR_IN(3), DATAIN(2) => DATA_WR_IN(2), DATAIN(1)
                           => DATA_WR_IN(1), DATAIN(0) => DATA_WR_IN(0), 
                           OUT1(31) => A_OUT(31), OUT1(30) => A_OUT(30), 
                           OUT1(29) => A_OUT(29), OUT1(28) => A_OUT(28), 
                           OUT1(27) => A_OUT(27), OUT1(26) => A_OUT(26), 
                           OUT1(25) => A_OUT(25), OUT1(24) => A_OUT(24), 
                           OUT1(23) => A_OUT(23), OUT1(22) => A_OUT(22), 
                           OUT1(21) => A_OUT(21), OUT1(20) => A_OUT(20), 
                           OUT1(19) => A_OUT(19), OUT1(18) => A_OUT(18), 
                           OUT1(17) => A_OUT(17), OUT1(16) => A_OUT(16), 
                           OUT1(15) => A_OUT(15), OUT1(14) => A_OUT(14), 
                           OUT1(13) => A_OUT(13), OUT1(12) => A_OUT(12), 
                           OUT1(11) => A_OUT(11), OUT1(10) => A_OUT(10), 
                           OUT1(9) => A_OUT(9), OUT1(8) => A_OUT(8), OUT1(7) =>
                           A_OUT(7), OUT1(6) => A_OUT(6), OUT1(5) => A_OUT(5), 
                           OUT1(4) => A_OUT(4), OUT1(3) => A_OUT(3), OUT1(2) =>
                           A_OUT(2), OUT1(1) => A_OUT(1), OUT1(0) => A_OUT(0), 
                           OUT2(31) => B_OUT(31), OUT2(30) => B_OUT(30), 
                           OUT2(29) => B_OUT(29), OUT2(28) => B_OUT(28), 
                           OUT2(27) => B_OUT(27), OUT2(26) => B_OUT(26), 
                           OUT2(25) => B_OUT(25), OUT2(24) => B_OUT(24), 
                           OUT2(23) => B_OUT(23), OUT2(22) => B_OUT(22), 
                           OUT2(21) => B_OUT(21), OUT2(20) => B_OUT(20), 
                           OUT2(19) => B_OUT(19), OUT2(18) => B_OUT(18), 
                           OUT2(17) => B_OUT(17), OUT2(16) => B_OUT(16), 
                           OUT2(15) => B_OUT(15), OUT2(14) => B_OUT(14), 
                           OUT2(13) => B_OUT(13), OUT2(12) => B_OUT(12), 
                           OUT2(11) => B_OUT(11), OUT2(10) => B_OUT(10), 
                           OUT2(9) => B_OUT(9), OUT2(8) => B_OUT(8), OUT2(7) =>
                           B_OUT(7), OUT2(6) => B_OUT(6), OUT2(5) => B_OUT(5), 
                           OUT2(4) => B_OUT(4), OUT2(3) => B_OUT(3), OUT2(2) =>
                           B_OUT(2), OUT2(1) => B_OUT(1), OUT2(0) => B_OUT(0));
   U3 : INV_X1 port map( A => RST, ZN => n1);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Fetch is

   port( CLK, RST, ZERO_FLAG : in std_logic;  PC_EXT, INS_IN : in 
         std_logic_vector (31 downto 0);  Bubble_in : in std_logic;  HDU_INS_IN
         , HDU_PC_IN, HDU_NPC_IN : in std_logic_vector (31 downto 0);  PC_OUT, 
         ADDR_OUT, NPC_OUT, INS_OUT : out std_logic_vector (31 downto 0));

end Fetch;

architecture SYN_struct of Fetch is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component Fetch_DW01_add_3
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component regn_N32_9
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_10
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_0
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, ADDR_OUT_31_port, ADDR_OUT_30_port, ADDR_OUT_29_port, 
      ADDR_OUT_28_port, n27, n28, ADDR_OUT_25_port, ADDR_OUT_24_port, n29, n30,
      n31, ADDR_OUT_20_port, n32, n33, n34, n35, n36, n37, n38, 
      ADDR_OUT_12_port, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      ADDR_OUT_1_port, ADDR_OUT_0_port, sig_RST, sig_NPC_31_port, 
      sig_NPC_30_port, sig_NPC_29_port, sig_NPC_28_port, sig_NPC_27_port, 
      sig_NPC_26_port, sig_NPC_25_port, sig_NPC_24_port, sig_NPC_23_port, 
      sig_NPC_22_port, sig_NPC_21_port, sig_NPC_20_port, sig_NPC_19_port, 
      sig_NPC_18_port, sig_NPC_17_port, sig_NPC_16_port, sig_NPC_15_port, 
      sig_NPC_14_port, sig_NPC_13_port, sig_NPC_12_port, sig_NPC_11_port, 
      sig_NPC_10_port, sig_NPC_9_port, sig_NPC_8_port, sig_NPC_7_port, 
      sig_NPC_6_port, sig_NPC_5_port, sig_NPC_4_port, sig_NPC_3_port, 
      sig_NPC_2_port, sig_NPC_1_port, sig_NPC_0_port, PC_MUX_OUT_31_port, 
      PC_MUX_OUT_30_port, PC_MUX_OUT_29_port, PC_MUX_OUT_28_port, 
      PC_MUX_OUT_27_port, PC_MUX_OUT_26_port, PC_MUX_OUT_25_port, 
      PC_MUX_OUT_24_port, PC_MUX_OUT_23_port, PC_MUX_OUT_22_port, 
      PC_MUX_OUT_21_port, PC_MUX_OUT_20_port, PC_MUX_OUT_19_port, 
      PC_MUX_OUT_18_port, PC_MUX_OUT_17_port, PC_MUX_OUT_16_port, 
      PC_MUX_OUT_15_port, PC_MUX_OUT_14_port, PC_MUX_OUT_13_port, 
      PC_MUX_OUT_12_port, PC_MUX_OUT_11_port, PC_MUX_OUT_10_port, 
      PC_MUX_OUT_9_port, PC_MUX_OUT_8_port, PC_MUX_OUT_7_port, 
      PC_MUX_OUT_6_port, PC_MUX_OUT_5_port, PC_MUX_OUT_4_port, 
      PC_MUX_OUT_3_port, PC_MUX_OUT_2_port, PC_MUX_OUT_1_port, 
      PC_MUX_OUT_0_port, sig_INS_31_port, sig_INS_30_port, sig_INS_29_port, 
      sig_INS_28_port, sig_INS_27_port, sig_INS_26_port, sig_INS_25_port, 
      sig_INS_24_port, sig_INS_23_port, sig_INS_22_port, sig_INS_21_port, 
      sig_INS_20_port, sig_INS_19_port, sig_INS_18_port, sig_INS_17_port, 
      sig_INS_16_port, sig_INS_15_port, sig_INS_14_port, sig_INS_13_port, 
      sig_INS_12_port, sig_INS_11_port, sig_INS_10_port, sig_INS_9_port, 
      sig_INS_8_port, sig_INS_7_port, sig_INS_6_port, sig_INS_5_port, 
      sig_INS_4_port, sig_INS_3_port, sig_INS_2_port, sig_INS_1_port, 
      sig_INS_0_port, n1, n2, n3, ADDR_OUT_23_port, ADDR_OUT_22_port, 
      ADDR_OUT_26_port, ADDR_OUT_4_port, ADDR_OUT_9_port, ADDR_OUT_8_port, 
      ADDR_OUT_2_port, ADDR_OUT_3_port, ADDR_OUT_21_port, ADDR_OUT_19_port, 
      ADDR_OUT_18_port, ADDR_OUT_16_port, ADDR_OUT_27_port, ADDR_OUT_7_port, 
      ADDR_OUT_15_port, ADDR_OUT_14_port, ADDR_OUT_5_port, ADDR_OUT_10_port, 
      ADDR_OUT_17_port, ADDR_OUT_11_port, ADDR_OUT_13_port, ADDR_OUT_6_port, 
      n26, n_1828 : std_logic;

begin
   ADDR_OUT <= ( ADDR_OUT_31_port, ADDR_OUT_30_port, ADDR_OUT_29_port, 
      ADDR_OUT_28_port, ADDR_OUT_27_port, ADDR_OUT_26_port, ADDR_OUT_25_port, 
      ADDR_OUT_24_port, ADDR_OUT_23_port, ADDR_OUT_22_port, ADDR_OUT_21_port, 
      ADDR_OUT_20_port, ADDR_OUT_19_port, ADDR_OUT_18_port, ADDR_OUT_17_port, 
      ADDR_OUT_16_port, ADDR_OUT_15_port, ADDR_OUT_14_port, ADDR_OUT_13_port, 
      ADDR_OUT_12_port, ADDR_OUT_11_port, ADDR_OUT_10_port, ADDR_OUT_9_port, 
      ADDR_OUT_8_port, ADDR_OUT_7_port, ADDR_OUT_6_port, ADDR_OUT_5_port, 
      ADDR_OUT_4_port, ADDR_OUT_3_port, ADDR_OUT_2_port, ADDR_OUT_1_port, 
      ADDR_OUT_0_port );
   
   X_Logic1_port <= '1';
   n1 <= '0';
   n2 <= '1';
   n3 <= '0';
   NPC_or_NPC_HDU : mux21_NBIT32_0 port map( A(31) => PC_EXT(31), A(30) => 
                           PC_EXT(30), A(29) => PC_EXT(29), A(28) => PC_EXT(28)
                           , A(27) => PC_EXT(27), A(26) => PC_EXT(26), A(25) =>
                           PC_EXT(25), A(24) => PC_EXT(24), A(23) => PC_EXT(23)
                           , A(22) => PC_EXT(22), A(21) => PC_EXT(21), A(20) =>
                           PC_EXT(20), A(19) => PC_EXT(19), A(18) => PC_EXT(18)
                           , A(17) => PC_EXT(17), A(16) => PC_EXT(16), A(15) =>
                           PC_EXT(15), A(14) => PC_EXT(14), A(13) => PC_EXT(13)
                           , A(12) => PC_EXT(12), A(11) => PC_EXT(11), A(10) =>
                           PC_EXT(10), A(9) => PC_EXT(9), A(8) => PC_EXT(8), 
                           A(7) => PC_EXT(7), A(6) => PC_EXT(6), A(5) => 
                           PC_EXT(5), A(4) => PC_EXT(4), A(3) => PC_EXT(3), 
                           A(2) => PC_EXT(2), A(1) => PC_EXT(1), A(0) => 
                           PC_EXT(0), B(31) => HDU_NPC_IN(31), B(30) => 
                           HDU_NPC_IN(30), B(29) => HDU_NPC_IN(29), B(28) => 
                           HDU_NPC_IN(28), B(27) => HDU_NPC_IN(27), B(26) => 
                           HDU_NPC_IN(26), B(25) => HDU_NPC_IN(25), B(24) => 
                           HDU_NPC_IN(24), B(23) => HDU_NPC_IN(23), B(22) => 
                           HDU_NPC_IN(22), B(21) => HDU_NPC_IN(21), B(20) => 
                           HDU_NPC_IN(20), B(19) => HDU_NPC_IN(19), B(18) => 
                           HDU_NPC_IN(18), B(17) => HDU_NPC_IN(17), B(16) => 
                           HDU_NPC_IN(16), B(15) => HDU_NPC_IN(15), B(14) => 
                           HDU_NPC_IN(14), B(13) => HDU_NPC_IN(13), B(12) => 
                           HDU_NPC_IN(12), B(11) => HDU_NPC_IN(11), B(10) => 
                           HDU_NPC_IN(10), B(9) => HDU_NPC_IN(9), B(8) => 
                           HDU_NPC_IN(8), B(7) => HDU_NPC_IN(7), B(6) => 
                           HDU_NPC_IN(6), B(5) => HDU_NPC_IN(5), B(4) => 
                           HDU_NPC_IN(4), B(3) => HDU_NPC_IN(3), B(2) => 
                           HDU_NPC_IN(2), B(1) => HDU_NPC_IN(1), B(0) => 
                           HDU_NPC_IN(0), S => Bubble_in, Z(31) => 
                           sig_NPC_31_port, Z(30) => sig_NPC_30_port, Z(29) => 
                           sig_NPC_29_port, Z(28) => sig_NPC_28_port, Z(27) => 
                           sig_NPC_27_port, Z(26) => sig_NPC_26_port, Z(25) => 
                           sig_NPC_25_port, Z(24) => sig_NPC_24_port, Z(23) => 
                           sig_NPC_23_port, Z(22) => sig_NPC_22_port, Z(21) => 
                           sig_NPC_21_port, Z(20) => sig_NPC_20_port, Z(19) => 
                           sig_NPC_19_port, Z(18) => sig_NPC_18_port, Z(17) => 
                           sig_NPC_17_port, Z(16) => sig_NPC_16_port, Z(15) => 
                           sig_NPC_15_port, Z(14) => sig_NPC_14_port, Z(13) => 
                           sig_NPC_13_port, Z(12) => sig_NPC_12_port, Z(11) => 
                           sig_NPC_11_port, Z(10) => sig_NPC_10_port, Z(9) => 
                           sig_NPC_9_port, Z(8) => sig_NPC_8_port, Z(7) => 
                           sig_NPC_7_port, Z(6) => sig_NPC_6_port, Z(5) => 
                           sig_NPC_5_port, Z(4) => sig_NPC_4_port, Z(3) => 
                           sig_NPC_3_port, Z(2) => sig_NPC_2_port, Z(1) => 
                           sig_NPC_1_port, Z(0) => sig_NPC_0_port);
   PC_or_PC_HDU : mux21_NBIT32_5 port map( A(31) => ADDR_OUT_31_port, A(30) => 
                           ADDR_OUT_30_port, A(29) => ADDR_OUT_29_port, A(28) 
                           => ADDR_OUT_28_port, A(27) => ADDR_OUT_27_port, 
                           A(26) => ADDR_OUT_26_port, A(25) => ADDR_OUT_25_port
                           , A(24) => ADDR_OUT_24_port, A(23) => 
                           ADDR_OUT_23_port, A(22) => ADDR_OUT_22_port, A(21) 
                           => ADDR_OUT_21_port, A(20) => ADDR_OUT_20_port, 
                           A(19) => ADDR_OUT_19_port, A(18) => ADDR_OUT_18_port
                           , A(17) => ADDR_OUT_17_port, A(16) => 
                           ADDR_OUT_16_port, A(15) => ADDR_OUT_15_port, A(14) 
                           => ADDR_OUT_14_port, A(13) => ADDR_OUT_13_port, 
                           A(12) => ADDR_OUT_12_port, A(11) => ADDR_OUT_11_port
                           , A(10) => ADDR_OUT_10_port, A(9) => ADDR_OUT_9_port
                           , A(8) => ADDR_OUT_8_port, A(7) => ADDR_OUT_7_port, 
                           A(6) => ADDR_OUT_6_port, A(5) => ADDR_OUT_5_port, 
                           A(4) => ADDR_OUT_4_port, A(3) => ADDR_OUT_3_port, 
                           A(2) => ADDR_OUT_2_port, A(1) => ADDR_OUT_1_port, 
                           A(0) => ADDR_OUT_0_port, B(31) => HDU_PC_IN(31), 
                           B(30) => HDU_PC_IN(30), B(29) => HDU_PC_IN(29), 
                           B(28) => HDU_PC_IN(28), B(27) => HDU_PC_IN(27), 
                           B(26) => HDU_PC_IN(26), B(25) => HDU_PC_IN(25), 
                           B(24) => HDU_PC_IN(24), B(23) => HDU_PC_IN(23), 
                           B(22) => HDU_PC_IN(22), B(21) => HDU_PC_IN(21), 
                           B(20) => HDU_PC_IN(20), B(19) => HDU_PC_IN(19), 
                           B(18) => HDU_PC_IN(18), B(17) => HDU_PC_IN(17), 
                           B(16) => HDU_PC_IN(16), B(15) => HDU_PC_IN(15), 
                           B(14) => HDU_PC_IN(14), B(13) => HDU_PC_IN(13), 
                           B(12) => HDU_PC_IN(12), B(11) => HDU_PC_IN(11), 
                           B(10) => HDU_PC_IN(10), B(9) => HDU_PC_IN(9), B(8) 
                           => HDU_PC_IN(8), B(7) => HDU_PC_IN(7), B(6) => 
                           HDU_PC_IN(6), B(5) => HDU_PC_IN(5), B(4) => 
                           HDU_PC_IN(4), B(3) => HDU_PC_IN(3), B(2) => 
                           HDU_PC_IN(2), B(1) => HDU_PC_IN(1), B(0) => 
                           HDU_PC_IN(0), S => Bubble_in, Z(31) => 
                           PC_MUX_OUT_31_port, Z(30) => PC_MUX_OUT_30_port, 
                           Z(29) => PC_MUX_OUT_29_port, Z(28) => 
                           PC_MUX_OUT_28_port, Z(27) => PC_MUX_OUT_27_port, 
                           Z(26) => PC_MUX_OUT_26_port, Z(25) => 
                           PC_MUX_OUT_25_port, Z(24) => PC_MUX_OUT_24_port, 
                           Z(23) => PC_MUX_OUT_23_port, Z(22) => 
                           PC_MUX_OUT_22_port, Z(21) => PC_MUX_OUT_21_port, 
                           Z(20) => PC_MUX_OUT_20_port, Z(19) => 
                           PC_MUX_OUT_19_port, Z(18) => PC_MUX_OUT_18_port, 
                           Z(17) => PC_MUX_OUT_17_port, Z(16) => 
                           PC_MUX_OUT_16_port, Z(15) => PC_MUX_OUT_15_port, 
                           Z(14) => PC_MUX_OUT_14_port, Z(13) => 
                           PC_MUX_OUT_13_port, Z(12) => PC_MUX_OUT_12_port, 
                           Z(11) => PC_MUX_OUT_11_port, Z(10) => 
                           PC_MUX_OUT_10_port, Z(9) => PC_MUX_OUT_9_port, Z(8) 
                           => PC_MUX_OUT_8_port, Z(7) => PC_MUX_OUT_7_port, 
                           Z(6) => PC_MUX_OUT_6_port, Z(5) => PC_MUX_OUT_5_port
                           , Z(4) => PC_MUX_OUT_4_port, Z(3) => 
                           PC_MUX_OUT_3_port, Z(2) => PC_MUX_OUT_2_port, Z(1) 
                           => PC_MUX_OUT_1_port, Z(0) => PC_MUX_OUT_0_port);
   INS_or_HDU_INS : mux21_NBIT32_4 port map( A(31) => INS_IN(31), A(30) => 
                           INS_IN(30), A(29) => INS_IN(29), A(28) => INS_IN(28)
                           , A(27) => INS_IN(27), A(26) => INS_IN(26), A(25) =>
                           INS_IN(25), A(24) => INS_IN(24), A(23) => INS_IN(23)
                           , A(22) => INS_IN(22), A(21) => INS_IN(21), A(20) =>
                           INS_IN(20), A(19) => INS_IN(19), A(18) => INS_IN(18)
                           , A(17) => INS_IN(17), A(16) => INS_IN(16), A(15) =>
                           INS_IN(15), A(14) => INS_IN(14), A(13) => INS_IN(13)
                           , A(12) => INS_IN(12), A(11) => INS_IN(11), A(10) =>
                           INS_IN(10), A(9) => INS_IN(9), A(8) => INS_IN(8), 
                           A(7) => INS_IN(7), A(6) => INS_IN(6), A(5) => 
                           INS_IN(5), A(4) => INS_IN(4), A(3) => INS_IN(3), 
                           A(2) => INS_IN(2), A(1) => INS_IN(1), A(0) => 
                           INS_IN(0), B(31) => HDU_INS_IN(31), B(30) => 
                           HDU_INS_IN(30), B(29) => HDU_INS_IN(29), B(28) => 
                           HDU_INS_IN(28), B(27) => HDU_INS_IN(27), B(26) => 
                           HDU_INS_IN(26), B(25) => HDU_INS_IN(25), B(24) => 
                           HDU_INS_IN(24), B(23) => HDU_INS_IN(23), B(22) => 
                           HDU_INS_IN(22), B(21) => HDU_INS_IN(21), B(20) => 
                           HDU_INS_IN(20), B(19) => HDU_INS_IN(19), B(18) => 
                           HDU_INS_IN(18), B(17) => HDU_INS_IN(17), B(16) => 
                           HDU_INS_IN(16), B(15) => HDU_INS_IN(15), B(14) => 
                           HDU_INS_IN(14), B(13) => HDU_INS_IN(13), B(12) => 
                           HDU_INS_IN(12), B(11) => HDU_INS_IN(11), B(10) => 
                           HDU_INS_IN(10), B(9) => HDU_INS_IN(9), B(8) => 
                           HDU_INS_IN(8), B(7) => HDU_INS_IN(7), B(6) => 
                           HDU_INS_IN(6), B(5) => HDU_INS_IN(5), B(4) => 
                           HDU_INS_IN(4), B(3) => HDU_INS_IN(3), B(2) => 
                           HDU_INS_IN(2), B(1) => HDU_INS_IN(1), B(0) => 
                           HDU_INS_IN(0), S => Bubble_in, Z(31) => 
                           sig_INS_31_port, Z(30) => sig_INS_30_port, Z(29) => 
                           sig_INS_29_port, Z(28) => sig_INS_28_port, Z(27) => 
                           sig_INS_27_port, Z(26) => sig_INS_26_port, Z(25) => 
                           sig_INS_25_port, Z(24) => sig_INS_24_port, Z(23) => 
                           sig_INS_23_port, Z(22) => sig_INS_22_port, Z(21) => 
                           sig_INS_21_port, Z(20) => sig_INS_20_port, Z(19) => 
                           sig_INS_19_port, Z(18) => sig_INS_18_port, Z(17) => 
                           sig_INS_17_port, Z(16) => sig_INS_16_port, Z(15) => 
                           sig_INS_15_port, Z(14) => sig_INS_14_port, Z(13) => 
                           sig_INS_13_port, Z(12) => sig_INS_12_port, Z(11) => 
                           sig_INS_11_port, Z(10) => sig_INS_10_port, Z(9) => 
                           sig_INS_9_port, Z(8) => sig_INS_8_port, Z(7) => 
                           sig_INS_7_port, Z(6) => sig_INS_6_port, Z(5) => 
                           sig_INS_5_port, Z(4) => sig_INS_4_port, Z(3) => 
                           sig_INS_3_port, Z(2) => sig_INS_2_port, Z(1) => 
                           sig_INS_1_port, Z(0) => sig_INS_0_port);
   PC : regn_N32_0 port map( DIN(31) => sig_NPC_31_port, DIN(30) => 
                           sig_NPC_30_port, DIN(29) => sig_NPC_29_port, DIN(28)
                           => sig_NPC_28_port, DIN(27) => sig_NPC_27_port, 
                           DIN(26) => sig_NPC_26_port, DIN(25) => 
                           sig_NPC_25_port, DIN(24) => sig_NPC_24_port, DIN(23)
                           => sig_NPC_23_port, DIN(22) => sig_NPC_22_port, 
                           DIN(21) => sig_NPC_21_port, DIN(20) => 
                           sig_NPC_20_port, DIN(19) => sig_NPC_19_port, DIN(18)
                           => sig_NPC_18_port, DIN(17) => sig_NPC_17_port, 
                           DIN(16) => sig_NPC_16_port, DIN(15) => 
                           sig_NPC_15_port, DIN(14) => sig_NPC_14_port, DIN(13)
                           => sig_NPC_13_port, DIN(12) => sig_NPC_12_port, 
                           DIN(11) => sig_NPC_11_port, DIN(10) => 
                           sig_NPC_10_port, DIN(9) => sig_NPC_9_port, DIN(8) =>
                           sig_NPC_8_port, DIN(7) => sig_NPC_7_port, DIN(6) => 
                           sig_NPC_6_port, DIN(5) => sig_NPC_5_port, DIN(4) => 
                           sig_NPC_4_port, DIN(3) => sig_NPC_3_port, DIN(2) => 
                           sig_NPC_2_port, DIN(1) => sig_NPC_1_port, DIN(0) => 
                           sig_NPC_0_port, CLK => CLK, EN => X_Logic1_port, RST
                           => RST, DOUT(31) => ADDR_OUT_31_port, DOUT(30) => 
                           ADDR_OUT_30_port, DOUT(29) => ADDR_OUT_29_port, 
                           DOUT(28) => ADDR_OUT_28_port, DOUT(27) => n27, 
                           DOUT(26) => n28, DOUT(25) => ADDR_OUT_25_port, 
                           DOUT(24) => ADDR_OUT_24_port, DOUT(23) => n29, 
                           DOUT(22) => n30, DOUT(21) => n31, DOUT(20) => 
                           ADDR_OUT_20_port, DOUT(19) => n32, DOUT(18) => n33, 
                           DOUT(17) => n34, DOUT(16) => n35, DOUT(15) => n36, 
                           DOUT(14) => n37, DOUT(13) => n38, DOUT(12) => 
                           ADDR_OUT_12_port, DOUT(11) => n39, DOUT(10) => n40, 
                           DOUT(9) => n41, DOUT(8) => n42, DOUT(7) => n43, 
                           DOUT(6) => n44, DOUT(5) => n45, DOUT(4) => n46, 
                           DOUT(3) => n47, DOUT(2) => n48, DOUT(1) => 
                           ADDR_OUT_1_port, DOUT(0) => ADDR_OUT_0_port);
   PC_reg : regn_N32_10 port map( DIN(31) => PC_MUX_OUT_31_port, DIN(30) => 
                           PC_MUX_OUT_30_port, DIN(29) => PC_MUX_OUT_29_port, 
                           DIN(28) => PC_MUX_OUT_28_port, DIN(27) => 
                           PC_MUX_OUT_27_port, DIN(26) => PC_MUX_OUT_26_port, 
                           DIN(25) => PC_MUX_OUT_25_port, DIN(24) => 
                           PC_MUX_OUT_24_port, DIN(23) => PC_MUX_OUT_23_port, 
                           DIN(22) => PC_MUX_OUT_22_port, DIN(21) => 
                           PC_MUX_OUT_21_port, DIN(20) => PC_MUX_OUT_20_port, 
                           DIN(19) => PC_MUX_OUT_19_port, DIN(18) => 
                           PC_MUX_OUT_18_port, DIN(17) => PC_MUX_OUT_17_port, 
                           DIN(16) => PC_MUX_OUT_16_port, DIN(15) => 
                           PC_MUX_OUT_15_port, DIN(14) => PC_MUX_OUT_14_port, 
                           DIN(13) => PC_MUX_OUT_13_port, DIN(12) => 
                           PC_MUX_OUT_12_port, DIN(11) => PC_MUX_OUT_11_port, 
                           DIN(10) => PC_MUX_OUT_10_port, DIN(9) => 
                           PC_MUX_OUT_9_port, DIN(8) => PC_MUX_OUT_8_port, 
                           DIN(7) => PC_MUX_OUT_7_port, DIN(6) => 
                           PC_MUX_OUT_6_port, DIN(5) => PC_MUX_OUT_5_port, 
                           DIN(4) => PC_MUX_OUT_4_port, DIN(3) => 
                           PC_MUX_OUT_3_port, DIN(2) => PC_MUX_OUT_2_port, 
                           DIN(1) => PC_MUX_OUT_1_port, DIN(0) => 
                           PC_MUX_OUT_0_port, CLK => CLK, EN => X_Logic1_port, 
                           RST => sig_RST, DOUT(31) => PC_OUT(31), DOUT(30) => 
                           PC_OUT(30), DOUT(29) => PC_OUT(29), DOUT(28) => 
                           PC_OUT(28), DOUT(27) => PC_OUT(27), DOUT(26) => 
                           PC_OUT(26), DOUT(25) => PC_OUT(25), DOUT(24) => 
                           PC_OUT(24), DOUT(23) => PC_OUT(23), DOUT(22) => 
                           PC_OUT(22), DOUT(21) => PC_OUT(21), DOUT(20) => 
                           PC_OUT(20), DOUT(19) => PC_OUT(19), DOUT(18) => 
                           PC_OUT(18), DOUT(17) => PC_OUT(17), DOUT(16) => 
                           PC_OUT(16), DOUT(15) => PC_OUT(15), DOUT(14) => 
                           PC_OUT(14), DOUT(13) => PC_OUT(13), DOUT(12) => 
                           PC_OUT(12), DOUT(11) => PC_OUT(11), DOUT(10) => 
                           PC_OUT(10), DOUT(9) => PC_OUT(9), DOUT(8) => 
                           PC_OUT(8), DOUT(7) => PC_OUT(7), DOUT(6) => 
                           PC_OUT(6), DOUT(5) => PC_OUT(5), DOUT(4) => 
                           PC_OUT(4), DOUT(3) => PC_OUT(3), DOUT(2) => 
                           PC_OUT(2), DOUT(1) => PC_OUT(1), DOUT(0) => 
                           PC_OUT(0));
   IR : regn_N32_9 port map( DIN(31) => sig_INS_31_port, DIN(30) => 
                           sig_INS_30_port, DIN(29) => sig_INS_29_port, DIN(28)
                           => sig_INS_28_port, DIN(27) => sig_INS_27_port, 
                           DIN(26) => sig_INS_26_port, DIN(25) => 
                           sig_INS_25_port, DIN(24) => sig_INS_24_port, DIN(23)
                           => sig_INS_23_port, DIN(22) => sig_INS_22_port, 
                           DIN(21) => sig_INS_21_port, DIN(20) => 
                           sig_INS_20_port, DIN(19) => sig_INS_19_port, DIN(18)
                           => sig_INS_18_port, DIN(17) => sig_INS_17_port, 
                           DIN(16) => sig_INS_16_port, DIN(15) => 
                           sig_INS_15_port, DIN(14) => sig_INS_14_port, DIN(13)
                           => sig_INS_13_port, DIN(12) => sig_INS_12_port, 
                           DIN(11) => sig_INS_11_port, DIN(10) => 
                           sig_INS_10_port, DIN(9) => sig_INS_9_port, DIN(8) =>
                           sig_INS_8_port, DIN(7) => sig_INS_7_port, DIN(6) => 
                           sig_INS_6_port, DIN(5) => sig_INS_5_port, DIN(4) => 
                           sig_INS_4_port, DIN(3) => sig_INS_3_port, DIN(2) => 
                           sig_INS_2_port, DIN(1) => sig_INS_1_port, DIN(0) => 
                           sig_INS_0_port, CLK => CLK, EN => X_Logic1_port, RST
                           => sig_RST, DOUT(31) => INS_OUT(31), DOUT(30) => 
                           INS_OUT(30), DOUT(29) => INS_OUT(29), DOUT(28) => 
                           INS_OUT(28), DOUT(27) => INS_OUT(27), DOUT(26) => 
                           INS_OUT(26), DOUT(25) => INS_OUT(25), DOUT(24) => 
                           INS_OUT(24), DOUT(23) => INS_OUT(23), DOUT(22) => 
                           INS_OUT(22), DOUT(21) => INS_OUT(21), DOUT(20) => 
                           INS_OUT(20), DOUT(19) => INS_OUT(19), DOUT(18) => 
                           INS_OUT(18), DOUT(17) => INS_OUT(17), DOUT(16) => 
                           INS_OUT(16), DOUT(15) => INS_OUT(15), DOUT(14) => 
                           INS_OUT(14), DOUT(13) => INS_OUT(13), DOUT(12) => 
                           INS_OUT(12), DOUT(11) => INS_OUT(11), DOUT(10) => 
                           INS_OUT(10), DOUT(9) => INS_OUT(9), DOUT(8) => 
                           INS_OUT(8), DOUT(7) => INS_OUT(7), DOUT(6) => 
                           INS_OUT(6), DOUT(5) => INS_OUT(5), DOUT(4) => 
                           INS_OUT(4), DOUT(3) => INS_OUT(3), DOUT(2) => 
                           INS_OUT(2), DOUT(1) => INS_OUT(1), DOUT(0) => 
                           INS_OUT(0));
   add_54 : Fetch_DW01_add_3 port map( A(31) => ADDR_OUT_31_port, A(30) => 
                           ADDR_OUT_30_port, A(29) => ADDR_OUT_29_port, A(28) 
                           => ADDR_OUT_28_port, A(27) => n27, A(26) => n28, 
                           A(25) => ADDR_OUT_25_port, A(24) => ADDR_OUT_24_port
                           , A(23) => n29, A(22) => n30, A(21) => n31, A(20) =>
                           ADDR_OUT_20_port, A(19) => n32, A(18) => n33, A(17) 
                           => n34, A(16) => n35, A(15) => n36, A(14) => n37, 
                           A(13) => n38, A(12) => ADDR_OUT_12_port, A(11) => 
                           n39, A(10) => n40, A(9) => n41, A(8) => n42, A(7) =>
                           n43, A(6) => n44, A(5) => n45, A(4) => n46, A(3) => 
                           n47, A(2) => n48, A(1) => ADDR_OUT_1_port, A(0) => 
                           ADDR_OUT_0_port, B(31) => n1, B(30) => n1, B(29) => 
                           n1, B(28) => n1, B(27) => n1, B(26) => n1, B(25) => 
                           n1, B(24) => n1, B(23) => n1, B(22) => n1, B(21) => 
                           n1, B(20) => n1, B(19) => n1, B(18) => n1, B(17) => 
                           n1, B(16) => n1, B(15) => n1, B(14) => n1, B(13) => 
                           n1, B(12) => n1, B(11) => n1, B(10) => n1, B(9) => 
                           n1, B(8) => n1, B(7) => n1, B(6) => n1, B(5) => n1, 
                           B(4) => n1, B(3) => n1, B(2) => n2, B(1) => n1, B(0)
                           => n1, CI => n3, SUM(31) => NPC_OUT(31), SUM(30) => 
                           NPC_OUT(30), SUM(29) => NPC_OUT(29), SUM(28) => 
                           NPC_OUT(28), SUM(27) => NPC_OUT(27), SUM(26) => 
                           NPC_OUT(26), SUM(25) => NPC_OUT(25), SUM(24) => 
                           NPC_OUT(24), SUM(23) => NPC_OUT(23), SUM(22) => 
                           NPC_OUT(22), SUM(21) => NPC_OUT(21), SUM(20) => 
                           NPC_OUT(20), SUM(19) => NPC_OUT(19), SUM(18) => 
                           NPC_OUT(18), SUM(17) => NPC_OUT(17), SUM(16) => 
                           NPC_OUT(16), SUM(15) => NPC_OUT(15), SUM(14) => 
                           NPC_OUT(14), SUM(13) => NPC_OUT(13), SUM(12) => 
                           NPC_OUT(12), SUM(11) => NPC_OUT(11), SUM(10) => 
                           NPC_OUT(10), SUM(9) => NPC_OUT(9), SUM(8) => 
                           NPC_OUT(8), SUM(7) => NPC_OUT(7), SUM(6) => 
                           NPC_OUT(6), SUM(5) => NPC_OUT(5), SUM(4) => 
                           NPC_OUT(4), SUM(3) => NPC_OUT(3), SUM(2) => 
                           NPC_OUT(2), SUM(1) => NPC_OUT(1), SUM(0) => 
                           NPC_OUT(0), CO => n_1828);
   U6 : BUF_X1 port map( A => n46, Z => ADDR_OUT_4_port);
   U7 : CLKBUF_X1 port map( A => n29, Z => ADDR_OUT_23_port);
   U8 : CLKBUF_X1 port map( A => n30, Z => ADDR_OUT_22_port);
   U9 : CLKBUF_X1 port map( A => n28, Z => ADDR_OUT_26_port);
   U10 : CLKBUF_X1 port map( A => n41, Z => ADDR_OUT_9_port);
   U11 : CLKBUF_X1 port map( A => n42, Z => ADDR_OUT_8_port);
   U12 : CLKBUF_X1 port map( A => n48, Z => ADDR_OUT_2_port);
   U13 : CLKBUF_X1 port map( A => n47, Z => ADDR_OUT_3_port);
   U14 : CLKBUF_X1 port map( A => n31, Z => ADDR_OUT_21_port);
   U15 : CLKBUF_X1 port map( A => n32, Z => ADDR_OUT_19_port);
   U16 : CLKBUF_X1 port map( A => n33, Z => ADDR_OUT_18_port);
   U17 : CLKBUF_X1 port map( A => n35, Z => ADDR_OUT_16_port);
   U18 : CLKBUF_X1 port map( A => n27, Z => ADDR_OUT_27_port);
   U19 : CLKBUF_X1 port map( A => n43, Z => ADDR_OUT_7_port);
   U20 : NOR2_X1 port map( A1 => ZERO_FLAG, A2 => n26, ZN => sig_RST);
   U21 : CLKBUF_X1 port map( A => n36, Z => ADDR_OUT_15_port);
   U22 : CLKBUF_X1 port map( A => n37, Z => ADDR_OUT_14_port);
   U23 : CLKBUF_X1 port map( A => n45, Z => ADDR_OUT_5_port);
   U24 : CLKBUF_X1 port map( A => n40, Z => ADDR_OUT_10_port);
   U25 : CLKBUF_X1 port map( A => n34, Z => ADDR_OUT_17_port);
   U26 : CLKBUF_X1 port map( A => n39, Z => ADDR_OUT_11_port);
   U27 : CLKBUF_X1 port map( A => n38, Z => ADDR_OUT_13_port);
   U28 : CLKBUF_X1 port map( A => n44, Z => ADDR_OUT_6_port);
   U29 : INV_X1 port map( A => RST, ZN => n26);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity hardwired_cu_NBIT32 is

   port( REG_LATCH_EN, RD1, RD2, MUX_A_SEL : out std_logic;  MUX_B_SEL : out 
         std_logic_vector (1 downto 0);  ALU_OPC : out std_logic_vector (0 to 
         3);  ALU_OUTREG_EN, DRAM_R_IN : out std_logic;  JUMP_TYPE : out 
         std_logic_vector (1 downto 0);  MEM_EN_IN, DRAM_W_IN, RF_WE, 
         DRAM_EN_IN, WB_MUX_SEL : out std_logic;  INS_IN : in std_logic_vector 
         (31 downto 0);  Bubble, Clk, Rst : in std_logic);

end hardwired_cu_NBIT32;

architecture SYN_bhv of hardwired_cu_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal AluOP_E_3_port, AluOP_E_2_port, AluOP_E_1_port, AluOP_E_0_port, N24, 
      N25, N26, N27, n19, n20, n21, n22, n23, n24_port, n25_port, n26_port, 
      n27_port, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40
      , n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, 
      n55, n56, n58, n59, n60, n61, n62, n63, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n_1829, n_1830, n_1831, 
      n_1832, n_1833, n_1834, n_1835, n_1836 : std_logic;

begin
   
   AluOP_E_reg_3_inst : DFFR_X1 port map( D => N27, CK => Clk, RN => Rst, Q => 
                           AluOP_E_3_port, QN => n_1829);
   ALU_OPC_reg_3_inst : DFFR_X1 port map( D => AluOP_E_3_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(0), QN => n_1830);
   AluOP_E_reg_2_inst : DFFR_X1 port map( D => N26, CK => Clk, RN => Rst, Q => 
                           AluOP_E_2_port, QN => n_1831);
   ALU_OPC_reg_2_inst : DFFR_X1 port map( D => AluOP_E_2_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(1), QN => n_1832);
   AluOP_E_reg_1_inst : DFFR_X1 port map( D => N25, CK => Clk, RN => Rst, Q => 
                           AluOP_E_1_port, QN => n_1833);
   ALU_OPC_reg_1_inst : DFFR_X1 port map( D => AluOP_E_1_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(2), QN => n_1834);
   AluOP_E_reg_0_inst : DFFR_X1 port map( D => N24, CK => Clk, RN => Rst, Q => 
                           AluOP_E_0_port, QN => n_1835);
   ALU_OPC_reg_0_inst : DFFR_X1 port map( D => AluOP_E_0_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(3), QN => n_1836);
   WB_MUX_SEL <= '0';
   DRAM_EN_IN <= '0';
   RF_WE <= '0';
   DRAM_W_IN <= '0';
   MEM_EN_IN <= '0';
   JUMP_TYPE(0) <= '0';
   JUMP_TYPE(1) <= '0';
   DRAM_R_IN <= '0';
   ALU_OUTREG_EN <= '0';
   MUX_B_SEL(0) <= '0';
   MUX_B_SEL(1) <= '0';
   MUX_A_SEL <= '0';
   RD2 <= '0';
   RD1 <= '0';
   REG_LATCH_EN <= '0';
   U74 : XOR2_X1 port map( A => n2, B => INS_IN(1), Z => n33);
   U75 : NAND3_X1 port map( A1 => n16, A2 => n13, A3 => INS_IN(30), ZN => n37);
   U76 : OAI33_X1 port map( A1 => n26_port, A2 => n13, A3 => n17, B1 => n46, B2
                           => INS_IN(30), B3 => INS_IN(28), ZN => n43);
   U77 : OAI33_X1 port map( A1 => n24_port, A2 => n25_port, A3 => n17, B1 => n3
                           , B2 => n8, B3 => n34, ZN => n50);
   U78 : OAI33_X1 port map( A1 => n12, A2 => n56, A3 => n11, B1 => n27_port, B2
                           => INS_IN(30), B3 => n25_port, ZN => n55);
   U79 : NAND3_X1 port map( A1 => n51, A2 => n7, A3 => INS_IN(5), ZN => n35);
   U80 : OAI33_X1 port map( A1 => n58, A2 => n13, A3 => n17, B1 => n59, B2 => 
                           n39, B3 => n6, ZN => n48);
   U81 : NAND3_X1 port map( A1 => INS_IN(3), A2 => n51, A3 => INS_IN(5), ZN => 
                           n39);
   U82 : NAND3_X1 port map( A1 => n15, A2 => n18, A3 => INS_IN(28), ZN => 
                           n24_port);
   U83 : NAND3_X1 port map( A1 => n10, A2 => n13, A3 => n63, ZN => n34);
   U84 : NAND3_X1 port map( A1 => n16, A2 => n17, A3 => INS_IN(28), ZN => n36);
   U18 : INV_X1 port map( A => n25_port, ZN => n10);
   U19 : NAND2_X1 port map( A1 => n12, A2 => n11, ZN => n25_port);
   U20 : AOI21_X1 port map( B1 => n40, B2 => n41, A => Bubble, ZN => N25);
   U21 : AOI211_X1 port map( C1 => n14, C2 => n10, A => n38, B => n48, ZN => 
                           n40);
   U22 : AOI221_X1 port map( B1 => n42, B2 => n5, C1 => n16, C2 => n43, A => 
                           n44, ZN => n41);
   U23 : INV_X1 port map( A => n47, ZN => n5);
   U24 : AOI21_X1 port map( B1 => n28, B2 => n29, A => Bubble, ZN => N26);
   U25 : AOI21_X1 port map( B1 => n20, B2 => n6, A => n38, ZN => n28);
   U26 : NOR3_X1 port map( A1 => n30, A2 => n31, A3 => n32, ZN => n29);
   U27 : AOI21_X1 port map( B1 => n36, B2 => n37, A => n26_port, ZN => n30);
   U28 : INV_X1 port map( A => n36, ZN => n14);
   U29 : INV_X1 port map( A => n27_port, ZN => n16);
   U30 : OR2_X1 port map( A1 => n49, A2 => n50, ZN => n38);
   U31 : INV_X1 port map( A => n52, ZN => n3);
   U32 : INV_X1 port map( A => n51, ZN => n8);
   U33 : NAND2_X1 port map( A1 => n16, A2 => n10, ZN => n58);
   U34 : OR3_X1 port map( A1 => INS_IN(0), A2 => INS_IN(1), A3 => n34, ZN => 
                           n59);
   U35 : NOR4_X1 port map( A1 => INS_IN(6), A2 => INS_IN(4), A3 => INS_IN(10), 
                           A4 => n62, ZN => n51);
   U36 : OR3_X1 port map( A1 => INS_IN(9), A2 => INS_IN(8), A3 => INS_IN(7), ZN
                           => n62);
   U37 : NAND2_X1 port map( A1 => INS_IN(27), A2 => n11, ZN => n46);
   U38 : NOR3_X1 port map( A1 => INS_IN(29), A2 => INS_IN(31), A3 => INS_IN(30)
                           , ZN => n63);
   U39 : NOR4_X1 port map( A1 => n2, A2 => n39, A3 => n34, A4 => INS_IN(1), ZN 
                           => n20);
   U40 : NOR4_X1 port map( A1 => n6, A2 => INS_IN(0), A3 => INS_IN(3), A4 => 
                           INS_IN(5), ZN => n52);
   U41 : NOR4_X1 port map( A1 => n33, A2 => n34, A3 => n6, A4 => n35, ZN => n32
                           );
   U42 : NOR4_X1 port map( A1 => INS_IN(1), A2 => n4, A3 => n34, A4 => n6, ZN 
                           => n44);
   U43 : INV_X1 port map( A => n45, ZN => n4);
   U44 : OAI21_X1 port map( B1 => n35, B2 => INS_IN(0), A => n39, ZN => n45);
   U45 : NOR3_X1 port map( A1 => n34, A2 => INS_IN(0), A3 => n35, ZN => n42);
   U46 : INV_X1 port map( A => INS_IN(3), ZN => n7);
   U47 : NOR3_X1 port map( A1 => n36, A2 => INS_IN(26), A3 => n12, ZN => n31);
   U48 : INV_X1 port map( A => INS_IN(2), ZN => n6);
   U49 : INV_X1 port map( A => INS_IN(30), ZN => n17);
   U50 : AOI22_X1 port map( A1 => n15, A2 => n18, B1 => INS_IN(31), B2 => n17, 
                           ZN => n56);
   U51 : NAND2_X1 port map( A1 => INS_IN(26), A2 => n12, ZN => n26_port);
   U52 : INV_X1 port map( A => INS_IN(27), ZN => n12);
   U53 : AOI21_X1 port map( B1 => n53, B2 => n54, A => Bubble, ZN => N24);
   U54 : AOI211_X1 port map( C1 => n14, C2 => n10, A => n49, B => n23, ZN => 
                           n53);
   U55 : AOI221_X1 port map( B1 => n42, B2 => n47, C1 => n55, C2 => n13, A => 
                           n31, ZN => n54);
   U56 : INV_X1 port map( A => INS_IN(28), ZN => n13);
   U57 : NAND2_X1 port map( A1 => INS_IN(29), A2 => n18, ZN => n27_port);
   U58 : OR2_X1 port map( A1 => n48, A2 => n1, ZN => n23);
   U59 : NOR3_X1 port map( A1 => n26_port, A2 => INS_IN(30), A3 => n24_port, ZN
                           => n1);
   U60 : NAND2_X1 port map( A1 => INS_IN(1), A2 => n6, ZN => n47);
   U61 : INV_X1 port map( A => INS_IN(31), ZN => n18);
   U62 : INV_X1 port map( A => INS_IN(26), ZN => n11);
   U63 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => n49);
   U64 : OR4_X1 port map( A1 => n12, A2 => n24_port, A3 => n17, A4 => 
                           INS_IN(26), ZN => n61);
   U65 : NAND4_X1 port map( A1 => INS_IN(1), A2 => n52, A3 => n9, A4 => n51, ZN
                           => n60);
   U66 : INV_X1 port map( A => n34, ZN => n9);
   U67 : NOR2_X1 port map( A1 => Bubble, A2 => n19, ZN => N27);
   U68 : NOR4_X1 port map( A1 => n20, A2 => n21, A3 => n22, A4 => n23, ZN => 
                           n19);
   U69 : NOR3_X1 port map( A1 => n26_port, A2 => n27_port, A3 => n17, ZN => n21
                           );
   U70 : NOR3_X1 port map( A1 => n24_port, A2 => INS_IN(30), A3 => n25_port, ZN
                           => n22);
   U71 : INV_X1 port map( A => INS_IN(0), ZN => n2);
   U72 : INV_X1 port map( A => INS_IN(29), ZN => n15);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Datapath is

   port( CLK, RST : in std_logic;  INS_IN, DATA_IN : in std_logic_vector (31 
         downto 0);  REG_LATCH_EN, RD1, RD2, MUX_A_SEL : in std_logic;  
         MUX_B_SEL : in std_logic_vector (1 downto 0);  ALU_OPC : in 
         std_logic_vector (0 to 3);  ALU_OUTREG_EN : in std_logic;  JUMP_TYPE :
         in std_logic_vector (1 downto 0);  DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, 
         RF_WE, DRAM_EN_IN, WB_MUX_SEL : in std_logic;  INS_OUT, IRAM_ADDR_OUT,
         DRAM_ADDR_OUT, DATA_OUT : out std_logic_vector (31 downto 0);  
         DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble_out : out std_logic);

end Datapath;

architecture SYN_struct of Datapath is

   component HazardDetection
      port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : in std_logic_vector
            (4 downto 0);  DRAM_R : in std_logic;  INS_IN, PC_IN : in 
            std_logic_vector (31 downto 0);  Bubble : out std_logic;  
            HDU_INS_OUT, HDU_PC_OUT, HDU_NPC_OUT : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Writeback
      port( WB_MUX_SEL : in std_logic;  DATA_IN, ALU_RES_IN : in 
            std_logic_vector (31 downto 0);  ADD_WR_IN : in std_logic_vector (4
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0);  
            ADD_WR_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component ff_2
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Memory
      port( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, DRAM_EN_IN : in 
            std_logic;  PC_SEL : in std_logic_vector (1 downto 0);  NPC_IN, 
            NPC_ABS, NPC_REL, ALU_RES_IN, B_IN : in std_logic_vector (31 downto
            0);  ADD_WR_IN : in std_logic_vector (4 downto 0);  DRAM_DATA_IN : 
            in std_logic_vector (31 downto 0);  PC_OUT : out std_logic_vector 
            (31 downto 0);  DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT : out std_logic
            ;  DRAM_ADDR_OUT, DRAM_DATA_OUT, DATA_OUT, ALU_RES_OUT, OP_MEM : 
            out std_logic_vector (31 downto 0);  ADD_WR_MEM, ADD_WR_OUT : out 
            std_logic_vector (4 downto 0));
   end component;
   
   component ff_0
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Execute
      port( CLK, RST, MUX_A_SEL : in std_logic;  MUX_B_SEL : in 
            std_logic_vector (1 downto 0);  ALU_OPC : in std_logic_vector (0 to
            3);  ALU_OUTREG_EN : in std_logic;  JUMP_TYPE : in std_logic_vector
            (1 downto 0);  PC_IN, A_IN, B_IN, IMM_IN : in std_logic_vector (31 
            downto 0);  ADD_WR_IN, ADD_RS1_IN, ADD_RS2_IN, ADD_WR_MEM, 
            ADD_WR_WB : in std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB 
            : in std_logic;  OP_MEM, OP_WB : in std_logic_vector (31 downto 0);
            PC_SEL : out std_logic_vector (1 downto 0);  ZERO_FLAG : out 
            std_logic;  NPC_ABS, NPC_REL, ALU_RES, B_OUT : out std_logic_vector
            (31 downto 0);  ADD_WR_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component Decode
      port( CLK, RST, REG_LATCH_EN, RD1, RD2, RF_WE, ZERO_FLAG : in std_logic; 
            PC_IN, INS_IN : in std_logic_vector (31 downto 0);  ADD_WR : in 
            std_logic_vector (4 downto 0);  DATA_WR_IN : in std_logic_vector 
            (31 downto 0);  PC_OUT, A_OUT, B_OUT, IMM_OUT : out 
            std_logic_vector (31 downto 0);  ADD_RS1_HDU, ADD_RS2_HDU, 
            ADD_WR_OUT, ADD_RS1_OUT, ADD_RS2_OUT : out std_logic_vector (4 
            downto 0));
   end component;
   
   component Fetch
      port( CLK, RST, ZERO_FLAG : in std_logic;  PC_EXT, INS_IN : in 
            std_logic_vector (31 downto 0);  Bubble_in : in std_logic;  
            HDU_INS_IN, HDU_PC_IN, HDU_NPC_IN : in std_logic_vector (31 downto 
            0);  PC_OUT, ADDR_OUT, NPC_OUT, INS_OUT : out std_logic_vector (31 
            downto 0));
   end component;
   
   signal X_Logic1_port, INS_OUT_31_port, INS_OUT_30_port, INS_OUT_29_port, 
      INS_OUT_28_port, INS_OUT_27_port, INS_OUT_26_port, INS_OUT_25_port, 
      INS_OUT_24_port, INS_OUT_23_port, INS_OUT_22_port, INS_OUT_21_port, 
      INS_OUT_20_port, INS_OUT_19_port, INS_OUT_18_port, INS_OUT_17_port, 
      INS_OUT_16_port, INS_OUT_15_port, INS_OUT_14_port, INS_OUT_13_port, 
      INS_OUT_12_port, INS_OUT_11_port, INS_OUT_10_port, INS_OUT_9_port, 
      INS_OUT_8_port, INS_OUT_7_port, INS_OUT_6_port, INS_OUT_5_port, 
      INS_OUT_4_port, INS_OUT_3_port, INS_OUT_2_port, INS_OUT_1_port, 
      INS_OUT_0_port, Bubble_out_port, ZERO_FLAG_EX, PC_MEM_OUT_31_port, 
      PC_MEM_OUT_30_port, PC_MEM_OUT_29_port, PC_MEM_OUT_28_port, 
      PC_MEM_OUT_27_port, PC_MEM_OUT_26_port, PC_MEM_OUT_25_port, 
      PC_MEM_OUT_24_port, PC_MEM_OUT_23_port, PC_MEM_OUT_22_port, 
      PC_MEM_OUT_21_port, PC_MEM_OUT_20_port, PC_MEM_OUT_19_port, 
      PC_MEM_OUT_18_port, PC_MEM_OUT_17_port, PC_MEM_OUT_16_port, 
      PC_MEM_OUT_15_port, PC_MEM_OUT_14_port, PC_MEM_OUT_13_port, 
      PC_MEM_OUT_12_port, PC_MEM_OUT_11_port, PC_MEM_OUT_10_port, 
      PC_MEM_OUT_9_port, PC_MEM_OUT_8_port, PC_MEM_OUT_7_port, 
      PC_MEM_OUT_6_port, PC_MEM_OUT_5_port, PC_MEM_OUT_4_port, 
      PC_MEM_OUT_3_port, PC_MEM_OUT_2_port, PC_MEM_OUT_1_port, 
      PC_MEM_OUT_0_port, sig_HDU_INS_OUT_31_port, sig_HDU_INS_OUT_30_port, 
      sig_HDU_INS_OUT_29_port, sig_HDU_INS_OUT_28_port, sig_HDU_INS_OUT_27_port
      , sig_HDU_INS_OUT_26_port, sig_HDU_INS_OUT_25_port, 
      sig_HDU_INS_OUT_24_port, sig_HDU_INS_OUT_23_port, sig_HDU_INS_OUT_22_port
      , sig_HDU_INS_OUT_21_port, sig_HDU_INS_OUT_20_port, 
      sig_HDU_INS_OUT_19_port, sig_HDU_INS_OUT_18_port, sig_HDU_INS_OUT_17_port
      , sig_HDU_INS_OUT_16_port, sig_HDU_INS_OUT_15_port, 
      sig_HDU_INS_OUT_14_port, sig_HDU_INS_OUT_13_port, sig_HDU_INS_OUT_12_port
      , sig_HDU_INS_OUT_11_port, sig_HDU_INS_OUT_10_port, 
      sig_HDU_INS_OUT_9_port, sig_HDU_INS_OUT_8_port, sig_HDU_INS_OUT_7_port, 
      sig_HDU_INS_OUT_6_port, sig_HDU_INS_OUT_5_port, sig_HDU_INS_OUT_4_port, 
      sig_HDU_INS_OUT_3_port, sig_HDU_INS_OUT_2_port, sig_HDU_INS_OUT_1_port, 
      sig_HDU_INS_OUT_0_port, sig_HDU_PC_OUT_31_port, sig_HDU_PC_OUT_30_port, 
      sig_HDU_PC_OUT_29_port, sig_HDU_PC_OUT_28_port, sig_HDU_PC_OUT_27_port, 
      sig_HDU_PC_OUT_26_port, sig_HDU_PC_OUT_25_port, sig_HDU_PC_OUT_24_port, 
      sig_HDU_PC_OUT_23_port, sig_HDU_PC_OUT_22_port, sig_HDU_PC_OUT_21_port, 
      sig_HDU_PC_OUT_20_port, sig_HDU_PC_OUT_19_port, sig_HDU_PC_OUT_18_port, 
      sig_HDU_PC_OUT_17_port, sig_HDU_PC_OUT_16_port, sig_HDU_PC_OUT_15_port, 
      sig_HDU_PC_OUT_14_port, sig_HDU_PC_OUT_13_port, sig_HDU_PC_OUT_12_port, 
      sig_HDU_PC_OUT_11_port, sig_HDU_PC_OUT_10_port, sig_HDU_PC_OUT_9_port, 
      sig_HDU_PC_OUT_8_port, sig_HDU_PC_OUT_7_port, sig_HDU_PC_OUT_6_port, 
      sig_HDU_PC_OUT_5_port, sig_HDU_PC_OUT_4_port, sig_HDU_PC_OUT_3_port, 
      sig_HDU_PC_OUT_2_port, sig_HDU_PC_OUT_1_port, sig_HDU_PC_OUT_0_port, 
      sig_HDU_NPC_OUT_31_port, sig_HDU_NPC_OUT_30_port, sig_HDU_NPC_OUT_29_port
      , sig_HDU_NPC_OUT_28_port, sig_HDU_NPC_OUT_27_port, 
      sig_HDU_NPC_OUT_26_port, sig_HDU_NPC_OUT_25_port, sig_HDU_NPC_OUT_24_port
      , sig_HDU_NPC_OUT_23_port, sig_HDU_NPC_OUT_22_port, 
      sig_HDU_NPC_OUT_21_port, sig_HDU_NPC_OUT_20_port, sig_HDU_NPC_OUT_19_port
      , sig_HDU_NPC_OUT_18_port, sig_HDU_NPC_OUT_17_port, 
      sig_HDU_NPC_OUT_16_port, sig_HDU_NPC_OUT_15_port, sig_HDU_NPC_OUT_14_port
      , sig_HDU_NPC_OUT_13_port, sig_HDU_NPC_OUT_12_port, 
      sig_HDU_NPC_OUT_11_port, sig_HDU_NPC_OUT_10_port, sig_HDU_NPC_OUT_9_port,
      sig_HDU_NPC_OUT_8_port, sig_HDU_NPC_OUT_7_port, sig_HDU_NPC_OUT_6_port, 
      sig_HDU_NPC_OUT_5_port, sig_HDU_NPC_OUT_4_port, sig_HDU_NPC_OUT_3_port, 
      sig_HDU_NPC_OUT_2_port, sig_HDU_NPC_OUT_1_port, sig_HDU_NPC_OUT_0_port, 
      PC_FETCH_OUT_31_port, PC_FETCH_OUT_30_port, PC_FETCH_OUT_29_port, 
      PC_FETCH_OUT_28_port, PC_FETCH_OUT_27_port, PC_FETCH_OUT_26_port, 
      PC_FETCH_OUT_25_port, PC_FETCH_OUT_24_port, PC_FETCH_OUT_23_port, 
      PC_FETCH_OUT_22_port, PC_FETCH_OUT_21_port, PC_FETCH_OUT_20_port, 
      PC_FETCH_OUT_19_port, PC_FETCH_OUT_18_port, PC_FETCH_OUT_17_port, 
      PC_FETCH_OUT_16_port, PC_FETCH_OUT_15_port, PC_FETCH_OUT_14_port, 
      PC_FETCH_OUT_13_port, PC_FETCH_OUT_12_port, PC_FETCH_OUT_11_port, 
      PC_FETCH_OUT_10_port, PC_FETCH_OUT_9_port, PC_FETCH_OUT_8_port, 
      PC_FETCH_OUT_7_port, PC_FETCH_OUT_6_port, PC_FETCH_OUT_5_port, 
      PC_FETCH_OUT_4_port, PC_FETCH_OUT_3_port, PC_FETCH_OUT_2_port, 
      PC_FETCH_OUT_1_port, PC_FETCH_OUT_0_port, NPC_FETCH_OUT_31_port, 
      NPC_FETCH_OUT_30_port, NPC_FETCH_OUT_29_port, NPC_FETCH_OUT_28_port, 
      NPC_FETCH_OUT_27_port, NPC_FETCH_OUT_26_port, NPC_FETCH_OUT_25_port, 
      NPC_FETCH_OUT_24_port, NPC_FETCH_OUT_23_port, NPC_FETCH_OUT_22_port, 
      NPC_FETCH_OUT_21_port, NPC_FETCH_OUT_20_port, NPC_FETCH_OUT_19_port, 
      NPC_FETCH_OUT_18_port, NPC_FETCH_OUT_17_port, NPC_FETCH_OUT_16_port, 
      NPC_FETCH_OUT_15_port, NPC_FETCH_OUT_14_port, NPC_FETCH_OUT_13_port, 
      NPC_FETCH_OUT_12_port, NPC_FETCH_OUT_11_port, NPC_FETCH_OUT_10_port, 
      NPC_FETCH_OUT_9_port, NPC_FETCH_OUT_8_port, NPC_FETCH_OUT_7_port, 
      NPC_FETCH_OUT_6_port, NPC_FETCH_OUT_5_port, NPC_FETCH_OUT_4_port, 
      NPC_FETCH_OUT_3_port, NPC_FETCH_OUT_2_port, NPC_FETCH_OUT_1_port, 
      NPC_FETCH_OUT_0_port, RF_WE_WB, ADD_WR_WB_4_port, ADD_WR_WB_3_port, 
      ADD_WR_WB_2_port, ADD_WR_WB_1_port, ADD_WR_WB_0_port, OP_WB_31_port, 
      OP_WB_30_port, OP_WB_29_port, OP_WB_28_port, OP_WB_27_port, OP_WB_26_port
      , OP_WB_25_port, OP_WB_24_port, OP_WB_23_port, OP_WB_22_port, 
      OP_WB_21_port, OP_WB_20_port, OP_WB_19_port, OP_WB_18_port, OP_WB_17_port
      , OP_WB_16_port, OP_WB_15_port, OP_WB_14_port, OP_WB_13_port, 
      OP_WB_12_port, OP_WB_11_port, OP_WB_10_port, OP_WB_9_port, OP_WB_8_port, 
      OP_WB_7_port, OP_WB_6_port, OP_WB_5_port, OP_WB_4_port, OP_WB_3_port, 
      OP_WB_2_port, OP_WB_1_port, OP_WB_0_port, PC_DECODE_OUT_31_port, 
      PC_DECODE_OUT_30_port, PC_DECODE_OUT_29_port, PC_DECODE_OUT_28_port, 
      PC_DECODE_OUT_27_port, PC_DECODE_OUT_26_port, PC_DECODE_OUT_25_port, 
      PC_DECODE_OUT_24_port, PC_DECODE_OUT_23_port, PC_DECODE_OUT_22_port, 
      PC_DECODE_OUT_21_port, PC_DECODE_OUT_20_port, PC_DECODE_OUT_19_port, 
      PC_DECODE_OUT_18_port, PC_DECODE_OUT_17_port, PC_DECODE_OUT_16_port, 
      PC_DECODE_OUT_15_port, PC_DECODE_OUT_14_port, PC_DECODE_OUT_13_port, 
      PC_DECODE_OUT_12_port, PC_DECODE_OUT_11_port, PC_DECODE_OUT_10_port, 
      PC_DECODE_OUT_9_port, PC_DECODE_OUT_8_port, PC_DECODE_OUT_7_port, 
      PC_DECODE_OUT_6_port, PC_DECODE_OUT_5_port, PC_DECODE_OUT_4_port, 
      PC_DECODE_OUT_3_port, PC_DECODE_OUT_2_port, PC_DECODE_OUT_1_port, 
      PC_DECODE_OUT_0_port, A_DECODE_OUT_31_port, A_DECODE_OUT_30_port, 
      A_DECODE_OUT_29_port, A_DECODE_OUT_28_port, A_DECODE_OUT_27_port, 
      A_DECODE_OUT_26_port, A_DECODE_OUT_25_port, A_DECODE_OUT_24_port, 
      A_DECODE_OUT_23_port, A_DECODE_OUT_22_port, A_DECODE_OUT_21_port, 
      A_DECODE_OUT_20_port, A_DECODE_OUT_19_port, A_DECODE_OUT_18_port, 
      A_DECODE_OUT_17_port, A_DECODE_OUT_16_port, A_DECODE_OUT_15_port, 
      A_DECODE_OUT_14_port, A_DECODE_OUT_13_port, A_DECODE_OUT_12_port, 
      A_DECODE_OUT_11_port, A_DECODE_OUT_10_port, A_DECODE_OUT_9_port, 
      A_DECODE_OUT_8_port, A_DECODE_OUT_7_port, A_DECODE_OUT_6_port, 
      A_DECODE_OUT_5_port, A_DECODE_OUT_4_port, A_DECODE_OUT_3_port, 
      A_DECODE_OUT_2_port, A_DECODE_OUT_1_port, A_DECODE_OUT_0_port, 
      B_DECODE_OUT_31_port, B_DECODE_OUT_30_port, B_DECODE_OUT_29_port, 
      B_DECODE_OUT_28_port, B_DECODE_OUT_27_port, B_DECODE_OUT_26_port, 
      B_DECODE_OUT_25_port, B_DECODE_OUT_24_port, B_DECODE_OUT_23_port, 
      B_DECODE_OUT_22_port, B_DECODE_OUT_21_port, B_DECODE_OUT_20_port, 
      B_DECODE_OUT_19_port, B_DECODE_OUT_18_port, B_DECODE_OUT_17_port, 
      B_DECODE_OUT_16_port, B_DECODE_OUT_15_port, B_DECODE_OUT_14_port, 
      B_DECODE_OUT_13_port, B_DECODE_OUT_12_port, B_DECODE_OUT_11_port, 
      B_DECODE_OUT_10_port, B_DECODE_OUT_9_port, B_DECODE_OUT_8_port, 
      B_DECODE_OUT_7_port, B_DECODE_OUT_6_port, B_DECODE_OUT_5_port, 
      B_DECODE_OUT_4_port, B_DECODE_OUT_3_port, B_DECODE_OUT_2_port, 
      B_DECODE_OUT_1_port, B_DECODE_OUT_0_port, IMM_DECODE_OUT_31_port, 
      IMM_DECODE_OUT_30_port, IMM_DECODE_OUT_29_port, IMM_DECODE_OUT_28_port, 
      IMM_DECODE_OUT_27_port, IMM_DECODE_OUT_26_port, IMM_DECODE_OUT_25_port, 
      IMM_DECODE_OUT_24_port, IMM_DECODE_OUT_23_port, IMM_DECODE_OUT_22_port, 
      IMM_DECODE_OUT_21_port, IMM_DECODE_OUT_20_port, IMM_DECODE_OUT_19_port, 
      IMM_DECODE_OUT_18_port, IMM_DECODE_OUT_17_port, IMM_DECODE_OUT_16_port, 
      IMM_DECODE_OUT_15_port, IMM_DECODE_OUT_14_port, IMM_DECODE_OUT_13_port, 
      IMM_DECODE_OUT_12_port, IMM_DECODE_OUT_11_port, IMM_DECODE_OUT_10_port, 
      IMM_DECODE_OUT_9_port, IMM_DECODE_OUT_8_port, IMM_DECODE_OUT_7_port, 
      IMM_DECODE_OUT_6_port, IMM_DECODE_OUT_5_port, IMM_DECODE_OUT_4_port, 
      IMM_DECODE_OUT_3_port, IMM_DECODE_OUT_2_port, IMM_DECODE_OUT_1_port, 
      IMM_DECODE_OUT_0_port, ADD_RS1_HDU_4_port, ADD_RS1_HDU_3_port, 
      ADD_RS1_HDU_2_port, ADD_RS1_HDU_1_port, ADD_RS1_HDU_0_port, 
      ADD_RS2_HDU_4_port, ADD_RS2_HDU_3_port, ADD_RS2_HDU_2_port, 
      ADD_RS2_HDU_1_port, ADD_RS2_HDU_0_port, ADD_WR_DECODE_OUT_4_port, 
      ADD_WR_DECODE_OUT_3_port, ADD_WR_DECODE_OUT_2_port, 
      ADD_WR_DECODE_OUT_1_port, ADD_WR_DECODE_OUT_0_port, 
      ADD_RS1_DECODE_OUT_4_port, ADD_RS1_DECODE_OUT_3_port, 
      ADD_RS1_DECODE_OUT_2_port, ADD_RS1_DECODE_OUT_1_port, 
      ADD_RS1_DECODE_OUT_0_port, ADD_RS2_DECODE_OUT_4_port, 
      ADD_RS2_DECODE_OUT_3_port, ADD_RS2_DECODE_OUT_2_port, 
      ADD_RS2_DECODE_OUT_1_port, ADD_RS2_DECODE_OUT_0_port, ADD_WR_MEM_4_port, 
      ADD_WR_MEM_3_port, ADD_WR_MEM_2_port, ADD_WR_MEM_1_port, 
      ADD_WR_MEM_0_port, OP_MEM_31_port, OP_MEM_30_port, OP_MEM_29_port, 
      OP_MEM_28_port, OP_MEM_27_port, OP_MEM_26_port, OP_MEM_25_port, 
      OP_MEM_24_port, OP_MEM_23_port, OP_MEM_22_port, OP_MEM_21_port, 
      OP_MEM_20_port, OP_MEM_19_port, OP_MEM_18_port, OP_MEM_17_port, 
      OP_MEM_16_port, OP_MEM_15_port, OP_MEM_14_port, OP_MEM_13_port, 
      OP_MEM_12_port, OP_MEM_11_port, OP_MEM_10_port, OP_MEM_9_port, 
      OP_MEM_8_port, OP_MEM_7_port, OP_MEM_6_port, OP_MEM_5_port, OP_MEM_4_port
      , OP_MEM_3_port, OP_MEM_2_port, OP_MEM_1_port, OP_MEM_0_port, 
      PC_SEL_EX_1_port, PC_SEL_EX_0_port, NPC_ABS_EX_31_port, 
      NPC_ABS_EX_30_port, NPC_ABS_EX_29_port, NPC_ABS_EX_28_port, 
      NPC_ABS_EX_27_port, NPC_ABS_EX_26_port, NPC_ABS_EX_25_port, 
      NPC_ABS_EX_24_port, NPC_ABS_EX_23_port, NPC_ABS_EX_22_port, 
      NPC_ABS_EX_21_port, NPC_ABS_EX_20_port, NPC_ABS_EX_19_port, 
      NPC_ABS_EX_18_port, NPC_ABS_EX_17_port, NPC_ABS_EX_16_port, 
      NPC_ABS_EX_15_port, NPC_ABS_EX_14_port, NPC_ABS_EX_13_port, 
      NPC_ABS_EX_12_port, NPC_ABS_EX_11_port, NPC_ABS_EX_10_port, 
      NPC_ABS_EX_9_port, NPC_ABS_EX_8_port, NPC_ABS_EX_7_port, 
      NPC_ABS_EX_6_port, NPC_ABS_EX_5_port, NPC_ABS_EX_4_port, 
      NPC_ABS_EX_3_port, NPC_ABS_EX_2_port, NPC_ABS_EX_1_port, 
      NPC_ABS_EX_0_port, NPC_REL_EX_31_port, NPC_REL_EX_30_port, 
      NPC_REL_EX_29_port, NPC_REL_EX_28_port, NPC_REL_EX_27_port, 
      NPC_REL_EX_26_port, NPC_REL_EX_25_port, NPC_REL_EX_24_port, 
      NPC_REL_EX_23_port, NPC_REL_EX_22_port, NPC_REL_EX_21_port, 
      NPC_REL_EX_20_port, NPC_REL_EX_19_port, NPC_REL_EX_18_port, 
      NPC_REL_EX_17_port, NPC_REL_EX_16_port, NPC_REL_EX_15_port, 
      NPC_REL_EX_14_port, NPC_REL_EX_13_port, NPC_REL_EX_12_port, 
      NPC_REL_EX_11_port, NPC_REL_EX_10_port, NPC_REL_EX_9_port, 
      NPC_REL_EX_8_port, NPC_REL_EX_7_port, NPC_REL_EX_6_port, 
      NPC_REL_EX_5_port, NPC_REL_EX_4_port, NPC_REL_EX_3_port, 
      NPC_REL_EX_2_port, NPC_REL_EX_1_port, NPC_REL_EX_0_port, 
      ALU_RES_EX_31_port, ALU_RES_EX_30_port, ALU_RES_EX_29_port, 
      ALU_RES_EX_28_port, ALU_RES_EX_27_port, ALU_RES_EX_26_port, 
      ALU_RES_EX_25_port, ALU_RES_EX_24_port, ALU_RES_EX_23_port, 
      ALU_RES_EX_22_port, ALU_RES_EX_21_port, ALU_RES_EX_20_port, 
      ALU_RES_EX_19_port, ALU_RES_EX_18_port, ALU_RES_EX_17_port, 
      ALU_RES_EX_16_port, ALU_RES_EX_15_port, ALU_RES_EX_14_port, 
      ALU_RES_EX_13_port, ALU_RES_EX_12_port, ALU_RES_EX_11_port, 
      ALU_RES_EX_10_port, ALU_RES_EX_9_port, ALU_RES_EX_8_port, 
      ALU_RES_EX_7_port, ALU_RES_EX_6_port, ALU_RES_EX_5_port, 
      ALU_RES_EX_4_port, ALU_RES_EX_3_port, ALU_RES_EX_2_port, 
      ALU_RES_EX_1_port, ALU_RES_EX_0_port, B_EX_OUT_31_port, B_EX_OUT_30_port,
      B_EX_OUT_29_port, B_EX_OUT_28_port, B_EX_OUT_27_port, B_EX_OUT_26_port, 
      B_EX_OUT_25_port, B_EX_OUT_24_port, B_EX_OUT_23_port, B_EX_OUT_22_port, 
      B_EX_OUT_21_port, B_EX_OUT_20_port, B_EX_OUT_19_port, B_EX_OUT_18_port, 
      B_EX_OUT_17_port, B_EX_OUT_16_port, B_EX_OUT_15_port, B_EX_OUT_14_port, 
      B_EX_OUT_13_port, B_EX_OUT_12_port, B_EX_OUT_11_port, B_EX_OUT_10_port, 
      B_EX_OUT_9_port, B_EX_OUT_8_port, B_EX_OUT_7_port, B_EX_OUT_6_port, 
      B_EX_OUT_5_port, B_EX_OUT_4_port, B_EX_OUT_3_port, B_EX_OUT_2_port, 
      B_EX_OUT_1_port, B_EX_OUT_0_port, ADD_WR_EX_OUT_4_port, 
      ADD_WR_EX_OUT_3_port, ADD_WR_EX_OUT_2_port, ADD_WR_EX_OUT_1_port, 
      ADD_WR_EX_OUT_0_port, DRAM_R_MEM, DATA_MEM_OUT_31_port, 
      DATA_MEM_OUT_30_port, DATA_MEM_OUT_29_port, DATA_MEM_OUT_28_port, 
      DATA_MEM_OUT_27_port, DATA_MEM_OUT_26_port, DATA_MEM_OUT_25_port, 
      DATA_MEM_OUT_24_port, DATA_MEM_OUT_23_port, DATA_MEM_OUT_22_port, 
      DATA_MEM_OUT_21_port, DATA_MEM_OUT_20_port, DATA_MEM_OUT_19_port, 
      DATA_MEM_OUT_18_port, DATA_MEM_OUT_17_port, DATA_MEM_OUT_16_port, 
      DATA_MEM_OUT_15_port, DATA_MEM_OUT_14_port, DATA_MEM_OUT_13_port, 
      DATA_MEM_OUT_12_port, DATA_MEM_OUT_11_port, DATA_MEM_OUT_10_port, 
      DATA_MEM_OUT_9_port, DATA_MEM_OUT_8_port, DATA_MEM_OUT_7_port, 
      DATA_MEM_OUT_6_port, DATA_MEM_OUT_5_port, DATA_MEM_OUT_4_port, 
      DATA_MEM_OUT_3_port, DATA_MEM_OUT_2_port, DATA_MEM_OUT_1_port, 
      DATA_MEM_OUT_0_port, ALU_RES_MEM_31_port, ALU_RES_MEM_30_port, 
      ALU_RES_MEM_29_port, ALU_RES_MEM_28_port, ALU_RES_MEM_27_port, 
      ALU_RES_MEM_26_port, ALU_RES_MEM_25_port, ALU_RES_MEM_24_port, 
      ALU_RES_MEM_23_port, ALU_RES_MEM_22_port, ALU_RES_MEM_21_port, 
      ALU_RES_MEM_20_port, ALU_RES_MEM_19_port, ALU_RES_MEM_18_port, 
      ALU_RES_MEM_17_port, ALU_RES_MEM_16_port, ALU_RES_MEM_15_port, 
      ALU_RES_MEM_14_port, ALU_RES_MEM_13_port, ALU_RES_MEM_12_port, 
      ALU_RES_MEM_11_port, ALU_RES_MEM_10_port, ALU_RES_MEM_9_port, 
      ALU_RES_MEM_8_port, ALU_RES_MEM_7_port, ALU_RES_MEM_6_port, 
      ALU_RES_MEM_5_port, ALU_RES_MEM_4_port, ALU_RES_MEM_3_port, 
      ALU_RES_MEM_2_port, ALU_RES_MEM_1_port, ALU_RES_MEM_0_port, 
      ADD_WR_MEM_OUT_4_port, ADD_WR_MEM_OUT_3_port, ADD_WR_MEM_OUT_2_port, 
      ADD_WR_MEM_OUT_1_port, ADD_WR_MEM_OUT_0_port : std_logic;

begin
   INS_OUT <= ( INS_OUT_31_port, INS_OUT_30_port, INS_OUT_29_port, 
      INS_OUT_28_port, INS_OUT_27_port, INS_OUT_26_port, INS_OUT_25_port, 
      INS_OUT_24_port, INS_OUT_23_port, INS_OUT_22_port, INS_OUT_21_port, 
      INS_OUT_20_port, INS_OUT_19_port, INS_OUT_18_port, INS_OUT_17_port, 
      INS_OUT_16_port, INS_OUT_15_port, INS_OUT_14_port, INS_OUT_13_port, 
      INS_OUT_12_port, INS_OUT_11_port, INS_OUT_10_port, INS_OUT_9_port, 
      INS_OUT_8_port, INS_OUT_7_port, INS_OUT_6_port, INS_OUT_5_port, 
      INS_OUT_4_port, INS_OUT_3_port, INS_OUT_2_port, INS_OUT_1_port, 
      INS_OUT_0_port );
   Bubble_out <= Bubble_out_port;
   
   X_Logic1_port <= '1';
   FetchStage : Fetch port map( CLK => CLK, RST => RST, ZERO_FLAG => 
                           ZERO_FLAG_EX, PC_EXT(31) => PC_MEM_OUT_31_port, 
                           PC_EXT(30) => PC_MEM_OUT_30_port, PC_EXT(29) => 
                           PC_MEM_OUT_29_port, PC_EXT(28) => PC_MEM_OUT_28_port
                           , PC_EXT(27) => PC_MEM_OUT_27_port, PC_EXT(26) => 
                           PC_MEM_OUT_26_port, PC_EXT(25) => PC_MEM_OUT_25_port
                           , PC_EXT(24) => PC_MEM_OUT_24_port, PC_EXT(23) => 
                           PC_MEM_OUT_23_port, PC_EXT(22) => PC_MEM_OUT_22_port
                           , PC_EXT(21) => PC_MEM_OUT_21_port, PC_EXT(20) => 
                           PC_MEM_OUT_20_port, PC_EXT(19) => PC_MEM_OUT_19_port
                           , PC_EXT(18) => PC_MEM_OUT_18_port, PC_EXT(17) => 
                           PC_MEM_OUT_17_port, PC_EXT(16) => PC_MEM_OUT_16_port
                           , PC_EXT(15) => PC_MEM_OUT_15_port, PC_EXT(14) => 
                           PC_MEM_OUT_14_port, PC_EXT(13) => PC_MEM_OUT_13_port
                           , PC_EXT(12) => PC_MEM_OUT_12_port, PC_EXT(11) => 
                           PC_MEM_OUT_11_port, PC_EXT(10) => PC_MEM_OUT_10_port
                           , PC_EXT(9) => PC_MEM_OUT_9_port, PC_EXT(8) => 
                           PC_MEM_OUT_8_port, PC_EXT(7) => PC_MEM_OUT_7_port, 
                           PC_EXT(6) => PC_MEM_OUT_6_port, PC_EXT(5) => 
                           PC_MEM_OUT_5_port, PC_EXT(4) => PC_MEM_OUT_4_port, 
                           PC_EXT(3) => PC_MEM_OUT_3_port, PC_EXT(2) => 
                           PC_MEM_OUT_2_port, PC_EXT(1) => PC_MEM_OUT_1_port, 
                           PC_EXT(0) => PC_MEM_OUT_0_port, INS_IN(31) => 
                           INS_IN(31), INS_IN(30) => INS_IN(30), INS_IN(29) => 
                           INS_IN(29), INS_IN(28) => INS_IN(28), INS_IN(27) => 
                           INS_IN(27), INS_IN(26) => INS_IN(26), INS_IN(25) => 
                           INS_IN(25), INS_IN(24) => INS_IN(24), INS_IN(23) => 
                           INS_IN(23), INS_IN(22) => INS_IN(22), INS_IN(21) => 
                           INS_IN(21), INS_IN(20) => INS_IN(20), INS_IN(19) => 
                           INS_IN(19), INS_IN(18) => INS_IN(18), INS_IN(17) => 
                           INS_IN(17), INS_IN(16) => INS_IN(16), INS_IN(15) => 
                           INS_IN(15), INS_IN(14) => INS_IN(14), INS_IN(13) => 
                           INS_IN(13), INS_IN(12) => INS_IN(12), INS_IN(11) => 
                           INS_IN(11), INS_IN(10) => INS_IN(10), INS_IN(9) => 
                           INS_IN(9), INS_IN(8) => INS_IN(8), INS_IN(7) => 
                           INS_IN(7), INS_IN(6) => INS_IN(6), INS_IN(5) => 
                           INS_IN(5), INS_IN(4) => INS_IN(4), INS_IN(3) => 
                           INS_IN(3), INS_IN(2) => INS_IN(2), INS_IN(1) => 
                           INS_IN(1), INS_IN(0) => INS_IN(0), Bubble_in => 
                           Bubble_out_port, HDU_INS_IN(31) => 
                           sig_HDU_INS_OUT_31_port, HDU_INS_IN(30) => 
                           sig_HDU_INS_OUT_30_port, HDU_INS_IN(29) => 
                           sig_HDU_INS_OUT_29_port, HDU_INS_IN(28) => 
                           sig_HDU_INS_OUT_28_port, HDU_INS_IN(27) => 
                           sig_HDU_INS_OUT_27_port, HDU_INS_IN(26) => 
                           sig_HDU_INS_OUT_26_port, HDU_INS_IN(25) => 
                           sig_HDU_INS_OUT_25_port, HDU_INS_IN(24) => 
                           sig_HDU_INS_OUT_24_port, HDU_INS_IN(23) => 
                           sig_HDU_INS_OUT_23_port, HDU_INS_IN(22) => 
                           sig_HDU_INS_OUT_22_port, HDU_INS_IN(21) => 
                           sig_HDU_INS_OUT_21_port, HDU_INS_IN(20) => 
                           sig_HDU_INS_OUT_20_port, HDU_INS_IN(19) => 
                           sig_HDU_INS_OUT_19_port, HDU_INS_IN(18) => 
                           sig_HDU_INS_OUT_18_port, HDU_INS_IN(17) => 
                           sig_HDU_INS_OUT_17_port, HDU_INS_IN(16) => 
                           sig_HDU_INS_OUT_16_port, HDU_INS_IN(15) => 
                           sig_HDU_INS_OUT_15_port, HDU_INS_IN(14) => 
                           sig_HDU_INS_OUT_14_port, HDU_INS_IN(13) => 
                           sig_HDU_INS_OUT_13_port, HDU_INS_IN(12) => 
                           sig_HDU_INS_OUT_12_port, HDU_INS_IN(11) => 
                           sig_HDU_INS_OUT_11_port, HDU_INS_IN(10) => 
                           sig_HDU_INS_OUT_10_port, HDU_INS_IN(9) => 
                           sig_HDU_INS_OUT_9_port, HDU_INS_IN(8) => 
                           sig_HDU_INS_OUT_8_port, HDU_INS_IN(7) => 
                           sig_HDU_INS_OUT_7_port, HDU_INS_IN(6) => 
                           sig_HDU_INS_OUT_6_port, HDU_INS_IN(5) => 
                           sig_HDU_INS_OUT_5_port, HDU_INS_IN(4) => 
                           sig_HDU_INS_OUT_4_port, HDU_INS_IN(3) => 
                           sig_HDU_INS_OUT_3_port, HDU_INS_IN(2) => 
                           sig_HDU_INS_OUT_2_port, HDU_INS_IN(1) => 
                           sig_HDU_INS_OUT_1_port, HDU_INS_IN(0) => 
                           sig_HDU_INS_OUT_0_port, HDU_PC_IN(31) => 
                           sig_HDU_PC_OUT_31_port, HDU_PC_IN(30) => 
                           sig_HDU_PC_OUT_30_port, HDU_PC_IN(29) => 
                           sig_HDU_PC_OUT_29_port, HDU_PC_IN(28) => 
                           sig_HDU_PC_OUT_28_port, HDU_PC_IN(27) => 
                           sig_HDU_PC_OUT_27_port, HDU_PC_IN(26) => 
                           sig_HDU_PC_OUT_26_port, HDU_PC_IN(25) => 
                           sig_HDU_PC_OUT_25_port, HDU_PC_IN(24) => 
                           sig_HDU_PC_OUT_24_port, HDU_PC_IN(23) => 
                           sig_HDU_PC_OUT_23_port, HDU_PC_IN(22) => 
                           sig_HDU_PC_OUT_22_port, HDU_PC_IN(21) => 
                           sig_HDU_PC_OUT_21_port, HDU_PC_IN(20) => 
                           sig_HDU_PC_OUT_20_port, HDU_PC_IN(19) => 
                           sig_HDU_PC_OUT_19_port, HDU_PC_IN(18) => 
                           sig_HDU_PC_OUT_18_port, HDU_PC_IN(17) => 
                           sig_HDU_PC_OUT_17_port, HDU_PC_IN(16) => 
                           sig_HDU_PC_OUT_16_port, HDU_PC_IN(15) => 
                           sig_HDU_PC_OUT_15_port, HDU_PC_IN(14) => 
                           sig_HDU_PC_OUT_14_port, HDU_PC_IN(13) => 
                           sig_HDU_PC_OUT_13_port, HDU_PC_IN(12) => 
                           sig_HDU_PC_OUT_12_port, HDU_PC_IN(11) => 
                           sig_HDU_PC_OUT_11_port, HDU_PC_IN(10) => 
                           sig_HDU_PC_OUT_10_port, HDU_PC_IN(9) => 
                           sig_HDU_PC_OUT_9_port, HDU_PC_IN(8) => 
                           sig_HDU_PC_OUT_8_port, HDU_PC_IN(7) => 
                           sig_HDU_PC_OUT_7_port, HDU_PC_IN(6) => 
                           sig_HDU_PC_OUT_6_port, HDU_PC_IN(5) => 
                           sig_HDU_PC_OUT_5_port, HDU_PC_IN(4) => 
                           sig_HDU_PC_OUT_4_port, HDU_PC_IN(3) => 
                           sig_HDU_PC_OUT_3_port, HDU_PC_IN(2) => 
                           sig_HDU_PC_OUT_2_port, HDU_PC_IN(1) => 
                           sig_HDU_PC_OUT_1_port, HDU_PC_IN(0) => 
                           sig_HDU_PC_OUT_0_port, HDU_NPC_IN(31) => 
                           sig_HDU_NPC_OUT_31_port, HDU_NPC_IN(30) => 
                           sig_HDU_NPC_OUT_30_port, HDU_NPC_IN(29) => 
                           sig_HDU_NPC_OUT_29_port, HDU_NPC_IN(28) => 
                           sig_HDU_NPC_OUT_28_port, HDU_NPC_IN(27) => 
                           sig_HDU_NPC_OUT_27_port, HDU_NPC_IN(26) => 
                           sig_HDU_NPC_OUT_26_port, HDU_NPC_IN(25) => 
                           sig_HDU_NPC_OUT_25_port, HDU_NPC_IN(24) => 
                           sig_HDU_NPC_OUT_24_port, HDU_NPC_IN(23) => 
                           sig_HDU_NPC_OUT_23_port, HDU_NPC_IN(22) => 
                           sig_HDU_NPC_OUT_22_port, HDU_NPC_IN(21) => 
                           sig_HDU_NPC_OUT_21_port, HDU_NPC_IN(20) => 
                           sig_HDU_NPC_OUT_20_port, HDU_NPC_IN(19) => 
                           sig_HDU_NPC_OUT_19_port, HDU_NPC_IN(18) => 
                           sig_HDU_NPC_OUT_18_port, HDU_NPC_IN(17) => 
                           sig_HDU_NPC_OUT_17_port, HDU_NPC_IN(16) => 
                           sig_HDU_NPC_OUT_16_port, HDU_NPC_IN(15) => 
                           sig_HDU_NPC_OUT_15_port, HDU_NPC_IN(14) => 
                           sig_HDU_NPC_OUT_14_port, HDU_NPC_IN(13) => 
                           sig_HDU_NPC_OUT_13_port, HDU_NPC_IN(12) => 
                           sig_HDU_NPC_OUT_12_port, HDU_NPC_IN(11) => 
                           sig_HDU_NPC_OUT_11_port, HDU_NPC_IN(10) => 
                           sig_HDU_NPC_OUT_10_port, HDU_NPC_IN(9) => 
                           sig_HDU_NPC_OUT_9_port, HDU_NPC_IN(8) => 
                           sig_HDU_NPC_OUT_8_port, HDU_NPC_IN(7) => 
                           sig_HDU_NPC_OUT_7_port, HDU_NPC_IN(6) => 
                           sig_HDU_NPC_OUT_6_port, HDU_NPC_IN(5) => 
                           sig_HDU_NPC_OUT_5_port, HDU_NPC_IN(4) => 
                           sig_HDU_NPC_OUT_4_port, HDU_NPC_IN(3) => 
                           sig_HDU_NPC_OUT_3_port, HDU_NPC_IN(2) => 
                           sig_HDU_NPC_OUT_2_port, HDU_NPC_IN(1) => 
                           sig_HDU_NPC_OUT_1_port, HDU_NPC_IN(0) => 
                           sig_HDU_NPC_OUT_0_port, PC_OUT(31) => 
                           PC_FETCH_OUT_31_port, PC_OUT(30) => 
                           PC_FETCH_OUT_30_port, PC_OUT(29) => 
                           PC_FETCH_OUT_29_port, PC_OUT(28) => 
                           PC_FETCH_OUT_28_port, PC_OUT(27) => 
                           PC_FETCH_OUT_27_port, PC_OUT(26) => 
                           PC_FETCH_OUT_26_port, PC_OUT(25) => 
                           PC_FETCH_OUT_25_port, PC_OUT(24) => 
                           PC_FETCH_OUT_24_port, PC_OUT(23) => 
                           PC_FETCH_OUT_23_port, PC_OUT(22) => 
                           PC_FETCH_OUT_22_port, PC_OUT(21) => 
                           PC_FETCH_OUT_21_port, PC_OUT(20) => 
                           PC_FETCH_OUT_20_port, PC_OUT(19) => 
                           PC_FETCH_OUT_19_port, PC_OUT(18) => 
                           PC_FETCH_OUT_18_port, PC_OUT(17) => 
                           PC_FETCH_OUT_17_port, PC_OUT(16) => 
                           PC_FETCH_OUT_16_port, PC_OUT(15) => 
                           PC_FETCH_OUT_15_port, PC_OUT(14) => 
                           PC_FETCH_OUT_14_port, PC_OUT(13) => 
                           PC_FETCH_OUT_13_port, PC_OUT(12) => 
                           PC_FETCH_OUT_12_port, PC_OUT(11) => 
                           PC_FETCH_OUT_11_port, PC_OUT(10) => 
                           PC_FETCH_OUT_10_port, PC_OUT(9) => 
                           PC_FETCH_OUT_9_port, PC_OUT(8) => 
                           PC_FETCH_OUT_8_port, PC_OUT(7) => 
                           PC_FETCH_OUT_7_port, PC_OUT(6) => 
                           PC_FETCH_OUT_6_port, PC_OUT(5) => 
                           PC_FETCH_OUT_5_port, PC_OUT(4) => 
                           PC_FETCH_OUT_4_port, PC_OUT(3) => 
                           PC_FETCH_OUT_3_port, PC_OUT(2) => 
                           PC_FETCH_OUT_2_port, PC_OUT(1) => 
                           PC_FETCH_OUT_1_port, PC_OUT(0) => 
                           PC_FETCH_OUT_0_port, ADDR_OUT(31) => 
                           IRAM_ADDR_OUT(31), ADDR_OUT(30) => IRAM_ADDR_OUT(30)
                           , ADDR_OUT(29) => IRAM_ADDR_OUT(29), ADDR_OUT(28) =>
                           IRAM_ADDR_OUT(28), ADDR_OUT(27) => IRAM_ADDR_OUT(27)
                           , ADDR_OUT(26) => IRAM_ADDR_OUT(26), ADDR_OUT(25) =>
                           IRAM_ADDR_OUT(25), ADDR_OUT(24) => IRAM_ADDR_OUT(24)
                           , ADDR_OUT(23) => IRAM_ADDR_OUT(23), ADDR_OUT(22) =>
                           IRAM_ADDR_OUT(22), ADDR_OUT(21) => IRAM_ADDR_OUT(21)
                           , ADDR_OUT(20) => IRAM_ADDR_OUT(20), ADDR_OUT(19) =>
                           IRAM_ADDR_OUT(19), ADDR_OUT(18) => IRAM_ADDR_OUT(18)
                           , ADDR_OUT(17) => IRAM_ADDR_OUT(17), ADDR_OUT(16) =>
                           IRAM_ADDR_OUT(16), ADDR_OUT(15) => IRAM_ADDR_OUT(15)
                           , ADDR_OUT(14) => IRAM_ADDR_OUT(14), ADDR_OUT(13) =>
                           IRAM_ADDR_OUT(13), ADDR_OUT(12) => IRAM_ADDR_OUT(12)
                           , ADDR_OUT(11) => IRAM_ADDR_OUT(11), ADDR_OUT(10) =>
                           IRAM_ADDR_OUT(10), ADDR_OUT(9) => IRAM_ADDR_OUT(9), 
                           ADDR_OUT(8) => IRAM_ADDR_OUT(8), ADDR_OUT(7) => 
                           IRAM_ADDR_OUT(7), ADDR_OUT(6) => IRAM_ADDR_OUT(6), 
                           ADDR_OUT(5) => IRAM_ADDR_OUT(5), ADDR_OUT(4) => 
                           IRAM_ADDR_OUT(4), ADDR_OUT(3) => IRAM_ADDR_OUT(3), 
                           ADDR_OUT(2) => IRAM_ADDR_OUT(2), ADDR_OUT(1) => 
                           IRAM_ADDR_OUT(1), ADDR_OUT(0) => IRAM_ADDR_OUT(0), 
                           NPC_OUT(31) => NPC_FETCH_OUT_31_port, NPC_OUT(30) =>
                           NPC_FETCH_OUT_30_port, NPC_OUT(29) => 
                           NPC_FETCH_OUT_29_port, NPC_OUT(28) => 
                           NPC_FETCH_OUT_28_port, NPC_OUT(27) => 
                           NPC_FETCH_OUT_27_port, NPC_OUT(26) => 
                           NPC_FETCH_OUT_26_port, NPC_OUT(25) => 
                           NPC_FETCH_OUT_25_port, NPC_OUT(24) => 
                           NPC_FETCH_OUT_24_port, NPC_OUT(23) => 
                           NPC_FETCH_OUT_23_port, NPC_OUT(22) => 
                           NPC_FETCH_OUT_22_port, NPC_OUT(21) => 
                           NPC_FETCH_OUT_21_port, NPC_OUT(20) => 
                           NPC_FETCH_OUT_20_port, NPC_OUT(19) => 
                           NPC_FETCH_OUT_19_port, NPC_OUT(18) => 
                           NPC_FETCH_OUT_18_port, NPC_OUT(17) => 
                           NPC_FETCH_OUT_17_port, NPC_OUT(16) => 
                           NPC_FETCH_OUT_16_port, NPC_OUT(15) => 
                           NPC_FETCH_OUT_15_port, NPC_OUT(14) => 
                           NPC_FETCH_OUT_14_port, NPC_OUT(13) => 
                           NPC_FETCH_OUT_13_port, NPC_OUT(12) => 
                           NPC_FETCH_OUT_12_port, NPC_OUT(11) => 
                           NPC_FETCH_OUT_11_port, NPC_OUT(10) => 
                           NPC_FETCH_OUT_10_port, NPC_OUT(9) => 
                           NPC_FETCH_OUT_9_port, NPC_OUT(8) => 
                           NPC_FETCH_OUT_8_port, NPC_OUT(7) => 
                           NPC_FETCH_OUT_7_port, NPC_OUT(6) => 
                           NPC_FETCH_OUT_6_port, NPC_OUT(5) => 
                           NPC_FETCH_OUT_5_port, NPC_OUT(4) => 
                           NPC_FETCH_OUT_4_port, NPC_OUT(3) => 
                           NPC_FETCH_OUT_3_port, NPC_OUT(2) => 
                           NPC_FETCH_OUT_2_port, NPC_OUT(1) => 
                           NPC_FETCH_OUT_1_port, NPC_OUT(0) => 
                           NPC_FETCH_OUT_0_port, INS_OUT(31) => INS_OUT_31_port
                           , INS_OUT(30) => INS_OUT_30_port, INS_OUT(29) => 
                           INS_OUT_29_port, INS_OUT(28) => INS_OUT_28_port, 
                           INS_OUT(27) => INS_OUT_27_port, INS_OUT(26) => 
                           INS_OUT_26_port, INS_OUT(25) => INS_OUT_25_port, 
                           INS_OUT(24) => INS_OUT_24_port, INS_OUT(23) => 
                           INS_OUT_23_port, INS_OUT(22) => INS_OUT_22_port, 
                           INS_OUT(21) => INS_OUT_21_port, INS_OUT(20) => 
                           INS_OUT_20_port, INS_OUT(19) => INS_OUT_19_port, 
                           INS_OUT(18) => INS_OUT_18_port, INS_OUT(17) => 
                           INS_OUT_17_port, INS_OUT(16) => INS_OUT_16_port, 
                           INS_OUT(15) => INS_OUT_15_port, INS_OUT(14) => 
                           INS_OUT_14_port, INS_OUT(13) => INS_OUT_13_port, 
                           INS_OUT(12) => INS_OUT_12_port, INS_OUT(11) => 
                           INS_OUT_11_port, INS_OUT(10) => INS_OUT_10_port, 
                           INS_OUT(9) => INS_OUT_9_port, INS_OUT(8) => 
                           INS_OUT_8_port, INS_OUT(7) => INS_OUT_7_port, 
                           INS_OUT(6) => INS_OUT_6_port, INS_OUT(5) => 
                           INS_OUT_5_port, INS_OUT(4) => INS_OUT_4_port, 
                           INS_OUT(3) => INS_OUT_3_port, INS_OUT(2) => 
                           INS_OUT_2_port, INS_OUT(1) => INS_OUT_1_port, 
                           INS_OUT(0) => INS_OUT_0_port);
   DecodeStage : Decode port map( CLK => CLK, RST => RST, REG_LATCH_EN => 
                           REG_LATCH_EN, RD1 => RD1, RD2 => RD2, RF_WE => 
                           RF_WE_WB, ZERO_FLAG => ZERO_FLAG_EX, PC_IN(31) => 
                           PC_FETCH_OUT_31_port, PC_IN(30) => 
                           PC_FETCH_OUT_30_port, PC_IN(29) => 
                           PC_FETCH_OUT_29_port, PC_IN(28) => 
                           PC_FETCH_OUT_28_port, PC_IN(27) => 
                           PC_FETCH_OUT_27_port, PC_IN(26) => 
                           PC_FETCH_OUT_26_port, PC_IN(25) => 
                           PC_FETCH_OUT_25_port, PC_IN(24) => 
                           PC_FETCH_OUT_24_port, PC_IN(23) => 
                           PC_FETCH_OUT_23_port, PC_IN(22) => 
                           PC_FETCH_OUT_22_port, PC_IN(21) => 
                           PC_FETCH_OUT_21_port, PC_IN(20) => 
                           PC_FETCH_OUT_20_port, PC_IN(19) => 
                           PC_FETCH_OUT_19_port, PC_IN(18) => 
                           PC_FETCH_OUT_18_port, PC_IN(17) => 
                           PC_FETCH_OUT_17_port, PC_IN(16) => 
                           PC_FETCH_OUT_16_port, PC_IN(15) => 
                           PC_FETCH_OUT_15_port, PC_IN(14) => 
                           PC_FETCH_OUT_14_port, PC_IN(13) => 
                           PC_FETCH_OUT_13_port, PC_IN(12) => 
                           PC_FETCH_OUT_12_port, PC_IN(11) => 
                           PC_FETCH_OUT_11_port, PC_IN(10) => 
                           PC_FETCH_OUT_10_port, PC_IN(9) => 
                           PC_FETCH_OUT_9_port, PC_IN(8) => PC_FETCH_OUT_8_port
                           , PC_IN(7) => PC_FETCH_OUT_7_port, PC_IN(6) => 
                           PC_FETCH_OUT_6_port, PC_IN(5) => PC_FETCH_OUT_5_port
                           , PC_IN(4) => PC_FETCH_OUT_4_port, PC_IN(3) => 
                           PC_FETCH_OUT_3_port, PC_IN(2) => PC_FETCH_OUT_2_port
                           , PC_IN(1) => PC_FETCH_OUT_1_port, PC_IN(0) => 
                           PC_FETCH_OUT_0_port, INS_IN(31) => INS_OUT_31_port, 
                           INS_IN(30) => INS_OUT_30_port, INS_IN(29) => 
                           INS_OUT_29_port, INS_IN(28) => INS_OUT_28_port, 
                           INS_IN(27) => INS_OUT_27_port, INS_IN(26) => 
                           INS_OUT_26_port, INS_IN(25) => INS_OUT_25_port, 
                           INS_IN(24) => INS_OUT_24_port, INS_IN(23) => 
                           INS_OUT_23_port, INS_IN(22) => INS_OUT_22_port, 
                           INS_IN(21) => INS_OUT_21_port, INS_IN(20) => 
                           INS_OUT_20_port, INS_IN(19) => INS_OUT_19_port, 
                           INS_IN(18) => INS_OUT_18_port, INS_IN(17) => 
                           INS_OUT_17_port, INS_IN(16) => INS_OUT_16_port, 
                           INS_IN(15) => INS_OUT_15_port, INS_IN(14) => 
                           INS_OUT_14_port, INS_IN(13) => INS_OUT_13_port, 
                           INS_IN(12) => INS_OUT_12_port, INS_IN(11) => 
                           INS_OUT_11_port, INS_IN(10) => INS_OUT_10_port, 
                           INS_IN(9) => INS_OUT_9_port, INS_IN(8) => 
                           INS_OUT_8_port, INS_IN(7) => INS_OUT_7_port, 
                           INS_IN(6) => INS_OUT_6_port, INS_IN(5) => 
                           INS_OUT_5_port, INS_IN(4) => INS_OUT_4_port, 
                           INS_IN(3) => INS_OUT_3_port, INS_IN(2) => 
                           INS_OUT_2_port, INS_IN(1) => INS_OUT_1_port, 
                           INS_IN(0) => INS_OUT_0_port, ADD_WR(4) => 
                           ADD_WR_WB_4_port, ADD_WR(3) => ADD_WR_WB_3_port, 
                           ADD_WR(2) => ADD_WR_WB_2_port, ADD_WR(1) => 
                           ADD_WR_WB_1_port, ADD_WR(0) => ADD_WR_WB_0_port, 
                           DATA_WR_IN(31) => OP_WB_31_port, DATA_WR_IN(30) => 
                           OP_WB_30_port, DATA_WR_IN(29) => OP_WB_29_port, 
                           DATA_WR_IN(28) => OP_WB_28_port, DATA_WR_IN(27) => 
                           OP_WB_27_port, DATA_WR_IN(26) => OP_WB_26_port, 
                           DATA_WR_IN(25) => OP_WB_25_port, DATA_WR_IN(24) => 
                           OP_WB_24_port, DATA_WR_IN(23) => OP_WB_23_port, 
                           DATA_WR_IN(22) => OP_WB_22_port, DATA_WR_IN(21) => 
                           OP_WB_21_port, DATA_WR_IN(20) => OP_WB_20_port, 
                           DATA_WR_IN(19) => OP_WB_19_port, DATA_WR_IN(18) => 
                           OP_WB_18_port, DATA_WR_IN(17) => OP_WB_17_port, 
                           DATA_WR_IN(16) => OP_WB_16_port, DATA_WR_IN(15) => 
                           OP_WB_15_port, DATA_WR_IN(14) => OP_WB_14_port, 
                           DATA_WR_IN(13) => OP_WB_13_port, DATA_WR_IN(12) => 
                           OP_WB_12_port, DATA_WR_IN(11) => OP_WB_11_port, 
                           DATA_WR_IN(10) => OP_WB_10_port, DATA_WR_IN(9) => 
                           OP_WB_9_port, DATA_WR_IN(8) => OP_WB_8_port, 
                           DATA_WR_IN(7) => OP_WB_7_port, DATA_WR_IN(6) => 
                           OP_WB_6_port, DATA_WR_IN(5) => OP_WB_5_port, 
                           DATA_WR_IN(4) => OP_WB_4_port, DATA_WR_IN(3) => 
                           OP_WB_3_port, DATA_WR_IN(2) => OP_WB_2_port, 
                           DATA_WR_IN(1) => OP_WB_1_port, DATA_WR_IN(0) => 
                           OP_WB_0_port, PC_OUT(31) => PC_DECODE_OUT_31_port, 
                           PC_OUT(30) => PC_DECODE_OUT_30_port, PC_OUT(29) => 
                           PC_DECODE_OUT_29_port, PC_OUT(28) => 
                           PC_DECODE_OUT_28_port, PC_OUT(27) => 
                           PC_DECODE_OUT_27_port, PC_OUT(26) => 
                           PC_DECODE_OUT_26_port, PC_OUT(25) => 
                           PC_DECODE_OUT_25_port, PC_OUT(24) => 
                           PC_DECODE_OUT_24_port, PC_OUT(23) => 
                           PC_DECODE_OUT_23_port, PC_OUT(22) => 
                           PC_DECODE_OUT_22_port, PC_OUT(21) => 
                           PC_DECODE_OUT_21_port, PC_OUT(20) => 
                           PC_DECODE_OUT_20_port, PC_OUT(19) => 
                           PC_DECODE_OUT_19_port, PC_OUT(18) => 
                           PC_DECODE_OUT_18_port, PC_OUT(17) => 
                           PC_DECODE_OUT_17_port, PC_OUT(16) => 
                           PC_DECODE_OUT_16_port, PC_OUT(15) => 
                           PC_DECODE_OUT_15_port, PC_OUT(14) => 
                           PC_DECODE_OUT_14_port, PC_OUT(13) => 
                           PC_DECODE_OUT_13_port, PC_OUT(12) => 
                           PC_DECODE_OUT_12_port, PC_OUT(11) => 
                           PC_DECODE_OUT_11_port, PC_OUT(10) => 
                           PC_DECODE_OUT_10_port, PC_OUT(9) => 
                           PC_DECODE_OUT_9_port, PC_OUT(8) => 
                           PC_DECODE_OUT_8_port, PC_OUT(7) => 
                           PC_DECODE_OUT_7_port, PC_OUT(6) => 
                           PC_DECODE_OUT_6_port, PC_OUT(5) => 
                           PC_DECODE_OUT_5_port, PC_OUT(4) => 
                           PC_DECODE_OUT_4_port, PC_OUT(3) => 
                           PC_DECODE_OUT_3_port, PC_OUT(2) => 
                           PC_DECODE_OUT_2_port, PC_OUT(1) => 
                           PC_DECODE_OUT_1_port, PC_OUT(0) => 
                           PC_DECODE_OUT_0_port, A_OUT(31) => 
                           A_DECODE_OUT_31_port, A_OUT(30) => 
                           A_DECODE_OUT_30_port, A_OUT(29) => 
                           A_DECODE_OUT_29_port, A_OUT(28) => 
                           A_DECODE_OUT_28_port, A_OUT(27) => 
                           A_DECODE_OUT_27_port, A_OUT(26) => 
                           A_DECODE_OUT_26_port, A_OUT(25) => 
                           A_DECODE_OUT_25_port, A_OUT(24) => 
                           A_DECODE_OUT_24_port, A_OUT(23) => 
                           A_DECODE_OUT_23_port, A_OUT(22) => 
                           A_DECODE_OUT_22_port, A_OUT(21) => 
                           A_DECODE_OUT_21_port, A_OUT(20) => 
                           A_DECODE_OUT_20_port, A_OUT(19) => 
                           A_DECODE_OUT_19_port, A_OUT(18) => 
                           A_DECODE_OUT_18_port, A_OUT(17) => 
                           A_DECODE_OUT_17_port, A_OUT(16) => 
                           A_DECODE_OUT_16_port, A_OUT(15) => 
                           A_DECODE_OUT_15_port, A_OUT(14) => 
                           A_DECODE_OUT_14_port, A_OUT(13) => 
                           A_DECODE_OUT_13_port, A_OUT(12) => 
                           A_DECODE_OUT_12_port, A_OUT(11) => 
                           A_DECODE_OUT_11_port, A_OUT(10) => 
                           A_DECODE_OUT_10_port, A_OUT(9) => 
                           A_DECODE_OUT_9_port, A_OUT(8) => A_DECODE_OUT_8_port
                           , A_OUT(7) => A_DECODE_OUT_7_port, A_OUT(6) => 
                           A_DECODE_OUT_6_port, A_OUT(5) => A_DECODE_OUT_5_port
                           , A_OUT(4) => A_DECODE_OUT_4_port, A_OUT(3) => 
                           A_DECODE_OUT_3_port, A_OUT(2) => A_DECODE_OUT_2_port
                           , A_OUT(1) => A_DECODE_OUT_1_port, A_OUT(0) => 
                           A_DECODE_OUT_0_port, B_OUT(31) => 
                           B_DECODE_OUT_31_port, B_OUT(30) => 
                           B_DECODE_OUT_30_port, B_OUT(29) => 
                           B_DECODE_OUT_29_port, B_OUT(28) => 
                           B_DECODE_OUT_28_port, B_OUT(27) => 
                           B_DECODE_OUT_27_port, B_OUT(26) => 
                           B_DECODE_OUT_26_port, B_OUT(25) => 
                           B_DECODE_OUT_25_port, B_OUT(24) => 
                           B_DECODE_OUT_24_port, B_OUT(23) => 
                           B_DECODE_OUT_23_port, B_OUT(22) => 
                           B_DECODE_OUT_22_port, B_OUT(21) => 
                           B_DECODE_OUT_21_port, B_OUT(20) => 
                           B_DECODE_OUT_20_port, B_OUT(19) => 
                           B_DECODE_OUT_19_port, B_OUT(18) => 
                           B_DECODE_OUT_18_port, B_OUT(17) => 
                           B_DECODE_OUT_17_port, B_OUT(16) => 
                           B_DECODE_OUT_16_port, B_OUT(15) => 
                           B_DECODE_OUT_15_port, B_OUT(14) => 
                           B_DECODE_OUT_14_port, B_OUT(13) => 
                           B_DECODE_OUT_13_port, B_OUT(12) => 
                           B_DECODE_OUT_12_port, B_OUT(11) => 
                           B_DECODE_OUT_11_port, B_OUT(10) => 
                           B_DECODE_OUT_10_port, B_OUT(9) => 
                           B_DECODE_OUT_9_port, B_OUT(8) => B_DECODE_OUT_8_port
                           , B_OUT(7) => B_DECODE_OUT_7_port, B_OUT(6) => 
                           B_DECODE_OUT_6_port, B_OUT(5) => B_DECODE_OUT_5_port
                           , B_OUT(4) => B_DECODE_OUT_4_port, B_OUT(3) => 
                           B_DECODE_OUT_3_port, B_OUT(2) => B_DECODE_OUT_2_port
                           , B_OUT(1) => B_DECODE_OUT_1_port, B_OUT(0) => 
                           B_DECODE_OUT_0_port, IMM_OUT(31) => 
                           IMM_DECODE_OUT_31_port, IMM_OUT(30) => 
                           IMM_DECODE_OUT_30_port, IMM_OUT(29) => 
                           IMM_DECODE_OUT_29_port, IMM_OUT(28) => 
                           IMM_DECODE_OUT_28_port, IMM_OUT(27) => 
                           IMM_DECODE_OUT_27_port, IMM_OUT(26) => 
                           IMM_DECODE_OUT_26_port, IMM_OUT(25) => 
                           IMM_DECODE_OUT_25_port, IMM_OUT(24) => 
                           IMM_DECODE_OUT_24_port, IMM_OUT(23) => 
                           IMM_DECODE_OUT_23_port, IMM_OUT(22) => 
                           IMM_DECODE_OUT_22_port, IMM_OUT(21) => 
                           IMM_DECODE_OUT_21_port, IMM_OUT(20) => 
                           IMM_DECODE_OUT_20_port, IMM_OUT(19) => 
                           IMM_DECODE_OUT_19_port, IMM_OUT(18) => 
                           IMM_DECODE_OUT_18_port, IMM_OUT(17) => 
                           IMM_DECODE_OUT_17_port, IMM_OUT(16) => 
                           IMM_DECODE_OUT_16_port, IMM_OUT(15) => 
                           IMM_DECODE_OUT_15_port, IMM_OUT(14) => 
                           IMM_DECODE_OUT_14_port, IMM_OUT(13) => 
                           IMM_DECODE_OUT_13_port, IMM_OUT(12) => 
                           IMM_DECODE_OUT_12_port, IMM_OUT(11) => 
                           IMM_DECODE_OUT_11_port, IMM_OUT(10) => 
                           IMM_DECODE_OUT_10_port, IMM_OUT(9) => 
                           IMM_DECODE_OUT_9_port, IMM_OUT(8) => 
                           IMM_DECODE_OUT_8_port, IMM_OUT(7) => 
                           IMM_DECODE_OUT_7_port, IMM_OUT(6) => 
                           IMM_DECODE_OUT_6_port, IMM_OUT(5) => 
                           IMM_DECODE_OUT_5_port, IMM_OUT(4) => 
                           IMM_DECODE_OUT_4_port, IMM_OUT(3) => 
                           IMM_DECODE_OUT_3_port, IMM_OUT(2) => 
                           IMM_DECODE_OUT_2_port, IMM_OUT(1) => 
                           IMM_DECODE_OUT_1_port, IMM_OUT(0) => 
                           IMM_DECODE_OUT_0_port, ADD_RS1_HDU(4) => 
                           ADD_RS1_HDU_4_port, ADD_RS1_HDU(3) => 
                           ADD_RS1_HDU_3_port, ADD_RS1_HDU(2) => 
                           ADD_RS1_HDU_2_port, ADD_RS1_HDU(1) => 
                           ADD_RS1_HDU_1_port, ADD_RS1_HDU(0) => 
                           ADD_RS1_HDU_0_port, ADD_RS2_HDU(4) => 
                           ADD_RS2_HDU_4_port, ADD_RS2_HDU(3) => 
                           ADD_RS2_HDU_3_port, ADD_RS2_HDU(2) => 
                           ADD_RS2_HDU_2_port, ADD_RS2_HDU(1) => 
                           ADD_RS2_HDU_1_port, ADD_RS2_HDU(0) => 
                           ADD_RS2_HDU_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_DECODE_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_DECODE_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_DECODE_OUT_0_port, ADD_RS1_OUT(4) => 
                           ADD_RS1_DECODE_OUT_4_port, ADD_RS1_OUT(3) => 
                           ADD_RS1_DECODE_OUT_3_port, ADD_RS1_OUT(2) => 
                           ADD_RS1_DECODE_OUT_2_port, ADD_RS1_OUT(1) => 
                           ADD_RS1_DECODE_OUT_1_port, ADD_RS1_OUT(0) => 
                           ADD_RS1_DECODE_OUT_0_port, ADD_RS2_OUT(4) => 
                           ADD_RS2_DECODE_OUT_4_port, ADD_RS2_OUT(3) => 
                           ADD_RS2_DECODE_OUT_3_port, ADD_RS2_OUT(2) => 
                           ADD_RS2_DECODE_OUT_2_port, ADD_RS2_OUT(1) => 
                           ADD_RS2_DECODE_OUT_1_port, ADD_RS2_OUT(0) => 
                           ADD_RS2_DECODE_OUT_0_port);
   ExecuteStage : Execute port map( CLK => CLK, RST => RST, MUX_A_SEL => 
                           MUX_A_SEL, MUX_B_SEL(1) => MUX_B_SEL(1), 
                           MUX_B_SEL(0) => MUX_B_SEL(0), ALU_OPC(0) => 
                           ALU_OPC(0), ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => 
                           ALU_OPC(2), ALU_OPC(3) => ALU_OPC(3), ALU_OUTREG_EN 
                           => ALU_OUTREG_EN, JUMP_TYPE(1) => JUMP_TYPE(1), 
                           JUMP_TYPE(0) => JUMP_TYPE(0), PC_IN(31) => 
                           PC_DECODE_OUT_31_port, PC_IN(30) => 
                           PC_DECODE_OUT_30_port, PC_IN(29) => 
                           PC_DECODE_OUT_29_port, PC_IN(28) => 
                           PC_DECODE_OUT_28_port, PC_IN(27) => 
                           PC_DECODE_OUT_27_port, PC_IN(26) => 
                           PC_DECODE_OUT_26_port, PC_IN(25) => 
                           PC_DECODE_OUT_25_port, PC_IN(24) => 
                           PC_DECODE_OUT_24_port, PC_IN(23) => 
                           PC_DECODE_OUT_23_port, PC_IN(22) => 
                           PC_DECODE_OUT_22_port, PC_IN(21) => 
                           PC_DECODE_OUT_21_port, PC_IN(20) => 
                           PC_DECODE_OUT_20_port, PC_IN(19) => 
                           PC_DECODE_OUT_19_port, PC_IN(18) => 
                           PC_DECODE_OUT_18_port, PC_IN(17) => 
                           PC_DECODE_OUT_17_port, PC_IN(16) => 
                           PC_DECODE_OUT_16_port, PC_IN(15) => 
                           PC_DECODE_OUT_15_port, PC_IN(14) => 
                           PC_DECODE_OUT_14_port, PC_IN(13) => 
                           PC_DECODE_OUT_13_port, PC_IN(12) => 
                           PC_DECODE_OUT_12_port, PC_IN(11) => 
                           PC_DECODE_OUT_11_port, PC_IN(10) => 
                           PC_DECODE_OUT_10_port, PC_IN(9) => 
                           PC_DECODE_OUT_9_port, PC_IN(8) => 
                           PC_DECODE_OUT_8_port, PC_IN(7) => 
                           PC_DECODE_OUT_7_port, PC_IN(6) => 
                           PC_DECODE_OUT_6_port, PC_IN(5) => 
                           PC_DECODE_OUT_5_port, PC_IN(4) => 
                           PC_DECODE_OUT_4_port, PC_IN(3) => 
                           PC_DECODE_OUT_3_port, PC_IN(2) => 
                           PC_DECODE_OUT_2_port, PC_IN(1) => 
                           PC_DECODE_OUT_1_port, PC_IN(0) => 
                           PC_DECODE_OUT_0_port, A_IN(31) => 
                           A_DECODE_OUT_31_port, A_IN(30) => 
                           A_DECODE_OUT_30_port, A_IN(29) => 
                           A_DECODE_OUT_29_port, A_IN(28) => 
                           A_DECODE_OUT_28_port, A_IN(27) => 
                           A_DECODE_OUT_27_port, A_IN(26) => 
                           A_DECODE_OUT_26_port, A_IN(25) => 
                           A_DECODE_OUT_25_port, A_IN(24) => 
                           A_DECODE_OUT_24_port, A_IN(23) => 
                           A_DECODE_OUT_23_port, A_IN(22) => 
                           A_DECODE_OUT_22_port, A_IN(21) => 
                           A_DECODE_OUT_21_port, A_IN(20) => 
                           A_DECODE_OUT_20_port, A_IN(19) => 
                           A_DECODE_OUT_19_port, A_IN(18) => 
                           A_DECODE_OUT_18_port, A_IN(17) => 
                           A_DECODE_OUT_17_port, A_IN(16) => 
                           A_DECODE_OUT_16_port, A_IN(15) => 
                           A_DECODE_OUT_15_port, A_IN(14) => 
                           A_DECODE_OUT_14_port, A_IN(13) => 
                           A_DECODE_OUT_13_port, A_IN(12) => 
                           A_DECODE_OUT_12_port, A_IN(11) => 
                           A_DECODE_OUT_11_port, A_IN(10) => 
                           A_DECODE_OUT_10_port, A_IN(9) => A_DECODE_OUT_9_port
                           , A_IN(8) => A_DECODE_OUT_8_port, A_IN(7) => 
                           A_DECODE_OUT_7_port, A_IN(6) => A_DECODE_OUT_6_port,
                           A_IN(5) => A_DECODE_OUT_5_port, A_IN(4) => 
                           A_DECODE_OUT_4_port, A_IN(3) => A_DECODE_OUT_3_port,
                           A_IN(2) => A_DECODE_OUT_2_port, A_IN(1) => 
                           A_DECODE_OUT_1_port, A_IN(0) => A_DECODE_OUT_0_port,
                           B_IN(31) => B_DECODE_OUT_31_port, B_IN(30) => 
                           B_DECODE_OUT_30_port, B_IN(29) => 
                           B_DECODE_OUT_29_port, B_IN(28) => 
                           B_DECODE_OUT_28_port, B_IN(27) => 
                           B_DECODE_OUT_27_port, B_IN(26) => 
                           B_DECODE_OUT_26_port, B_IN(25) => 
                           B_DECODE_OUT_25_port, B_IN(24) => 
                           B_DECODE_OUT_24_port, B_IN(23) => 
                           B_DECODE_OUT_23_port, B_IN(22) => 
                           B_DECODE_OUT_22_port, B_IN(21) => 
                           B_DECODE_OUT_21_port, B_IN(20) => 
                           B_DECODE_OUT_20_port, B_IN(19) => 
                           B_DECODE_OUT_19_port, B_IN(18) => 
                           B_DECODE_OUT_18_port, B_IN(17) => 
                           B_DECODE_OUT_17_port, B_IN(16) => 
                           B_DECODE_OUT_16_port, B_IN(15) => 
                           B_DECODE_OUT_15_port, B_IN(14) => 
                           B_DECODE_OUT_14_port, B_IN(13) => 
                           B_DECODE_OUT_13_port, B_IN(12) => 
                           B_DECODE_OUT_12_port, B_IN(11) => 
                           B_DECODE_OUT_11_port, B_IN(10) => 
                           B_DECODE_OUT_10_port, B_IN(9) => B_DECODE_OUT_9_port
                           , B_IN(8) => B_DECODE_OUT_8_port, B_IN(7) => 
                           B_DECODE_OUT_7_port, B_IN(6) => B_DECODE_OUT_6_port,
                           B_IN(5) => B_DECODE_OUT_5_port, B_IN(4) => 
                           B_DECODE_OUT_4_port, B_IN(3) => B_DECODE_OUT_3_port,
                           B_IN(2) => B_DECODE_OUT_2_port, B_IN(1) => 
                           B_DECODE_OUT_1_port, B_IN(0) => B_DECODE_OUT_0_port,
                           IMM_IN(31) => IMM_DECODE_OUT_31_port, IMM_IN(30) => 
                           IMM_DECODE_OUT_30_port, IMM_IN(29) => 
                           IMM_DECODE_OUT_29_port, IMM_IN(28) => 
                           IMM_DECODE_OUT_28_port, IMM_IN(27) => 
                           IMM_DECODE_OUT_27_port, IMM_IN(26) => 
                           IMM_DECODE_OUT_26_port, IMM_IN(25) => 
                           IMM_DECODE_OUT_25_port, IMM_IN(24) => 
                           IMM_DECODE_OUT_24_port, IMM_IN(23) => 
                           IMM_DECODE_OUT_23_port, IMM_IN(22) => 
                           IMM_DECODE_OUT_22_port, IMM_IN(21) => 
                           IMM_DECODE_OUT_21_port, IMM_IN(20) => 
                           IMM_DECODE_OUT_20_port, IMM_IN(19) => 
                           IMM_DECODE_OUT_19_port, IMM_IN(18) => 
                           IMM_DECODE_OUT_18_port, IMM_IN(17) => 
                           IMM_DECODE_OUT_17_port, IMM_IN(16) => 
                           IMM_DECODE_OUT_16_port, IMM_IN(15) => 
                           IMM_DECODE_OUT_15_port, IMM_IN(14) => 
                           IMM_DECODE_OUT_14_port, IMM_IN(13) => 
                           IMM_DECODE_OUT_13_port, IMM_IN(12) => 
                           IMM_DECODE_OUT_12_port, IMM_IN(11) => 
                           IMM_DECODE_OUT_11_port, IMM_IN(10) => 
                           IMM_DECODE_OUT_10_port, IMM_IN(9) => 
                           IMM_DECODE_OUT_9_port, IMM_IN(8) => 
                           IMM_DECODE_OUT_8_port, IMM_IN(7) => 
                           IMM_DECODE_OUT_7_port, IMM_IN(6) => 
                           IMM_DECODE_OUT_6_port, IMM_IN(5) => 
                           IMM_DECODE_OUT_5_port, IMM_IN(4) => 
                           IMM_DECODE_OUT_4_port, IMM_IN(3) => 
                           IMM_DECODE_OUT_3_port, IMM_IN(2) => 
                           IMM_DECODE_OUT_2_port, IMM_IN(1) => 
                           IMM_DECODE_OUT_1_port, IMM_IN(0) => 
                           IMM_DECODE_OUT_0_port, ADD_WR_IN(4) => 
                           ADD_WR_DECODE_OUT_4_port, ADD_WR_IN(3) => 
                           ADD_WR_DECODE_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_DECODE_OUT_0_port, ADD_RS1_IN(4) => 
                           ADD_RS1_DECODE_OUT_4_port, ADD_RS1_IN(3) => 
                           ADD_RS1_DECODE_OUT_3_port, ADD_RS1_IN(2) => 
                           ADD_RS1_DECODE_OUT_2_port, ADD_RS1_IN(1) => 
                           ADD_RS1_DECODE_OUT_1_port, ADD_RS1_IN(0) => 
                           ADD_RS1_DECODE_OUT_0_port, ADD_RS2_IN(4) => 
                           ADD_RS2_DECODE_OUT_4_port, ADD_RS2_IN(3) => 
                           ADD_RS2_DECODE_OUT_3_port, ADD_RS2_IN(2) => 
                           ADD_RS2_DECODE_OUT_2_port, ADD_RS2_IN(1) => 
                           ADD_RS2_DECODE_OUT_1_port, ADD_RS2_IN(0) => 
                           ADD_RS2_DECODE_OUT_0_port, ADD_WR_MEM(4) => 
                           ADD_WR_MEM_4_port, ADD_WR_MEM(3) => 
                           ADD_WR_MEM_3_port, ADD_WR_MEM(2) => 
                           ADD_WR_MEM_2_port, ADD_WR_MEM(1) => 
                           ADD_WR_MEM_1_port, ADD_WR_MEM(0) => 
                           ADD_WR_MEM_0_port, ADD_WR_WB(4) => ADD_WR_WB_4_port,
                           ADD_WR_WB(3) => ADD_WR_WB_3_port, ADD_WR_WB(2) => 
                           ADD_WR_WB_2_port, ADD_WR_WB(1) => ADD_WR_WB_1_port, 
                           ADD_WR_WB(0) => ADD_WR_WB_0_port, RF_WE_MEM => RF_WE
                           , RF_WE_WB => RF_WE_WB, OP_MEM(31) => OP_MEM_31_port
                           , OP_MEM(30) => OP_MEM_30_port, OP_MEM(29) => 
                           OP_MEM_29_port, OP_MEM(28) => OP_MEM_28_port, 
                           OP_MEM(27) => OP_MEM_27_port, OP_MEM(26) => 
                           OP_MEM_26_port, OP_MEM(25) => OP_MEM_25_port, 
                           OP_MEM(24) => OP_MEM_24_port, OP_MEM(23) => 
                           OP_MEM_23_port, OP_MEM(22) => OP_MEM_22_port, 
                           OP_MEM(21) => OP_MEM_21_port, OP_MEM(20) => 
                           OP_MEM_20_port, OP_MEM(19) => OP_MEM_19_port, 
                           OP_MEM(18) => OP_MEM_18_port, OP_MEM(17) => 
                           OP_MEM_17_port, OP_MEM(16) => OP_MEM_16_port, 
                           OP_MEM(15) => OP_MEM_15_port, OP_MEM(14) => 
                           OP_MEM_14_port, OP_MEM(13) => OP_MEM_13_port, 
                           OP_MEM(12) => OP_MEM_12_port, OP_MEM(11) => 
                           OP_MEM_11_port, OP_MEM(10) => OP_MEM_10_port, 
                           OP_MEM(9) => OP_MEM_9_port, OP_MEM(8) => 
                           OP_MEM_8_port, OP_MEM(7) => OP_MEM_7_port, OP_MEM(6)
                           => OP_MEM_6_port, OP_MEM(5) => OP_MEM_5_port, 
                           OP_MEM(4) => OP_MEM_4_port, OP_MEM(3) => 
                           OP_MEM_3_port, OP_MEM(2) => OP_MEM_2_port, OP_MEM(1)
                           => OP_MEM_1_port, OP_MEM(0) => OP_MEM_0_port, 
                           OP_WB(31) => OP_WB_31_port, OP_WB(30) => 
                           OP_WB_30_port, OP_WB(29) => OP_WB_29_port, OP_WB(28)
                           => OP_WB_28_port, OP_WB(27) => OP_WB_27_port, 
                           OP_WB(26) => OP_WB_26_port, OP_WB(25) => 
                           OP_WB_25_port, OP_WB(24) => OP_WB_24_port, OP_WB(23)
                           => OP_WB_23_port, OP_WB(22) => OP_WB_22_port, 
                           OP_WB(21) => OP_WB_21_port, OP_WB(20) => 
                           OP_WB_20_port, OP_WB(19) => OP_WB_19_port, OP_WB(18)
                           => OP_WB_18_port, OP_WB(17) => OP_WB_17_port, 
                           OP_WB(16) => OP_WB_16_port, OP_WB(15) => 
                           OP_WB_15_port, OP_WB(14) => OP_WB_14_port, OP_WB(13)
                           => OP_WB_13_port, OP_WB(12) => OP_WB_12_port, 
                           OP_WB(11) => OP_WB_11_port, OP_WB(10) => 
                           OP_WB_10_port, OP_WB(9) => OP_WB_9_port, OP_WB(8) =>
                           OP_WB_8_port, OP_WB(7) => OP_WB_7_port, OP_WB(6) => 
                           OP_WB_6_port, OP_WB(5) => OP_WB_5_port, OP_WB(4) => 
                           OP_WB_4_port, OP_WB(3) => OP_WB_3_port, OP_WB(2) => 
                           OP_WB_2_port, OP_WB(1) => OP_WB_1_port, OP_WB(0) => 
                           OP_WB_0_port, PC_SEL(1) => PC_SEL_EX_1_port, 
                           PC_SEL(0) => PC_SEL_EX_0_port, ZERO_FLAG => 
                           ZERO_FLAG_EX, NPC_ABS(31) => NPC_ABS_EX_31_port, 
                           NPC_ABS(30) => NPC_ABS_EX_30_port, NPC_ABS(29) => 
                           NPC_ABS_EX_29_port, NPC_ABS(28) => 
                           NPC_ABS_EX_28_port, NPC_ABS(27) => 
                           NPC_ABS_EX_27_port, NPC_ABS(26) => 
                           NPC_ABS_EX_26_port, NPC_ABS(25) => 
                           NPC_ABS_EX_25_port, NPC_ABS(24) => 
                           NPC_ABS_EX_24_port, NPC_ABS(23) => 
                           NPC_ABS_EX_23_port, NPC_ABS(22) => 
                           NPC_ABS_EX_22_port, NPC_ABS(21) => 
                           NPC_ABS_EX_21_port, NPC_ABS(20) => 
                           NPC_ABS_EX_20_port, NPC_ABS(19) => 
                           NPC_ABS_EX_19_port, NPC_ABS(18) => 
                           NPC_ABS_EX_18_port, NPC_ABS(17) => 
                           NPC_ABS_EX_17_port, NPC_ABS(16) => 
                           NPC_ABS_EX_16_port, NPC_ABS(15) => 
                           NPC_ABS_EX_15_port, NPC_ABS(14) => 
                           NPC_ABS_EX_14_port, NPC_ABS(13) => 
                           NPC_ABS_EX_13_port, NPC_ABS(12) => 
                           NPC_ABS_EX_12_port, NPC_ABS(11) => 
                           NPC_ABS_EX_11_port, NPC_ABS(10) => 
                           NPC_ABS_EX_10_port, NPC_ABS(9) => NPC_ABS_EX_9_port,
                           NPC_ABS(8) => NPC_ABS_EX_8_port, NPC_ABS(7) => 
                           NPC_ABS_EX_7_port, NPC_ABS(6) => NPC_ABS_EX_6_port, 
                           NPC_ABS(5) => NPC_ABS_EX_5_port, NPC_ABS(4) => 
                           NPC_ABS_EX_4_port, NPC_ABS(3) => NPC_ABS_EX_3_port, 
                           NPC_ABS(2) => NPC_ABS_EX_2_port, NPC_ABS(1) => 
                           NPC_ABS_EX_1_port, NPC_ABS(0) => NPC_ABS_EX_0_port, 
                           NPC_REL(31) => NPC_REL_EX_31_port, NPC_REL(30) => 
                           NPC_REL_EX_30_port, NPC_REL(29) => 
                           NPC_REL_EX_29_port, NPC_REL(28) => 
                           NPC_REL_EX_28_port, NPC_REL(27) => 
                           NPC_REL_EX_27_port, NPC_REL(26) => 
                           NPC_REL_EX_26_port, NPC_REL(25) => 
                           NPC_REL_EX_25_port, NPC_REL(24) => 
                           NPC_REL_EX_24_port, NPC_REL(23) => 
                           NPC_REL_EX_23_port, NPC_REL(22) => 
                           NPC_REL_EX_22_port, NPC_REL(21) => 
                           NPC_REL_EX_21_port, NPC_REL(20) => 
                           NPC_REL_EX_20_port, NPC_REL(19) => 
                           NPC_REL_EX_19_port, NPC_REL(18) => 
                           NPC_REL_EX_18_port, NPC_REL(17) => 
                           NPC_REL_EX_17_port, NPC_REL(16) => 
                           NPC_REL_EX_16_port, NPC_REL(15) => 
                           NPC_REL_EX_15_port, NPC_REL(14) => 
                           NPC_REL_EX_14_port, NPC_REL(13) => 
                           NPC_REL_EX_13_port, NPC_REL(12) => 
                           NPC_REL_EX_12_port, NPC_REL(11) => 
                           NPC_REL_EX_11_port, NPC_REL(10) => 
                           NPC_REL_EX_10_port, NPC_REL(9) => NPC_REL_EX_9_port,
                           NPC_REL(8) => NPC_REL_EX_8_port, NPC_REL(7) => 
                           NPC_REL_EX_7_port, NPC_REL(6) => NPC_REL_EX_6_port, 
                           NPC_REL(5) => NPC_REL_EX_5_port, NPC_REL(4) => 
                           NPC_REL_EX_4_port, NPC_REL(3) => NPC_REL_EX_3_port, 
                           NPC_REL(2) => NPC_REL_EX_2_port, NPC_REL(1) => 
                           NPC_REL_EX_1_port, NPC_REL(0) => NPC_REL_EX_0_port, 
                           ALU_RES(31) => ALU_RES_EX_31_port, ALU_RES(30) => 
                           ALU_RES_EX_30_port, ALU_RES(29) => 
                           ALU_RES_EX_29_port, ALU_RES(28) => 
                           ALU_RES_EX_28_port, ALU_RES(27) => 
                           ALU_RES_EX_27_port, ALU_RES(26) => 
                           ALU_RES_EX_26_port, ALU_RES(25) => 
                           ALU_RES_EX_25_port, ALU_RES(24) => 
                           ALU_RES_EX_24_port, ALU_RES(23) => 
                           ALU_RES_EX_23_port, ALU_RES(22) => 
                           ALU_RES_EX_22_port, ALU_RES(21) => 
                           ALU_RES_EX_21_port, ALU_RES(20) => 
                           ALU_RES_EX_20_port, ALU_RES(19) => 
                           ALU_RES_EX_19_port, ALU_RES(18) => 
                           ALU_RES_EX_18_port, ALU_RES(17) => 
                           ALU_RES_EX_17_port, ALU_RES(16) => 
                           ALU_RES_EX_16_port, ALU_RES(15) => 
                           ALU_RES_EX_15_port, ALU_RES(14) => 
                           ALU_RES_EX_14_port, ALU_RES(13) => 
                           ALU_RES_EX_13_port, ALU_RES(12) => 
                           ALU_RES_EX_12_port, ALU_RES(11) => 
                           ALU_RES_EX_11_port, ALU_RES(10) => 
                           ALU_RES_EX_10_port, ALU_RES(9) => ALU_RES_EX_9_port,
                           ALU_RES(8) => ALU_RES_EX_8_port, ALU_RES(7) => 
                           ALU_RES_EX_7_port, ALU_RES(6) => ALU_RES_EX_6_port, 
                           ALU_RES(5) => ALU_RES_EX_5_port, ALU_RES(4) => 
                           ALU_RES_EX_4_port, ALU_RES(3) => ALU_RES_EX_3_port, 
                           ALU_RES(2) => ALU_RES_EX_2_port, ALU_RES(1) => 
                           ALU_RES_EX_1_port, ALU_RES(0) => ALU_RES_EX_0_port, 
                           B_OUT(31) => B_EX_OUT_31_port, B_OUT(30) => 
                           B_EX_OUT_30_port, B_OUT(29) => B_EX_OUT_29_port, 
                           B_OUT(28) => B_EX_OUT_28_port, B_OUT(27) => 
                           B_EX_OUT_27_port, B_OUT(26) => B_EX_OUT_26_port, 
                           B_OUT(25) => B_EX_OUT_25_port, B_OUT(24) => 
                           B_EX_OUT_24_port, B_OUT(23) => B_EX_OUT_23_port, 
                           B_OUT(22) => B_EX_OUT_22_port, B_OUT(21) => 
                           B_EX_OUT_21_port, B_OUT(20) => B_EX_OUT_20_port, 
                           B_OUT(19) => B_EX_OUT_19_port, B_OUT(18) => 
                           B_EX_OUT_18_port, B_OUT(17) => B_EX_OUT_17_port, 
                           B_OUT(16) => B_EX_OUT_16_port, B_OUT(15) => 
                           B_EX_OUT_15_port, B_OUT(14) => B_EX_OUT_14_port, 
                           B_OUT(13) => B_EX_OUT_13_port, B_OUT(12) => 
                           B_EX_OUT_12_port, B_OUT(11) => B_EX_OUT_11_port, 
                           B_OUT(10) => B_EX_OUT_10_port, B_OUT(9) => 
                           B_EX_OUT_9_port, B_OUT(8) => B_EX_OUT_8_port, 
                           B_OUT(7) => B_EX_OUT_7_port, B_OUT(6) => 
                           B_EX_OUT_6_port, B_OUT(5) => B_EX_OUT_5_port, 
                           B_OUT(4) => B_EX_OUT_4_port, B_OUT(3) => 
                           B_EX_OUT_3_port, B_OUT(2) => B_EX_OUT_2_port, 
                           B_OUT(1) => B_EX_OUT_1_port, B_OUT(0) => 
                           B_EX_OUT_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_EX_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_EX_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_EX_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_EX_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_EX_OUT_0_port);
   DRAM_R_ff : ff_0 port map( D => DRAM_R_IN, CLK => CLK, EN => X_Logic1_port, 
                           RST => RST, Q => DRAM_R_MEM);
   MemoryStage : Memory port map( CLK => CLK, RST => RST, MEM_EN_IN => 
                           MEM_EN_IN, DRAM_R_IN => DRAM_R_MEM, DRAM_W_IN => 
                           DRAM_W_IN, DRAM_EN_IN => DRAM_EN_IN, PC_SEL(1) => 
                           PC_SEL_EX_1_port, PC_SEL(0) => PC_SEL_EX_0_port, 
                           NPC_IN(31) => NPC_FETCH_OUT_31_port, NPC_IN(30) => 
                           NPC_FETCH_OUT_30_port, NPC_IN(29) => 
                           NPC_FETCH_OUT_29_port, NPC_IN(28) => 
                           NPC_FETCH_OUT_28_port, NPC_IN(27) => 
                           NPC_FETCH_OUT_27_port, NPC_IN(26) => 
                           NPC_FETCH_OUT_26_port, NPC_IN(25) => 
                           NPC_FETCH_OUT_25_port, NPC_IN(24) => 
                           NPC_FETCH_OUT_24_port, NPC_IN(23) => 
                           NPC_FETCH_OUT_23_port, NPC_IN(22) => 
                           NPC_FETCH_OUT_22_port, NPC_IN(21) => 
                           NPC_FETCH_OUT_21_port, NPC_IN(20) => 
                           NPC_FETCH_OUT_20_port, NPC_IN(19) => 
                           NPC_FETCH_OUT_19_port, NPC_IN(18) => 
                           NPC_FETCH_OUT_18_port, NPC_IN(17) => 
                           NPC_FETCH_OUT_17_port, NPC_IN(16) => 
                           NPC_FETCH_OUT_16_port, NPC_IN(15) => 
                           NPC_FETCH_OUT_15_port, NPC_IN(14) => 
                           NPC_FETCH_OUT_14_port, NPC_IN(13) => 
                           NPC_FETCH_OUT_13_port, NPC_IN(12) => 
                           NPC_FETCH_OUT_12_port, NPC_IN(11) => 
                           NPC_FETCH_OUT_11_port, NPC_IN(10) => 
                           NPC_FETCH_OUT_10_port, NPC_IN(9) => 
                           NPC_FETCH_OUT_9_port, NPC_IN(8) => 
                           NPC_FETCH_OUT_8_port, NPC_IN(7) => 
                           NPC_FETCH_OUT_7_port, NPC_IN(6) => 
                           NPC_FETCH_OUT_6_port, NPC_IN(5) => 
                           NPC_FETCH_OUT_5_port, NPC_IN(4) => 
                           NPC_FETCH_OUT_4_port, NPC_IN(3) => 
                           NPC_FETCH_OUT_3_port, NPC_IN(2) => 
                           NPC_FETCH_OUT_2_port, NPC_IN(1) => 
                           NPC_FETCH_OUT_1_port, NPC_IN(0) => 
                           NPC_FETCH_OUT_0_port, NPC_ABS(31) => 
                           NPC_ABS_EX_31_port, NPC_ABS(30) => 
                           NPC_ABS_EX_30_port, NPC_ABS(29) => 
                           NPC_ABS_EX_29_port, NPC_ABS(28) => 
                           NPC_ABS_EX_28_port, NPC_ABS(27) => 
                           NPC_ABS_EX_27_port, NPC_ABS(26) => 
                           NPC_ABS_EX_26_port, NPC_ABS(25) => 
                           NPC_ABS_EX_25_port, NPC_ABS(24) => 
                           NPC_ABS_EX_24_port, NPC_ABS(23) => 
                           NPC_ABS_EX_23_port, NPC_ABS(22) => 
                           NPC_ABS_EX_22_port, NPC_ABS(21) => 
                           NPC_ABS_EX_21_port, NPC_ABS(20) => 
                           NPC_ABS_EX_20_port, NPC_ABS(19) => 
                           NPC_ABS_EX_19_port, NPC_ABS(18) => 
                           NPC_ABS_EX_18_port, NPC_ABS(17) => 
                           NPC_ABS_EX_17_port, NPC_ABS(16) => 
                           NPC_ABS_EX_16_port, NPC_ABS(15) => 
                           NPC_ABS_EX_15_port, NPC_ABS(14) => 
                           NPC_ABS_EX_14_port, NPC_ABS(13) => 
                           NPC_ABS_EX_13_port, NPC_ABS(12) => 
                           NPC_ABS_EX_12_port, NPC_ABS(11) => 
                           NPC_ABS_EX_11_port, NPC_ABS(10) => 
                           NPC_ABS_EX_10_port, NPC_ABS(9) => NPC_ABS_EX_9_port,
                           NPC_ABS(8) => NPC_ABS_EX_8_port, NPC_ABS(7) => 
                           NPC_ABS_EX_7_port, NPC_ABS(6) => NPC_ABS_EX_6_port, 
                           NPC_ABS(5) => NPC_ABS_EX_5_port, NPC_ABS(4) => 
                           NPC_ABS_EX_4_port, NPC_ABS(3) => NPC_ABS_EX_3_port, 
                           NPC_ABS(2) => NPC_ABS_EX_2_port, NPC_ABS(1) => 
                           NPC_ABS_EX_1_port, NPC_ABS(0) => NPC_ABS_EX_0_port, 
                           NPC_REL(31) => NPC_REL_EX_31_port, NPC_REL(30) => 
                           NPC_REL_EX_30_port, NPC_REL(29) => 
                           NPC_REL_EX_29_port, NPC_REL(28) => 
                           NPC_REL_EX_28_port, NPC_REL(27) => 
                           NPC_REL_EX_27_port, NPC_REL(26) => 
                           NPC_REL_EX_26_port, NPC_REL(25) => 
                           NPC_REL_EX_25_port, NPC_REL(24) => 
                           NPC_REL_EX_24_port, NPC_REL(23) => 
                           NPC_REL_EX_23_port, NPC_REL(22) => 
                           NPC_REL_EX_22_port, NPC_REL(21) => 
                           NPC_REL_EX_21_port, NPC_REL(20) => 
                           NPC_REL_EX_20_port, NPC_REL(19) => 
                           NPC_REL_EX_19_port, NPC_REL(18) => 
                           NPC_REL_EX_18_port, NPC_REL(17) => 
                           NPC_REL_EX_17_port, NPC_REL(16) => 
                           NPC_REL_EX_16_port, NPC_REL(15) => 
                           NPC_REL_EX_15_port, NPC_REL(14) => 
                           NPC_REL_EX_14_port, NPC_REL(13) => 
                           NPC_REL_EX_13_port, NPC_REL(12) => 
                           NPC_REL_EX_12_port, NPC_REL(11) => 
                           NPC_REL_EX_11_port, NPC_REL(10) => 
                           NPC_REL_EX_10_port, NPC_REL(9) => NPC_REL_EX_9_port,
                           NPC_REL(8) => NPC_REL_EX_8_port, NPC_REL(7) => 
                           NPC_REL_EX_7_port, NPC_REL(6) => NPC_REL_EX_6_port, 
                           NPC_REL(5) => NPC_REL_EX_5_port, NPC_REL(4) => 
                           NPC_REL_EX_4_port, NPC_REL(3) => NPC_REL_EX_3_port, 
                           NPC_REL(2) => NPC_REL_EX_2_port, NPC_REL(1) => 
                           NPC_REL_EX_1_port, NPC_REL(0) => NPC_REL_EX_0_port, 
                           ALU_RES_IN(31) => ALU_RES_EX_31_port, ALU_RES_IN(30)
                           => ALU_RES_EX_30_port, ALU_RES_IN(29) => 
                           ALU_RES_EX_29_port, ALU_RES_IN(28) => 
                           ALU_RES_EX_28_port, ALU_RES_IN(27) => 
                           ALU_RES_EX_27_port, ALU_RES_IN(26) => 
                           ALU_RES_EX_26_port, ALU_RES_IN(25) => 
                           ALU_RES_EX_25_port, ALU_RES_IN(24) => 
                           ALU_RES_EX_24_port, ALU_RES_IN(23) => 
                           ALU_RES_EX_23_port, ALU_RES_IN(22) => 
                           ALU_RES_EX_22_port, ALU_RES_IN(21) => 
                           ALU_RES_EX_21_port, ALU_RES_IN(20) => 
                           ALU_RES_EX_20_port, ALU_RES_IN(19) => 
                           ALU_RES_EX_19_port, ALU_RES_IN(18) => 
                           ALU_RES_EX_18_port, ALU_RES_IN(17) => 
                           ALU_RES_EX_17_port, ALU_RES_IN(16) => 
                           ALU_RES_EX_16_port, ALU_RES_IN(15) => 
                           ALU_RES_EX_15_port, ALU_RES_IN(14) => 
                           ALU_RES_EX_14_port, ALU_RES_IN(13) => 
                           ALU_RES_EX_13_port, ALU_RES_IN(12) => 
                           ALU_RES_EX_12_port, ALU_RES_IN(11) => 
                           ALU_RES_EX_11_port, ALU_RES_IN(10) => 
                           ALU_RES_EX_10_port, ALU_RES_IN(9) => 
                           ALU_RES_EX_9_port, ALU_RES_IN(8) => 
                           ALU_RES_EX_8_port, ALU_RES_IN(7) => 
                           ALU_RES_EX_7_port, ALU_RES_IN(6) => 
                           ALU_RES_EX_6_port, ALU_RES_IN(5) => 
                           ALU_RES_EX_5_port, ALU_RES_IN(4) => 
                           ALU_RES_EX_4_port, ALU_RES_IN(3) => 
                           ALU_RES_EX_3_port, ALU_RES_IN(2) => 
                           ALU_RES_EX_2_port, ALU_RES_IN(1) => 
                           ALU_RES_EX_1_port, ALU_RES_IN(0) => 
                           ALU_RES_EX_0_port, B_IN(31) => B_EX_OUT_31_port, 
                           B_IN(30) => B_EX_OUT_30_port, B_IN(29) => 
                           B_EX_OUT_29_port, B_IN(28) => B_EX_OUT_28_port, 
                           B_IN(27) => B_EX_OUT_27_port, B_IN(26) => 
                           B_EX_OUT_26_port, B_IN(25) => B_EX_OUT_25_port, 
                           B_IN(24) => B_EX_OUT_24_port, B_IN(23) => 
                           B_EX_OUT_23_port, B_IN(22) => B_EX_OUT_22_port, 
                           B_IN(21) => B_EX_OUT_21_port, B_IN(20) => 
                           B_EX_OUT_20_port, B_IN(19) => B_EX_OUT_19_port, 
                           B_IN(18) => B_EX_OUT_18_port, B_IN(17) => 
                           B_EX_OUT_17_port, B_IN(16) => B_EX_OUT_16_port, 
                           B_IN(15) => B_EX_OUT_15_port, B_IN(14) => 
                           B_EX_OUT_14_port, B_IN(13) => B_EX_OUT_13_port, 
                           B_IN(12) => B_EX_OUT_12_port, B_IN(11) => 
                           B_EX_OUT_11_port, B_IN(10) => B_EX_OUT_10_port, 
                           B_IN(9) => B_EX_OUT_9_port, B_IN(8) => 
                           B_EX_OUT_8_port, B_IN(7) => B_EX_OUT_7_port, B_IN(6)
                           => B_EX_OUT_6_port, B_IN(5) => B_EX_OUT_5_port, 
                           B_IN(4) => B_EX_OUT_4_port, B_IN(3) => 
                           B_EX_OUT_3_port, B_IN(2) => B_EX_OUT_2_port, B_IN(1)
                           => B_EX_OUT_1_port, B_IN(0) => B_EX_OUT_0_port, 
                           ADD_WR_IN(4) => ADD_WR_EX_OUT_4_port, ADD_WR_IN(3) 
                           => ADD_WR_EX_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_EX_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_EX_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_EX_OUT_0_port, DRAM_DATA_IN(31) => 
                           DATA_IN(31), DRAM_DATA_IN(30) => DATA_IN(30), 
                           DRAM_DATA_IN(29) => DATA_IN(29), DRAM_DATA_IN(28) =>
                           DATA_IN(28), DRAM_DATA_IN(27) => DATA_IN(27), 
                           DRAM_DATA_IN(26) => DATA_IN(26), DRAM_DATA_IN(25) =>
                           DATA_IN(25), DRAM_DATA_IN(24) => DATA_IN(24), 
                           DRAM_DATA_IN(23) => DATA_IN(23), DRAM_DATA_IN(22) =>
                           DATA_IN(22), DRAM_DATA_IN(21) => DATA_IN(21), 
                           DRAM_DATA_IN(20) => DATA_IN(20), DRAM_DATA_IN(19) =>
                           DATA_IN(19), DRAM_DATA_IN(18) => DATA_IN(18), 
                           DRAM_DATA_IN(17) => DATA_IN(17), DRAM_DATA_IN(16) =>
                           DATA_IN(16), DRAM_DATA_IN(15) => DATA_IN(15), 
                           DRAM_DATA_IN(14) => DATA_IN(14), DRAM_DATA_IN(13) =>
                           DATA_IN(13), DRAM_DATA_IN(12) => DATA_IN(12), 
                           DRAM_DATA_IN(11) => DATA_IN(11), DRAM_DATA_IN(10) =>
                           DATA_IN(10), DRAM_DATA_IN(9) => DATA_IN(9), 
                           DRAM_DATA_IN(8) => DATA_IN(8), DRAM_DATA_IN(7) => 
                           DATA_IN(7), DRAM_DATA_IN(6) => DATA_IN(6), 
                           DRAM_DATA_IN(5) => DATA_IN(5), DRAM_DATA_IN(4) => 
                           DATA_IN(4), DRAM_DATA_IN(3) => DATA_IN(3), 
                           DRAM_DATA_IN(2) => DATA_IN(2), DRAM_DATA_IN(1) => 
                           DATA_IN(1), DRAM_DATA_IN(0) => DATA_IN(0), 
                           PC_OUT(31) => PC_MEM_OUT_31_port, PC_OUT(30) => 
                           PC_MEM_OUT_30_port, PC_OUT(29) => PC_MEM_OUT_29_port
                           , PC_OUT(28) => PC_MEM_OUT_28_port, PC_OUT(27) => 
                           PC_MEM_OUT_27_port, PC_OUT(26) => PC_MEM_OUT_26_port
                           , PC_OUT(25) => PC_MEM_OUT_25_port, PC_OUT(24) => 
                           PC_MEM_OUT_24_port, PC_OUT(23) => PC_MEM_OUT_23_port
                           , PC_OUT(22) => PC_MEM_OUT_22_port, PC_OUT(21) => 
                           PC_MEM_OUT_21_port, PC_OUT(20) => PC_MEM_OUT_20_port
                           , PC_OUT(19) => PC_MEM_OUT_19_port, PC_OUT(18) => 
                           PC_MEM_OUT_18_port, PC_OUT(17) => PC_MEM_OUT_17_port
                           , PC_OUT(16) => PC_MEM_OUT_16_port, PC_OUT(15) => 
                           PC_MEM_OUT_15_port, PC_OUT(14) => PC_MEM_OUT_14_port
                           , PC_OUT(13) => PC_MEM_OUT_13_port, PC_OUT(12) => 
                           PC_MEM_OUT_12_port, PC_OUT(11) => PC_MEM_OUT_11_port
                           , PC_OUT(10) => PC_MEM_OUT_10_port, PC_OUT(9) => 
                           PC_MEM_OUT_9_port, PC_OUT(8) => PC_MEM_OUT_8_port, 
                           PC_OUT(7) => PC_MEM_OUT_7_port, PC_OUT(6) => 
                           PC_MEM_OUT_6_port, PC_OUT(5) => PC_MEM_OUT_5_port, 
                           PC_OUT(4) => PC_MEM_OUT_4_port, PC_OUT(3) => 
                           PC_MEM_OUT_3_port, PC_OUT(2) => PC_MEM_OUT_2_port, 
                           PC_OUT(1) => PC_MEM_OUT_1_port, PC_OUT(0) => 
                           PC_MEM_OUT_0_port, DRAM_EN_OUT => DRAM_EN_OUT, 
                           DRAM_R_OUT => DRAM_R_OUT, DRAM_W_OUT => DRAM_W_OUT, 
                           DRAM_ADDR_OUT(31) => DRAM_ADDR_OUT(31), 
                           DRAM_ADDR_OUT(30) => DRAM_ADDR_OUT(30), 
                           DRAM_ADDR_OUT(29) => DRAM_ADDR_OUT(29), 
                           DRAM_ADDR_OUT(28) => DRAM_ADDR_OUT(28), 
                           DRAM_ADDR_OUT(27) => DRAM_ADDR_OUT(27), 
                           DRAM_ADDR_OUT(26) => DRAM_ADDR_OUT(26), 
                           DRAM_ADDR_OUT(25) => DRAM_ADDR_OUT(25), 
                           DRAM_ADDR_OUT(24) => DRAM_ADDR_OUT(24), 
                           DRAM_ADDR_OUT(23) => DRAM_ADDR_OUT(23), 
                           DRAM_ADDR_OUT(22) => DRAM_ADDR_OUT(22), 
                           DRAM_ADDR_OUT(21) => DRAM_ADDR_OUT(21), 
                           DRAM_ADDR_OUT(20) => DRAM_ADDR_OUT(20), 
                           DRAM_ADDR_OUT(19) => DRAM_ADDR_OUT(19), 
                           DRAM_ADDR_OUT(18) => DRAM_ADDR_OUT(18), 
                           DRAM_ADDR_OUT(17) => DRAM_ADDR_OUT(17), 
                           DRAM_ADDR_OUT(16) => DRAM_ADDR_OUT(16), 
                           DRAM_ADDR_OUT(15) => DRAM_ADDR_OUT(15), 
                           DRAM_ADDR_OUT(14) => DRAM_ADDR_OUT(14), 
                           DRAM_ADDR_OUT(13) => DRAM_ADDR_OUT(13), 
                           DRAM_ADDR_OUT(12) => DRAM_ADDR_OUT(12), 
                           DRAM_ADDR_OUT(11) => DRAM_ADDR_OUT(11), 
                           DRAM_ADDR_OUT(10) => DRAM_ADDR_OUT(10), 
                           DRAM_ADDR_OUT(9) => DRAM_ADDR_OUT(9), 
                           DRAM_ADDR_OUT(8) => DRAM_ADDR_OUT(8), 
                           DRAM_ADDR_OUT(7) => DRAM_ADDR_OUT(7), 
                           DRAM_ADDR_OUT(6) => DRAM_ADDR_OUT(6), 
                           DRAM_ADDR_OUT(5) => DRAM_ADDR_OUT(5), 
                           DRAM_ADDR_OUT(4) => DRAM_ADDR_OUT(4), 
                           DRAM_ADDR_OUT(3) => DRAM_ADDR_OUT(3), 
                           DRAM_ADDR_OUT(2) => DRAM_ADDR_OUT(2), 
                           DRAM_ADDR_OUT(1) => DRAM_ADDR_OUT(1), 
                           DRAM_ADDR_OUT(0) => DRAM_ADDR_OUT(0), 
                           DRAM_DATA_OUT(31) => DATA_OUT(31), DRAM_DATA_OUT(30)
                           => DATA_OUT(30), DRAM_DATA_OUT(29) => DATA_OUT(29), 
                           DRAM_DATA_OUT(28) => DATA_OUT(28), DRAM_DATA_OUT(27)
                           => DATA_OUT(27), DRAM_DATA_OUT(26) => DATA_OUT(26), 
                           DRAM_DATA_OUT(25) => DATA_OUT(25), DRAM_DATA_OUT(24)
                           => DATA_OUT(24), DRAM_DATA_OUT(23) => DATA_OUT(23), 
                           DRAM_DATA_OUT(22) => DATA_OUT(22), DRAM_DATA_OUT(21)
                           => DATA_OUT(21), DRAM_DATA_OUT(20) => DATA_OUT(20), 
                           DRAM_DATA_OUT(19) => DATA_OUT(19), DRAM_DATA_OUT(18)
                           => DATA_OUT(18), DRAM_DATA_OUT(17) => DATA_OUT(17), 
                           DRAM_DATA_OUT(16) => DATA_OUT(16), DRAM_DATA_OUT(15)
                           => DATA_OUT(15), DRAM_DATA_OUT(14) => DATA_OUT(14), 
                           DRAM_DATA_OUT(13) => DATA_OUT(13), DRAM_DATA_OUT(12)
                           => DATA_OUT(12), DRAM_DATA_OUT(11) => DATA_OUT(11), 
                           DRAM_DATA_OUT(10) => DATA_OUT(10), DRAM_DATA_OUT(9) 
                           => DATA_OUT(9), DRAM_DATA_OUT(8) => DATA_OUT(8), 
                           DRAM_DATA_OUT(7) => DATA_OUT(7), DRAM_DATA_OUT(6) =>
                           DATA_OUT(6), DRAM_DATA_OUT(5) => DATA_OUT(5), 
                           DRAM_DATA_OUT(4) => DATA_OUT(4), DRAM_DATA_OUT(3) =>
                           DATA_OUT(3), DRAM_DATA_OUT(2) => DATA_OUT(2), 
                           DRAM_DATA_OUT(1) => DATA_OUT(1), DRAM_DATA_OUT(0) =>
                           DATA_OUT(0), DATA_OUT(31) => DATA_MEM_OUT_31_port, 
                           DATA_OUT(30) => DATA_MEM_OUT_30_port, DATA_OUT(29) 
                           => DATA_MEM_OUT_29_port, DATA_OUT(28) => 
                           DATA_MEM_OUT_28_port, DATA_OUT(27) => 
                           DATA_MEM_OUT_27_port, DATA_OUT(26) => 
                           DATA_MEM_OUT_26_port, DATA_OUT(25) => 
                           DATA_MEM_OUT_25_port, DATA_OUT(24) => 
                           DATA_MEM_OUT_24_port, DATA_OUT(23) => 
                           DATA_MEM_OUT_23_port, DATA_OUT(22) => 
                           DATA_MEM_OUT_22_port, DATA_OUT(21) => 
                           DATA_MEM_OUT_21_port, DATA_OUT(20) => 
                           DATA_MEM_OUT_20_port, DATA_OUT(19) => 
                           DATA_MEM_OUT_19_port, DATA_OUT(18) => 
                           DATA_MEM_OUT_18_port, DATA_OUT(17) => 
                           DATA_MEM_OUT_17_port, DATA_OUT(16) => 
                           DATA_MEM_OUT_16_port, DATA_OUT(15) => 
                           DATA_MEM_OUT_15_port, DATA_OUT(14) => 
                           DATA_MEM_OUT_14_port, DATA_OUT(13) => 
                           DATA_MEM_OUT_13_port, DATA_OUT(12) => 
                           DATA_MEM_OUT_12_port, DATA_OUT(11) => 
                           DATA_MEM_OUT_11_port, DATA_OUT(10) => 
                           DATA_MEM_OUT_10_port, DATA_OUT(9) => 
                           DATA_MEM_OUT_9_port, DATA_OUT(8) => 
                           DATA_MEM_OUT_8_port, DATA_OUT(7) => 
                           DATA_MEM_OUT_7_port, DATA_OUT(6) => 
                           DATA_MEM_OUT_6_port, DATA_OUT(5) => 
                           DATA_MEM_OUT_5_port, DATA_OUT(4) => 
                           DATA_MEM_OUT_4_port, DATA_OUT(3) => 
                           DATA_MEM_OUT_3_port, DATA_OUT(2) => 
                           DATA_MEM_OUT_2_port, DATA_OUT(1) => 
                           DATA_MEM_OUT_1_port, DATA_OUT(0) => 
                           DATA_MEM_OUT_0_port, ALU_RES_OUT(31) => 
                           ALU_RES_MEM_31_port, ALU_RES_OUT(30) => 
                           ALU_RES_MEM_30_port, ALU_RES_OUT(29) => 
                           ALU_RES_MEM_29_port, ALU_RES_OUT(28) => 
                           ALU_RES_MEM_28_port, ALU_RES_OUT(27) => 
                           ALU_RES_MEM_27_port, ALU_RES_OUT(26) => 
                           ALU_RES_MEM_26_port, ALU_RES_OUT(25) => 
                           ALU_RES_MEM_25_port, ALU_RES_OUT(24) => 
                           ALU_RES_MEM_24_port, ALU_RES_OUT(23) => 
                           ALU_RES_MEM_23_port, ALU_RES_OUT(22) => 
                           ALU_RES_MEM_22_port, ALU_RES_OUT(21) => 
                           ALU_RES_MEM_21_port, ALU_RES_OUT(20) => 
                           ALU_RES_MEM_20_port, ALU_RES_OUT(19) => 
                           ALU_RES_MEM_19_port, ALU_RES_OUT(18) => 
                           ALU_RES_MEM_18_port, ALU_RES_OUT(17) => 
                           ALU_RES_MEM_17_port, ALU_RES_OUT(16) => 
                           ALU_RES_MEM_16_port, ALU_RES_OUT(15) => 
                           ALU_RES_MEM_15_port, ALU_RES_OUT(14) => 
                           ALU_RES_MEM_14_port, ALU_RES_OUT(13) => 
                           ALU_RES_MEM_13_port, ALU_RES_OUT(12) => 
                           ALU_RES_MEM_12_port, ALU_RES_OUT(11) => 
                           ALU_RES_MEM_11_port, ALU_RES_OUT(10) => 
                           ALU_RES_MEM_10_port, ALU_RES_OUT(9) => 
                           ALU_RES_MEM_9_port, ALU_RES_OUT(8) => 
                           ALU_RES_MEM_8_port, ALU_RES_OUT(7) => 
                           ALU_RES_MEM_7_port, ALU_RES_OUT(6) => 
                           ALU_RES_MEM_6_port, ALU_RES_OUT(5) => 
                           ALU_RES_MEM_5_port, ALU_RES_OUT(4) => 
                           ALU_RES_MEM_4_port, ALU_RES_OUT(3) => 
                           ALU_RES_MEM_3_port, ALU_RES_OUT(2) => 
                           ALU_RES_MEM_2_port, ALU_RES_OUT(1) => 
                           ALU_RES_MEM_1_port, ALU_RES_OUT(0) => 
                           ALU_RES_MEM_0_port, OP_MEM(31) => OP_MEM_31_port, 
                           OP_MEM(30) => OP_MEM_30_port, OP_MEM(29) => 
                           OP_MEM_29_port, OP_MEM(28) => OP_MEM_28_port, 
                           OP_MEM(27) => OP_MEM_27_port, OP_MEM(26) => 
                           OP_MEM_26_port, OP_MEM(25) => OP_MEM_25_port, 
                           OP_MEM(24) => OP_MEM_24_port, OP_MEM(23) => 
                           OP_MEM_23_port, OP_MEM(22) => OP_MEM_22_port, 
                           OP_MEM(21) => OP_MEM_21_port, OP_MEM(20) => 
                           OP_MEM_20_port, OP_MEM(19) => OP_MEM_19_port, 
                           OP_MEM(18) => OP_MEM_18_port, OP_MEM(17) => 
                           OP_MEM_17_port, OP_MEM(16) => OP_MEM_16_port, 
                           OP_MEM(15) => OP_MEM_15_port, OP_MEM(14) => 
                           OP_MEM_14_port, OP_MEM(13) => OP_MEM_13_port, 
                           OP_MEM(12) => OP_MEM_12_port, OP_MEM(11) => 
                           OP_MEM_11_port, OP_MEM(10) => OP_MEM_10_port, 
                           OP_MEM(9) => OP_MEM_9_port, OP_MEM(8) => 
                           OP_MEM_8_port, OP_MEM(7) => OP_MEM_7_port, OP_MEM(6)
                           => OP_MEM_6_port, OP_MEM(5) => OP_MEM_5_port, 
                           OP_MEM(4) => OP_MEM_4_port, OP_MEM(3) => 
                           OP_MEM_3_port, OP_MEM(2) => OP_MEM_2_port, OP_MEM(1)
                           => OP_MEM_1_port, OP_MEM(0) => OP_MEM_0_port, 
                           ADD_WR_MEM(4) => ADD_WR_MEM_4_port, ADD_WR_MEM(3) =>
                           ADD_WR_MEM_3_port, ADD_WR_MEM(2) => 
                           ADD_WR_MEM_2_port, ADD_WR_MEM(1) => 
                           ADD_WR_MEM_1_port, ADD_WR_MEM(0) => 
                           ADD_WR_MEM_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_MEM_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_MEM_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_MEM_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_MEM_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_MEM_OUT_0_port);
   RF_WE_ff : ff_2 port map( D => RF_WE, CLK => CLK, EN => X_Logic1_port, RST 
                           => RST, Q => RF_WE_WB);
   WritebackStage : Writeback port map( WB_MUX_SEL => WB_MUX_SEL, DATA_IN(31) 
                           => DATA_MEM_OUT_31_port, DATA_IN(30) => 
                           DATA_MEM_OUT_30_port, DATA_IN(29) => 
                           DATA_MEM_OUT_29_port, DATA_IN(28) => 
                           DATA_MEM_OUT_28_port, DATA_IN(27) => 
                           DATA_MEM_OUT_27_port, DATA_IN(26) => 
                           DATA_MEM_OUT_26_port, DATA_IN(25) => 
                           DATA_MEM_OUT_25_port, DATA_IN(24) => 
                           DATA_MEM_OUT_24_port, DATA_IN(23) => 
                           DATA_MEM_OUT_23_port, DATA_IN(22) => 
                           DATA_MEM_OUT_22_port, DATA_IN(21) => 
                           DATA_MEM_OUT_21_port, DATA_IN(20) => 
                           DATA_MEM_OUT_20_port, DATA_IN(19) => 
                           DATA_MEM_OUT_19_port, DATA_IN(18) => 
                           DATA_MEM_OUT_18_port, DATA_IN(17) => 
                           DATA_MEM_OUT_17_port, DATA_IN(16) => 
                           DATA_MEM_OUT_16_port, DATA_IN(15) => 
                           DATA_MEM_OUT_15_port, DATA_IN(14) => 
                           DATA_MEM_OUT_14_port, DATA_IN(13) => 
                           DATA_MEM_OUT_13_port, DATA_IN(12) => 
                           DATA_MEM_OUT_12_port, DATA_IN(11) => 
                           DATA_MEM_OUT_11_port, DATA_IN(10) => 
                           DATA_MEM_OUT_10_port, DATA_IN(9) => 
                           DATA_MEM_OUT_9_port, DATA_IN(8) => 
                           DATA_MEM_OUT_8_port, DATA_IN(7) => 
                           DATA_MEM_OUT_7_port, DATA_IN(6) => 
                           DATA_MEM_OUT_6_port, DATA_IN(5) => 
                           DATA_MEM_OUT_5_port, DATA_IN(4) => 
                           DATA_MEM_OUT_4_port, DATA_IN(3) => 
                           DATA_MEM_OUT_3_port, DATA_IN(2) => 
                           DATA_MEM_OUT_2_port, DATA_IN(1) => 
                           DATA_MEM_OUT_1_port, DATA_IN(0) => 
                           DATA_MEM_OUT_0_port, ALU_RES_IN(31) => 
                           ALU_RES_MEM_31_port, ALU_RES_IN(30) => 
                           ALU_RES_MEM_30_port, ALU_RES_IN(29) => 
                           ALU_RES_MEM_29_port, ALU_RES_IN(28) => 
                           ALU_RES_MEM_28_port, ALU_RES_IN(27) => 
                           ALU_RES_MEM_27_port, ALU_RES_IN(26) => 
                           ALU_RES_MEM_26_port, ALU_RES_IN(25) => 
                           ALU_RES_MEM_25_port, ALU_RES_IN(24) => 
                           ALU_RES_MEM_24_port, ALU_RES_IN(23) => 
                           ALU_RES_MEM_23_port, ALU_RES_IN(22) => 
                           ALU_RES_MEM_22_port, ALU_RES_IN(21) => 
                           ALU_RES_MEM_21_port, ALU_RES_IN(20) => 
                           ALU_RES_MEM_20_port, ALU_RES_IN(19) => 
                           ALU_RES_MEM_19_port, ALU_RES_IN(18) => 
                           ALU_RES_MEM_18_port, ALU_RES_IN(17) => 
                           ALU_RES_MEM_17_port, ALU_RES_IN(16) => 
                           ALU_RES_MEM_16_port, ALU_RES_IN(15) => 
                           ALU_RES_MEM_15_port, ALU_RES_IN(14) => 
                           ALU_RES_MEM_14_port, ALU_RES_IN(13) => 
                           ALU_RES_MEM_13_port, ALU_RES_IN(12) => 
                           ALU_RES_MEM_12_port, ALU_RES_IN(11) => 
                           ALU_RES_MEM_11_port, ALU_RES_IN(10) => 
                           ALU_RES_MEM_10_port, ALU_RES_IN(9) => 
                           ALU_RES_MEM_9_port, ALU_RES_IN(8) => 
                           ALU_RES_MEM_8_port, ALU_RES_IN(7) => 
                           ALU_RES_MEM_7_port, ALU_RES_IN(6) => 
                           ALU_RES_MEM_6_port, ALU_RES_IN(5) => 
                           ALU_RES_MEM_5_port, ALU_RES_IN(4) => 
                           ALU_RES_MEM_4_port, ALU_RES_IN(3) => 
                           ALU_RES_MEM_3_port, ALU_RES_IN(2) => 
                           ALU_RES_MEM_2_port, ALU_RES_IN(1) => 
                           ALU_RES_MEM_1_port, ALU_RES_IN(0) => 
                           ALU_RES_MEM_0_port, ADD_WR_IN(4) => 
                           ADD_WR_MEM_OUT_4_port, ADD_WR_IN(3) => 
                           ADD_WR_MEM_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_MEM_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_MEM_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_MEM_OUT_0_port, DATA_OUT(31) => OP_WB_31_port
                           , DATA_OUT(30) => OP_WB_30_port, DATA_OUT(29) => 
                           OP_WB_29_port, DATA_OUT(28) => OP_WB_28_port, 
                           DATA_OUT(27) => OP_WB_27_port, DATA_OUT(26) => 
                           OP_WB_26_port, DATA_OUT(25) => OP_WB_25_port, 
                           DATA_OUT(24) => OP_WB_24_port, DATA_OUT(23) => 
                           OP_WB_23_port, DATA_OUT(22) => OP_WB_22_port, 
                           DATA_OUT(21) => OP_WB_21_port, DATA_OUT(20) => 
                           OP_WB_20_port, DATA_OUT(19) => OP_WB_19_port, 
                           DATA_OUT(18) => OP_WB_18_port, DATA_OUT(17) => 
                           OP_WB_17_port, DATA_OUT(16) => OP_WB_16_port, 
                           DATA_OUT(15) => OP_WB_15_port, DATA_OUT(14) => 
                           OP_WB_14_port, DATA_OUT(13) => OP_WB_13_port, 
                           DATA_OUT(12) => OP_WB_12_port, DATA_OUT(11) => 
                           OP_WB_11_port, DATA_OUT(10) => OP_WB_10_port, 
                           DATA_OUT(9) => OP_WB_9_port, DATA_OUT(8) => 
                           OP_WB_8_port, DATA_OUT(7) => OP_WB_7_port, 
                           DATA_OUT(6) => OP_WB_6_port, DATA_OUT(5) => 
                           OP_WB_5_port, DATA_OUT(4) => OP_WB_4_port, 
                           DATA_OUT(3) => OP_WB_3_port, DATA_OUT(2) => 
                           OP_WB_2_port, DATA_OUT(1) => OP_WB_1_port, 
                           DATA_OUT(0) => OP_WB_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_WB_4_port, ADD_WR_OUT(3) => ADD_WR_WB_3_port,
                           ADD_WR_OUT(2) => ADD_WR_WB_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_WB_1_port, ADD_WR_OUT(0) => ADD_WR_WB_0_port)
                           ;
   HDU : HazardDetection port map( RST => RST, ADD_RS1(4) => ADD_RS1_HDU_4_port
                           , ADD_RS1(3) => ADD_RS1_HDU_3_port, ADD_RS1(2) => 
                           ADD_RS1_HDU_2_port, ADD_RS1(1) => ADD_RS1_HDU_1_port
                           , ADD_RS1(0) => ADD_RS1_HDU_0_port, ADD_RS2(4) => 
                           ADD_RS2_HDU_4_port, ADD_RS2(3) => ADD_RS2_HDU_3_port
                           , ADD_RS2(2) => ADD_RS2_HDU_2_port, ADD_RS2(1) => 
                           ADD_RS2_HDU_1_port, ADD_RS2(0) => ADD_RS2_HDU_0_port
                           , ADD_WR(4) => ADD_WR_DECODE_OUT_4_port, ADD_WR(3) 
                           => ADD_WR_DECODE_OUT_3_port, ADD_WR(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR(0) => 
                           ADD_WR_DECODE_OUT_0_port, DRAM_R => DRAM_R_IN, 
                           INS_IN(31) => INS_OUT_31_port, INS_IN(30) => 
                           INS_OUT_30_port, INS_IN(29) => INS_OUT_29_port, 
                           INS_IN(28) => INS_OUT_28_port, INS_IN(27) => 
                           INS_OUT_27_port, INS_IN(26) => INS_OUT_26_port, 
                           INS_IN(25) => INS_OUT_25_port, INS_IN(24) => 
                           INS_OUT_24_port, INS_IN(23) => INS_OUT_23_port, 
                           INS_IN(22) => INS_OUT_22_port, INS_IN(21) => 
                           INS_OUT_21_port, INS_IN(20) => INS_OUT_20_port, 
                           INS_IN(19) => INS_OUT_19_port, INS_IN(18) => 
                           INS_OUT_18_port, INS_IN(17) => INS_OUT_17_port, 
                           INS_IN(16) => INS_OUT_16_port, INS_IN(15) => 
                           INS_OUT_15_port, INS_IN(14) => INS_OUT_14_port, 
                           INS_IN(13) => INS_OUT_13_port, INS_IN(12) => 
                           INS_OUT_12_port, INS_IN(11) => INS_OUT_11_port, 
                           INS_IN(10) => INS_OUT_10_port, INS_IN(9) => 
                           INS_OUT_9_port, INS_IN(8) => INS_OUT_8_port, 
                           INS_IN(7) => INS_OUT_7_port, INS_IN(6) => 
                           INS_OUT_6_port, INS_IN(5) => INS_OUT_5_port, 
                           INS_IN(4) => INS_OUT_4_port, INS_IN(3) => 
                           INS_OUT_3_port, INS_IN(2) => INS_OUT_2_port, 
                           INS_IN(1) => INS_OUT_1_port, INS_IN(0) => 
                           INS_OUT_0_port, PC_IN(31) => PC_FETCH_OUT_31_port, 
                           PC_IN(30) => PC_FETCH_OUT_30_port, PC_IN(29) => 
                           PC_FETCH_OUT_29_port, PC_IN(28) => 
                           PC_FETCH_OUT_28_port, PC_IN(27) => 
                           PC_FETCH_OUT_27_port, PC_IN(26) => 
                           PC_FETCH_OUT_26_port, PC_IN(25) => 
                           PC_FETCH_OUT_25_port, PC_IN(24) => 
                           PC_FETCH_OUT_24_port, PC_IN(23) => 
                           PC_FETCH_OUT_23_port, PC_IN(22) => 
                           PC_FETCH_OUT_22_port, PC_IN(21) => 
                           PC_FETCH_OUT_21_port, PC_IN(20) => 
                           PC_FETCH_OUT_20_port, PC_IN(19) => 
                           PC_FETCH_OUT_19_port, PC_IN(18) => 
                           PC_FETCH_OUT_18_port, PC_IN(17) => 
                           PC_FETCH_OUT_17_port, PC_IN(16) => 
                           PC_FETCH_OUT_16_port, PC_IN(15) => 
                           PC_FETCH_OUT_15_port, PC_IN(14) => 
                           PC_FETCH_OUT_14_port, PC_IN(13) => 
                           PC_FETCH_OUT_13_port, PC_IN(12) => 
                           PC_FETCH_OUT_12_port, PC_IN(11) => 
                           PC_FETCH_OUT_11_port, PC_IN(10) => 
                           PC_FETCH_OUT_10_port, PC_IN(9) => 
                           PC_FETCH_OUT_9_port, PC_IN(8) => PC_FETCH_OUT_8_port
                           , PC_IN(7) => PC_FETCH_OUT_7_port, PC_IN(6) => 
                           PC_FETCH_OUT_6_port, PC_IN(5) => PC_FETCH_OUT_5_port
                           , PC_IN(4) => PC_FETCH_OUT_4_port, PC_IN(3) => 
                           PC_FETCH_OUT_3_port, PC_IN(2) => PC_FETCH_OUT_2_port
                           , PC_IN(1) => PC_FETCH_OUT_1_port, PC_IN(0) => 
                           PC_FETCH_OUT_0_port, Bubble => Bubble_out_port, 
                           HDU_INS_OUT(31) => sig_HDU_INS_OUT_31_port, 
                           HDU_INS_OUT(30) => sig_HDU_INS_OUT_30_port, 
                           HDU_INS_OUT(29) => sig_HDU_INS_OUT_29_port, 
                           HDU_INS_OUT(28) => sig_HDU_INS_OUT_28_port, 
                           HDU_INS_OUT(27) => sig_HDU_INS_OUT_27_port, 
                           HDU_INS_OUT(26) => sig_HDU_INS_OUT_26_port, 
                           HDU_INS_OUT(25) => sig_HDU_INS_OUT_25_port, 
                           HDU_INS_OUT(24) => sig_HDU_INS_OUT_24_port, 
                           HDU_INS_OUT(23) => sig_HDU_INS_OUT_23_port, 
                           HDU_INS_OUT(22) => sig_HDU_INS_OUT_22_port, 
                           HDU_INS_OUT(21) => sig_HDU_INS_OUT_21_port, 
                           HDU_INS_OUT(20) => sig_HDU_INS_OUT_20_port, 
                           HDU_INS_OUT(19) => sig_HDU_INS_OUT_19_port, 
                           HDU_INS_OUT(18) => sig_HDU_INS_OUT_18_port, 
                           HDU_INS_OUT(17) => sig_HDU_INS_OUT_17_port, 
                           HDU_INS_OUT(16) => sig_HDU_INS_OUT_16_port, 
                           HDU_INS_OUT(15) => sig_HDU_INS_OUT_15_port, 
                           HDU_INS_OUT(14) => sig_HDU_INS_OUT_14_port, 
                           HDU_INS_OUT(13) => sig_HDU_INS_OUT_13_port, 
                           HDU_INS_OUT(12) => sig_HDU_INS_OUT_12_port, 
                           HDU_INS_OUT(11) => sig_HDU_INS_OUT_11_port, 
                           HDU_INS_OUT(10) => sig_HDU_INS_OUT_10_port, 
                           HDU_INS_OUT(9) => sig_HDU_INS_OUT_9_port, 
                           HDU_INS_OUT(8) => sig_HDU_INS_OUT_8_port, 
                           HDU_INS_OUT(7) => sig_HDU_INS_OUT_7_port, 
                           HDU_INS_OUT(6) => sig_HDU_INS_OUT_6_port, 
                           HDU_INS_OUT(5) => sig_HDU_INS_OUT_5_port, 
                           HDU_INS_OUT(4) => sig_HDU_INS_OUT_4_port, 
                           HDU_INS_OUT(3) => sig_HDU_INS_OUT_3_port, 
                           HDU_INS_OUT(2) => sig_HDU_INS_OUT_2_port, 
                           HDU_INS_OUT(1) => sig_HDU_INS_OUT_1_port, 
                           HDU_INS_OUT(0) => sig_HDU_INS_OUT_0_port, 
                           HDU_PC_OUT(31) => sig_HDU_PC_OUT_31_port, 
                           HDU_PC_OUT(30) => sig_HDU_PC_OUT_30_port, 
                           HDU_PC_OUT(29) => sig_HDU_PC_OUT_29_port, 
                           HDU_PC_OUT(28) => sig_HDU_PC_OUT_28_port, 
                           HDU_PC_OUT(27) => sig_HDU_PC_OUT_27_port, 
                           HDU_PC_OUT(26) => sig_HDU_PC_OUT_26_port, 
                           HDU_PC_OUT(25) => sig_HDU_PC_OUT_25_port, 
                           HDU_PC_OUT(24) => sig_HDU_PC_OUT_24_port, 
                           HDU_PC_OUT(23) => sig_HDU_PC_OUT_23_port, 
                           HDU_PC_OUT(22) => sig_HDU_PC_OUT_22_port, 
                           HDU_PC_OUT(21) => sig_HDU_PC_OUT_21_port, 
                           HDU_PC_OUT(20) => sig_HDU_PC_OUT_20_port, 
                           HDU_PC_OUT(19) => sig_HDU_PC_OUT_19_port, 
                           HDU_PC_OUT(18) => sig_HDU_PC_OUT_18_port, 
                           HDU_PC_OUT(17) => sig_HDU_PC_OUT_17_port, 
                           HDU_PC_OUT(16) => sig_HDU_PC_OUT_16_port, 
                           HDU_PC_OUT(15) => sig_HDU_PC_OUT_15_port, 
                           HDU_PC_OUT(14) => sig_HDU_PC_OUT_14_port, 
                           HDU_PC_OUT(13) => sig_HDU_PC_OUT_13_port, 
                           HDU_PC_OUT(12) => sig_HDU_PC_OUT_12_port, 
                           HDU_PC_OUT(11) => sig_HDU_PC_OUT_11_port, 
                           HDU_PC_OUT(10) => sig_HDU_PC_OUT_10_port, 
                           HDU_PC_OUT(9) => sig_HDU_PC_OUT_9_port, 
                           HDU_PC_OUT(8) => sig_HDU_PC_OUT_8_port, 
                           HDU_PC_OUT(7) => sig_HDU_PC_OUT_7_port, 
                           HDU_PC_OUT(6) => sig_HDU_PC_OUT_6_port, 
                           HDU_PC_OUT(5) => sig_HDU_PC_OUT_5_port, 
                           HDU_PC_OUT(4) => sig_HDU_PC_OUT_4_port, 
                           HDU_PC_OUT(3) => sig_HDU_PC_OUT_3_port, 
                           HDU_PC_OUT(2) => sig_HDU_PC_OUT_2_port, 
                           HDU_PC_OUT(1) => sig_HDU_PC_OUT_1_port, 
                           HDU_PC_OUT(0) => sig_HDU_PC_OUT_0_port, 
                           HDU_NPC_OUT(31) => sig_HDU_NPC_OUT_31_port, 
                           HDU_NPC_OUT(30) => sig_HDU_NPC_OUT_30_port, 
                           HDU_NPC_OUT(29) => sig_HDU_NPC_OUT_29_port, 
                           HDU_NPC_OUT(28) => sig_HDU_NPC_OUT_28_port, 
                           HDU_NPC_OUT(27) => sig_HDU_NPC_OUT_27_port, 
                           HDU_NPC_OUT(26) => sig_HDU_NPC_OUT_26_port, 
                           HDU_NPC_OUT(25) => sig_HDU_NPC_OUT_25_port, 
                           HDU_NPC_OUT(24) => sig_HDU_NPC_OUT_24_port, 
                           HDU_NPC_OUT(23) => sig_HDU_NPC_OUT_23_port, 
                           HDU_NPC_OUT(22) => sig_HDU_NPC_OUT_22_port, 
                           HDU_NPC_OUT(21) => sig_HDU_NPC_OUT_21_port, 
                           HDU_NPC_OUT(20) => sig_HDU_NPC_OUT_20_port, 
                           HDU_NPC_OUT(19) => sig_HDU_NPC_OUT_19_port, 
                           HDU_NPC_OUT(18) => sig_HDU_NPC_OUT_18_port, 
                           HDU_NPC_OUT(17) => sig_HDU_NPC_OUT_17_port, 
                           HDU_NPC_OUT(16) => sig_HDU_NPC_OUT_16_port, 
                           HDU_NPC_OUT(15) => sig_HDU_NPC_OUT_15_port, 
                           HDU_NPC_OUT(14) => sig_HDU_NPC_OUT_14_port, 
                           HDU_NPC_OUT(13) => sig_HDU_NPC_OUT_13_port, 
                           HDU_NPC_OUT(12) => sig_HDU_NPC_OUT_12_port, 
                           HDU_NPC_OUT(11) => sig_HDU_NPC_OUT_11_port, 
                           HDU_NPC_OUT(10) => sig_HDU_NPC_OUT_10_port, 
                           HDU_NPC_OUT(9) => sig_HDU_NPC_OUT_9_port, 
                           HDU_NPC_OUT(8) => sig_HDU_NPC_OUT_8_port, 
                           HDU_NPC_OUT(7) => sig_HDU_NPC_OUT_7_port, 
                           HDU_NPC_OUT(6) => sig_HDU_NPC_OUT_6_port, 
                           HDU_NPC_OUT(5) => sig_HDU_NPC_OUT_5_port, 
                           HDU_NPC_OUT(4) => sig_HDU_NPC_OUT_4_port, 
                           HDU_NPC_OUT(3) => sig_HDU_NPC_OUT_3_port, 
                           HDU_NPC_OUT(2) => sig_HDU_NPC_OUT_2_port, 
                           HDU_NPC_OUT(1) => sig_HDU_NPC_OUT_1_port, 
                           HDU_NPC_OUT(0) => sig_HDU_NPC_OUT_0_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( Clk, Rst : in std_logic);

end DLX;

architecture SYN_dlx_rtl of DLX is

   component DRAM
      port( En, Rst : in std_logic;  ADDR_IN, DATA_IN : in std_logic_vector (31
            downto 0);  DRAM_W, DRAM_R : in std_logic;  DATA_OUT : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component IRAM
      port( Rst : in std_logic;  Addr : in std_logic_vector (31 downto 0);  
            Iout : out std_logic_vector (31 downto 0));
   end component;
   
   component hardwired_cu_NBIT32
      port( REG_LATCH_EN, RD1, RD2, MUX_A_SEL : out std_logic;  MUX_B_SEL : out
            std_logic_vector (1 downto 0);  ALU_OPC : out std_logic_vector (0 
            to 3);  ALU_OUTREG_EN, DRAM_R_IN : out std_logic;  JUMP_TYPE : out 
            std_logic_vector (1 downto 0);  MEM_EN_IN, DRAM_W_IN, RF_WE, 
            DRAM_EN_IN, WB_MUX_SEL : out std_logic;  INS_IN : in 
            std_logic_vector (31 downto 0);  Bubble, Clk, Rst : in std_logic);
   end component;
   
   component Datapath
      port( CLK, RST : in std_logic;  INS_IN, DATA_IN : in std_logic_vector (31
            downto 0);  REG_LATCH_EN, RD1, RD2, MUX_A_SEL : in std_logic;  
            MUX_B_SEL : in std_logic_vector (1 downto 0);  ALU_OPC : in 
            std_logic_vector (0 to 3);  ALU_OUTREG_EN : in std_logic;  
            JUMP_TYPE : in std_logic_vector (1 downto 0);  DRAM_R_IN, MEM_EN_IN
            , DRAM_W_IN, RF_WE, DRAM_EN_IN, WB_MUX_SEL : in std_logic;  INS_OUT
            , IRAM_ADDR_OUT, DRAM_ADDR_OUT, DATA_OUT : out std_logic_vector (31
            downto 0);  DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble_out : out 
            std_logic);
   end component;
   
   signal INS_IN_31_port, INS_IN_30_port, INS_IN_29_port, INS_IN_28_port, 
      INS_IN_27_port, INS_IN_26_port, INS_IN_25_port, INS_IN_24_port, 
      INS_IN_23_port, INS_IN_22_port, INS_IN_21_port, INS_IN_20_port, 
      INS_IN_19_port, INS_IN_18_port, INS_IN_17_port, INS_IN_16_port, 
      INS_IN_15_port, INS_IN_14_port, INS_IN_13_port, INS_IN_12_port, 
      INS_IN_11_port, INS_IN_10_port, INS_IN_9_port, INS_IN_8_port, 
      INS_IN_7_port, INS_IN_6_port, INS_IN_5_port, INS_IN_4_port, INS_IN_3_port
      , INS_IN_2_port, INS_IN_1_port, INS_IN_0_port, DATA_IN_31_port, 
      DATA_IN_30_port, DATA_IN_29_port, DATA_IN_28_port, DATA_IN_27_port, 
      DATA_IN_26_port, DATA_IN_25_port, DATA_IN_24_port, DATA_IN_23_port, 
      DATA_IN_22_port, DATA_IN_21_port, DATA_IN_20_port, DATA_IN_19_port, 
      DATA_IN_18_port, DATA_IN_17_port, DATA_IN_16_port, DATA_IN_15_port, 
      DATA_IN_14_port, DATA_IN_13_port, DATA_IN_12_port, DATA_IN_11_port, 
      DATA_IN_10_port, DATA_IN_9_port, DATA_IN_8_port, DATA_IN_7_port, 
      DATA_IN_6_port, DATA_IN_5_port, DATA_IN_4_port, DATA_IN_3_port, 
      DATA_IN_2_port, DATA_IN_1_port, DATA_IN_0_port, REG_LATCH_EN, RD1, RD2, 
      MUX_A_SEL, MUX_B_SEL_1_port, MUX_B_SEL_0_port, ALU_OPC_3_port, 
      ALU_OPC_2_port, ALU_OPC_1_port, ALU_OPC_0_port, ALU_OUTREG_EN, 
      JUMP_TYPE_1_port, JUMP_TYPE_0_port, DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, 
      RF_WE, DRAM_EN_IN, WB_MUX_SEL, IRAM_ADDR_OUT_31_port, 
      IRAM_ADDR_OUT_30_port, IRAM_ADDR_OUT_29_port, IRAM_ADDR_OUT_28_port, 
      IRAM_ADDR_OUT_27_port, IRAM_ADDR_OUT_26_port, IRAM_ADDR_OUT_25_port, 
      IRAM_ADDR_OUT_24_port, IRAM_ADDR_OUT_23_port, IRAM_ADDR_OUT_22_port, 
      IRAM_ADDR_OUT_21_port, IRAM_ADDR_OUT_20_port, IRAM_ADDR_OUT_19_port, 
      IRAM_ADDR_OUT_18_port, IRAM_ADDR_OUT_17_port, IRAM_ADDR_OUT_16_port, 
      IRAM_ADDR_OUT_15_port, IRAM_ADDR_OUT_14_port, IRAM_ADDR_OUT_13_port, 
      IRAM_ADDR_OUT_12_port, IRAM_ADDR_OUT_11_port, IRAM_ADDR_OUT_10_port, 
      IRAM_ADDR_OUT_9_port, IRAM_ADDR_OUT_8_port, IRAM_ADDR_OUT_7_port, 
      IRAM_ADDR_OUT_6_port, IRAM_ADDR_OUT_5_port, IRAM_ADDR_OUT_4_port, 
      IRAM_ADDR_OUT_3_port, IRAM_ADDR_OUT_2_port, IRAM_ADDR_OUT_1_port, 
      IRAM_ADDR_OUT_0_port, DRAM_ADDR_OUT_31_port, DRAM_ADDR_OUT_30_port, 
      DRAM_ADDR_OUT_29_port, DRAM_ADDR_OUT_28_port, DRAM_ADDR_OUT_27_port, 
      DRAM_ADDR_OUT_26_port, DRAM_ADDR_OUT_25_port, DRAM_ADDR_OUT_24_port, 
      DRAM_ADDR_OUT_23_port, DRAM_ADDR_OUT_22_port, DRAM_ADDR_OUT_21_port, 
      DRAM_ADDR_OUT_20_port, DRAM_ADDR_OUT_19_port, DRAM_ADDR_OUT_18_port, 
      DRAM_ADDR_OUT_17_port, DRAM_ADDR_OUT_16_port, DRAM_ADDR_OUT_15_port, 
      DRAM_ADDR_OUT_14_port, DRAM_ADDR_OUT_13_port, DRAM_ADDR_OUT_12_port, 
      DRAM_ADDR_OUT_11_port, DRAM_ADDR_OUT_10_port, DRAM_ADDR_OUT_9_port, 
      DRAM_ADDR_OUT_8_port, DRAM_ADDR_OUT_7_port, DRAM_ADDR_OUT_6_port, 
      DRAM_ADDR_OUT_5_port, DRAM_ADDR_OUT_4_port, DRAM_ADDR_OUT_3_port, 
      DRAM_ADDR_OUT_2_port, DRAM_ADDR_OUT_1_port, DRAM_ADDR_OUT_0_port, 
      DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, DATA_OUT_28_port, 
      DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, DATA_OUT_24_port, 
      DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, DATA_OUT_20_port, 
      DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, DATA_OUT_16_port, 
      DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, DATA_OUT_12_port, 
      DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, DATA_OUT_8_port, 
      DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, DATA_OUT_4_port, 
      DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, DATA_OUT_0_port, 
      DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble, n_1837, n_1838, n_1839, 
      n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, 
      n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, 
      n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, 
      n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, 
      n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883 : 
      std_logic;

begin
   
   DP : Datapath port map( CLK => Clk, RST => Rst, INS_IN(31) => INS_IN_31_port
                           , INS_IN(30) => INS_IN_30_port, INS_IN(29) => 
                           INS_IN_29_port, INS_IN(28) => INS_IN_28_port, 
                           INS_IN(27) => INS_IN_27_port, INS_IN(26) => 
                           INS_IN_26_port, INS_IN(25) => INS_IN_25_port, 
                           INS_IN(24) => INS_IN_24_port, INS_IN(23) => 
                           INS_IN_23_port, INS_IN(22) => INS_IN_22_port, 
                           INS_IN(21) => INS_IN_21_port, INS_IN(20) => 
                           INS_IN_20_port, INS_IN(19) => INS_IN_19_port, 
                           INS_IN(18) => INS_IN_18_port, INS_IN(17) => 
                           INS_IN_17_port, INS_IN(16) => INS_IN_16_port, 
                           INS_IN(15) => INS_IN_15_port, INS_IN(14) => 
                           INS_IN_14_port, INS_IN(13) => INS_IN_13_port, 
                           INS_IN(12) => INS_IN_12_port, INS_IN(11) => 
                           INS_IN_11_port, INS_IN(10) => INS_IN_10_port, 
                           INS_IN(9) => INS_IN_9_port, INS_IN(8) => 
                           INS_IN_8_port, INS_IN(7) => INS_IN_7_port, INS_IN(6)
                           => INS_IN_6_port, INS_IN(5) => INS_IN_5_port, 
                           INS_IN(4) => INS_IN_4_port, INS_IN(3) => 
                           INS_IN_3_port, INS_IN(2) => INS_IN_2_port, INS_IN(1)
                           => INS_IN_1_port, INS_IN(0) => INS_IN_0_port, 
                           DATA_IN(31) => DATA_IN_31_port, DATA_IN(30) => 
                           DATA_IN_30_port, DATA_IN(29) => DATA_IN_29_port, 
                           DATA_IN(28) => DATA_IN_28_port, DATA_IN(27) => 
                           DATA_IN_27_port, DATA_IN(26) => DATA_IN_26_port, 
                           DATA_IN(25) => DATA_IN_25_port, DATA_IN(24) => 
                           DATA_IN_24_port, DATA_IN(23) => DATA_IN_23_port, 
                           DATA_IN(22) => DATA_IN_22_port, DATA_IN(21) => 
                           DATA_IN_21_port, DATA_IN(20) => DATA_IN_20_port, 
                           DATA_IN(19) => DATA_IN_19_port, DATA_IN(18) => 
                           DATA_IN_18_port, DATA_IN(17) => DATA_IN_17_port, 
                           DATA_IN(16) => DATA_IN_16_port, DATA_IN(15) => 
                           DATA_IN_15_port, DATA_IN(14) => DATA_IN_14_port, 
                           DATA_IN(13) => DATA_IN_13_port, DATA_IN(12) => 
                           DATA_IN_12_port, DATA_IN(11) => DATA_IN_11_port, 
                           DATA_IN(10) => DATA_IN_10_port, DATA_IN(9) => 
                           DATA_IN_9_port, DATA_IN(8) => DATA_IN_8_port, 
                           DATA_IN(7) => DATA_IN_7_port, DATA_IN(6) => 
                           DATA_IN_6_port, DATA_IN(5) => DATA_IN_5_port, 
                           DATA_IN(4) => DATA_IN_4_port, DATA_IN(3) => 
                           DATA_IN_3_port, DATA_IN(2) => DATA_IN_2_port, 
                           DATA_IN(1) => DATA_IN_1_port, DATA_IN(0) => 
                           DATA_IN_0_port, REG_LATCH_EN => REG_LATCH_EN, RD1 =>
                           RD1, RD2 => RD2, MUX_A_SEL => MUX_A_SEL, 
                           MUX_B_SEL(1) => MUX_B_SEL_1_port, MUX_B_SEL(0) => 
                           MUX_B_SEL_0_port, ALU_OPC(0) => ALU_OPC_3_port, 
                           ALU_OPC(1) => ALU_OPC_2_port, ALU_OPC(2) => 
                           ALU_OPC_1_port, ALU_OPC(3) => ALU_OPC_0_port, 
                           ALU_OUTREG_EN => ALU_OUTREG_EN, JUMP_TYPE(1) => 
                           JUMP_TYPE_1_port, JUMP_TYPE(0) => JUMP_TYPE_0_port, 
                           DRAM_R_IN => DRAM_R_IN, MEM_EN_IN => MEM_EN_IN, 
                           DRAM_W_IN => DRAM_W_IN, RF_WE => RF_WE, DRAM_EN_IN 
                           => DRAM_EN_IN, WB_MUX_SEL => WB_MUX_SEL, INS_OUT(31)
                           => n_1837, INS_OUT(30) => n_1838, INS_OUT(29) => 
                           n_1839, INS_OUT(28) => n_1840, INS_OUT(27) => n_1841
                           , INS_OUT(26) => n_1842, INS_OUT(25) => n_1843, 
                           INS_OUT(24) => n_1844, INS_OUT(23) => n_1845, 
                           INS_OUT(22) => n_1846, INS_OUT(21) => n_1847, 
                           INS_OUT(20) => n_1848, INS_OUT(19) => n_1849, 
                           INS_OUT(18) => n_1850, INS_OUT(17) => n_1851, 
                           INS_OUT(16) => n_1852, INS_OUT(15) => n_1853, 
                           INS_OUT(14) => n_1854, INS_OUT(13) => n_1855, 
                           INS_OUT(12) => n_1856, INS_OUT(11) => n_1857, 
                           INS_OUT(10) => n_1858, INS_OUT(9) => n_1859, 
                           INS_OUT(8) => n_1860, INS_OUT(7) => n_1861, 
                           INS_OUT(6) => n_1862, INS_OUT(5) => n_1863, 
                           INS_OUT(4) => n_1864, INS_OUT(3) => n_1865, 
                           INS_OUT(2) => n_1866, INS_OUT(1) => n_1867, 
                           INS_OUT(0) => n_1868, IRAM_ADDR_OUT(31) => 
                           IRAM_ADDR_OUT_31_port, IRAM_ADDR_OUT(30) => 
                           IRAM_ADDR_OUT_30_port, IRAM_ADDR_OUT(29) => 
                           IRAM_ADDR_OUT_29_port, IRAM_ADDR_OUT(28) => 
                           IRAM_ADDR_OUT_28_port, IRAM_ADDR_OUT(27) => 
                           IRAM_ADDR_OUT_27_port, IRAM_ADDR_OUT(26) => 
                           IRAM_ADDR_OUT_26_port, IRAM_ADDR_OUT(25) => 
                           IRAM_ADDR_OUT_25_port, IRAM_ADDR_OUT(24) => 
                           IRAM_ADDR_OUT_24_port, IRAM_ADDR_OUT(23) => 
                           IRAM_ADDR_OUT_23_port, IRAM_ADDR_OUT(22) => 
                           IRAM_ADDR_OUT_22_port, IRAM_ADDR_OUT(21) => 
                           IRAM_ADDR_OUT_21_port, IRAM_ADDR_OUT(20) => 
                           IRAM_ADDR_OUT_20_port, IRAM_ADDR_OUT(19) => 
                           IRAM_ADDR_OUT_19_port, IRAM_ADDR_OUT(18) => 
                           IRAM_ADDR_OUT_18_port, IRAM_ADDR_OUT(17) => 
                           IRAM_ADDR_OUT_17_port, IRAM_ADDR_OUT(16) => 
                           IRAM_ADDR_OUT_16_port, IRAM_ADDR_OUT(15) => 
                           IRAM_ADDR_OUT_15_port, IRAM_ADDR_OUT(14) => 
                           IRAM_ADDR_OUT_14_port, IRAM_ADDR_OUT(13) => 
                           IRAM_ADDR_OUT_13_port, IRAM_ADDR_OUT(12) => 
                           IRAM_ADDR_OUT_12_port, IRAM_ADDR_OUT(11) => 
                           IRAM_ADDR_OUT_11_port, IRAM_ADDR_OUT(10) => 
                           IRAM_ADDR_OUT_10_port, IRAM_ADDR_OUT(9) => 
                           IRAM_ADDR_OUT_9_port, IRAM_ADDR_OUT(8) => 
                           IRAM_ADDR_OUT_8_port, IRAM_ADDR_OUT(7) => 
                           IRAM_ADDR_OUT_7_port, IRAM_ADDR_OUT(6) => 
                           IRAM_ADDR_OUT_6_port, IRAM_ADDR_OUT(5) => 
                           IRAM_ADDR_OUT_5_port, IRAM_ADDR_OUT(4) => 
                           IRAM_ADDR_OUT_4_port, IRAM_ADDR_OUT(3) => 
                           IRAM_ADDR_OUT_3_port, IRAM_ADDR_OUT(2) => 
                           IRAM_ADDR_OUT_2_port, IRAM_ADDR_OUT(1) => 
                           IRAM_ADDR_OUT_1_port, IRAM_ADDR_OUT(0) => 
                           IRAM_ADDR_OUT_0_port, DRAM_ADDR_OUT(31) => 
                           DRAM_ADDR_OUT_31_port, DRAM_ADDR_OUT(30) => 
                           DRAM_ADDR_OUT_30_port, DRAM_ADDR_OUT(29) => 
                           DRAM_ADDR_OUT_29_port, DRAM_ADDR_OUT(28) => 
                           DRAM_ADDR_OUT_28_port, DRAM_ADDR_OUT(27) => 
                           DRAM_ADDR_OUT_27_port, DRAM_ADDR_OUT(26) => 
                           DRAM_ADDR_OUT_26_port, DRAM_ADDR_OUT(25) => 
                           DRAM_ADDR_OUT_25_port, DRAM_ADDR_OUT(24) => 
                           DRAM_ADDR_OUT_24_port, DRAM_ADDR_OUT(23) => 
                           DRAM_ADDR_OUT_23_port, DRAM_ADDR_OUT(22) => 
                           DRAM_ADDR_OUT_22_port, DRAM_ADDR_OUT(21) => 
                           DRAM_ADDR_OUT_21_port, DRAM_ADDR_OUT(20) => 
                           DRAM_ADDR_OUT_20_port, DRAM_ADDR_OUT(19) => 
                           DRAM_ADDR_OUT_19_port, DRAM_ADDR_OUT(18) => 
                           DRAM_ADDR_OUT_18_port, DRAM_ADDR_OUT(17) => 
                           DRAM_ADDR_OUT_17_port, DRAM_ADDR_OUT(16) => 
                           DRAM_ADDR_OUT_16_port, DRAM_ADDR_OUT(15) => 
                           DRAM_ADDR_OUT_15_port, DRAM_ADDR_OUT(14) => 
                           DRAM_ADDR_OUT_14_port, DRAM_ADDR_OUT(13) => 
                           DRAM_ADDR_OUT_13_port, DRAM_ADDR_OUT(12) => 
                           DRAM_ADDR_OUT_12_port, DRAM_ADDR_OUT(11) => 
                           DRAM_ADDR_OUT_11_port, DRAM_ADDR_OUT(10) => 
                           DRAM_ADDR_OUT_10_port, DRAM_ADDR_OUT(9) => 
                           DRAM_ADDR_OUT_9_port, DRAM_ADDR_OUT(8) => 
                           DRAM_ADDR_OUT_8_port, DRAM_ADDR_OUT(7) => 
                           DRAM_ADDR_OUT_7_port, DRAM_ADDR_OUT(6) => 
                           DRAM_ADDR_OUT_6_port, DRAM_ADDR_OUT(5) => 
                           DRAM_ADDR_OUT_5_port, DRAM_ADDR_OUT(4) => 
                           DRAM_ADDR_OUT_4_port, DRAM_ADDR_OUT(3) => 
                           DRAM_ADDR_OUT_3_port, DRAM_ADDR_OUT(2) => 
                           DRAM_ADDR_OUT_2_port, DRAM_ADDR_OUT(1) => 
                           DRAM_ADDR_OUT_1_port, DRAM_ADDR_OUT(0) => 
                           DRAM_ADDR_OUT_0_port, DATA_OUT(31) => 
                           DATA_OUT_31_port, DATA_OUT(30) => DATA_OUT_30_port, 
                           DATA_OUT(29) => DATA_OUT_29_port, DATA_OUT(28) => 
                           DATA_OUT_28_port, DATA_OUT(27) => DATA_OUT_27_port, 
                           DATA_OUT(26) => DATA_OUT_26_port, DATA_OUT(25) => 
                           DATA_OUT_25_port, DATA_OUT(24) => DATA_OUT_24_port, 
                           DATA_OUT(23) => DATA_OUT_23_port, DATA_OUT(22) => 
                           DATA_OUT_22_port, DATA_OUT(21) => DATA_OUT_21_port, 
                           DATA_OUT(20) => DATA_OUT_20_port, DATA_OUT(19) => 
                           DATA_OUT_19_port, DATA_OUT(18) => DATA_OUT_18_port, 
                           DATA_OUT(17) => DATA_OUT_17_port, DATA_OUT(16) => 
                           DATA_OUT_16_port, DATA_OUT(15) => DATA_OUT_15_port, 
                           DATA_OUT(14) => DATA_OUT_14_port, DATA_OUT(13) => 
                           DATA_OUT_13_port, DATA_OUT(12) => DATA_OUT_12_port, 
                           DATA_OUT(11) => DATA_OUT_11_port, DATA_OUT(10) => 
                           DATA_OUT_10_port, DATA_OUT(9) => DATA_OUT_9_port, 
                           DATA_OUT(8) => DATA_OUT_8_port, DATA_OUT(7) => 
                           DATA_OUT_7_port, DATA_OUT(6) => DATA_OUT_6_port, 
                           DATA_OUT(5) => DATA_OUT_5_port, DATA_OUT(4) => 
                           DATA_OUT_4_port, DATA_OUT(3) => DATA_OUT_3_port, 
                           DATA_OUT(2) => DATA_OUT_2_port, DATA_OUT(1) => 
                           DATA_OUT_1_port, DATA_OUT(0) => DATA_OUT_0_port, 
                           DRAM_EN_OUT => DRAM_EN_OUT, DRAM_R_OUT => DRAM_R_OUT
                           , DRAM_W_OUT => DRAM_W_OUT, Bubble_out => Bubble);
   CU : hardwired_cu_NBIT32 port map( REG_LATCH_EN => n_1869, RD1 => n_1870, 
                           RD2 => n_1871, MUX_A_SEL => n_1872, MUX_B_SEL(1) => 
                           n_1873, MUX_B_SEL(0) => n_1874, ALU_OPC(0) => 
                           ALU_OPC_3_port, ALU_OPC(1) => ALU_OPC_2_port, 
                           ALU_OPC(2) => ALU_OPC_1_port, ALU_OPC(3) => 
                           ALU_OPC_0_port, ALU_OUTREG_EN => n_1875, DRAM_R_IN 
                           => n_1876, JUMP_TYPE(1) => n_1877, JUMP_TYPE(0) => 
                           n_1878, MEM_EN_IN => n_1879, DRAM_W_IN => n_1880, 
                           RF_WE => n_1881, DRAM_EN_IN => n_1882, WB_MUX_SEL =>
                           n_1883, INS_IN(31) => INS_IN_31_port, INS_IN(30) => 
                           INS_IN_30_port, INS_IN(29) => INS_IN_29_port, 
                           INS_IN(28) => INS_IN_28_port, INS_IN(27) => 
                           INS_IN_27_port, INS_IN(26) => INS_IN_26_port, 
                           INS_IN(25) => INS_IN_25_port, INS_IN(24) => 
                           INS_IN_24_port, INS_IN(23) => INS_IN_23_port, 
                           INS_IN(22) => INS_IN_22_port, INS_IN(21) => 
                           INS_IN_21_port, INS_IN(20) => INS_IN_20_port, 
                           INS_IN(19) => INS_IN_19_port, INS_IN(18) => 
                           INS_IN_18_port, INS_IN(17) => INS_IN_17_port, 
                           INS_IN(16) => INS_IN_16_port, INS_IN(15) => 
                           INS_IN_15_port, INS_IN(14) => INS_IN_14_port, 
                           INS_IN(13) => INS_IN_13_port, INS_IN(12) => 
                           INS_IN_12_port, INS_IN(11) => INS_IN_11_port, 
                           INS_IN(10) => INS_IN_10_port, INS_IN(9) => 
                           INS_IN_9_port, INS_IN(8) => INS_IN_8_port, INS_IN(7)
                           => INS_IN_7_port, INS_IN(6) => INS_IN_6_port, 
                           INS_IN(5) => INS_IN_5_port, INS_IN(4) => 
                           INS_IN_4_port, INS_IN(3) => INS_IN_3_port, INS_IN(2)
                           => INS_IN_2_port, INS_IN(1) => INS_IN_1_port, 
                           INS_IN(0) => INS_IN_0_port, Bubble => Bubble, Clk =>
                           Clk, Rst => Rst);
   IRAM_I : IRAM port map( Rst => Rst, Addr(31) => IRAM_ADDR_OUT_31_port, 
                           Addr(30) => IRAM_ADDR_OUT_30_port, Addr(29) => 
                           IRAM_ADDR_OUT_29_port, Addr(28) => 
                           IRAM_ADDR_OUT_28_port, Addr(27) => 
                           IRAM_ADDR_OUT_27_port, Addr(26) => 
                           IRAM_ADDR_OUT_26_port, Addr(25) => 
                           IRAM_ADDR_OUT_25_port, Addr(24) => 
                           IRAM_ADDR_OUT_24_port, Addr(23) => 
                           IRAM_ADDR_OUT_23_port, Addr(22) => 
                           IRAM_ADDR_OUT_22_port, Addr(21) => 
                           IRAM_ADDR_OUT_21_port, Addr(20) => 
                           IRAM_ADDR_OUT_20_port, Addr(19) => 
                           IRAM_ADDR_OUT_19_port, Addr(18) => 
                           IRAM_ADDR_OUT_18_port, Addr(17) => 
                           IRAM_ADDR_OUT_17_port, Addr(16) => 
                           IRAM_ADDR_OUT_16_port, Addr(15) => 
                           IRAM_ADDR_OUT_15_port, Addr(14) => 
                           IRAM_ADDR_OUT_14_port, Addr(13) => 
                           IRAM_ADDR_OUT_13_port, Addr(12) => 
                           IRAM_ADDR_OUT_12_port, Addr(11) => 
                           IRAM_ADDR_OUT_11_port, Addr(10) => 
                           IRAM_ADDR_OUT_10_port, Addr(9) => 
                           IRAM_ADDR_OUT_9_port, Addr(8) => 
                           IRAM_ADDR_OUT_8_port, Addr(7) => 
                           IRAM_ADDR_OUT_7_port, Addr(6) => 
                           IRAM_ADDR_OUT_6_port, Addr(5) => 
                           IRAM_ADDR_OUT_5_port, Addr(4) => 
                           IRAM_ADDR_OUT_4_port, Addr(3) => 
                           IRAM_ADDR_OUT_3_port, Addr(2) => 
                           IRAM_ADDR_OUT_2_port, Addr(1) => 
                           IRAM_ADDR_OUT_1_port, Addr(0) => 
                           IRAM_ADDR_OUT_0_port, Iout(31) => INS_IN_31_port, 
                           Iout(30) => INS_IN_30_port, Iout(29) => 
                           INS_IN_29_port, Iout(28) => INS_IN_28_port, Iout(27)
                           => INS_IN_27_port, Iout(26) => INS_IN_26_port, 
                           Iout(25) => INS_IN_25_port, Iout(24) => 
                           INS_IN_24_port, Iout(23) => INS_IN_23_port, Iout(22)
                           => INS_IN_22_port, Iout(21) => INS_IN_21_port, 
                           Iout(20) => INS_IN_20_port, Iout(19) => 
                           INS_IN_19_port, Iout(18) => INS_IN_18_port, Iout(17)
                           => INS_IN_17_port, Iout(16) => INS_IN_16_port, 
                           Iout(15) => INS_IN_15_port, Iout(14) => 
                           INS_IN_14_port, Iout(13) => INS_IN_13_port, Iout(12)
                           => INS_IN_12_port, Iout(11) => INS_IN_11_port, 
                           Iout(10) => INS_IN_10_port, Iout(9) => INS_IN_9_port
                           , Iout(8) => INS_IN_8_port, Iout(7) => INS_IN_7_port
                           , Iout(6) => INS_IN_6_port, Iout(5) => INS_IN_5_port
                           , Iout(4) => INS_IN_4_port, Iout(3) => INS_IN_3_port
                           , Iout(2) => INS_IN_2_port, Iout(1) => INS_IN_1_port
                           , Iout(0) => INS_IN_0_port);
   DRAM_I : DRAM port map( En => DRAM_EN_OUT, Rst => Rst, ADDR_IN(31) => 
                           DRAM_ADDR_OUT_31_port, ADDR_IN(30) => 
                           DRAM_ADDR_OUT_30_port, ADDR_IN(29) => 
                           DRAM_ADDR_OUT_29_port, ADDR_IN(28) => 
                           DRAM_ADDR_OUT_28_port, ADDR_IN(27) => 
                           DRAM_ADDR_OUT_27_port, ADDR_IN(26) => 
                           DRAM_ADDR_OUT_26_port, ADDR_IN(25) => 
                           DRAM_ADDR_OUT_25_port, ADDR_IN(24) => 
                           DRAM_ADDR_OUT_24_port, ADDR_IN(23) => 
                           DRAM_ADDR_OUT_23_port, ADDR_IN(22) => 
                           DRAM_ADDR_OUT_22_port, ADDR_IN(21) => 
                           DRAM_ADDR_OUT_21_port, ADDR_IN(20) => 
                           DRAM_ADDR_OUT_20_port, ADDR_IN(19) => 
                           DRAM_ADDR_OUT_19_port, ADDR_IN(18) => 
                           DRAM_ADDR_OUT_18_port, ADDR_IN(17) => 
                           DRAM_ADDR_OUT_17_port, ADDR_IN(16) => 
                           DRAM_ADDR_OUT_16_port, ADDR_IN(15) => 
                           DRAM_ADDR_OUT_15_port, ADDR_IN(14) => 
                           DRAM_ADDR_OUT_14_port, ADDR_IN(13) => 
                           DRAM_ADDR_OUT_13_port, ADDR_IN(12) => 
                           DRAM_ADDR_OUT_12_port, ADDR_IN(11) => 
                           DRAM_ADDR_OUT_11_port, ADDR_IN(10) => 
                           DRAM_ADDR_OUT_10_port, ADDR_IN(9) => 
                           DRAM_ADDR_OUT_9_port, ADDR_IN(8) => 
                           DRAM_ADDR_OUT_8_port, ADDR_IN(7) => 
                           DRAM_ADDR_OUT_7_port, ADDR_IN(6) => 
                           DRAM_ADDR_OUT_6_port, ADDR_IN(5) => 
                           DRAM_ADDR_OUT_5_port, ADDR_IN(4) => 
                           DRAM_ADDR_OUT_4_port, ADDR_IN(3) => 
                           DRAM_ADDR_OUT_3_port, ADDR_IN(2) => 
                           DRAM_ADDR_OUT_2_port, ADDR_IN(1) => 
                           DRAM_ADDR_OUT_1_port, ADDR_IN(0) => 
                           DRAM_ADDR_OUT_0_port, DATA_IN(31) => 
                           DATA_OUT_31_port, DATA_IN(30) => DATA_OUT_30_port, 
                           DATA_IN(29) => DATA_OUT_29_port, DATA_IN(28) => 
                           DATA_OUT_28_port, DATA_IN(27) => DATA_OUT_27_port, 
                           DATA_IN(26) => DATA_OUT_26_port, DATA_IN(25) => 
                           DATA_OUT_25_port, DATA_IN(24) => DATA_OUT_24_port, 
                           DATA_IN(23) => DATA_OUT_23_port, DATA_IN(22) => 
                           DATA_OUT_22_port, DATA_IN(21) => DATA_OUT_21_port, 
                           DATA_IN(20) => DATA_OUT_20_port, DATA_IN(19) => 
                           DATA_OUT_19_port, DATA_IN(18) => DATA_OUT_18_port, 
                           DATA_IN(17) => DATA_OUT_17_port, DATA_IN(16) => 
                           DATA_OUT_16_port, DATA_IN(15) => DATA_OUT_15_port, 
                           DATA_IN(14) => DATA_OUT_14_port, DATA_IN(13) => 
                           DATA_OUT_13_port, DATA_IN(12) => DATA_OUT_12_port, 
                           DATA_IN(11) => DATA_OUT_11_port, DATA_IN(10) => 
                           DATA_OUT_10_port, DATA_IN(9) => DATA_OUT_9_port, 
                           DATA_IN(8) => DATA_OUT_8_port, DATA_IN(7) => 
                           DATA_OUT_7_port, DATA_IN(6) => DATA_OUT_6_port, 
                           DATA_IN(5) => DATA_OUT_5_port, DATA_IN(4) => 
                           DATA_OUT_4_port, DATA_IN(3) => DATA_OUT_3_port, 
                           DATA_IN(2) => DATA_OUT_2_port, DATA_IN(1) => 
                           DATA_OUT_1_port, DATA_IN(0) => DATA_OUT_0_port, 
                           DRAM_W => DRAM_W_OUT, DRAM_R => DRAM_R_OUT, 
                           DATA_OUT(31) => DATA_IN_31_port, DATA_OUT(30) => 
                           DATA_IN_30_port, DATA_OUT(29) => DATA_IN_29_port, 
                           DATA_OUT(28) => DATA_IN_28_port, DATA_OUT(27) => 
                           DATA_IN_27_port, DATA_OUT(26) => DATA_IN_26_port, 
                           DATA_OUT(25) => DATA_IN_25_port, DATA_OUT(24) => 
                           DATA_IN_24_port, DATA_OUT(23) => DATA_IN_23_port, 
                           DATA_OUT(22) => DATA_IN_22_port, DATA_OUT(21) => 
                           DATA_IN_21_port, DATA_OUT(20) => DATA_IN_20_port, 
                           DATA_OUT(19) => DATA_IN_19_port, DATA_OUT(18) => 
                           DATA_IN_18_port, DATA_OUT(17) => DATA_IN_17_port, 
                           DATA_OUT(16) => DATA_IN_16_port, DATA_OUT(15) => 
                           DATA_IN_15_port, DATA_OUT(14) => DATA_IN_14_port, 
                           DATA_OUT(13) => DATA_IN_13_port, DATA_OUT(12) => 
                           DATA_IN_12_port, DATA_OUT(11) => DATA_IN_11_port, 
                           DATA_OUT(10) => DATA_IN_10_port, DATA_OUT(9) => 
                           DATA_IN_9_port, DATA_OUT(8) => DATA_IN_8_port, 
                           DATA_OUT(7) => DATA_IN_7_port, DATA_OUT(6) => 
                           DATA_IN_6_port, DATA_OUT(5) => DATA_IN_5_port, 
                           DATA_OUT(4) => DATA_IN_4_port, DATA_OUT(3) => 
                           DATA_IN_3_port, DATA_OUT(2) => DATA_IN_2_port, 
                           DATA_OUT(1) => DATA_IN_1_port, DATA_OUT(0) => 
                           DATA_IN_0_port);
   WB_MUX_SEL <= '0';
   DRAM_EN_IN <= '0';
   RF_WE <= '0';
   DRAM_W_IN <= '0';
   MEM_EN_IN <= '0';
   JUMP_TYPE_0_port <= '0';
   JUMP_TYPE_1_port <= '0';
   DRAM_R_IN <= '0';
   ALU_OUTREG_EN <= '0';
   MUX_B_SEL_0_port <= '0';
   MUX_B_SEL_1_port <= '0';
   MUX_A_SEL <= '0';
   RD2 <= '0';
   RD1 <= '0';
   REG_LATCH_EN <= '0';

end SYN_dlx_rtl;
