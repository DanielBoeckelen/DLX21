
module mux21_NBIT32_0 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n36, n37, n38, n39, n40, n43, n54, n65, n1, n2, n3;

  INV_X2 U1 ( .A(n2), .ZN(n1) );
  INV_X1 U2 ( .A(n54), .ZN(Z[1]) );
  AOI22_X1 U3 ( .A1(A[1]), .A2(n2), .B1(B[1]), .B2(S), .ZN(n54) );
  INV_X1 U4 ( .A(n43), .ZN(Z[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(n3), .B1(B[2]), .B2(S), .ZN(n43) );
  INV_X1 U6 ( .A(n40), .ZN(Z[3]) );
  AOI22_X1 U7 ( .A1(A[3]), .A2(n2), .B1(B[3]), .B2(S), .ZN(n40) );
  INV_X1 U8 ( .A(n36), .ZN(Z[7]) );
  AOI22_X1 U9 ( .A1(A[7]), .A2(n3), .B1(B[7]), .B2(S), .ZN(n36) );
  INV_X1 U10 ( .A(n37), .ZN(Z[6]) );
  AOI22_X1 U11 ( .A1(A[6]), .A2(n3), .B1(B[6]), .B2(S), .ZN(n37) );
  INV_X1 U12 ( .A(n38), .ZN(Z[5]) );
  AOI22_X1 U13 ( .A1(A[5]), .A2(n2), .B1(B[5]), .B2(S), .ZN(n38) );
  INV_X1 U14 ( .A(n39), .ZN(Z[4]) );
  AOI22_X1 U15 ( .A1(A[4]), .A2(n2), .B1(B[4]), .B2(S), .ZN(n39) );
  INV_X1 U16 ( .A(n65), .ZN(Z[0]) );
  AOI22_X1 U17 ( .A1(A[0]), .A2(n3), .B1(B[0]), .B2(S), .ZN(n65) );
  INV_X1 U18 ( .A(S), .ZN(n2) );
  INV_X1 U19 ( .A(S), .ZN(n3) );
  MUX2_X1 U20 ( .A(A[8]), .B(B[8]), .S(n1), .Z(Z[8]) );
  MUX2_X1 U21 ( .A(A[9]), .B(B[9]), .S(n1), .Z(Z[9]) );
  MUX2_X1 U22 ( .A(A[10]), .B(B[10]), .S(n1), .Z(Z[10]) );
  MUX2_X1 U23 ( .A(A[11]), .B(B[11]), .S(n1), .Z(Z[11]) );
  MUX2_X1 U24 ( .A(A[12]), .B(B[12]), .S(n1), .Z(Z[12]) );
  MUX2_X1 U25 ( .A(A[13]), .B(B[13]), .S(n1), .Z(Z[13]) );
  MUX2_X1 U26 ( .A(A[14]), .B(B[14]), .S(n1), .Z(Z[14]) );
  MUX2_X1 U27 ( .A(A[15]), .B(B[15]), .S(n1), .Z(Z[15]) );
  MUX2_X1 U28 ( .A(A[16]), .B(B[16]), .S(n1), .Z(Z[16]) );
  MUX2_X1 U29 ( .A(A[17]), .B(B[17]), .S(n1), .Z(Z[17]) );
  MUX2_X1 U30 ( .A(A[18]), .B(B[18]), .S(n1), .Z(Z[18]) );
  MUX2_X1 U31 ( .A(A[19]), .B(B[19]), .S(n1), .Z(Z[19]) );
  MUX2_X1 U32 ( .A(A[20]), .B(B[20]), .S(n1), .Z(Z[20]) );
  MUX2_X1 U33 ( .A(A[21]), .B(B[21]), .S(n1), .Z(Z[21]) );
  MUX2_X1 U34 ( .A(A[22]), .B(B[22]), .S(n1), .Z(Z[22]) );
  MUX2_X1 U35 ( .A(A[23]), .B(B[23]), .S(n1), .Z(Z[23]) );
  MUX2_X1 U36 ( .A(A[24]), .B(B[24]), .S(n1), .Z(Z[24]) );
  MUX2_X1 U37 ( .A(A[25]), .B(B[25]), .S(n1), .Z(Z[25]) );
  MUX2_X1 U38 ( .A(A[26]), .B(B[26]), .S(n1), .Z(Z[26]) );
  MUX2_X1 U39 ( .A(A[27]), .B(B[27]), .S(n1), .Z(Z[27]) );
  MUX2_X1 U40 ( .A(A[28]), .B(B[28]), .S(n1), .Z(Z[28]) );
  MUX2_X1 U41 ( .A(A[29]), .B(B[29]), .S(n1), .Z(Z[29]) );
  MUX2_X1 U42 ( .A(A[30]), .B(B[30]), .S(n1), .Z(Z[30]) );
  MUX2_X1 U43 ( .A(A[31]), .B(B[31]), .S(n1), .Z(Z[31]) );
endmodule


module mux21_NBIT32_6 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104;

  BUF_X2 U1 ( .A(n2), .Z(n7) );
  INV_X2 U2 ( .A(S), .ZN(n3) );
  CLKBUF_X1 U3 ( .A(S), .Z(n2) );
  CLKBUF_X1 U4 ( .A(S), .Z(n1) );
  CLKBUF_X1 U5 ( .A(n4), .Z(n8) );
  CLKBUF_X1 U6 ( .A(n1), .Z(n4) );
  BUF_X1 U7 ( .A(n1), .Z(n6) );
  BUF_X1 U8 ( .A(n1), .Z(n5) );
  INV_X1 U9 ( .A(n95), .ZN(Z[2]) );
  AOI22_X1 U10 ( .A1(A[2]), .A2(n3), .B1(B[2]), .B2(n5), .ZN(n95) );
  INV_X1 U11 ( .A(n84), .ZN(Z[1]) );
  AOI22_X1 U12 ( .A1(A[1]), .A2(n3), .B1(B[1]), .B2(n7), .ZN(n84) );
  INV_X1 U13 ( .A(n73), .ZN(Z[0]) );
  AOI22_X1 U14 ( .A1(A[0]), .A2(n3), .B1(B[0]), .B2(n8), .ZN(n73) );
  INV_X1 U15 ( .A(n98), .ZN(Z[3]) );
  AOI22_X1 U16 ( .A1(A[3]), .A2(n3), .B1(B[3]), .B2(n5), .ZN(n98) );
  INV_X1 U17 ( .A(n99), .ZN(Z[4]) );
  AOI22_X1 U18 ( .A1(A[4]), .A2(n3), .B1(B[4]), .B2(n5), .ZN(n99) );
  INV_X1 U19 ( .A(n100), .ZN(Z[5]) );
  AOI22_X1 U20 ( .A1(A[5]), .A2(n3), .B1(B[5]), .B2(n4), .ZN(n100) );
  INV_X1 U21 ( .A(n101), .ZN(Z[6]) );
  AOI22_X1 U22 ( .A1(A[6]), .A2(n3), .B1(B[6]), .B2(n4), .ZN(n101) );
  INV_X1 U23 ( .A(n102), .ZN(Z[7]) );
  AOI22_X1 U24 ( .A1(A[7]), .A2(n3), .B1(B[7]), .B2(n4), .ZN(n102) );
  INV_X1 U25 ( .A(n103), .ZN(Z[8]) );
  AOI22_X1 U26 ( .A1(A[8]), .A2(n3), .B1(B[8]), .B2(n4), .ZN(n103) );
  INV_X1 U27 ( .A(n74), .ZN(Z[10]) );
  AOI22_X1 U28 ( .A1(A[10]), .A2(n3), .B1(B[10]), .B2(n8), .ZN(n74) );
  INV_X1 U29 ( .A(n75), .ZN(Z[11]) );
  AOI22_X1 U30 ( .A1(A[11]), .A2(n3), .B1(B[11]), .B2(n8), .ZN(n75) );
  INV_X1 U31 ( .A(n76), .ZN(Z[12]) );
  AOI22_X1 U32 ( .A1(A[12]), .A2(n3), .B1(B[12]), .B2(n8), .ZN(n76) );
  INV_X1 U33 ( .A(n77), .ZN(Z[13]) );
  AOI22_X1 U34 ( .A1(A[13]), .A2(n3), .B1(B[13]), .B2(n1), .ZN(n77) );
  INV_X1 U35 ( .A(n78), .ZN(Z[14]) );
  AOI22_X1 U36 ( .A1(A[14]), .A2(n3), .B1(B[14]), .B2(n2), .ZN(n78) );
  INV_X1 U37 ( .A(n79), .ZN(Z[15]) );
  AOI22_X1 U38 ( .A1(A[15]), .A2(n3), .B1(B[15]), .B2(n2), .ZN(n79) );
  INV_X1 U39 ( .A(n80), .ZN(Z[16]) );
  AOI22_X1 U40 ( .A1(A[16]), .A2(n3), .B1(B[16]), .B2(n2), .ZN(n80) );
  INV_X1 U41 ( .A(n81), .ZN(Z[17]) );
  AOI22_X1 U42 ( .A1(A[17]), .A2(n3), .B1(B[17]), .B2(n1), .ZN(n81) );
  INV_X1 U43 ( .A(n82), .ZN(Z[18]) );
  AOI22_X1 U44 ( .A1(A[18]), .A2(n3), .B1(B[18]), .B2(n2), .ZN(n82) );
  INV_X1 U45 ( .A(n83), .ZN(Z[19]) );
  AOI22_X1 U46 ( .A1(A[19]), .A2(n3), .B1(B[19]), .B2(n1), .ZN(n83) );
  INV_X1 U47 ( .A(n85), .ZN(Z[20]) );
  AOI22_X1 U48 ( .A1(A[20]), .A2(n3), .B1(B[20]), .B2(n2), .ZN(n85) );
  INV_X1 U49 ( .A(n86), .ZN(Z[21]) );
  AOI22_X1 U50 ( .A1(A[21]), .A2(n3), .B1(B[21]), .B2(n6), .ZN(n86) );
  INV_X1 U51 ( .A(n87), .ZN(Z[22]) );
  AOI22_X1 U52 ( .A1(A[22]), .A2(n3), .B1(B[22]), .B2(n7), .ZN(n87) );
  INV_X1 U53 ( .A(n88), .ZN(Z[23]) );
  AOI22_X1 U54 ( .A1(A[23]), .A2(n3), .B1(B[23]), .B2(n7), .ZN(n88) );
  INV_X1 U55 ( .A(n89), .ZN(Z[24]) );
  AOI22_X1 U56 ( .A1(A[24]), .A2(n3), .B1(B[24]), .B2(n7), .ZN(n89) );
  INV_X1 U57 ( .A(n90), .ZN(Z[25]) );
  AOI22_X1 U58 ( .A1(A[25]), .A2(n3), .B1(B[25]), .B2(n7), .ZN(n90) );
  INV_X1 U59 ( .A(n91), .ZN(Z[26]) );
  AOI22_X1 U60 ( .A1(A[26]), .A2(n3), .B1(B[26]), .B2(n6), .ZN(n91) );
  INV_X1 U61 ( .A(n92), .ZN(Z[27]) );
  AOI22_X1 U62 ( .A1(A[27]), .A2(n3), .B1(B[27]), .B2(n6), .ZN(n92) );
  INV_X1 U63 ( .A(n93), .ZN(Z[28]) );
  AOI22_X1 U64 ( .A1(A[28]), .A2(n3), .B1(B[28]), .B2(n6), .ZN(n93) );
  INV_X1 U65 ( .A(n94), .ZN(Z[29]) );
  AOI22_X1 U66 ( .A1(A[29]), .A2(n3), .B1(B[29]), .B2(n6), .ZN(n94) );
  INV_X1 U67 ( .A(n96), .ZN(Z[30]) );
  AOI22_X1 U68 ( .A1(A[30]), .A2(n3), .B1(B[30]), .B2(n5), .ZN(n96) );
  INV_X1 U69 ( .A(n97), .ZN(Z[31]) );
  AOI22_X1 U70 ( .A1(A[31]), .A2(n3), .B1(B[31]), .B2(n5), .ZN(n97) );
  INV_X1 U71 ( .A(n104), .ZN(Z[9]) );
  AOI22_X1 U72 ( .A1(A[9]), .A2(n3), .B1(n8), .B2(B[9]), .ZN(n104) );
endmodule


module mux21_NBIT32_5 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99;

  BUF_X2 U1 ( .A(S), .Z(n3) );
  INV_X2 U2 ( .A(n3), .ZN(n1) );
  BUF_X1 U3 ( .A(S), .Z(n2) );
  INV_X1 U4 ( .A(n86), .ZN(Z[26]) );
  INV_X1 U5 ( .A(n91), .ZN(Z[30]) );
  INV_X1 U6 ( .A(n88), .ZN(Z[28]) );
  INV_X1 U7 ( .A(n92), .ZN(Z[31]) );
  INV_X1 U8 ( .A(n87), .ZN(Z[27]) );
  INV_X1 U9 ( .A(n89), .ZN(Z[29]) );
  INV_X1 U10 ( .A(n79), .ZN(Z[1]) );
  AOI22_X1 U11 ( .A1(A[1]), .A2(n1), .B1(B[1]), .B2(n3), .ZN(n79) );
  INV_X1 U12 ( .A(n90), .ZN(Z[2]) );
  AOI22_X1 U13 ( .A1(A[2]), .A2(n1), .B1(B[2]), .B2(n2), .ZN(n90) );
  INV_X1 U14 ( .A(n93), .ZN(Z[3]) );
  AOI22_X1 U15 ( .A1(A[3]), .A2(n1), .B1(B[3]), .B2(n2), .ZN(n93) );
  INV_X1 U16 ( .A(n94), .ZN(Z[4]) );
  AOI22_X1 U17 ( .A1(A[4]), .A2(n1), .B1(B[4]), .B2(n2), .ZN(n94) );
  INV_X1 U18 ( .A(n95), .ZN(Z[5]) );
  AOI22_X1 U19 ( .A1(A[5]), .A2(n1), .B1(B[5]), .B2(n3), .ZN(n95) );
  INV_X1 U20 ( .A(n96), .ZN(Z[6]) );
  AOI22_X1 U21 ( .A1(A[6]), .A2(n1), .B1(B[6]), .B2(n3), .ZN(n96) );
  INV_X1 U22 ( .A(n97), .ZN(Z[7]) );
  AOI22_X1 U23 ( .A1(A[7]), .A2(n1), .B1(B[7]), .B2(n3), .ZN(n97) );
  INV_X1 U24 ( .A(n98), .ZN(Z[8]) );
  AOI22_X1 U25 ( .A1(A[8]), .A2(n1), .B1(B[8]), .B2(n3), .ZN(n98) );
  INV_X1 U26 ( .A(n69), .ZN(Z[10]) );
  AOI22_X1 U27 ( .A1(A[10]), .A2(n1), .B1(B[10]), .B2(n3), .ZN(n69) );
  INV_X1 U28 ( .A(n70), .ZN(Z[11]) );
  AOI22_X1 U29 ( .A1(A[11]), .A2(n1), .B1(B[11]), .B2(n3), .ZN(n70) );
  INV_X1 U30 ( .A(n71), .ZN(Z[12]) );
  AOI22_X1 U31 ( .A1(A[12]), .A2(n1), .B1(B[12]), .B2(n3), .ZN(n71) );
  INV_X1 U32 ( .A(n72), .ZN(Z[13]) );
  AOI22_X1 U33 ( .A1(A[13]), .A2(n1), .B1(B[13]), .B2(n3), .ZN(n72) );
  INV_X1 U34 ( .A(n73), .ZN(Z[14]) );
  AOI22_X1 U35 ( .A1(A[14]), .A2(n1), .B1(B[14]), .B2(n3), .ZN(n73) );
  INV_X1 U36 ( .A(n74), .ZN(Z[15]) );
  AOI22_X1 U37 ( .A1(A[15]), .A2(n1), .B1(B[15]), .B2(n3), .ZN(n74) );
  INV_X1 U38 ( .A(n75), .ZN(Z[16]) );
  AOI22_X1 U39 ( .A1(A[16]), .A2(n1), .B1(B[16]), .B2(n3), .ZN(n75) );
  INV_X1 U40 ( .A(n76), .ZN(Z[17]) );
  AOI22_X1 U41 ( .A1(A[17]), .A2(n1), .B1(B[17]), .B2(n3), .ZN(n76) );
  INV_X1 U42 ( .A(n77), .ZN(Z[18]) );
  AOI22_X1 U43 ( .A1(A[18]), .A2(n1), .B1(B[18]), .B2(n3), .ZN(n77) );
  INV_X1 U44 ( .A(n78), .ZN(Z[19]) );
  AOI22_X1 U45 ( .A1(A[19]), .A2(n1), .B1(B[19]), .B2(n3), .ZN(n78) );
  INV_X1 U46 ( .A(n80), .ZN(Z[20]) );
  AOI22_X1 U47 ( .A1(A[20]), .A2(n1), .B1(B[20]), .B2(n3), .ZN(n80) );
  INV_X1 U48 ( .A(n81), .ZN(Z[21]) );
  AOI22_X1 U49 ( .A1(A[21]), .A2(n1), .B1(B[21]), .B2(n3), .ZN(n81) );
  INV_X1 U50 ( .A(n82), .ZN(Z[22]) );
  AOI22_X1 U51 ( .A1(A[22]), .A2(n1), .B1(B[22]), .B2(n3), .ZN(n82) );
  INV_X1 U52 ( .A(n83), .ZN(Z[23]) );
  AOI22_X1 U53 ( .A1(A[23]), .A2(n1), .B1(B[23]), .B2(n3), .ZN(n83) );
  INV_X1 U54 ( .A(n84), .ZN(Z[24]) );
  AOI22_X1 U55 ( .A1(A[24]), .A2(n1), .B1(B[24]), .B2(n3), .ZN(n84) );
  INV_X1 U56 ( .A(n85), .ZN(Z[25]) );
  AOI22_X1 U57 ( .A1(A[25]), .A2(n1), .B1(B[25]), .B2(n3), .ZN(n85) );
  INV_X1 U58 ( .A(n99), .ZN(Z[9]) );
  AOI22_X1 U59 ( .A1(A[9]), .A2(n1), .B1(n3), .B2(B[9]), .ZN(n99) );
  INV_X1 U60 ( .A(n68), .ZN(Z[0]) );
  AOI22_X1 U61 ( .A1(A[0]), .A2(n1), .B1(B[0]), .B2(n3), .ZN(n68) );
  AOI22_X1 U62 ( .A1(A[29]), .A2(n1), .B1(B[29]), .B2(n3), .ZN(n89) );
  AOI22_X1 U63 ( .A1(A[30]), .A2(n1), .B1(B[30]), .B2(n3), .ZN(n91) );
  AOI22_X1 U64 ( .A1(A[27]), .A2(n1), .B1(B[27]), .B2(n3), .ZN(n87) );
  AOI22_X1 U65 ( .A1(A[28]), .A2(n1), .B1(B[28]), .B2(n3), .ZN(n88) );
  AOI22_X1 U66 ( .A1(A[26]), .A2(n1), .B1(B[26]), .B2(n3), .ZN(n86) );
  AOI22_X1 U67 ( .A1(A[31]), .A2(n1), .B1(B[31]), .B2(n2), .ZN(n92) );
endmodule


module regn_N32_0 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n9, n10, n11, n12, n13, n14, n16, n17, n18, n19, n20, n21, n22;

  DFFR_X1 \DOUT_reg[31]  ( .D(n96), .CK(CLK), .RN(n11), .Q(DOUT[31]) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n95), .CK(CLK), .RN(n11), .Q(DOUT[30]) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n94), .CK(CLK), .RN(n11), .Q(DOUT[29]) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n93), .CK(CLK), .RN(n11), .Q(DOUT[28]) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n92), .CK(CLK), .RN(n11), .Q(DOUT[27]) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n91), .CK(CLK), .RN(n11), .Q(DOUT[26]) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n90), .CK(CLK), .RN(n11), .Q(DOUT[25]) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n89), .CK(CLK), .RN(n11), .Q(DOUT[24]) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n88), .CK(CLK), .RN(n10), .Q(DOUT[23]) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n87), .CK(CLK), .RN(n10), .Q(DOUT[22]) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n86), .CK(CLK), .RN(n10), .Q(DOUT[21]) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n85), .CK(CLK), .RN(n10), .Q(DOUT[20]) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n84), .CK(CLK), .RN(n10), .Q(DOUT[19]) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n83), .CK(CLK), .RN(n10), .Q(DOUT[18]), .QN(n51)
         );
  DFFR_X1 \DOUT_reg[17]  ( .D(n82), .CK(CLK), .RN(n10), .Q(DOUT[17]), .QN(n50)
         );
  DFFR_X1 \DOUT_reg[16]  ( .D(n81), .CK(CLK), .RN(n10), .Q(DOUT[16]), .QN(n49)
         );
  DFFR_X1 \DOUT_reg[15]  ( .D(n80), .CK(CLK), .RN(n10), .Q(DOUT[15]), .QN(n48)
         );
  DFFR_X1 \DOUT_reg[14]  ( .D(n79), .CK(CLK), .RN(n10), .Q(DOUT[14]), .QN(n47)
         );
  DFFR_X1 \DOUT_reg[13]  ( .D(n78), .CK(CLK), .RN(n10), .Q(DOUT[13]), .QN(n46)
         );
  DFFR_X1 \DOUT_reg[12]  ( .D(n77), .CK(CLK), .RN(n10), .Q(DOUT[12]), .QN(n45)
         );
  DFFR_X1 \DOUT_reg[11]  ( .D(n76), .CK(CLK), .RN(n9), .Q(DOUT[11]) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n75), .CK(CLK), .RN(n9), .Q(DOUT[10]), .QN(n43)
         );
  DFFR_X1 \DOUT_reg[9]  ( .D(n74), .CK(CLK), .RN(n9), .Q(DOUT[9]), .QN(n42) );
  DFFR_X1 \DOUT_reg[8]  ( .D(n73), .CK(CLK), .RN(n9), .Q(DOUT[8]), .QN(n41) );
  DFFR_X1 \DOUT_reg[7]  ( .D(n72), .CK(CLK), .RN(n9), .Q(DOUT[7]), .QN(n40) );
  DFFR_X1 \DOUT_reg[6]  ( .D(n71), .CK(CLK), .RN(n9), .Q(DOUT[6]), .QN(n39) );
  DFFR_X1 \DOUT_reg[5]  ( .D(n70), .CK(CLK), .RN(n9), .Q(DOUT[5]), .QN(n38) );
  DFFR_X1 \DOUT_reg[4]  ( .D(n69), .CK(CLK), .RN(n9), .Q(DOUT[4]), .QN(n37) );
  DFFR_X1 \DOUT_reg[3]  ( .D(n68), .CK(CLK), .RN(n9), .Q(DOUT[3]), .QN(n36) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n67), .CK(CLK), .RN(n9), .Q(DOUT[2]), .QN(n35) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n66), .CK(CLK), .RN(n9), .Q(DOUT[1]), .QN(n34) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n65), .CK(CLK), .RN(n9), .Q(DOUT[0]), .QN(n33) );
  BUF_X1 U2 ( .A(RST), .Z(n9) );
  BUF_X1 U3 ( .A(RST), .Z(n10) );
  BUF_X1 U4 ( .A(RST), .Z(n11) );
  OAI21_X1 U5 ( .B1(n34), .B2(EN), .A(n2), .ZN(n66) );
  NAND2_X1 U6 ( .A1(DIN[1]), .A2(EN), .ZN(n2) );
  OAI21_X1 U7 ( .B1(n35), .B2(EN), .A(n3), .ZN(n67) );
  NAND2_X1 U8 ( .A1(DIN[2]), .A2(EN), .ZN(n3) );
  OAI21_X1 U9 ( .B1(n36), .B2(EN), .A(n4), .ZN(n68) );
  NAND2_X1 U10 ( .A1(DIN[3]), .A2(EN), .ZN(n4) );
  OAI21_X1 U11 ( .B1(n40), .B2(EN), .A(n8), .ZN(n72) );
  NAND2_X1 U12 ( .A1(DIN[7]), .A2(EN), .ZN(n8) );
  OAI21_X1 U13 ( .B1(n39), .B2(EN), .A(n7), .ZN(n71) );
  NAND2_X1 U14 ( .A1(DIN[6]), .A2(EN), .ZN(n7) );
  OAI21_X1 U15 ( .B1(n38), .B2(EN), .A(n6), .ZN(n70) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n6) );
  OAI21_X1 U17 ( .B1(n37), .B2(EN), .A(n5), .ZN(n69) );
  NAND2_X1 U18 ( .A1(DIN[4]), .A2(EN), .ZN(n5) );
  OAI21_X1 U19 ( .B1(n33), .B2(EN), .A(n1), .ZN(n65) );
  NAND2_X1 U20 ( .A1(EN), .A2(DIN[0]), .ZN(n1) );
  INV_X1 U21 ( .A(n41), .ZN(n12) );
  MUX2_X1 U22 ( .A(n12), .B(DIN[8]), .S(EN), .Z(n73) );
  INV_X1 U23 ( .A(n42), .ZN(n13) );
  MUX2_X1 U24 ( .A(n13), .B(DIN[9]), .S(EN), .Z(n74) );
  INV_X1 U25 ( .A(n43), .ZN(n14) );
  MUX2_X1 U26 ( .A(n14), .B(DIN[10]), .S(EN), .Z(n75) );
  MUX2_X1 U27 ( .A(DOUT[11]), .B(DIN[11]), .S(EN), .Z(n76) );
  INV_X1 U28 ( .A(n45), .ZN(n16) );
  MUX2_X1 U29 ( .A(n16), .B(DIN[12]), .S(EN), .Z(n77) );
  INV_X1 U30 ( .A(n46), .ZN(n17) );
  MUX2_X1 U31 ( .A(n17), .B(DIN[13]), .S(EN), .Z(n78) );
  INV_X1 U32 ( .A(n47), .ZN(n18) );
  MUX2_X1 U33 ( .A(n18), .B(DIN[14]), .S(EN), .Z(n79) );
  INV_X1 U34 ( .A(n48), .ZN(n19) );
  MUX2_X1 U35 ( .A(n19), .B(DIN[15]), .S(EN), .Z(n80) );
  INV_X1 U36 ( .A(n49), .ZN(n20) );
  MUX2_X1 U37 ( .A(n20), .B(DIN[16]), .S(EN), .Z(n81) );
  INV_X1 U38 ( .A(n50), .ZN(n21) );
  MUX2_X1 U39 ( .A(n21), .B(DIN[17]), .S(EN), .Z(n82) );
  INV_X1 U40 ( .A(n51), .ZN(n22) );
  MUX2_X1 U41 ( .A(n22), .B(DIN[18]), .S(EN), .Z(n83) );
  MUX2_X1 U42 ( .A(DOUT[19]), .B(DIN[19]), .S(EN), .Z(n84) );
  MUX2_X1 U43 ( .A(DOUT[20]), .B(DIN[20]), .S(EN), .Z(n85) );
  MUX2_X1 U44 ( .A(DOUT[21]), .B(DIN[21]), .S(EN), .Z(n86) );
  MUX2_X1 U45 ( .A(DOUT[22]), .B(DIN[22]), .S(EN), .Z(n87) );
  MUX2_X1 U46 ( .A(DOUT[23]), .B(DIN[23]), .S(EN), .Z(n88) );
  MUX2_X1 U47 ( .A(DOUT[24]), .B(DIN[24]), .S(EN), .Z(n89) );
  MUX2_X1 U48 ( .A(DOUT[25]), .B(DIN[25]), .S(EN), .Z(n90) );
  MUX2_X1 U49 ( .A(DOUT[26]), .B(DIN[26]), .S(EN), .Z(n91) );
  MUX2_X1 U50 ( .A(DOUT[27]), .B(DIN[27]), .S(EN), .Z(n92) );
  MUX2_X1 U51 ( .A(DOUT[28]), .B(DIN[28]), .S(EN), .Z(n93) );
  MUX2_X1 U52 ( .A(DOUT[29]), .B(DIN[29]), .S(EN), .Z(n94) );
  MUX2_X1 U53 ( .A(DOUT[30]), .B(DIN[30]), .S(EN), .Z(n95) );
  MUX2_X1 U54 ( .A(DOUT[31]), .B(DIN[31]), .S(EN), .Z(n96) );
endmodule


module regn_N32_9 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U6 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U7 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U10 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U11 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U24 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U25 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U26 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U27 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U28 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U29 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U30 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U31 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U32 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U33 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U34 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U35 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U36 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U37 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U38 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U39 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U40 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U41 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U42 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U43 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U44 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U45 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U46 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U47 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U48 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U49 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U50 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U51 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U52 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U53 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U54 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U55 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U56 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U57 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U58 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U59 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U60 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U61 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U62 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U63 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U64 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U65 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U66 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
  OAI21_X1 U67 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U68 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
endmodule


module regn_N32_8 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  DFFR_X2 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X2 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X2 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  NAND2_X1 U5 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  NAND2_X1 U6 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  NAND2_X1 U7 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  NAND2_X1 U8 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
  NAND2_X1 U9 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U10 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U11 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U12 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U13 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U14 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U15 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U16 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U17 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U18 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U19 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U20 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U21 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U22 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U23 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U24 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U25 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U26 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U27 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U28 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U29 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U30 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U31 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U32 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U33 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U34 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U35 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U36 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U37 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U38 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U39 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U40 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U41 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U42 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U43 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U44 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U45 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U46 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U47 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U48 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U49 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U50 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U51 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U52 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U53 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U54 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U55 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U56 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U57 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U58 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U59 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U60 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U61 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U62 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U63 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U64 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  OAI21_X1 U65 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  OAI21_X1 U66 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  OAI21_X1 U68 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
endmodule


module Fetch_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AND3_X1 U2 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n1) );
  AND2_X1 U3 ( .A1(n40), .A2(n53), .ZN(n2) );
  AND2_X1 U4 ( .A1(n40), .A2(n66), .ZN(n3) );
  AND2_X1 U5 ( .A1(n12), .A2(n25), .ZN(n23) );
  NOR2_X1 U6 ( .A1(n15), .A2(n17), .ZN(n108) );
  NOR2_X1 U7 ( .A1(n45), .A2(n47), .ZN(n49) );
  NOR2_X1 U8 ( .A1(n45), .A2(n41), .ZN(n44) );
  NAND2_X1 U9 ( .A1(n19), .A2(n20), .ZN(n15) );
  NOR2_X1 U10 ( .A1(n99), .A2(n5), .ZN(n4) );
  OR2_X1 U11 ( .A1(n97), .A2(n98), .ZN(n5) );
  AND2_X1 U12 ( .A1(n38), .A2(n40), .ZN(n6) );
  AND2_X1 U13 ( .A1(n59), .A2(n40), .ZN(n7) );
  OR2_X1 U14 ( .A1(n98), .A2(n99), .ZN(n100) );
  INV_X1 U15 ( .A(n34), .ZN(n33) );
  INV_X1 U16 ( .A(n97), .ZN(n101) );
  AND2_X1 U17 ( .A1(n22), .A2(n23), .ZN(n8) );
  AND2_X1 U18 ( .A1(n107), .A2(n108), .ZN(n9) );
  INV_X1 U19 ( .A(n29), .ZN(n31) );
  INV_X1 U20 ( .A(n22), .ZN(n24) );
  INV_X1 U21 ( .A(n25), .ZN(n27) );
  INV_X1 U22 ( .A(n17), .ZN(n16) );
  INV_X1 U23 ( .A(n20), .ZN(n18) );
  INV_X1 U24 ( .A(n107), .ZN(n109) );
  INV_X1 U25 ( .A(n80), .ZN(n40) );
  NOR2_X1 U26 ( .A1(n83), .A2(n84), .ZN(n82) );
  NOR2_X1 U27 ( .A1(n85), .A2(n86), .ZN(n81) );
  NAND4_X1 U28 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(A[19]), .ZN(n68) );
  AND2_X1 U29 ( .A1(n4), .A2(A[13]), .ZN(n94) );
  NOR2_X1 U30 ( .A1(n111), .A2(n103), .ZN(n19) );
  NAND4_X1 U31 ( .A1(A[24]), .A2(A[25]), .A3(A[26]), .A4(A[27]), .ZN(n47) );
  NAND4_X1 U32 ( .A1(A[4]), .A2(A[5]), .A3(n90), .A4(A[7]), .ZN(n103) );
  NAND4_X1 U33 ( .A1(n107), .A2(n110), .A3(n20), .A4(A[11]), .ZN(n98) );
  INV_X1 U34 ( .A(n105), .ZN(n110) );
  NAND4_X1 U35 ( .A1(A[14]), .A2(A[15]), .A3(A[3]), .A4(A[7]), .ZN(n83) );
  NOR2_X1 U36 ( .A1(n41), .A2(n43), .ZN(n39) );
  AND3_X1 U37 ( .A1(A[16]), .A2(A[17]), .A3(n40), .ZN(n10) );
  AND2_X1 U38 ( .A1(n40), .A2(A[16]), .ZN(n11) );
  NAND2_X1 U39 ( .A1(n58), .A2(n59), .ZN(n55) );
  NOR2_X1 U40 ( .A1(n60), .A2(n61), .ZN(n58) );
  NAND2_X1 U41 ( .A1(A[22]), .A2(A[23]), .ZN(n60) );
  NAND2_X1 U42 ( .A1(n62), .A2(A[21]), .ZN(n61) );
  NAND2_X1 U43 ( .A1(n102), .A2(n28), .ZN(n99) );
  NAND2_X1 U44 ( .A1(n46), .A2(A[28]), .ZN(n41) );
  NOR2_X1 U45 ( .A1(n54), .A2(n55), .ZN(n53) );
  NAND2_X1 U46 ( .A1(A[25]), .A2(A[24]), .ZN(n54) );
  AND2_X1 U47 ( .A1(n28), .A2(n29), .ZN(n12) );
  NOR2_X1 U48 ( .A1(n67), .A2(n68), .ZN(n66) );
  NAND2_X1 U49 ( .A1(A[21]), .A2(n62), .ZN(n67) );
  INV_X1 U50 ( .A(n32), .ZN(n29) );
  INV_X1 U51 ( .A(n104), .ZN(n20) );
  NAND2_X1 U52 ( .A1(n72), .A2(n40), .ZN(n69) );
  NOR2_X1 U53 ( .A1(n68), .A2(n73), .ZN(n72) );
  INV_X1 U54 ( .A(n26), .ZN(n22) );
  INV_X1 U55 ( .A(n89), .ZN(n107) );
  AND2_X1 U56 ( .A1(n10), .A2(A[18]), .ZN(n76) );
  AND2_X1 U57 ( .A1(n2), .A2(A[26]), .ZN(n51) );
  AND2_X1 U58 ( .A1(n3), .A2(A[22]), .ZN(n64) );
  NAND2_X1 U59 ( .A1(A[14]), .A2(n94), .ZN(n91) );
  AND2_X1 U60 ( .A1(n6), .A2(A[24]), .ZN(n13) );
  INV_X1 U61 ( .A(n26), .ZN(n90) );
  INV_X1 U62 ( .A(n30), .ZN(n25) );
  INV_X1 U63 ( .A(A[24]), .ZN(n57) );
  INV_X1 U64 ( .A(A[16]), .ZN(n79) );
  AND2_X1 U65 ( .A1(n1), .A2(A[30]), .ZN(n14) );
  INV_X1 U66 ( .A(n71), .ZN(n70) );
  INV_X1 U67 ( .A(n93), .ZN(n92) );
  INV_X1 U68 ( .A(n62), .ZN(n73) );
  INV_X1 U69 ( .A(A[7]), .ZN(n21) );
  INV_X1 U70 ( .A(A[25]), .ZN(n56) );
  INV_X1 U71 ( .A(A[11]), .ZN(n106) );
  INV_X1 U72 ( .A(A[18]), .ZN(n77) );
  INV_X1 U73 ( .A(A[26]), .ZN(n52) );
  INV_X1 U74 ( .A(A[17]), .ZN(n78) );
  INV_X1 U75 ( .A(A[22]), .ZN(n65) );
  INV_X1 U76 ( .A(A[13]), .ZN(n96) );
  INV_X1 U77 ( .A(A[28]), .ZN(n48) );
  INV_X1 U78 ( .A(A[29]), .ZN(n43) );
  INV_X1 U79 ( .A(A[14]), .ZN(n95) );
  INV_X1 U80 ( .A(A[19]), .ZN(n75) );
  INV_X1 U81 ( .A(A[27]), .ZN(n50) );
  INV_X1 U82 ( .A(A[23]), .ZN(n63) );
  NOR2_X1 U83 ( .A1(n34), .A2(n42), .ZN(n28) );
  INV_X1 U84 ( .A(A[2]), .ZN(n42) );
  XNOR2_X1 U85 ( .A(n106), .B(n9), .ZN(SUM[11]) );
  XNOR2_X1 U86 ( .A(n40), .B(n79), .ZN(SUM[16]) );
  XNOR2_X1 U87 ( .A(n21), .B(n8), .ZN(SUM[7]) );
  INV_X1 U88 ( .A(n74), .ZN(n62) );
  INV_X1 U89 ( .A(A[20]), .ZN(n74) );
  XNOR2_X1 U90 ( .A(n69), .B(n70), .ZN(SUM[21]) );
  XNOR2_X1 U91 ( .A(n91), .B(n92), .ZN(SUM[15]) );
  XNOR2_X1 U92 ( .A(n100), .B(n101), .ZN(SUM[12]) );
  XNOR2_X1 U93 ( .A(n1), .B(n37), .ZN(SUM[30]) );
  XNOR2_X1 U94 ( .A(n6), .B(n57), .ZN(SUM[24]) );
  XNOR2_X1 U95 ( .A(n73), .B(n7), .ZN(SUM[20]) );
  XNOR2_X1 U96 ( .A(n56), .B(n13), .ZN(SUM[25]) );
  XNOR2_X1 U97 ( .A(n77), .B(n10), .ZN(SUM[18]) );
  XNOR2_X1 U98 ( .A(n52), .B(n2), .ZN(SUM[26]) );
  XNOR2_X1 U99 ( .A(n48), .B(n49), .ZN(SUM[28]) );
  XNOR2_X1 U100 ( .A(n78), .B(n11), .ZN(SUM[17]) );
  XNOR2_X1 U101 ( .A(n43), .B(n44), .ZN(SUM[29]) );
  XNOR2_X1 U102 ( .A(n65), .B(n3), .ZN(SUM[22]) );
  XNOR2_X1 U103 ( .A(n96), .B(n4), .ZN(SUM[13]) );
  INV_X1 U104 ( .A(A[6]), .ZN(n26) );
  INV_X1 U105 ( .A(A[4]), .ZN(n32) );
  INV_X1 U106 ( .A(A[8]), .ZN(n104) );
  INV_X1 U107 ( .A(A[9]), .ZN(n105) );
  INV_X1 U108 ( .A(A[5]), .ZN(n30) );
  INV_X1 U109 ( .A(A[30]), .ZN(n37) );
  INV_X1 U110 ( .A(A[2]), .ZN(SUM[2]) );
  XNOR2_X1 U111 ( .A(SUM[2]), .B(n33), .ZN(SUM[3]) );
  XNOR2_X1 U112 ( .A(n24), .B(n23), .ZN(SUM[6]) );
  XNOR2_X1 U113 ( .A(n27), .B(n12), .ZN(SUM[5]) );
  XNOR2_X1 U114 ( .A(n31), .B(n28), .ZN(SUM[4]) );
  XNOR2_X1 U115 ( .A(n36), .B(n14), .ZN(SUM[31]) );
  INV_X1 U116 ( .A(A[15]), .ZN(n93) );
  INV_X1 U117 ( .A(A[31]), .ZN(n36) );
  XNOR2_X1 U118 ( .A(n15), .B(n16), .ZN(SUM[9]) );
  XNOR2_X1 U119 ( .A(n18), .B(n19), .ZN(SUM[8]) );
  INV_X1 U120 ( .A(n47), .ZN(n46) );
  INV_X1 U121 ( .A(n6), .ZN(n45) );
  XNOR2_X1 U122 ( .A(n50), .B(n51), .ZN(SUM[27]) );
  INV_X1 U123 ( .A(n55), .ZN(n38) );
  XNOR2_X1 U124 ( .A(n63), .B(n64), .ZN(SUM[23]) );
  INV_X1 U125 ( .A(A[21]), .ZN(n71) );
  INV_X1 U126 ( .A(n68), .ZN(n59) );
  XNOR2_X1 U127 ( .A(n75), .B(n76), .ZN(SUM[19]) );
  NAND2_X1 U128 ( .A1(n81), .A2(n82), .ZN(n80) );
  NAND3_X1 U129 ( .A1(A[11]), .A2(A[13]), .A3(A[12]), .ZN(n84) );
  NAND3_X1 U130 ( .A1(A[4]), .A2(A[5]), .A3(A[2]), .ZN(n86) );
  NAND2_X1 U131 ( .A1(n87), .A2(n88), .ZN(n85) );
  NOR2_X1 U132 ( .A1(n104), .A2(n105), .ZN(n88) );
  NOR2_X1 U133 ( .A1(n89), .A2(n26), .ZN(n87) );
  INV_X1 U134 ( .A(A[10]), .ZN(n89) );
  XNOR2_X1 U135 ( .A(n95), .B(n94), .ZN(SUM[14]) );
  INV_X1 U136 ( .A(A[12]), .ZN(n97) );
  INV_X1 U137 ( .A(n103), .ZN(n102) );
  XNOR2_X1 U138 ( .A(n109), .B(n108), .ZN(SUM[10]) );
  INV_X1 U139 ( .A(n110), .ZN(n17) );
  INV_X1 U140 ( .A(n28), .ZN(n111) );
  INV_X1 U141 ( .A(A[3]), .ZN(n34) );
endmodule


module Fetch ( CLK, RST, ZERO_FLAG, PC_EXT, INS_IN, Bubble_in, HDU_INS_IN, 
        HDU_PC_IN, HDU_NPC_IN, PC_OUT, ADDR_OUT, NPC_OUT, INS_OUT );
  input [31:0] PC_EXT;
  input [31:0] INS_IN;
  input [31:0] HDU_INS_IN;
  input [31:0] HDU_PC_IN;
  input [31:0] HDU_NPC_IN;
  output [31:0] PC_OUT;
  output [31:0] ADDR_OUT;
  output [31:0] NPC_OUT;
  output [31:0] INS_OUT;
  input CLK, RST, ZERO_FLAG, Bubble_in;
  wire   sig_RST, n4;
  wire   [31:0] sig_NPC;
  wire   [31:0] PC_MUX_OUT;
  wire   [31:0] sig_INS;

  mux21_NBIT32_0 NPC_or_NPC_HDU ( .A(PC_EXT), .B(HDU_NPC_IN), .S(Bubble_in), 
        .Z(sig_NPC) );
  mux21_NBIT32_6 PC_or_PC_HDU ( .A(ADDR_OUT), .B(HDU_PC_IN), .S(Bubble_in), 
        .Z(PC_MUX_OUT) );
  mux21_NBIT32_5 INS_or_HDU_INS ( .A(INS_IN), .B(HDU_INS_IN), .S(Bubble_in), 
        .Z(sig_INS) );
  regn_N32_0 PC ( .DIN(sig_NPC), .CLK(CLK), .EN(1'b1), .RST(RST), .DOUT(
        ADDR_OUT) );
  regn_N32_9 PC_reg ( .DIN(PC_MUX_OUT), .CLK(CLK), .EN(1'b1), .RST(sig_RST), 
        .DOUT(PC_OUT) );
  regn_N32_8 IR ( .DIN(sig_INS), .CLK(CLK), .EN(1'b1), .RST(sig_RST), .DOUT(
        INS_OUT) );
  Fetch_DW01_add_1 add_54 ( .A(ADDR_OUT), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(NPC_OUT) );
  NOR2_X1 U6 ( .A1(ZERO_FLAG), .A2(n4), .ZN(sig_RST) );
  INV_X1 U7 ( .A(RST), .ZN(n4) );
endmodule


module instruction_type ( INST_IN, Rtype, Itype, Jtype );
  input [31:0] INST_IN;
  output Rtype, Itype, Jtype;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;

  BUF_X1 U1 ( .A(INST_IN[30]), .Z(n5) );
  CLKBUF_X1 U2 ( .A(n9), .Z(n1) );
  BUF_X1 U3 ( .A(INST_IN[26]), .Z(n9) );
  INV_X1 U4 ( .A(INST_IN[30]), .ZN(n2) );
  INV_X1 U5 ( .A(INST_IN[30]), .ZN(n3) );
  CLKBUF_X1 U6 ( .A(INST_IN[27]), .Z(n4) );
  INV_X1 U7 ( .A(n15), .ZN(n6) );
  INV_X1 U8 ( .A(INST_IN[27]), .ZN(n7) );
  NAND4_X1 U9 ( .A1(n13), .A2(n11), .A3(n2), .A4(n18), .ZN(n8) );
  INV_X1 U10 ( .A(INST_IN[31]), .ZN(n10) );
  INV_X1 U11 ( .A(INST_IN[28]), .ZN(n13) );
  INV_X1 U12 ( .A(INST_IN[29]), .ZN(n11) );
  INV_X1 U13 ( .A(INST_IN[30]), .ZN(n24) );
  INV_X1 U14 ( .A(INST_IN[31]), .ZN(n18) );
  NAND4_X1 U15 ( .A1(n13), .A2(n11), .A3(n24), .A4(n18), .ZN(n28) );
  INV_X1 U16 ( .A(INST_IN[27]), .ZN(n15) );
  NOR2_X1 U17 ( .A1(n15), .A2(n8), .ZN(Jtype) );
  MUX2_X1 U18 ( .A(n2), .B(n10), .S(INST_IN[29]), .Z(n12) );
  NAND3_X1 U19 ( .A1(n15), .A2(INST_IN[28]), .A3(n12), .ZN(n27) );
  OAI211_X1 U20 ( .C1(n13), .C2(n24), .A(INST_IN[29]), .B(n10), .ZN(n26) );
  NAND3_X1 U21 ( .A1(n9), .A2(n7), .A3(INST_IN[28]), .ZN(n14) );
  OAI211_X1 U22 ( .C1(INST_IN[28]), .C2(n15), .A(n14), .B(INST_IN[29]), .ZN(
        n23) );
  XOR2_X1 U23 ( .A(INST_IN[27]), .B(INST_IN[26]), .Z(n16) );
  NOR3_X1 U24 ( .A1(n16), .A2(INST_IN[28]), .A3(n10), .ZN(n22) );
  INV_X1 U25 ( .A(INST_IN[26]), .ZN(n17) );
  NAND3_X1 U26 ( .A1(INST_IN[28]), .A2(n18), .A3(n17), .ZN(n20) );
  AOI21_X1 U27 ( .B1(n4), .B2(n18), .A(INST_IN[29]), .ZN(n19) );
  NAND3_X1 U28 ( .A1(n19), .A2(n20), .A3(n5), .ZN(n21) );
  OAI221_X1 U29 ( .B1(n23), .B2(n3), .C1(n22), .C2(n5), .A(n21), .ZN(n25) );
  NAND3_X1 U30 ( .A1(n25), .A2(n26), .A3(n27), .ZN(Itype) );
  NOR3_X1 U31 ( .A1(n28), .A2(n1), .A3(n6), .ZN(Rtype) );
endmodule


module instruction_decomposition ( INST_IN, Rtype, Itype, Jtype, ADD_RS1, 
        ADD_RS2, ADD_WR, IMM, RD1, RD2 );
  input [31:0] INST_IN;
  output [4:0] ADD_RS1;
  output [4:0] ADD_RS2;
  output [4:0] ADD_WR;
  output [31:0] IMM;
  input Rtype, Itype, Jtype;
  output RD1, RD2;
  wire   n56, n33, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, \IMM[31] , n50, n51, n52, n53, n54, n55;
  assign IMM[25] = \IMM[31] ;
  assign IMM[26] = \IMM[31] ;
  assign IMM[27] = \IMM[31] ;
  assign IMM[28] = \IMM[31] ;
  assign IMM[29] = \IMM[31] ;
  assign IMM[30] = \IMM[31] ;
  assign IMM[31] = \IMM[31] ;

  INV_X1 U3 ( .A(RD1), .ZN(n1) );
  CLKBUF_X1 U4 ( .A(n7), .Z(RD1) );
  CLKBUF_X1 U5 ( .A(n1), .Z(n3) );
  BUF_X1 U6 ( .A(n56), .Z(n7) );
  AND2_X1 U7 ( .A1(n56), .A2(INST_IN[23]), .ZN(ADD_RS1[2]) );
  NOR2_X1 U8 ( .A1(n17), .A2(n18), .ZN(n4) );
  NOR2_X1 U9 ( .A1(n19), .A2(n5), .ZN(n20) );
  INV_X1 U10 ( .A(n4), .ZN(n5) );
  BUF_X1 U11 ( .A(n31), .Z(n8) );
  AND2_X2 U12 ( .A1(n7), .A2(INST_IN[21]), .ZN(ADD_RS1[0]) );
  AND2_X2 U13 ( .A1(n41), .A2(n13), .ZN(n14) );
  AND2_X1 U14 ( .A1(n31), .A2(n12), .ZN(n6) );
  AND2_X1 U15 ( .A1(n31), .A2(n12), .ZN(n15) );
  INV_X1 U16 ( .A(n16), .ZN(n9) );
  AOI211_X4 U17 ( .C1(n16), .C2(n13), .A(n34), .B(n15), .ZN(ADD_RS2[1]) );
  CLKBUF_X1 U18 ( .A(n13), .Z(n10) );
  NAND2_X1 U19 ( .A1(INST_IN[15]), .A2(n24), .ZN(n25) );
  AND2_X1 U20 ( .A1(n29), .A2(n28), .ZN(n11) );
  INV_X1 U21 ( .A(INST_IN[15]), .ZN(n51) );
  INV_X1 U22 ( .A(INST_IN[11]), .ZN(n55) );
  INV_X1 U23 ( .A(INST_IN[12]), .ZN(n54) );
  INV_X1 U24 ( .A(INST_IN[13]), .ZN(n53) );
  INV_X1 U25 ( .A(INST_IN[14]), .ZN(n52) );
  CLKBUF_X1 U26 ( .A(n40), .Z(n12) );
  BUF_X2 U27 ( .A(n40), .Z(n13) );
  NAND2_X1 U28 ( .A1(n3), .A2(Jtype), .ZN(n28) );
  INV_X1 U29 ( .A(n56), .ZN(n45) );
  NOR2_X1 U30 ( .A1(n43), .A2(n14), .ZN(ADD_RS1[3]) );
  AND2_X2 U31 ( .A1(RD2), .A2(INST_IN[18]), .ZN(ADD_RS2[2]) );
  INV_X1 U32 ( .A(Itype), .ZN(n16) );
  NOR3_X1 U33 ( .A1(n14), .A2(n6), .A3(n36), .ZN(ADD_RS2[3]) );
  OR4_X1 U34 ( .A1(n50), .A2(INST_IN[28]), .A3(INST_IN[29]), .A4(INST_IN[31]), 
        .ZN(n33) );
  NOR3_X2 U35 ( .A1(n14), .A2(n6), .A3(n32), .ZN(ADD_RS2[0]) );
  INV_X1 U36 ( .A(INST_IN[28]), .ZN(n21) );
  INV_X1 U37 ( .A(INST_IN[30]), .ZN(n26) );
  XOR2_X1 U38 ( .A(INST_IN[26]), .B(INST_IN[27]), .Z(n19) );
  INV_X1 U39 ( .A(INST_IN[31]), .ZN(n18) );
  INV_X1 U40 ( .A(INST_IN[29]), .ZN(n17) );
  NAND3_X1 U41 ( .A1(n20), .A2(n26), .A3(n21), .ZN(n31) );
  INV_X1 U42 ( .A(Itype), .ZN(n41) );
  INV_X1 U43 ( .A(Rtype), .ZN(n40) );
  OAI21_X1 U44 ( .B1(n8), .B2(n16), .A(n13), .ZN(RD2) );
  NAND2_X1 U45 ( .A1(n41), .A2(n13), .ZN(n56) );
  OAI21_X1 U46 ( .B1(Jtype), .B2(n9), .A(n10), .ZN(n23) );
  INV_X1 U47 ( .A(n23), .ZN(n22) );
  AND2_X1 U48 ( .A1(INST_IN[0]), .A2(n22), .ZN(IMM[0]) );
  AND2_X1 U49 ( .A1(INST_IN[1]), .A2(n22), .ZN(IMM[1]) );
  AND2_X1 U50 ( .A1(INST_IN[2]), .A2(n22), .ZN(IMM[2]) );
  AND2_X1 U51 ( .A1(INST_IN[3]), .A2(n22), .ZN(IMM[3]) );
  AND2_X1 U52 ( .A1(INST_IN[4]), .A2(n22), .ZN(IMM[4]) );
  AND2_X1 U53 ( .A1(INST_IN[5]), .A2(n22), .ZN(IMM[5]) );
  AND2_X1 U54 ( .A1(INST_IN[6]), .A2(n22), .ZN(IMM[6]) );
  AND2_X1 U55 ( .A1(INST_IN[7]), .A2(n22), .ZN(IMM[7]) );
  AND2_X1 U56 ( .A1(INST_IN[8]), .A2(n22), .ZN(IMM[8]) );
  AND2_X1 U57 ( .A1(INST_IN[9]), .A2(n22), .ZN(IMM[9]) );
  AND2_X1 U58 ( .A1(INST_IN[10]), .A2(n22), .ZN(IMM[10]) );
  NOR2_X1 U59 ( .A1(n55), .A2(n23), .ZN(IMM[11]) );
  NOR2_X1 U60 ( .A1(n54), .A2(n23), .ZN(IMM[12]) );
  NOR2_X1 U61 ( .A1(n53), .A2(n23), .ZN(IMM[13]) );
  NOR2_X1 U62 ( .A1(n52), .A2(n23), .ZN(IMM[14]) );
  NOR2_X1 U63 ( .A1(n51), .A2(n23), .ZN(IMM[15]) );
  INV_X1 U64 ( .A(INST_IN[16]), .ZN(n32) );
  NAND2_X1 U65 ( .A1(n9), .A2(n13), .ZN(n30) );
  INV_X1 U66 ( .A(n30), .ZN(n24) );
  OAI21_X1 U67 ( .B1(n32), .B2(n28), .A(n25), .ZN(IMM[16]) );
  INV_X1 U68 ( .A(INST_IN[17]), .ZN(n34) );
  OAI21_X1 U69 ( .B1(n34), .B2(n28), .A(n25), .ZN(IMM[17]) );
  INV_X1 U70 ( .A(INST_IN[18]), .ZN(n35) );
  OAI21_X1 U71 ( .B1(n35), .B2(n28), .A(n25), .ZN(IMM[18]) );
  INV_X1 U72 ( .A(INST_IN[19]), .ZN(n36) );
  OAI21_X1 U73 ( .B1(n36), .B2(n28), .A(n25), .ZN(IMM[19]) );
  INV_X1 U74 ( .A(INST_IN[20]), .ZN(n37) );
  OAI21_X1 U75 ( .B1(n37), .B2(n28), .A(n25), .ZN(IMM[20]) );
  INV_X1 U76 ( .A(INST_IN[21]), .ZN(n38) );
  OAI21_X1 U77 ( .B1(n38), .B2(n28), .A(n25), .ZN(IMM[21]) );
  INV_X1 U78 ( .A(INST_IN[22]), .ZN(n39) );
  OAI21_X1 U79 ( .B1(n39), .B2(n28), .A(n25), .ZN(IMM[22]) );
  INV_X1 U80 ( .A(INST_IN[23]), .ZN(n42) );
  OAI21_X1 U81 ( .B1(n42), .B2(n28), .A(n25), .ZN(IMM[23]) );
  INV_X1 U82 ( .A(INST_IN[24]), .ZN(n43) );
  OAI21_X1 U83 ( .B1(n43), .B2(n28), .A(n25), .ZN(IMM[24]) );
  INV_X1 U84 ( .A(INST_IN[25]), .ZN(n44) );
  OAI22_X1 U85 ( .A1(n51), .A2(n30), .B1(n44), .B2(n28), .ZN(\IMM[31] ) );
  INV_X1 U86 ( .A(INST_IN[26]), .ZN(n27) );
  OR4_X1 U87 ( .A1(n27), .A2(n26), .A3(n33), .A4(n30), .ZN(n29) );
  OAI221_X1 U88 ( .B1(n32), .B2(n30), .C1(n55), .C2(n10), .A(n11), .ZN(
        ADD_WR[0]) );
  OAI221_X1 U89 ( .B1(n34), .B2(n30), .C1(n54), .C2(n10), .A(n11), .ZN(
        ADD_WR[1]) );
  OAI221_X1 U90 ( .B1(n35), .B2(n30), .C1(n53), .C2(n10), .A(n11), .ZN(
        ADD_WR[2]) );
  OAI221_X1 U91 ( .B1(n36), .B2(n30), .C1(n52), .C2(n10), .A(n11), .ZN(
        ADD_WR[3]) );
  OAI221_X1 U92 ( .B1(n37), .B2(n30), .C1(n51), .C2(n10), .A(n11), .ZN(
        ADD_WR[4]) );
  NOR3_X1 U93 ( .A1(n14), .A2(n6), .A3(n37), .ZN(ADD_RS2[4]) );
  AOI21_X1 U94 ( .B1(n16), .B2(n13), .A(n39), .ZN(ADD_RS1[1]) );
  NOR2_X1 U95 ( .A1(n45), .A2(n44), .ZN(ADD_RS1[4]) );
  INV_X1 U96 ( .A(INST_IN[27]), .ZN(n50) );
endmodule


module regn_N32_7 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U6 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U7 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U8 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U9 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U10 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U11 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U12 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U13 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U14 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U15 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U16 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U17 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U18 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U19 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U20 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U21 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U22 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U23 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U24 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U25 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U26 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U27 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U28 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U29 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U30 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U31 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U32 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U33 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U34 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U35 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U36 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U37 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U38 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U39 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U40 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U41 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U42 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U43 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U44 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U45 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U46 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U47 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U48 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U49 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U50 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U51 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U52 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U53 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U54 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U55 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U56 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U57 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U58 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U59 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U60 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U61 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U62 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
  OAI21_X1 U63 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U64 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U65 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U66 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U67 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U68 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
endmodule


module regn_N32_6 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U6 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U7 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U8 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U9 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U10 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U11 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U12 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U13 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U14 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U15 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U16 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U17 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U18 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U19 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U20 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U21 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U22 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U23 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U24 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U25 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U26 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U27 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U28 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U29 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U30 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U31 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U32 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U33 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U34 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U35 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U36 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
  OAI21_X1 U37 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U38 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U39 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U40 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U41 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U42 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U43 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U44 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U45 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U46 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U47 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U48 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U49 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U50 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U51 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U52 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U53 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U54 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U55 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U56 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U57 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U58 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U59 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U60 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U61 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U62 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U63 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U64 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U65 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U66 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U67 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U68 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
endmodule


module regn_N5_0 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  DFFR_X1 \DOUT_reg[4]  ( .D(n15), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n10)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n14), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n9) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n13), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n8) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n12), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n7) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n11), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n6) );
  OAI21_X1 U2 ( .B1(n7), .B2(EN), .A(n2), .ZN(n12) );
  NAND2_X1 U3 ( .A1(DIN[1]), .A2(EN), .ZN(n2) );
  OAI21_X1 U4 ( .B1(n8), .B2(EN), .A(n3), .ZN(n13) );
  NAND2_X1 U5 ( .A1(DIN[2]), .A2(EN), .ZN(n3) );
  OAI21_X1 U6 ( .B1(n9), .B2(EN), .A(n4), .ZN(n14) );
  NAND2_X1 U7 ( .A1(DIN[3]), .A2(EN), .ZN(n4) );
  OAI21_X1 U8 ( .B1(n10), .B2(EN), .A(n5), .ZN(n15) );
  NAND2_X1 U9 ( .A1(DIN[4]), .A2(EN), .ZN(n5) );
  OAI21_X1 U10 ( .B1(n6), .B2(EN), .A(n1), .ZN(n11) );
  NAND2_X1 U11 ( .A1(EN), .A2(DIN[0]), .ZN(n1) );
endmodule


module regn_N5_4 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 \DOUT_reg[4]  ( .D(n16), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n21)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n17), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n22)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n18), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n23)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n19), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n24)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n20), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n25)
         );
  OAI21_X1 U2 ( .B1(n24), .B2(EN), .A(n29), .ZN(n19) );
  NAND2_X1 U3 ( .A1(DIN[1]), .A2(EN), .ZN(n29) );
  OAI21_X1 U4 ( .B1(n23), .B2(EN), .A(n28), .ZN(n18) );
  NAND2_X1 U5 ( .A1(DIN[2]), .A2(EN), .ZN(n28) );
  OAI21_X1 U6 ( .B1(n21), .B2(EN), .A(n26), .ZN(n16) );
  NAND2_X1 U7 ( .A1(DIN[4]), .A2(EN), .ZN(n26) );
  OAI21_X1 U8 ( .B1(n25), .B2(EN), .A(n30), .ZN(n20) );
  NAND2_X1 U9 ( .A1(EN), .A2(DIN[0]), .ZN(n30) );
  OAI21_X1 U10 ( .B1(n22), .B2(EN), .A(n27), .ZN(n17) );
  NAND2_X1 U11 ( .A1(DIN[3]), .A2(EN), .ZN(n27) );
endmodule


module regn_N5_3 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 \DOUT_reg[4]  ( .D(n16), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n21)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n17), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n22)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n18), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n23)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n19), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n24)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n20), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n25)
         );
  OAI21_X1 U2 ( .B1(n22), .B2(EN), .A(n27), .ZN(n17) );
  NAND2_X1 U3 ( .A1(DIN[3]), .A2(EN), .ZN(n27) );
  OAI21_X1 U4 ( .B1(n21), .B2(EN), .A(n26), .ZN(n16) );
  NAND2_X1 U5 ( .A1(DIN[4]), .A2(EN), .ZN(n26) );
  OAI21_X1 U6 ( .B1(n24), .B2(EN), .A(n29), .ZN(n19) );
  NAND2_X1 U7 ( .A1(DIN[1]), .A2(EN), .ZN(n29) );
  OAI21_X1 U8 ( .B1(n23), .B2(EN), .A(n28), .ZN(n18) );
  NAND2_X1 U9 ( .A1(DIN[2]), .A2(EN), .ZN(n28) );
  OAI21_X1 U10 ( .B1(n25), .B2(EN), .A(n30), .ZN(n20) );
  NAND2_X1 U11 ( .A1(EN), .A2(DIN[0]), .ZN(n30) );
endmodule


module mux21_NBIT5_0 ( A, B, S, Z );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Z;
  input S;
  wire   n7, n8, n9, n10, n11, n1, n2;

  BUF_X1 U1 ( .A(S), .Z(n1) );
  INV_X1 U2 ( .A(n10), .ZN(Z[1]) );
  AOI22_X1 U3 ( .A1(A[1]), .A2(n2), .B1(B[1]), .B2(n1), .ZN(n10) );
  INV_X1 U4 ( .A(n9), .ZN(Z[2]) );
  INV_X1 U5 ( .A(n7), .ZN(Z[4]) );
  INV_X1 U6 ( .A(n11), .ZN(Z[0]) );
  INV_X1 U7 ( .A(n8), .ZN(Z[3]) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(n2), .B1(B[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U9 ( .A1(A[2]), .A2(n2), .B1(B[2]), .B2(n1), .ZN(n9) );
  AOI22_X1 U10 ( .A1(A[4]), .A2(n2), .B1(S), .B2(B[4]), .ZN(n7) );
  AOI22_X1 U11 ( .A1(A[0]), .A2(n2), .B1(B[0]), .B2(n1), .ZN(n11) );
  INV_X1 U12 ( .A(S), .ZN(n2) );
endmodule


module mux21_NBIT5_2 ( A, B, S, Z );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Z;
  input S;
  wire   n1, n2, n3, n14, n15, n16, n17, n18;

  BUF_X1 U1 ( .A(S), .Z(n1) );
  BUF_X1 U2 ( .A(S), .Z(n2) );
  INV_X1 U3 ( .A(n17), .ZN(Z[3]) );
  INV_X1 U4 ( .A(n18), .ZN(Z[4]) );
  INV_X1 U5 ( .A(n15), .ZN(Z[1]) );
  INV_X1 U6 ( .A(n16), .ZN(Z[2]) );
  INV_X1 U7 ( .A(n14), .ZN(Z[0]) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(n3), .B1(B[3]), .B2(n1), .ZN(n17) );
  AOI22_X1 U9 ( .A1(A[4]), .A2(n3), .B1(n2), .B2(B[4]), .ZN(n18) );
  AOI22_X1 U10 ( .A1(A[1]), .A2(n3), .B1(B[1]), .B2(n1), .ZN(n15) );
  AOI22_X1 U11 ( .A1(A[0]), .A2(n3), .B1(B[0]), .B2(n1), .ZN(n14) );
  AOI22_X1 U12 ( .A1(A[2]), .A2(n3), .B1(B[2]), .B2(n1), .ZN(n16) );
  INV_X1 U13 ( .A(n2), .ZN(n3) );
endmodule


module mux21_NBIT5_1 ( A, B, S, Z );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Z;
  input S;
  wire   n1, n2, n3, n14, n15, n16, n17, n18;

  BUF_X1 U1 ( .A(S), .Z(n1) );
  BUF_X1 U2 ( .A(S), .Z(n2) );
  INV_X1 U3 ( .A(n15), .ZN(Z[1]) );
  AOI22_X1 U4 ( .A1(A[1]), .A2(n3), .B1(B[1]), .B2(n1), .ZN(n15) );
  INV_X1 U5 ( .A(n16), .ZN(Z[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n3), .B1(B[2]), .B2(n1), .ZN(n16) );
  INV_X1 U7 ( .A(n17), .ZN(Z[3]) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(n3), .B1(B[3]), .B2(n1), .ZN(n17) );
  INV_X1 U9 ( .A(n18), .ZN(Z[4]) );
  AOI22_X1 U10 ( .A1(A[4]), .A2(n3), .B1(n2), .B2(B[4]), .ZN(n18) );
  INV_X1 U11 ( .A(n14), .ZN(Z[0]) );
  AOI22_X1 U12 ( .A1(A[0]), .A2(n3), .B1(B[0]), .B2(n1), .ZN(n14) );
  INV_X1 U13 ( .A(n2), .ZN(n3) );
endmodule


module register_file_NBIT_ADD5_NBIT_DATA32 ( CLK, RST, ENABLE, RD1, RD2, WR, 
        ADD_WR, ADD_RS1, ADD_RS2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RST, ENABLE, RD1, RD2, WR;
  wire   n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235;

  DFFR_X1 \REGISTERS_reg[2][31]  ( .D(n3529), .CK(CLK), .RN(n1458), .Q(n5235)
         );
  DFFR_X1 \REGISTERS_reg[2][30]  ( .D(n3528), .CK(CLK), .RN(n1458), .Q(n5234)
         );
  DFFR_X1 \REGISTERS_reg[2][29]  ( .D(n3527), .CK(CLK), .RN(n1458), .Q(n5233)
         );
  DFFR_X1 \REGISTERS_reg[2][28]  ( .D(n3526), .CK(CLK), .RN(n1458), .Q(n5232)
         );
  DFFR_X1 \REGISTERS_reg[2][27]  ( .D(n3525), .CK(CLK), .RN(n1459), .Q(n5231)
         );
  DFFR_X1 \REGISTERS_reg[2][26]  ( .D(n3524), .CK(CLK), .RN(n1459), .Q(n5230)
         );
  DFFR_X1 \REGISTERS_reg[2][25]  ( .D(n3523), .CK(CLK), .RN(n1459), .Q(n5229)
         );
  DFFR_X1 \REGISTERS_reg[2][24]  ( .D(n3522), .CK(CLK), .RN(n1459), .Q(n5228)
         );
  DFFR_X1 \REGISTERS_reg[2][23]  ( .D(n3521), .CK(CLK), .RN(n1459), .Q(n5227)
         );
  DFFR_X1 \REGISTERS_reg[2][22]  ( .D(n3520), .CK(CLK), .RN(n1459), .Q(n5226)
         );
  DFFR_X1 \REGISTERS_reg[2][21]  ( .D(n3519), .CK(CLK), .RN(n1459), .Q(n5225)
         );
  DFFR_X1 \REGISTERS_reg[2][20]  ( .D(n3518), .CK(CLK), .RN(n1459), .Q(n5224)
         );
  DFFR_X1 \REGISTERS_reg[2][19]  ( .D(n3517), .CK(CLK), .RN(n1459), .Q(n5223)
         );
  DFFR_X1 \REGISTERS_reg[2][18]  ( .D(n3516), .CK(CLK), .RN(n1459), .Q(n5222)
         );
  DFFR_X1 \REGISTERS_reg[2][17]  ( .D(n3515), .CK(CLK), .RN(n1459), .Q(n5221)
         );
  DFFR_X1 \REGISTERS_reg[2][16]  ( .D(n3514), .CK(CLK), .RN(n1459), .Q(n5220)
         );
  DFFR_X1 \REGISTERS_reg[2][15]  ( .D(n3513), .CK(CLK), .RN(n1460), .Q(n5219)
         );
  DFFR_X1 \REGISTERS_reg[2][14]  ( .D(n3512), .CK(CLK), .RN(n1460), .Q(n5218)
         );
  DFFR_X1 \REGISTERS_reg[2][13]  ( .D(n3511), .CK(CLK), .RN(n1460), .Q(n5217)
         );
  DFFR_X1 \REGISTERS_reg[2][12]  ( .D(n3510), .CK(CLK), .RN(n1460), .Q(n5216)
         );
  DFFR_X1 \REGISTERS_reg[2][11]  ( .D(n3509), .CK(CLK), .RN(n1460), .Q(n5215)
         );
  DFFR_X1 \REGISTERS_reg[2][10]  ( .D(n3508), .CK(CLK), .RN(n1460), .Q(n5214)
         );
  DFFR_X1 \REGISTERS_reg[2][9]  ( .D(n3507), .CK(CLK), .RN(n1460), .Q(n5213)
         );
  DFFR_X1 \REGISTERS_reg[2][8]  ( .D(n3506), .CK(CLK), .RN(n1460), .Q(n5212)
         );
  DFFR_X1 \REGISTERS_reg[2][7]  ( .D(n3505), .CK(CLK), .RN(n1460), .Q(n5211)
         );
  DFFR_X1 \REGISTERS_reg[2][6]  ( .D(n3504), .CK(CLK), .RN(n1460), .Q(n5210)
         );
  DFFR_X1 \REGISTERS_reg[2][5]  ( .D(n3503), .CK(CLK), .RN(n1460), .Q(n5209)
         );
  DFFR_X1 \REGISTERS_reg[2][4]  ( .D(n3502), .CK(CLK), .RN(n1460), .Q(n5208)
         );
  DFFR_X1 \REGISTERS_reg[2][3]  ( .D(n3501), .CK(CLK), .RN(n1461), .Q(n5207)
         );
  DFFR_X1 \REGISTERS_reg[2][2]  ( .D(n3500), .CK(CLK), .RN(n1461), .Q(n5206)
         );
  DFFR_X1 \REGISTERS_reg[2][1]  ( .D(n3499), .CK(CLK), .RN(n1461), .Q(n5205)
         );
  DFFR_X1 \REGISTERS_reg[2][0]  ( .D(n3498), .CK(CLK), .RN(n1461), .Q(n5204)
         );
  DFFR_X1 \REGISTERS_reg[3][31]  ( .D(n3497), .CK(CLK), .RN(n1461), .Q(n5203), 
        .QN(n2201) );
  DFFR_X1 \REGISTERS_reg[3][30]  ( .D(n3496), .CK(CLK), .RN(n1461), .Q(n5202), 
        .QN(n2179) );
  DFFR_X1 \REGISTERS_reg[3][29]  ( .D(n3495), .CK(CLK), .RN(n1461), .Q(n5201), 
        .QN(n2158) );
  DFFR_X1 \REGISTERS_reg[3][28]  ( .D(n3494), .CK(CLK), .RN(n1461), .Q(n5200), 
        .QN(n2137) );
  DFFR_X1 \REGISTERS_reg[3][27]  ( .D(n3493), .CK(CLK), .RN(n1461), .Q(n5199), 
        .QN(n2116) );
  DFFR_X1 \REGISTERS_reg[3][26]  ( .D(n3492), .CK(CLK), .RN(n1461), .Q(n5198), 
        .QN(n2095) );
  DFFR_X1 \REGISTERS_reg[3][25]  ( .D(n3491), .CK(CLK), .RN(n1461), .Q(n5197), 
        .QN(n2074) );
  DFFR_X1 \REGISTERS_reg[3][24]  ( .D(n3490), .CK(CLK), .RN(n1461), .Q(n5196), 
        .QN(n2053) );
  DFFR_X1 \REGISTERS_reg[3][23]  ( .D(n3489), .CK(CLK), .RN(n1462), .Q(n5195), 
        .QN(n2032) );
  DFFR_X1 \REGISTERS_reg[3][22]  ( .D(n3488), .CK(CLK), .RN(n1462), .Q(n5194), 
        .QN(n2011) );
  DFFR_X1 \REGISTERS_reg[3][21]  ( .D(n3487), .CK(CLK), .RN(n1462), .Q(n5193), 
        .QN(n1991) );
  DFFR_X1 \REGISTERS_reg[3][20]  ( .D(n3486), .CK(CLK), .RN(n1462), .Q(n5192), 
        .QN(n1970) );
  DFFR_X1 \REGISTERS_reg[3][19]  ( .D(n3485), .CK(CLK), .RN(n1462), .Q(n5191), 
        .QN(n1950) );
  DFFR_X1 \REGISTERS_reg[3][18]  ( .D(n3484), .CK(CLK), .RN(n1462), .Q(n5190), 
        .QN(n1930) );
  DFFR_X1 \REGISTERS_reg[3][17]  ( .D(n3483), .CK(CLK), .RN(n1462), .Q(n5189), 
        .QN(n1910) );
  DFFR_X1 \REGISTERS_reg[3][16]  ( .D(n3482), .CK(CLK), .RN(n1462), .Q(n5188), 
        .QN(n1889) );
  DFFR_X1 \REGISTERS_reg[3][15]  ( .D(n3481), .CK(CLK), .RN(n1462), .Q(n5187), 
        .QN(n1870) );
  DFFR_X1 \REGISTERS_reg[3][14]  ( .D(n3480), .CK(CLK), .RN(n1462), .Q(n5186), 
        .QN(n1849) );
  DFFR_X1 \REGISTERS_reg[3][13]  ( .D(n3479), .CK(CLK), .RN(n1462), .Q(n5185), 
        .QN(n1828) );
  DFFR_X1 \REGISTERS_reg[3][12]  ( .D(n3478), .CK(CLK), .RN(n1462), .Q(n5184), 
        .QN(n1808) );
  DFFR_X1 \REGISTERS_reg[3][11]  ( .D(n3477), .CK(CLK), .RN(n1463), .Q(n5183), 
        .QN(n1787) );
  DFFR_X1 \REGISTERS_reg[3][10]  ( .D(n3476), .CK(CLK), .RN(n1463), .Q(n5182), 
        .QN(n1766) );
  DFFR_X1 \REGISTERS_reg[3][9]  ( .D(n3475), .CK(CLK), .RN(n1463), .Q(n5181), 
        .QN(n1745) );
  DFFR_X1 \REGISTERS_reg[3][8]  ( .D(n3474), .CK(CLK), .RN(n1463), .Q(n5180), 
        .QN(n1724) );
  DFFR_X1 \REGISTERS_reg[3][7]  ( .D(n3473), .CK(CLK), .RN(n1463), .Q(n5179), 
        .QN(n1703) );
  DFFR_X1 \REGISTERS_reg[3][6]  ( .D(n3472), .CK(CLK), .RN(n1463), .Q(n5178), 
        .QN(n1682) );
  DFFR_X1 \REGISTERS_reg[3][5]  ( .D(n3471), .CK(CLK), .RN(n1463), .Q(n5177), 
        .QN(n1661) );
  DFFR_X1 \REGISTERS_reg[3][4]  ( .D(n3470), .CK(CLK), .RN(n1463), .Q(n5176), 
        .QN(n1640) );
  DFFR_X1 \REGISTERS_reg[3][3]  ( .D(n3469), .CK(CLK), .RN(n1463), .Q(n5175), 
        .QN(n1620) );
  DFFR_X1 \REGISTERS_reg[3][2]  ( .D(n3468), .CK(CLK), .RN(n1463), .Q(n5174), 
        .QN(n1601) );
  DFFR_X1 \REGISTERS_reg[3][1]  ( .D(n3467), .CK(CLK), .RN(n1463), .Q(n5173), 
        .QN(n1581) );
  DFFR_X1 \REGISTERS_reg[3][0]  ( .D(n3466), .CK(CLK), .RN(n1463), .Q(n5172), 
        .QN(n1556) );
  DFFR_X1 \REGISTERS_reg[6][31]  ( .D(n3401), .CK(CLK), .RN(n1469), .Q(n5171), 
        .QN(n2215) );
  DFFR_X1 \REGISTERS_reg[6][30]  ( .D(n3400), .CK(CLK), .RN(n1469), .Q(n5170), 
        .QN(n2185) );
  DFFR_X1 \REGISTERS_reg[6][29]  ( .D(n3399), .CK(CLK), .RN(n1469), .Q(n5169), 
        .QN(n2164) );
  DFFR_X1 \REGISTERS_reg[6][28]  ( .D(n3398), .CK(CLK), .RN(n1469), .Q(n5168), 
        .QN(n2143) );
  DFFR_X1 \REGISTERS_reg[6][27]  ( .D(n3397), .CK(CLK), .RN(n1469), .Q(n5167), 
        .QN(n2122) );
  DFFR_X1 \REGISTERS_reg[6][26]  ( .D(n3396), .CK(CLK), .RN(n1469), .Q(n5166), 
        .QN(n2101) );
  DFFR_X1 \REGISTERS_reg[6][25]  ( .D(n3395), .CK(CLK), .RN(n1469), .Q(n5165), 
        .QN(n2080) );
  DFFR_X1 \REGISTERS_reg[6][24]  ( .D(n3394), .CK(CLK), .RN(n1469), .Q(n5164), 
        .QN(n2059) );
  DFFR_X1 \REGISTERS_reg[6][23]  ( .D(n3393), .CK(CLK), .RN(n1470), .Q(n5163), 
        .QN(n2038) );
  DFFR_X1 \REGISTERS_reg[6][22]  ( .D(n3392), .CK(CLK), .RN(n1470), .Q(n5162), 
        .QN(n2017) );
  DFFR_X1 \REGISTERS_reg[6][21]  ( .D(n3391), .CK(CLK), .RN(n1470), .Q(n5161), 
        .QN(n1997) );
  DFFR_X1 \REGISTERS_reg[6][20]  ( .D(n3390), .CK(CLK), .RN(n1470), .Q(n5160), 
        .QN(n1976) );
  DFFR_X1 \REGISTERS_reg[6][19]  ( .D(n3389), .CK(CLK), .RN(n1470), .Q(n5159), 
        .QN(n1956) );
  DFFR_X1 \REGISTERS_reg[6][18]  ( .D(n3388), .CK(CLK), .RN(n1470), .Q(n5158), 
        .QN(n1936) );
  DFFR_X1 \REGISTERS_reg[6][17]  ( .D(n3387), .CK(CLK), .RN(n1470), .Q(n5157), 
        .QN(n1916) );
  DFFR_X1 \REGISTERS_reg[6][16]  ( .D(n3386), .CK(CLK), .RN(n1470), .Q(n5156), 
        .QN(n1895) );
  DFFR_X1 \REGISTERS_reg[6][15]  ( .D(n3385), .CK(CLK), .RN(n1470), .Q(n5155), 
        .QN(n1874) );
  DFFR_X1 \REGISTERS_reg[6][14]  ( .D(n3384), .CK(CLK), .RN(n1470), .Q(n5154), 
        .QN(n1855) );
  DFFR_X1 \REGISTERS_reg[6][13]  ( .D(n3383), .CK(CLK), .RN(n1470), .Q(n5153), 
        .QN(n1834) );
  DFFR_X1 \REGISTERS_reg[6][12]  ( .D(n3382), .CK(CLK), .RN(n1470), .Q(n5152), 
        .QN(n1814) );
  DFFR_X1 \REGISTERS_reg[6][11]  ( .D(n3381), .CK(CLK), .RN(n1471), .Q(n5151), 
        .QN(n1793) );
  DFFR_X1 \REGISTERS_reg[6][10]  ( .D(n3380), .CK(CLK), .RN(n1471), .Q(n5150), 
        .QN(n1772) );
  DFFR_X1 \REGISTERS_reg[6][9]  ( .D(n3379), .CK(CLK), .RN(n1471), .Q(n5149), 
        .QN(n1751) );
  DFFR_X1 \REGISTERS_reg[6][8]  ( .D(n3378), .CK(CLK), .RN(n1471), .Q(n5148), 
        .QN(n1730) );
  DFFR_X1 \REGISTERS_reg[6][7]  ( .D(n3377), .CK(CLK), .RN(n1471), .Q(n5147), 
        .QN(n1709) );
  DFFR_X1 \REGISTERS_reg[6][6]  ( .D(n3376), .CK(CLK), .RN(n1471), .Q(n5146), 
        .QN(n1688) );
  DFFR_X1 \REGISTERS_reg[6][5]  ( .D(n3375), .CK(CLK), .RN(n1471), .Q(n5145), 
        .QN(n1667) );
  DFFR_X1 \REGISTERS_reg[6][4]  ( .D(n3374), .CK(CLK), .RN(n1471), .Q(n5144), 
        .QN(n1646) );
  DFFR_X1 \REGISTERS_reg[6][3]  ( .D(n3373), .CK(CLK), .RN(n1471), .Q(n5143), 
        .QN(n1626) );
  DFFR_X1 \REGISTERS_reg[6][2]  ( .D(n3372), .CK(CLK), .RN(n1471), .Q(n5142), 
        .QN(n1605) );
  DFFR_X1 \REGISTERS_reg[6][1]  ( .D(n3371), .CK(CLK), .RN(n1471), .Q(n5141), 
        .QN(n1587) );
  DFFR_X1 \REGISTERS_reg[6][0]  ( .D(n3370), .CK(CLK), .RN(n1471), .Q(n5140), 
        .QN(n1564) );
  DFFR_X1 \REGISTERS_reg[7][31]  ( .D(n3369), .CK(CLK), .RN(n1472), .Q(n5139)
         );
  DFFR_X1 \REGISTERS_reg[7][30]  ( .D(n3368), .CK(CLK), .RN(n1472), .Q(n5138)
         );
  DFFR_X1 \REGISTERS_reg[7][29]  ( .D(n3367), .CK(CLK), .RN(n1472), .Q(n5137)
         );
  DFFR_X1 \REGISTERS_reg[7][28]  ( .D(n3366), .CK(CLK), .RN(n1472), .Q(n5136)
         );
  DFFR_X1 \REGISTERS_reg[7][27]  ( .D(n3365), .CK(CLK), .RN(n1472), .Q(n5135)
         );
  DFFR_X1 \REGISTERS_reg[7][26]  ( .D(n3364), .CK(CLK), .RN(n1472), .Q(n5134)
         );
  DFFR_X1 \REGISTERS_reg[7][25]  ( .D(n3363), .CK(CLK), .RN(n1472), .Q(n5133)
         );
  DFFR_X1 \REGISTERS_reg[7][24]  ( .D(n3362), .CK(CLK), .RN(n1472), .Q(n5132)
         );
  DFFR_X1 \REGISTERS_reg[7][23]  ( .D(n3361), .CK(CLK), .RN(n1472), .Q(n5131)
         );
  DFFR_X1 \REGISTERS_reg[7][22]  ( .D(n3360), .CK(CLK), .RN(n1472), .Q(n5130)
         );
  DFFR_X1 \REGISTERS_reg[7][21]  ( .D(n3359), .CK(CLK), .RN(n1472), .Q(n5129)
         );
  DFFR_X1 \REGISTERS_reg[7][20]  ( .D(n3358), .CK(CLK), .RN(n1472), .Q(n5128)
         );
  DFFR_X1 \REGISTERS_reg[7][19]  ( .D(n3357), .CK(CLK), .RN(n1473), .Q(n5127)
         );
  DFFR_X1 \REGISTERS_reg[7][18]  ( .D(n3356), .CK(CLK), .RN(n1473), .Q(n5126)
         );
  DFFR_X1 \REGISTERS_reg[7][17]  ( .D(n3355), .CK(CLK), .RN(n1473), .Q(n5125)
         );
  DFFR_X1 \REGISTERS_reg[7][16]  ( .D(n3354), .CK(CLK), .RN(n1473), .Q(n5124)
         );
  DFFR_X1 \REGISTERS_reg[7][15]  ( .D(n3353), .CK(CLK), .RN(n1473), .Q(n5123)
         );
  DFFR_X1 \REGISTERS_reg[7][14]  ( .D(n3352), .CK(CLK), .RN(n1473), .Q(n5122)
         );
  DFFR_X1 \REGISTERS_reg[7][13]  ( .D(n3351), .CK(CLK), .RN(n1473), .Q(n5121)
         );
  DFFR_X1 \REGISTERS_reg[7][12]  ( .D(n3350), .CK(CLK), .RN(n1473), .Q(n5120)
         );
  DFFR_X1 \REGISTERS_reg[7][11]  ( .D(n3349), .CK(CLK), .RN(n1473), .Q(n5119)
         );
  DFFR_X1 \REGISTERS_reg[7][10]  ( .D(n3348), .CK(CLK), .RN(n1473), .Q(n5118)
         );
  DFFR_X1 \REGISTERS_reg[7][9]  ( .D(n3347), .CK(CLK), .RN(n1473), .Q(n5117)
         );
  DFFR_X1 \REGISTERS_reg[7][8]  ( .D(n3346), .CK(CLK), .RN(n1473), .Q(n5116)
         );
  DFFR_X1 \REGISTERS_reg[7][7]  ( .D(n3345), .CK(CLK), .RN(n1474), .Q(n5115)
         );
  DFFR_X1 \REGISTERS_reg[7][6]  ( .D(n3344), .CK(CLK), .RN(n1474), .Q(n5114)
         );
  DFFR_X1 \REGISTERS_reg[7][5]  ( .D(n3343), .CK(CLK), .RN(n1474), .Q(n5113)
         );
  DFFR_X1 \REGISTERS_reg[7][4]  ( .D(n3342), .CK(CLK), .RN(n1474), .Q(n5112)
         );
  DFFR_X1 \REGISTERS_reg[7][3]  ( .D(n3341), .CK(CLK), .RN(n1474), .Q(n5111)
         );
  DFFR_X1 \REGISTERS_reg[7][2]  ( .D(n3340), .CK(CLK), .RN(n1474), .Q(n5110)
         );
  DFFR_X1 \REGISTERS_reg[7][1]  ( .D(n3339), .CK(CLK), .RN(n1474), .Q(n5109)
         );
  DFFR_X1 \REGISTERS_reg[7][0]  ( .D(n3338), .CK(CLK), .RN(n1474), .Q(n5108)
         );
  DFFR_X1 \REGISTERS_reg[8][23]  ( .D(n3329), .CK(CLK), .RN(n1475), .QN(n237)
         );
  DFFR_X1 \REGISTERS_reg[8][22]  ( .D(n3328), .CK(CLK), .RN(n1475), .QN(n238)
         );
  DFFR_X1 \REGISTERS_reg[8][20]  ( .D(n3326), .CK(CLK), .RN(n1475), .QN(n240)
         );
  DFFR_X1 \REGISTERS_reg[8][19]  ( .D(n3325), .CK(CLK), .RN(n1475), .QN(n241)
         );
  DFFR_X1 \REGISTERS_reg[8][18]  ( .D(n3324), .CK(CLK), .RN(n1475), .QN(n242)
         );
  DFFR_X1 \REGISTERS_reg[8][17]  ( .D(n3323), .CK(CLK), .RN(n1475), .QN(n243)
         );
  DFFR_X1 \REGISTERS_reg[8][16]  ( .D(n3322), .CK(CLK), .RN(n1475), .QN(n244)
         );
  DFFR_X1 \REGISTERS_reg[8][15]  ( .D(n3321), .CK(CLK), .RN(n1476), .QN(n245)
         );
  DFFR_X1 \REGISTERS_reg[8][14]  ( .D(n3320), .CK(CLK), .RN(n1476), .QN(n246)
         );
  DFFR_X1 \REGISTERS_reg[8][13]  ( .D(n3319), .CK(CLK), .RN(n1476), .QN(n247)
         );
  DFFR_X1 \REGISTERS_reg[8][12]  ( .D(n3318), .CK(CLK), .RN(n1476), .QN(n248)
         );
  DFFR_X1 \REGISTERS_reg[8][11]  ( .D(n3317), .CK(CLK), .RN(n1476), .QN(n249)
         );
  DFFR_X1 \REGISTERS_reg[8][10]  ( .D(n3316), .CK(CLK), .RN(n1476), .QN(n250)
         );
  DFFR_X1 \REGISTERS_reg[8][9]  ( .D(n3315), .CK(CLK), .RN(n1476), .QN(n251)
         );
  DFFR_X1 \REGISTERS_reg[8][8]  ( .D(n3314), .CK(CLK), .RN(n1476), .QN(n252)
         );
  DFFR_X1 \REGISTERS_reg[8][7]  ( .D(n3313), .CK(CLK), .RN(n1476), .QN(n253)
         );
  DFFR_X1 \REGISTERS_reg[8][5]  ( .D(n3311), .CK(CLK), .RN(n1476), .QN(n255)
         );
  DFFR_X1 \REGISTERS_reg[8][4]  ( .D(n3310), .CK(CLK), .RN(n1476), .QN(n256)
         );
  DFFR_X1 \REGISTERS_reg[8][3]  ( .D(n3309), .CK(CLK), .RN(n1477), .QN(n257)
         );
  DFFR_X1 \REGISTERS_reg[8][2]  ( .D(n3308), .CK(CLK), .RN(n1477), .QN(n258)
         );
  DFFR_X1 \REGISTERS_reg[8][1]  ( .D(n3307), .CK(CLK), .RN(n1477), .QN(n259)
         );
  DFFR_X1 \REGISTERS_reg[8][0]  ( .D(n3306), .CK(CLK), .RN(n1477), .QN(n260)
         );
  DFFR_X1 \REGISTERS_reg[9][23]  ( .D(n3297), .CK(CLK), .RN(n1478), .Q(n212), 
        .QN(n269) );
  DFFR_X1 \REGISTERS_reg[9][22]  ( .D(n3296), .CK(CLK), .RN(n1478), .Q(n211), 
        .QN(n270) );
  DFFR_X1 \REGISTERS_reg[9][21]  ( .D(n3295), .CK(CLK), .RN(n1478), .Q(n210), 
        .QN(n271) );
  DFFR_X1 \REGISTERS_reg[9][20]  ( .D(n3294), .CK(CLK), .RN(n1478), .Q(n209), 
        .QN(n272) );
  DFFR_X1 \REGISTERS_reg[9][19]  ( .D(n3293), .CK(CLK), .RN(n1478), .Q(n208), 
        .QN(n273) );
  DFFR_X1 \REGISTERS_reg[9][18]  ( .D(n3292), .CK(CLK), .RN(n1478), .Q(n207), 
        .QN(n274) );
  DFFR_X1 \REGISTERS_reg[9][17]  ( .D(n3291), .CK(CLK), .RN(n1478), .Q(n206), 
        .QN(n275) );
  DFFR_X1 \REGISTERS_reg[9][16]  ( .D(n3290), .CK(CLK), .RN(n1478), .Q(n205), 
        .QN(n276) );
  DFFR_X1 \REGISTERS_reg[9][15]  ( .D(n3289), .CK(CLK), .RN(n1478), .Q(n204), 
        .QN(n277) );
  DFFR_X1 \REGISTERS_reg[9][14]  ( .D(n3288), .CK(CLK), .RN(n1478), .Q(n217), 
        .QN(n278) );
  DFFR_X1 \REGISTERS_reg[9][13]  ( .D(n3287), .CK(CLK), .RN(n1478), .Q(n216), 
        .QN(n279) );
  DFFR_X1 \REGISTERS_reg[9][12]  ( .D(n3286), .CK(CLK), .RN(n1478), .Q(n215), 
        .QN(n280) );
  DFFR_X1 \REGISTERS_reg[9][11]  ( .D(n3285), .CK(CLK), .RN(n1479), .Q(n214), 
        .QN(n281) );
  DFFR_X1 \REGISTERS_reg[9][10]  ( .D(n3284), .CK(CLK), .RN(n1479), .Q(n203), 
        .QN(n282) );
  DFFR_X1 \REGISTERS_reg[9][9]  ( .D(n3283), .CK(CLK), .RN(n1479), .Q(n213), 
        .QN(n283) );
  DFFR_X1 \REGISTERS_reg[9][8]  ( .D(n3282), .CK(CLK), .RN(n1479), .Q(n202), 
        .QN(n284) );
  DFFR_X1 \REGISTERS_reg[9][7]  ( .D(n3281), .CK(CLK), .RN(n1479), .Q(n201), 
        .QN(n285) );
  DFFR_X1 \REGISTERS_reg[9][6]  ( .D(n3280), .CK(CLK), .RN(n1479), .Q(n200), 
        .QN(n286) );
  DFFR_X1 \REGISTERS_reg[9][5]  ( .D(n3279), .CK(CLK), .RN(n1479), .Q(n199), 
        .QN(n287) );
  DFFR_X1 \REGISTERS_reg[9][4]  ( .D(n3278), .CK(CLK), .RN(n1479), .Q(n198), 
        .QN(n288) );
  DFFR_X1 \REGISTERS_reg[9][3]  ( .D(n3277), .CK(CLK), .RN(n1479), .Q(n197), 
        .QN(n289) );
  DFFR_X1 \REGISTERS_reg[9][2]  ( .D(n3276), .CK(CLK), .RN(n1479), .Q(n196), 
        .QN(n290) );
  DFFR_X1 \REGISTERS_reg[9][1]  ( .D(n3275), .CK(CLK), .RN(n1479), .Q(n195), 
        .QN(n291) );
  DFFR_X1 \REGISTERS_reg[9][0]  ( .D(n3274), .CK(CLK), .RN(n1479), .Q(n194), 
        .QN(n292) );
  DFFR_X1 \REGISTERS_reg[10][31]  ( .D(n3273), .CK(CLK), .RN(n1480), .Q(n5107), 
        .QN(n193) );
  DFFR_X1 \REGISTERS_reg[10][30]  ( .D(n3272), .CK(CLK), .RN(n1480), .Q(n5106), 
        .QN(n192) );
  DFFR_X1 \REGISTERS_reg[10][29]  ( .D(n3271), .CK(CLK), .RN(n1480), .Q(n5105), 
        .QN(n191) );
  DFFR_X1 \REGISTERS_reg[10][28]  ( .D(n3270), .CK(CLK), .RN(n1480), .Q(n5104), 
        .QN(n190) );
  DFFR_X1 \REGISTERS_reg[10][27]  ( .D(n3269), .CK(CLK), .RN(n1480), .Q(n5103), 
        .QN(n189) );
  DFFR_X1 \REGISTERS_reg[10][26]  ( .D(n3268), .CK(CLK), .RN(n1480), .Q(n5102), 
        .QN(n188) );
  DFFR_X1 \REGISTERS_reg[10][25]  ( .D(n3267), .CK(CLK), .RN(n1480), .Q(n5101), 
        .QN(n187) );
  DFFR_X1 \REGISTERS_reg[10][24]  ( .D(n3266), .CK(CLK), .RN(n1480), .Q(n5100), 
        .QN(n186) );
  DFFR_X1 \REGISTERS_reg[10][23]  ( .D(n3265), .CK(CLK), .RN(n1480), .Q(n5099), 
        .QN(n185) );
  DFFR_X1 \REGISTERS_reg[10][22]  ( .D(n3264), .CK(CLK), .RN(n1480), .Q(n5098), 
        .QN(n441) );
  DFFR_X1 \REGISTERS_reg[10][21]  ( .D(n3263), .CK(CLK), .RN(n1480), .Q(n5097), 
        .QN(n443) );
  DFFR_X1 \REGISTERS_reg[10][20]  ( .D(n3262), .CK(CLK), .RN(n1480), .Q(n5096), 
        .QN(n453) );
  DFFR_X1 \REGISTERS_reg[10][19]  ( .D(n3261), .CK(CLK), .RN(n1481), .Q(n5095), 
        .QN(n455) );
  DFFR_X1 \REGISTERS_reg[10][18]  ( .D(n3260), .CK(CLK), .RN(n1481), .Q(n5094), 
        .QN(n184) );
  DFFR_X1 \REGISTERS_reg[10][17]  ( .D(n3259), .CK(CLK), .RN(n1481), .Q(n5093), 
        .QN(n445) );
  DFFR_X1 \REGISTERS_reg[10][16]  ( .D(n3258), .CK(CLK), .RN(n1481), .Q(n5092), 
        .QN(n447) );
  DFFR_X1 \REGISTERS_reg[10][15]  ( .D(n3257), .CK(CLK), .RN(n1481), .Q(n5091), 
        .QN(n183) );
  DFFR_X1 \REGISTERS_reg[10][14]  ( .D(n3256), .CK(CLK), .RN(n1481), .Q(n5090), 
        .QN(n182) );
  DFFR_X1 \REGISTERS_reg[10][13]  ( .D(n3255), .CK(CLK), .RN(n1481), .Q(n5089), 
        .QN(n457) );
  DFFR_X1 \REGISTERS_reg[10][12]  ( .D(n3254), .CK(CLK), .RN(n1481), .Q(n5088), 
        .QN(n181) );
  DFFR_X1 \REGISTERS_reg[10][11]  ( .D(n3253), .CK(CLK), .RN(n1481), .Q(n5087), 
        .QN(n459) );
  DFFR_X1 \REGISTERS_reg[10][10]  ( .D(n3252), .CK(CLK), .RN(n1481), .Q(n5086), 
        .QN(n180) );
  DFFR_X1 \REGISTERS_reg[10][9]  ( .D(n3251), .CK(CLK), .RN(n1481), .Q(n5085), 
        .QN(n179) );
  DFFR_X1 \REGISTERS_reg[10][8]  ( .D(n3250), .CK(CLK), .RN(n1481), .Q(n5084), 
        .QN(n178) );
  DFFR_X1 \REGISTERS_reg[10][7]  ( .D(n3249), .CK(CLK), .RN(n1482), .Q(n5083), 
        .QN(n177) );
  DFFR_X1 \REGISTERS_reg[10][6]  ( .D(n3248), .CK(CLK), .RN(n1482), .Q(n5082), 
        .QN(n176) );
  DFFR_X1 \REGISTERS_reg[10][5]  ( .D(n3247), .CK(CLK), .RN(n1482), .Q(n5081), 
        .QN(n175) );
  DFFR_X1 \REGISTERS_reg[10][4]  ( .D(n3246), .CK(CLK), .RN(n1482), .Q(n5080), 
        .QN(n449) );
  DFFR_X1 \REGISTERS_reg[10][3]  ( .D(n3245), .CK(CLK), .RN(n1482), .Q(n5079), 
        .QN(n174) );
  DFFR_X1 \REGISTERS_reg[10][2]  ( .D(n3244), .CK(CLK), .RN(n1482), .Q(n5078), 
        .QN(n173) );
  DFFR_X1 \REGISTERS_reg[10][1]  ( .D(n3243), .CK(CLK), .RN(n1482), .Q(n5077), 
        .QN(n439) );
  DFFR_X1 \REGISTERS_reg[10][0]  ( .D(n3242), .CK(CLK), .RN(n1482), .Q(n5076), 
        .QN(n451) );
  DFFR_X1 \REGISTERS_reg[11][31]  ( .D(n3241), .CK(CLK), .RN(n1482), .Q(n5075), 
        .QN(n342) );
  DFFR_X1 \REGISTERS_reg[11][30]  ( .D(n3240), .CK(CLK), .RN(n1482), .Q(n5074), 
        .QN(n341) );
  DFFR_X1 \REGISTERS_reg[11][29]  ( .D(n3239), .CK(CLK), .RN(n1482), .Q(n5073), 
        .QN(n340) );
  DFFR_X1 \REGISTERS_reg[11][28]  ( .D(n3238), .CK(CLK), .RN(n1482), .Q(n5072), 
        .QN(n339) );
  DFFR_X1 \REGISTERS_reg[11][27]  ( .D(n3237), .CK(CLK), .RN(n1483), .Q(n5071), 
        .QN(n338) );
  DFFR_X1 \REGISTERS_reg[11][26]  ( .D(n3236), .CK(CLK), .RN(n1483), .Q(n5070), 
        .QN(n337) );
  DFFR_X1 \REGISTERS_reg[11][25]  ( .D(n3235), .CK(CLK), .RN(n1483), .Q(n5069), 
        .QN(n336) );
  DFFR_X1 \REGISTERS_reg[11][24]  ( .D(n3234), .CK(CLK), .RN(n1483), .Q(n5068), 
        .QN(n335) );
  DFFR_X1 \REGISTERS_reg[11][23]  ( .D(n3233), .CK(CLK), .RN(n1483), .Q(n5067), 
        .QN(n334) );
  DFFR_X1 \REGISTERS_reg[11][22]  ( .D(n3232), .CK(CLK), .RN(n1483), .Q(n5066), 
        .QN(n442) );
  DFFR_X1 \REGISTERS_reg[11][21]  ( .D(n3231), .CK(CLK), .RN(n1483), .Q(n5065), 
        .QN(n444) );
  DFFR_X1 \REGISTERS_reg[11][20]  ( .D(n3230), .CK(CLK), .RN(n1483), .Q(n5064), 
        .QN(n454) );
  DFFR_X1 \REGISTERS_reg[11][19]  ( .D(n3229), .CK(CLK), .RN(n1483), .Q(n5063), 
        .QN(n456) );
  DFFR_X1 \REGISTERS_reg[11][18]  ( .D(n3228), .CK(CLK), .RN(n1483), .Q(n5062), 
        .QN(n333) );
  DFFR_X1 \REGISTERS_reg[11][17]  ( .D(n3227), .CK(CLK), .RN(n1483), .Q(n5061), 
        .QN(n446) );
  DFFR_X1 \REGISTERS_reg[11][16]  ( .D(n3226), .CK(CLK), .RN(n1483), .Q(n5060), 
        .QN(n448) );
  DFFR_X1 \REGISTERS_reg[11][15]  ( .D(n3225), .CK(CLK), .RN(n1484), .Q(n5059), 
        .QN(n332) );
  DFFR_X1 \REGISTERS_reg[11][14]  ( .D(n3224), .CK(CLK), .RN(n1484), .Q(n5058), 
        .QN(n331) );
  DFFR_X1 \REGISTERS_reg[11][13]  ( .D(n3223), .CK(CLK), .RN(n1484), .Q(n5057), 
        .QN(n458) );
  DFFR_X1 \REGISTERS_reg[11][12]  ( .D(n3222), .CK(CLK), .RN(n1484), .Q(n5056), 
        .QN(n330) );
  DFFR_X1 \REGISTERS_reg[11][11]  ( .D(n3221), .CK(CLK), .RN(n1484), .Q(n5055), 
        .QN(n460) );
  DFFR_X1 \REGISTERS_reg[11][10]  ( .D(n3220), .CK(CLK), .RN(n1484), .Q(n5054), 
        .QN(n329) );
  DFFR_X1 \REGISTERS_reg[11][9]  ( .D(n3219), .CK(CLK), .RN(n1484), .Q(n5053), 
        .QN(n328) );
  DFFR_X1 \REGISTERS_reg[11][8]  ( .D(n3218), .CK(CLK), .RN(n1484), .Q(n5052), 
        .QN(n327) );
  DFFR_X1 \REGISTERS_reg[11][7]  ( .D(n3217), .CK(CLK), .RN(n1484), .Q(n5051), 
        .QN(n326) );
  DFFR_X1 \REGISTERS_reg[11][6]  ( .D(n3216), .CK(CLK), .RN(n1484), .Q(n5050), 
        .QN(n325) );
  DFFR_X1 \REGISTERS_reg[11][5]  ( .D(n3215), .CK(CLK), .RN(n1484), .Q(n5049), 
        .QN(n324) );
  DFFR_X1 \REGISTERS_reg[11][4]  ( .D(n3214), .CK(CLK), .RN(n1484), .Q(n5048), 
        .QN(n450) );
  DFFR_X1 \REGISTERS_reg[11][3]  ( .D(n3213), .CK(CLK), .RN(n1485), .Q(n5047), 
        .QN(n323) );
  DFFR_X1 \REGISTERS_reg[11][2]  ( .D(n3212), .CK(CLK), .RN(n1485), .Q(n5046), 
        .QN(n322) );
  DFFR_X1 \REGISTERS_reg[11][1]  ( .D(n3211), .CK(CLK), .RN(n1485), .Q(n5045), 
        .QN(n440) );
  DFFR_X1 \REGISTERS_reg[11][0]  ( .D(n3210), .CK(CLK), .RN(n1485), .Q(n5044), 
        .QN(n452) );
  DFFR_X1 \REGISTERS_reg[12][23]  ( .D(n3201), .CK(CLK), .RN(n1486), .Q(n2036), 
        .QN(n365) );
  DFFR_X1 \REGISTERS_reg[12][22]  ( .D(n3200), .CK(CLK), .RN(n1486), .Q(n2015), 
        .QN(n366) );
  DFFR_X1 \REGISTERS_reg[12][21]  ( .D(n3199), .CK(CLK), .RN(n1486), .Q(n1995), 
        .QN(n367) );
  DFFR_X1 \REGISTERS_reg[12][20]  ( .D(n3198), .CK(CLK), .RN(n1486), .Q(n1974), 
        .QN(n368) );
  DFFR_X1 \REGISTERS_reg[12][19]  ( .D(n3197), .CK(CLK), .RN(n1486), .Q(n1954), 
        .QN(n369) );
  DFFR_X1 \REGISTERS_reg[12][18]  ( .D(n3196), .CK(CLK), .RN(n1486), .Q(n1934), 
        .QN(n370) );
  DFFR_X1 \REGISTERS_reg[12][17]  ( .D(n3195), .CK(CLK), .RN(n1486), .Q(n1914), 
        .QN(n371) );
  DFFR_X1 \REGISTERS_reg[12][16]  ( .D(n3194), .CK(CLK), .RN(n1486), .Q(n1893), 
        .QN(n372) );
  DFFR_X1 \REGISTERS_reg[12][15]  ( .D(n3193), .CK(CLK), .RN(n1486), .Q(n221), 
        .QN(n373) );
  DFFR_X1 \REGISTERS_reg[12][14]  ( .D(n3192), .CK(CLK), .RN(n1486), .Q(n1853), 
        .QN(n374) );
  DFFR_X1 \REGISTERS_reg[12][13]  ( .D(n3191), .CK(CLK), .RN(n1486), .Q(n1832), 
        .QN(n375) );
  DFFR_X1 \REGISTERS_reg[12][12]  ( .D(n3190), .CK(CLK), .RN(n1486), .Q(n1812), 
        .QN(n376) );
  DFFR_X1 \REGISTERS_reg[12][11]  ( .D(n3189), .CK(CLK), .RN(n1487), .Q(n1791), 
        .QN(n377) );
  DFFR_X1 \REGISTERS_reg[12][10]  ( .D(n3188), .CK(CLK), .RN(n1487), .Q(n1770), 
        .QN(n378) );
  DFFR_X1 \REGISTERS_reg[12][9]  ( .D(n3187), .CK(CLK), .RN(n1487), .Q(n1749), 
        .QN(n379) );
  DFFR_X1 \REGISTERS_reg[12][8]  ( .D(n3186), .CK(CLK), .RN(n1487), .Q(n1728), 
        .QN(n380) );
  DFFR_X1 \REGISTERS_reg[12][7]  ( .D(n3185), .CK(CLK), .RN(n1487), .Q(n1707), 
        .QN(n381) );
  DFFR_X1 \REGISTERS_reg[12][6]  ( .D(n3184), .CK(CLK), .RN(n1487), .Q(n1686), 
        .QN(n382) );
  DFFR_X1 \REGISTERS_reg[12][5]  ( .D(n3183), .CK(CLK), .RN(n1487), .Q(n1665), 
        .QN(n383) );
  DFFR_X1 \REGISTERS_reg[12][4]  ( .D(n3182), .CK(CLK), .RN(n1487), .Q(n1644), 
        .QN(n384) );
  DFFR_X1 \REGISTERS_reg[12][3]  ( .D(n3181), .CK(CLK), .RN(n1487), .Q(n1624), 
        .QN(n385) );
  DFFR_X1 \REGISTERS_reg[12][2]  ( .D(n3180), .CK(CLK), .RN(n1487), .Q(n219), 
        .QN(n386) );
  DFFR_X1 \REGISTERS_reg[12][1]  ( .D(n3179), .CK(CLK), .RN(n1487), .Q(n1585), 
        .QN(n387) );
  DFFR_X1 \REGISTERS_reg[12][0]  ( .D(n3178), .CK(CLK), .RN(n1487), .Q(n1562), 
        .QN(n388) );
  DFFR_X1 \REGISTERS_reg[13][23]  ( .D(n3169), .CK(CLK), .RN(n1488), .Q(n2034), 
        .QN(n397) );
  DFFR_X1 \REGISTERS_reg[13][22]  ( .D(n3168), .CK(CLK), .RN(n1488), .Q(n2013), 
        .QN(n398) );
  DFFR_X1 \REGISTERS_reg[13][21]  ( .D(n3167), .CK(CLK), .RN(n1488), .Q(n1993), 
        .QN(n399) );
  DFFR_X1 \REGISTERS_reg[13][20]  ( .D(n3166), .CK(CLK), .RN(n1488), .Q(n1972), 
        .QN(n400) );
  DFFR_X1 \REGISTERS_reg[13][19]  ( .D(n3165), .CK(CLK), .RN(n1489), .Q(n1952), 
        .QN(n401) );
  DFFR_X1 \REGISTERS_reg[13][18]  ( .D(n3164), .CK(CLK), .RN(n1489), .Q(n1932), 
        .QN(n402) );
  DFFR_X1 \REGISTERS_reg[13][17]  ( .D(n3163), .CK(CLK), .RN(n1489), .Q(n1912), 
        .QN(n403) );
  DFFR_X1 \REGISTERS_reg[13][16]  ( .D(n3162), .CK(CLK), .RN(n1489), .Q(n1891), 
        .QN(n404) );
  DFFR_X1 \REGISTERS_reg[13][15]  ( .D(n3161), .CK(CLK), .RN(n1489), .Q(n220), 
        .QN(n405) );
  DFFR_X1 \REGISTERS_reg[13][14]  ( .D(n3160), .CK(CLK), .RN(n1489), .Q(n1851), 
        .QN(n406) );
  DFFR_X1 \REGISTERS_reg[13][13]  ( .D(n3159), .CK(CLK), .RN(n1489), .Q(n1830), 
        .QN(n407) );
  DFFR_X1 \REGISTERS_reg[13][12]  ( .D(n3158), .CK(CLK), .RN(n1489), .Q(n1810), 
        .QN(n408) );
  DFFR_X1 \REGISTERS_reg[13][11]  ( .D(n3157), .CK(CLK), .RN(n1489), .Q(n1789), 
        .QN(n409) );
  DFFR_X1 \REGISTERS_reg[13][10]  ( .D(n3156), .CK(CLK), .RN(n1489), .Q(n1768), 
        .QN(n410) );
  DFFR_X1 \REGISTERS_reg[13][9]  ( .D(n3155), .CK(CLK), .RN(n1489), .Q(n1747), 
        .QN(n411) );
  DFFR_X1 \REGISTERS_reg[13][8]  ( .D(n3154), .CK(CLK), .RN(n1489), .Q(n1726), 
        .QN(n412) );
  DFFR_X1 \REGISTERS_reg[13][7]  ( .D(n3153), .CK(CLK), .RN(n1490), .Q(n1705), 
        .QN(n413) );
  DFFR_X1 \REGISTERS_reg[13][6]  ( .D(n3152), .CK(CLK), .RN(n1490), .Q(n1684), 
        .QN(n414) );
  DFFR_X1 \REGISTERS_reg[13][5]  ( .D(n3151), .CK(CLK), .RN(n1490), .Q(n1663), 
        .QN(n415) );
  DFFR_X1 \REGISTERS_reg[13][4]  ( .D(n3150), .CK(CLK), .RN(n1490), .Q(n1642), 
        .QN(n416) );
  DFFR_X1 \REGISTERS_reg[13][3]  ( .D(n3149), .CK(CLK), .RN(n1490), .Q(n1622), 
        .QN(n417) );
  DFFR_X1 \REGISTERS_reg[13][2]  ( .D(n3148), .CK(CLK), .RN(n1490), .Q(n218), 
        .QN(n418) );
  DFFR_X1 \REGISTERS_reg[13][1]  ( .D(n3147), .CK(CLK), .RN(n1490), .Q(n1583), 
        .QN(n419) );
  DFFR_X1 \REGISTERS_reg[13][0]  ( .D(n3146), .CK(CLK), .RN(n1490), .Q(n1558), 
        .QN(n420) );
  DFFR_X1 \REGISTERS_reg[14][31]  ( .D(n3145), .CK(CLK), .RN(n1490), .Q(n5043), 
        .QN(n4095) );
  DFFR_X1 \REGISTERS_reg[14][30]  ( .D(n3144), .CK(CLK), .RN(n1490), .Q(n5042), 
        .QN(n4064) );
  DFFR_X1 \REGISTERS_reg[14][29]  ( .D(n3143), .CK(CLK), .RN(n1490), .Q(n5041), 
        .QN(n4038) );
  DFFR_X1 \REGISTERS_reg[14][28]  ( .D(n3142), .CK(CLK), .RN(n1490), .Q(n5040), 
        .QN(n4012) );
  DFFR_X1 \REGISTERS_reg[14][27]  ( .D(n3141), .CK(CLK), .RN(n1491), .Q(n5039), 
        .QN(n3986) );
  DFFR_X1 \REGISTERS_reg[14][26]  ( .D(n3140), .CK(CLK), .RN(n1491), .Q(n5038), 
        .QN(n3960) );
  DFFR_X1 \REGISTERS_reg[14][25]  ( .D(n3139), .CK(CLK), .RN(n1491), .Q(n5037), 
        .QN(n3934) );
  DFFR_X1 \REGISTERS_reg[14][24]  ( .D(n3138), .CK(CLK), .RN(n1491), .Q(n5036), 
        .QN(n3908) );
  DFFR_X1 \REGISTERS_reg[14][23]  ( .D(n3137), .CK(CLK), .RN(n1491), .Q(n5035), 
        .QN(n3882) );
  DFFR_X1 \REGISTERS_reg[14][22]  ( .D(n3136), .CK(CLK), .RN(n1491), .Q(n5034), 
        .QN(n3857) );
  DFFR_X1 \REGISTERS_reg[14][21]  ( .D(n3135), .CK(CLK), .RN(n1491), .Q(n5033), 
        .QN(n3832) );
  DFFR_X1 \REGISTERS_reg[14][20]  ( .D(n3134), .CK(CLK), .RN(n1491), .Q(n5032), 
        .QN(n3807) );
  DFFR_X1 \REGISTERS_reg[14][19]  ( .D(n3133), .CK(CLK), .RN(n1491), .Q(n5031), 
        .QN(n3782) );
  DFFR_X1 \REGISTERS_reg[14][18]  ( .D(n3132), .CK(CLK), .RN(n1491), .Q(n5030), 
        .QN(n3757) );
  DFFR_X1 \REGISTERS_reg[14][17]  ( .D(n3131), .CK(CLK), .RN(n1491), .Q(n5029), 
        .QN(n3732) );
  DFFR_X1 \REGISTERS_reg[14][16]  ( .D(n3130), .CK(CLK), .RN(n1491), .Q(n5028), 
        .QN(n3707) );
  DFFR_X1 \REGISTERS_reg[14][15]  ( .D(n3129), .CK(CLK), .RN(n1492), .Q(n5027), 
        .QN(n3682) );
  DFFR_X1 \REGISTERS_reg[14][14]  ( .D(n3128), .CK(CLK), .RN(n1492), .Q(n5026), 
        .QN(n3657) );
  DFFR_X1 \REGISTERS_reg[14][13]  ( .D(n3127), .CK(CLK), .RN(n1492), .Q(n5025), 
        .QN(n3632) );
  DFFR_X1 \REGISTERS_reg[14][12]  ( .D(n3126), .CK(CLK), .RN(n1492), .Q(n5024), 
        .QN(n3607) );
  DFFR_X1 \REGISTERS_reg[14][11]  ( .D(n3125), .CK(CLK), .RN(n1492), .Q(n5023), 
        .QN(n3582) );
  DFFR_X1 \REGISTERS_reg[14][10]  ( .D(n3124), .CK(CLK), .RN(n1492), .Q(n5022), 
        .QN(n2501) );
  DFFR_X1 \REGISTERS_reg[14][9]  ( .D(n3123), .CK(CLK), .RN(n1492), .Q(n5021), 
        .QN(n2476) );
  DFFR_X1 \REGISTERS_reg[14][8]  ( .D(n3122), .CK(CLK), .RN(n1492), .Q(n5020), 
        .QN(n2451) );
  DFFR_X1 \REGISTERS_reg[14][7]  ( .D(n3121), .CK(CLK), .RN(n1492), .Q(n5019), 
        .QN(n2426) );
  DFFR_X1 \REGISTERS_reg[14][6]  ( .D(n3120), .CK(CLK), .RN(n1492), .Q(n5018), 
        .QN(n2401) );
  DFFR_X1 \REGISTERS_reg[14][5]  ( .D(n3119), .CK(CLK), .RN(n1492), .Q(n5017), 
        .QN(n2376) );
  DFFR_X1 \REGISTERS_reg[14][4]  ( .D(n3118), .CK(CLK), .RN(n1492), .Q(n5016), 
        .QN(n2351) );
  DFFR_X1 \REGISTERS_reg[14][3]  ( .D(n3117), .CK(CLK), .RN(n1493), .Q(n5015), 
        .QN(n2326) );
  DFFR_X1 \REGISTERS_reg[14][2]  ( .D(n3116), .CK(CLK), .RN(n1493), .Q(n5014), 
        .QN(n2301) );
  DFFR_X1 \REGISTERS_reg[14][1]  ( .D(n3115), .CK(CLK), .RN(n1493), .Q(n5013), 
        .QN(n2276) );
  DFFR_X1 \REGISTERS_reg[14][0]  ( .D(n3114), .CK(CLK), .RN(n1493), .Q(n5012), 
        .QN(n2247) );
  DFFR_X1 \REGISTERS_reg[15][31]  ( .D(n3113), .CK(CLK), .RN(n1493), .Q(n5011), 
        .QN(n4093) );
  DFFR_X1 \REGISTERS_reg[15][30]  ( .D(n3112), .CK(CLK), .RN(n1493), .Q(n5010), 
        .QN(n4063) );
  DFFR_X1 \REGISTERS_reg[15][29]  ( .D(n3111), .CK(CLK), .RN(n1493), .Q(n5009), 
        .QN(n4037) );
  DFFR_X1 \REGISTERS_reg[15][28]  ( .D(n3110), .CK(CLK), .RN(n1493), .Q(n5008), 
        .QN(n4011) );
  DFFR_X1 \REGISTERS_reg[15][27]  ( .D(n3109), .CK(CLK), .RN(n1493), .Q(n5007), 
        .QN(n3985) );
  DFFR_X1 \REGISTERS_reg[15][26]  ( .D(n3108), .CK(CLK), .RN(n1493), .Q(n5006), 
        .QN(n3959) );
  DFFR_X1 \REGISTERS_reg[15][25]  ( .D(n3107), .CK(CLK), .RN(n1493), .Q(n5005), 
        .QN(n3933) );
  DFFR_X1 \REGISTERS_reg[15][24]  ( .D(n3106), .CK(CLK), .RN(n1493), .Q(n5004), 
        .QN(n3907) );
  DFFR_X1 \REGISTERS_reg[15][23]  ( .D(n3105), .CK(CLK), .RN(n1494), .Q(n5003), 
        .QN(n3881) );
  DFFR_X1 \REGISTERS_reg[15][22]  ( .D(n3104), .CK(CLK), .RN(n1494), .Q(n5002), 
        .QN(n3856) );
  DFFR_X1 \REGISTERS_reg[15][21]  ( .D(n3103), .CK(CLK), .RN(n1494), .Q(n5001), 
        .QN(n3831) );
  DFFR_X1 \REGISTERS_reg[15][20]  ( .D(n3102), .CK(CLK), .RN(n1494), .Q(n5000), 
        .QN(n3806) );
  DFFR_X1 \REGISTERS_reg[15][19]  ( .D(n3101), .CK(CLK), .RN(n1494), .Q(n4999), 
        .QN(n3781) );
  DFFR_X1 \REGISTERS_reg[15][18]  ( .D(n3100), .CK(CLK), .RN(n1494), .Q(n4998), 
        .QN(n3756) );
  DFFR_X1 \REGISTERS_reg[15][17]  ( .D(n3099), .CK(CLK), .RN(n1494), .Q(n4997), 
        .QN(n3731) );
  DFFR_X1 \REGISTERS_reg[15][16]  ( .D(n3098), .CK(CLK), .RN(n1494), .Q(n4996), 
        .QN(n3706) );
  DFFR_X1 \REGISTERS_reg[15][15]  ( .D(n3097), .CK(CLK), .RN(n1494), .Q(n4995), 
        .QN(n3681) );
  DFFR_X1 \REGISTERS_reg[15][14]  ( .D(n3096), .CK(CLK), .RN(n1494), .Q(n4994), 
        .QN(n3656) );
  DFFR_X1 \REGISTERS_reg[15][13]  ( .D(n3095), .CK(CLK), .RN(n1494), .Q(n4993), 
        .QN(n3631) );
  DFFR_X1 \REGISTERS_reg[15][12]  ( .D(n3094), .CK(CLK), .RN(n1494), .Q(n4992), 
        .QN(n3606) );
  DFFR_X1 \REGISTERS_reg[15][11]  ( .D(n3093), .CK(CLK), .RN(n1495), .Q(n4991), 
        .QN(n3581) );
  DFFR_X1 \REGISTERS_reg[15][10]  ( .D(n3092), .CK(CLK), .RN(n1495), .Q(n4990), 
        .QN(n2500) );
  DFFR_X1 \REGISTERS_reg[15][9]  ( .D(n3091), .CK(CLK), .RN(n1495), .Q(n4989), 
        .QN(n2475) );
  DFFR_X1 \REGISTERS_reg[15][8]  ( .D(n3090), .CK(CLK), .RN(n1495), .Q(n4988), 
        .QN(n2450) );
  DFFR_X1 \REGISTERS_reg[15][7]  ( .D(n3089), .CK(CLK), .RN(n1495), .Q(n4987), 
        .QN(n2425) );
  DFFR_X1 \REGISTERS_reg[15][6]  ( .D(n3088), .CK(CLK), .RN(n1495), .Q(n4986), 
        .QN(n2400) );
  DFFR_X1 \REGISTERS_reg[15][5]  ( .D(n3087), .CK(CLK), .RN(n1495), .Q(n4985), 
        .QN(n2375) );
  DFFR_X1 \REGISTERS_reg[15][4]  ( .D(n3086), .CK(CLK), .RN(n1495), .Q(n4984), 
        .QN(n2350) );
  DFFR_X1 \REGISTERS_reg[15][3]  ( .D(n3085), .CK(CLK), .RN(n1495), .Q(n4983), 
        .QN(n2325) );
  DFFR_X1 \REGISTERS_reg[15][2]  ( .D(n3084), .CK(CLK), .RN(n1495), .Q(n4982), 
        .QN(n2300) );
  DFFR_X1 \REGISTERS_reg[15][1]  ( .D(n3083), .CK(CLK), .RN(n1495), .Q(n4981), 
        .QN(n2275) );
  DFFR_X1 \REGISTERS_reg[15][0]  ( .D(n3082), .CK(CLK), .RN(n1495), .Q(n4980), 
        .QN(n2246) );
  DFFR_X1 \REGISTERS_reg[16][23]  ( .D(n3073), .CK(CLK), .RN(n1496), .Q(n4232)
         );
  DFFR_X1 \REGISTERS_reg[16][22]  ( .D(n3072), .CK(CLK), .RN(n1496), .Q(n4233)
         );
  DFFR_X1 \REGISTERS_reg[16][21]  ( .D(n3071), .CK(CLK), .RN(n1496), .Q(n4234)
         );
  DFFR_X1 \REGISTERS_reg[16][20]  ( .D(n3070), .CK(CLK), .RN(n1496), .Q(n4235)
         );
  DFFR_X1 \REGISTERS_reg[16][19]  ( .D(n3069), .CK(CLK), .RN(n1497), .Q(n4236)
         );
  DFFR_X1 \REGISTERS_reg[16][18]  ( .D(n3068), .CK(CLK), .RN(n1497), .Q(n4237)
         );
  DFFR_X1 \REGISTERS_reg[16][17]  ( .D(n3067), .CK(CLK), .RN(n1497), .Q(n4238)
         );
  DFFR_X1 \REGISTERS_reg[16][16]  ( .D(n3066), .CK(CLK), .RN(n1497), .Q(n4239)
         );
  DFFR_X1 \REGISTERS_reg[16][15]  ( .D(n3065), .CK(CLK), .RN(n1497), .Q(n4240)
         );
  DFFR_X1 \REGISTERS_reg[16][14]  ( .D(n3064), .CK(CLK), .RN(n1497), .Q(n4241)
         );
  DFFR_X1 \REGISTERS_reg[16][13]  ( .D(n3063), .CK(CLK), .RN(n1497), .Q(n4242)
         );
  DFFR_X1 \REGISTERS_reg[16][12]  ( .D(n3062), .CK(CLK), .RN(n1497), .Q(n4243)
         );
  DFFR_X1 \REGISTERS_reg[16][11]  ( .D(n3061), .CK(CLK), .RN(n1497), .Q(n4244)
         );
  DFFR_X1 \REGISTERS_reg[16][10]  ( .D(n3060), .CK(CLK), .RN(n1497), .Q(n4245)
         );
  DFFR_X1 \REGISTERS_reg[16][9]  ( .D(n3059), .CK(CLK), .RN(n1497), .Q(n4246)
         );
  DFFR_X1 \REGISTERS_reg[16][8]  ( .D(n3058), .CK(CLK), .RN(n1497), .Q(n4247)
         );
  DFFR_X1 \REGISTERS_reg[16][7]  ( .D(n3057), .CK(CLK), .RN(n1498), .Q(n4248)
         );
  DFFR_X1 \REGISTERS_reg[16][6]  ( .D(n3056), .CK(CLK), .RN(n1498), .Q(n4249)
         );
  DFFR_X1 \REGISTERS_reg[16][5]  ( .D(n3055), .CK(CLK), .RN(n1498), .Q(n4250)
         );
  DFFR_X1 \REGISTERS_reg[16][4]  ( .D(n3054), .CK(CLK), .RN(n1498), .Q(n4251)
         );
  DFFR_X1 \REGISTERS_reg[16][3]  ( .D(n3053), .CK(CLK), .RN(n1498), .Q(n4252)
         );
  DFFR_X1 \REGISTERS_reg[16][2]  ( .D(n3052), .CK(CLK), .RN(n1498), .Q(n4253)
         );
  DFFR_X1 \REGISTERS_reg[16][1]  ( .D(n3051), .CK(CLK), .RN(n1498), .Q(n4254)
         );
  DFFR_X1 \REGISTERS_reg[16][0]  ( .D(n3050), .CK(CLK), .RN(n1498), .Q(n4255)
         );
  DFFR_X1 \REGISTERS_reg[17][23]  ( .D(n3041), .CK(CLK), .RN(n1499), .Q(n3898), 
        .QN(n525) );
  DFFR_X1 \REGISTERS_reg[17][22]  ( .D(n3040), .CK(CLK), .RN(n1499), .Q(n3873), 
        .QN(n526) );
  DFFR_X1 \REGISTERS_reg[17][21]  ( .D(n3039), .CK(CLK), .RN(n1499), .Q(n3848), 
        .QN(n527) );
  DFFR_X1 \REGISTERS_reg[17][20]  ( .D(n3038), .CK(CLK), .RN(n1499), .Q(n3823), 
        .QN(n528) );
  DFFR_X1 \REGISTERS_reg[17][19]  ( .D(n3037), .CK(CLK), .RN(n1499), .Q(n3798), 
        .QN(n529) );
  DFFR_X1 \REGISTERS_reg[17][18]  ( .D(n3036), .CK(CLK), .RN(n1499), .Q(n3773), 
        .QN(n530) );
  DFFR_X1 \REGISTERS_reg[17][17]  ( .D(n3035), .CK(CLK), .RN(n1499), .Q(n3748), 
        .QN(n531) );
  DFFR_X1 \REGISTERS_reg[17][16]  ( .D(n3034), .CK(CLK), .RN(n1499), .Q(n3723), 
        .QN(n532) );
  DFFR_X1 \REGISTERS_reg[17][15]  ( .D(n3033), .CK(CLK), .RN(n1500), .Q(n3698), 
        .QN(n533) );
  DFFR_X1 \REGISTERS_reg[17][14]  ( .D(n3032), .CK(CLK), .RN(n1500), .Q(n3673), 
        .QN(n534) );
  DFFR_X1 \REGISTERS_reg[17][13]  ( .D(n3031), .CK(CLK), .RN(n1500), .Q(n3648), 
        .QN(n535) );
  DFFR_X1 \REGISTERS_reg[17][12]  ( .D(n3030), .CK(CLK), .RN(n1500), .Q(n3623), 
        .QN(n536) );
  DFFR_X1 \REGISTERS_reg[17][11]  ( .D(n3029), .CK(CLK), .RN(n1500), .Q(n3598), 
        .QN(n537) );
  DFFR_X1 \REGISTERS_reg[17][10]  ( .D(n3028), .CK(CLK), .RN(n1500), .Q(n3573), 
        .QN(n538) );
  DFFR_X1 \REGISTERS_reg[17][9]  ( .D(n3027), .CK(CLK), .RN(n1500), .Q(n2492), 
        .QN(n539) );
  DFFR_X1 \REGISTERS_reg[17][8]  ( .D(n3026), .CK(CLK), .RN(n1500), .Q(n2467), 
        .QN(n540) );
  DFFR_X1 \REGISTERS_reg[17][7]  ( .D(n3025), .CK(CLK), .RN(n1500), .Q(n2442), 
        .QN(n541) );
  DFFR_X1 \REGISTERS_reg[17][6]  ( .D(n3024), .CK(CLK), .RN(n1500), .Q(n2417), 
        .QN(n542) );
  DFFR_X1 \REGISTERS_reg[17][5]  ( .D(n3023), .CK(CLK), .RN(n1500), .Q(n2392), 
        .QN(n543) );
  DFFR_X1 \REGISTERS_reg[17][4]  ( .D(n3022), .CK(CLK), .RN(n1500), .Q(n2367), 
        .QN(n544) );
  DFFR_X1 \REGISTERS_reg[17][3]  ( .D(n3021), .CK(CLK), .RN(n1501), .Q(n2342), 
        .QN(n545) );
  DFFR_X1 \REGISTERS_reg[17][2]  ( .D(n3020), .CK(CLK), .RN(n1501), .Q(n2317), 
        .QN(n546) );
  DFFR_X1 \REGISTERS_reg[17][1]  ( .D(n3019), .CK(CLK), .RN(n1501), .Q(n2292), 
        .QN(n547) );
  DFFR_X1 \REGISTERS_reg[17][0]  ( .D(n3018), .CK(CLK), .RN(n1501), .Q(n2267), 
        .QN(n548) );
  DFFR_X1 \REGISTERS_reg[18][31]  ( .D(n3017), .CK(CLK), .RN(n1501), .Q(n4979)
         );
  DFFR_X1 \REGISTERS_reg[18][30]  ( .D(n3016), .CK(CLK), .RN(n1501), .Q(n4978)
         );
  DFFR_X1 \REGISTERS_reg[18][29]  ( .D(n3015), .CK(CLK), .RN(n1501), .Q(n4977)
         );
  DFFR_X1 \REGISTERS_reg[18][28]  ( .D(n3014), .CK(CLK), .RN(n1501), .Q(n4976)
         );
  DFFR_X1 \REGISTERS_reg[18][27]  ( .D(n3013), .CK(CLK), .RN(n1501), .Q(n4975)
         );
  DFFR_X1 \REGISTERS_reg[18][26]  ( .D(n3012), .CK(CLK), .RN(n1501), .Q(n4974)
         );
  DFFR_X1 \REGISTERS_reg[18][25]  ( .D(n3011), .CK(CLK), .RN(n1501), .Q(n4973)
         );
  DFFR_X1 \REGISTERS_reg[18][24]  ( .D(n3010), .CK(CLK), .RN(n1501), .Q(n4972)
         );
  DFFR_X1 \REGISTERS_reg[18][23]  ( .D(n3009), .CK(CLK), .RN(n1502), .Q(n4971)
         );
  DFFR_X1 \REGISTERS_reg[18][22]  ( .D(n3008), .CK(CLK), .RN(n1502), .Q(n4970)
         );
  DFFR_X1 \REGISTERS_reg[18][21]  ( .D(n3007), .CK(CLK), .RN(n1502), .Q(n4969)
         );
  DFFR_X1 \REGISTERS_reg[18][20]  ( .D(n3006), .CK(CLK), .RN(n1502), .Q(n4968)
         );
  DFFR_X1 \REGISTERS_reg[18][19]  ( .D(n3005), .CK(CLK), .RN(n1502), .Q(n4967)
         );
  DFFR_X1 \REGISTERS_reg[18][18]  ( .D(n3004), .CK(CLK), .RN(n1502), .Q(n4966)
         );
  DFFR_X1 \REGISTERS_reg[18][17]  ( .D(n3003), .CK(CLK), .RN(n1502), .Q(n4965)
         );
  DFFR_X1 \REGISTERS_reg[18][16]  ( .D(n3002), .CK(CLK), .RN(n1502), .Q(n4964)
         );
  DFFR_X1 \REGISTERS_reg[18][15]  ( .D(n3001), .CK(CLK), .RN(n1502), .Q(n4963)
         );
  DFFR_X1 \REGISTERS_reg[18][14]  ( .D(n3000), .CK(CLK), .RN(n1502), .Q(n4962)
         );
  DFFR_X1 \REGISTERS_reg[18][13]  ( .D(n2999), .CK(CLK), .RN(n1502), .Q(n4961)
         );
  DFFR_X1 \REGISTERS_reg[18][12]  ( .D(n2998), .CK(CLK), .RN(n1502), .Q(n4960)
         );
  DFFR_X1 \REGISTERS_reg[18][11]  ( .D(n2997), .CK(CLK), .RN(n1503), .Q(n4959)
         );
  DFFR_X1 \REGISTERS_reg[18][10]  ( .D(n2996), .CK(CLK), .RN(n1503), .Q(n4958)
         );
  DFFR_X1 \REGISTERS_reg[18][9]  ( .D(n2995), .CK(CLK), .RN(n1503), .Q(n4957)
         );
  DFFR_X1 \REGISTERS_reg[18][8]  ( .D(n2994), .CK(CLK), .RN(n1503), .Q(n4956)
         );
  DFFR_X1 \REGISTERS_reg[18][7]  ( .D(n2993), .CK(CLK), .RN(n1503), .Q(n4955)
         );
  DFFR_X1 \REGISTERS_reg[18][6]  ( .D(n2992), .CK(CLK), .RN(n1503), .Q(n4954)
         );
  DFFR_X1 \REGISTERS_reg[18][5]  ( .D(n2991), .CK(CLK), .RN(n1503), .Q(n4953)
         );
  DFFR_X1 \REGISTERS_reg[18][4]  ( .D(n2990), .CK(CLK), .RN(n1503), .Q(n4952)
         );
  DFFR_X1 \REGISTERS_reg[18][3]  ( .D(n2989), .CK(CLK), .RN(n1503), .Q(n4951)
         );
  DFFR_X1 \REGISTERS_reg[18][2]  ( .D(n2988), .CK(CLK), .RN(n1503), .Q(n4950)
         );
  DFFR_X1 \REGISTERS_reg[18][1]  ( .D(n2987), .CK(CLK), .RN(n1503), .Q(n4949)
         );
  DFFR_X1 \REGISTERS_reg[18][0]  ( .D(n2986), .CK(CLK), .RN(n1503), .Q(n4948)
         );
  DFFR_X1 \REGISTERS_reg[19][31]  ( .D(n2985), .CK(CLK), .RN(n1504), .Q(n4947), 
        .QN(n4115) );
  DFFR_X1 \REGISTERS_reg[19][30]  ( .D(n2984), .CK(CLK), .RN(n1504), .Q(n4946), 
        .QN(n4076) );
  DFFR_X1 \REGISTERS_reg[19][29]  ( .D(n2983), .CK(CLK), .RN(n1504), .Q(n4945), 
        .QN(n4050) );
  DFFR_X1 \REGISTERS_reg[19][28]  ( .D(n2982), .CK(CLK), .RN(n1504), .Q(n4944), 
        .QN(n4024) );
  DFFR_X1 \REGISTERS_reg[19][27]  ( .D(n2981), .CK(CLK), .RN(n1504), .Q(n4943), 
        .QN(n3998) );
  DFFR_X1 \REGISTERS_reg[19][26]  ( .D(n2980), .CK(CLK), .RN(n1504), .Q(n4942), 
        .QN(n3972) );
  DFFR_X1 \REGISTERS_reg[19][25]  ( .D(n2979), .CK(CLK), .RN(n1504), .Q(n4941), 
        .QN(n3946) );
  DFFR_X1 \REGISTERS_reg[19][24]  ( .D(n2978), .CK(CLK), .RN(n1504), .Q(n4940), 
        .QN(n3920) );
  DFFR_X1 \REGISTERS_reg[19][23]  ( .D(n2977), .CK(CLK), .RN(n1504), .Q(n4939), 
        .QN(n3894) );
  DFFR_X1 \REGISTERS_reg[19][22]  ( .D(n2976), .CK(CLK), .RN(n1504), .Q(n4938), 
        .QN(n3869) );
  DFFR_X1 \REGISTERS_reg[19][21]  ( .D(n2975), .CK(CLK), .RN(n1504), .Q(n4937), 
        .QN(n3844) );
  DFFR_X1 \REGISTERS_reg[19][20]  ( .D(n2974), .CK(CLK), .RN(n1504), .Q(n4936), 
        .QN(n3819) );
  DFFR_X1 \REGISTERS_reg[19][19]  ( .D(n2973), .CK(CLK), .RN(n1505), .Q(n4935), 
        .QN(n3794) );
  DFFR_X1 \REGISTERS_reg[19][18]  ( .D(n2972), .CK(CLK), .RN(n1505), .Q(n4934), 
        .QN(n3769) );
  DFFR_X1 \REGISTERS_reg[19][17]  ( .D(n2971), .CK(CLK), .RN(n1505), .Q(n4933), 
        .QN(n3744) );
  DFFR_X1 \REGISTERS_reg[19][16]  ( .D(n2970), .CK(CLK), .RN(n1505), .Q(n4932), 
        .QN(n3719) );
  DFFR_X1 \REGISTERS_reg[19][15]  ( .D(n2969), .CK(CLK), .RN(n1505), .Q(n4931), 
        .QN(n3694) );
  DFFR_X1 \REGISTERS_reg[19][14]  ( .D(n2968), .CK(CLK), .RN(n1505), .Q(n4930), 
        .QN(n3669) );
  DFFR_X1 \REGISTERS_reg[19][13]  ( .D(n2967), .CK(CLK), .RN(n1505), .Q(n4929), 
        .QN(n3644) );
  DFFR_X1 \REGISTERS_reg[19][12]  ( .D(n2966), .CK(CLK), .RN(n1505), .Q(n4928), 
        .QN(n3619) );
  DFFR_X1 \REGISTERS_reg[19][11]  ( .D(n2965), .CK(CLK), .RN(n1505), .Q(n4927), 
        .QN(n3594) );
  DFFR_X1 \REGISTERS_reg[19][10]  ( .D(n2964), .CK(CLK), .RN(n1505), .Q(n4926), 
        .QN(n3569) );
  DFFR_X1 \REGISTERS_reg[19][9]  ( .D(n2963), .CK(CLK), .RN(n1505), .Q(n4925), 
        .QN(n2488) );
  DFFR_X1 \REGISTERS_reg[19][8]  ( .D(n2962), .CK(CLK), .RN(n1505), .Q(n4924), 
        .QN(n2463) );
  DFFR_X1 \REGISTERS_reg[19][7]  ( .D(n2961), .CK(CLK), .RN(n1506), .Q(n4923), 
        .QN(n2438) );
  DFFR_X1 \REGISTERS_reg[19][6]  ( .D(n2960), .CK(CLK), .RN(n1506), .Q(n4922), 
        .QN(n2413) );
  DFFR_X1 \REGISTERS_reg[19][5]  ( .D(n2959), .CK(CLK), .RN(n1506), .Q(n4921), 
        .QN(n2388) );
  DFFR_X1 \REGISTERS_reg[19][4]  ( .D(n2958), .CK(CLK), .RN(n1506), .Q(n4920), 
        .QN(n2363) );
  DFFR_X1 \REGISTERS_reg[19][3]  ( .D(n2957), .CK(CLK), .RN(n1506), .Q(n4919), 
        .QN(n2338) );
  DFFR_X1 \REGISTERS_reg[19][2]  ( .D(n2956), .CK(CLK), .RN(n1506), .Q(n4918), 
        .QN(n2313) );
  DFFR_X1 \REGISTERS_reg[19][1]  ( .D(n2955), .CK(CLK), .RN(n1506), .Q(n4917), 
        .QN(n2288) );
  DFFR_X1 \REGISTERS_reg[19][0]  ( .D(n2954), .CK(CLK), .RN(n1506), .Q(n4916), 
        .QN(n2261) );
  DFFR_X1 \REGISTERS_reg[20][23]  ( .D(n2945), .CK(CLK), .RN(n1507), .QN(n621)
         );
  DFFR_X1 \REGISTERS_reg[20][22]  ( .D(n2944), .CK(CLK), .RN(n1507), .QN(n622)
         );
  DFFR_X1 \REGISTERS_reg[20][21]  ( .D(n2943), .CK(CLK), .RN(n1507), .QN(n623)
         );
  DFFR_X1 \REGISTERS_reg[20][20]  ( .D(n2942), .CK(CLK), .RN(n1507), .QN(n624)
         );
  DFFR_X1 \REGISTERS_reg[20][19]  ( .D(n2941), .CK(CLK), .RN(n1507), .QN(n625)
         );
  DFFR_X1 \REGISTERS_reg[20][18]  ( .D(n2940), .CK(CLK), .RN(n1507), .QN(n626)
         );
  DFFR_X1 \REGISTERS_reg[20][17]  ( .D(n2939), .CK(CLK), .RN(n1507), .QN(n627)
         );
  DFFR_X1 \REGISTERS_reg[20][16]  ( .D(n2938), .CK(CLK), .RN(n1507), .QN(n628)
         );
  DFFR_X1 \REGISTERS_reg[20][15]  ( .D(n2937), .CK(CLK), .RN(n1508), .QN(n629)
         );
  DFFR_X1 \REGISTERS_reg[20][14]  ( .D(n2936), .CK(CLK), .RN(n1508), .QN(n630)
         );
  DFFR_X1 \REGISTERS_reg[20][13]  ( .D(n2935), .CK(CLK), .RN(n1508), .QN(n631)
         );
  DFFR_X1 \REGISTERS_reg[20][12]  ( .D(n2934), .CK(CLK), .RN(n1508), .QN(n632)
         );
  DFFR_X1 \REGISTERS_reg[20][11]  ( .D(n2933), .CK(CLK), .RN(n1508), .QN(n633)
         );
  DFFR_X1 \REGISTERS_reg[20][10]  ( .D(n2932), .CK(CLK), .RN(n1508), .QN(n634)
         );
  DFFR_X1 \REGISTERS_reg[20][9]  ( .D(n2931), .CK(CLK), .RN(n1508), .QN(n635)
         );
  DFFR_X1 \REGISTERS_reg[20][8]  ( .D(n2930), .CK(CLK), .RN(n1508), .QN(n636)
         );
  DFFR_X1 \REGISTERS_reg[20][7]  ( .D(n2929), .CK(CLK), .RN(n1508), .QN(n637)
         );
  DFFR_X1 \REGISTERS_reg[20][6]  ( .D(n2928), .CK(CLK), .RN(n1508), .QN(n638)
         );
  DFFR_X1 \REGISTERS_reg[20][5]  ( .D(n2927), .CK(CLK), .RN(n1508), .QN(n639)
         );
  DFFR_X1 \REGISTERS_reg[20][4]  ( .D(n2926), .CK(CLK), .RN(n1508), .QN(n640)
         );
  DFFR_X1 \REGISTERS_reg[20][3]  ( .D(n2925), .CK(CLK), .RN(n1509), .QN(n641)
         );
  DFFR_X1 \REGISTERS_reg[20][2]  ( .D(n2924), .CK(CLK), .RN(n1509), .QN(n642)
         );
  DFFR_X1 \REGISTERS_reg[20][1]  ( .D(n2923), .CK(CLK), .RN(n1509), .QN(n643)
         );
  DFFR_X1 \REGISTERS_reg[20][0]  ( .D(n2922), .CK(CLK), .RN(n1509), .QN(n644)
         );
  DFFR_X1 \REGISTERS_reg[21][23]  ( .D(n2913), .CK(CLK), .RN(n1510), .Q(n4264)
         );
  DFFR_X1 \REGISTERS_reg[21][22]  ( .D(n2912), .CK(CLK), .RN(n1510), .Q(n4265)
         );
  DFFR_X1 \REGISTERS_reg[21][21]  ( .D(n2911), .CK(CLK), .RN(n1510), .Q(n4266)
         );
  DFFR_X1 \REGISTERS_reg[21][20]  ( .D(n2910), .CK(CLK), .RN(n1510), .Q(n4267)
         );
  DFFR_X1 \REGISTERS_reg[21][19]  ( .D(n2909), .CK(CLK), .RN(n1510), .Q(n4268)
         );
  DFFR_X1 \REGISTERS_reg[21][18]  ( .D(n2908), .CK(CLK), .RN(n1510), .Q(n4269)
         );
  DFFR_X1 \REGISTERS_reg[21][17]  ( .D(n2907), .CK(CLK), .RN(n1510), .Q(n4270)
         );
  DFFR_X1 \REGISTERS_reg[21][16]  ( .D(n2906), .CK(CLK), .RN(n1510), .Q(n4271)
         );
  DFFR_X1 \REGISTERS_reg[21][15]  ( .D(n2905), .CK(CLK), .RN(n1510), .Q(n4272)
         );
  DFFR_X1 \REGISTERS_reg[21][14]  ( .D(n2904), .CK(CLK), .RN(n1510), .Q(n4273)
         );
  DFFR_X1 \REGISTERS_reg[21][13]  ( .D(n2903), .CK(CLK), .RN(n1510), .Q(n4274)
         );
  DFFR_X1 \REGISTERS_reg[21][12]  ( .D(n2902), .CK(CLK), .RN(n1510), .Q(n4275)
         );
  DFFR_X1 \REGISTERS_reg[21][11]  ( .D(n2901), .CK(CLK), .RN(n1511), .Q(n4276)
         );
  DFFR_X1 \REGISTERS_reg[21][10]  ( .D(n2900), .CK(CLK), .RN(n1511), .Q(n4277)
         );
  DFFR_X1 \REGISTERS_reg[21][9]  ( .D(n2899), .CK(CLK), .RN(n1511), .Q(n4278)
         );
  DFFR_X1 \REGISTERS_reg[21][8]  ( .D(n2898), .CK(CLK), .RN(n1511), .Q(n4279)
         );
  DFFR_X1 \REGISTERS_reg[21][7]  ( .D(n2897), .CK(CLK), .RN(n1511), .Q(n4280)
         );
  DFFR_X1 \REGISTERS_reg[21][6]  ( .D(n2896), .CK(CLK), .RN(n1511), .Q(n4281)
         );
  DFFR_X1 \REGISTERS_reg[21][5]  ( .D(n2895), .CK(CLK), .RN(n1511), .Q(n4282)
         );
  DFFR_X1 \REGISTERS_reg[21][4]  ( .D(n2894), .CK(CLK), .RN(n1511), .Q(n4283)
         );
  DFFR_X1 \REGISTERS_reg[21][3]  ( .D(n2893), .CK(CLK), .RN(n1511), .Q(n4284)
         );
  DFFR_X1 \REGISTERS_reg[21][2]  ( .D(n2892), .CK(CLK), .RN(n1511), .Q(n4285)
         );
  DFFR_X1 \REGISTERS_reg[21][1]  ( .D(n2891), .CK(CLK), .RN(n1511), .Q(n4286)
         );
  DFFR_X1 \REGISTERS_reg[21][0]  ( .D(n2890), .CK(CLK), .RN(n1511), .Q(n4287)
         );
  DFFR_X1 \REGISTERS_reg[22][31]  ( .D(n2889), .CK(CLK), .RN(n1512), .Q(n4915), 
        .QN(n4117) );
  DFFR_X1 \REGISTERS_reg[22][30]  ( .D(n2888), .CK(CLK), .RN(n1512), .Q(n4914), 
        .QN(n4077) );
  DFFR_X1 \REGISTERS_reg[22][29]  ( .D(n2887), .CK(CLK), .RN(n1512), .Q(n4913), 
        .QN(n4051) );
  DFFR_X1 \REGISTERS_reg[22][28]  ( .D(n2886), .CK(CLK), .RN(n1512), .Q(n4912), 
        .QN(n4025) );
  DFFR_X1 \REGISTERS_reg[22][27]  ( .D(n2885), .CK(CLK), .RN(n1512), .Q(n4911), 
        .QN(n3999) );
  DFFR_X1 \REGISTERS_reg[22][26]  ( .D(n2884), .CK(CLK), .RN(n1512), .Q(n4910), 
        .QN(n3973) );
  DFFR_X1 \REGISTERS_reg[22][25]  ( .D(n2883), .CK(CLK), .RN(n1512), .Q(n4909), 
        .QN(n3947) );
  DFFR_X1 \REGISTERS_reg[22][24]  ( .D(n2882), .CK(CLK), .RN(n1512), .Q(n4908), 
        .QN(n3921) );
  DFFR_X1 \REGISTERS_reg[22][23]  ( .D(n2881), .CK(CLK), .RN(n1512), .Q(n4907), 
        .QN(n3895) );
  DFFR_X1 \REGISTERS_reg[22][22]  ( .D(n2880), .CK(CLK), .RN(n1512), .Q(n4906), 
        .QN(n3870) );
  DFFR_X1 \REGISTERS_reg[22][21]  ( .D(n2879), .CK(CLK), .RN(n1512), .Q(n4905), 
        .QN(n3845) );
  DFFR_X1 \REGISTERS_reg[22][20]  ( .D(n2878), .CK(CLK), .RN(n1512), .Q(n4904), 
        .QN(n3820) );
  DFFR_X1 \REGISTERS_reg[22][19]  ( .D(n2877), .CK(CLK), .RN(n1513), .Q(n4903), 
        .QN(n3795) );
  DFFR_X1 \REGISTERS_reg[22][18]  ( .D(n2876), .CK(CLK), .RN(n1513), .Q(n4902), 
        .QN(n3770) );
  DFFR_X1 \REGISTERS_reg[22][17]  ( .D(n2875), .CK(CLK), .RN(n1513), .Q(n4901), 
        .QN(n3745) );
  DFFR_X1 \REGISTERS_reg[22][16]  ( .D(n2874), .CK(CLK), .RN(n1513), .Q(n4900), 
        .QN(n3720) );
  DFFR_X1 \REGISTERS_reg[22][15]  ( .D(n2873), .CK(CLK), .RN(n1513), .Q(n4899), 
        .QN(n3695) );
  DFFR_X1 \REGISTERS_reg[22][14]  ( .D(n2872), .CK(CLK), .RN(n1513), .Q(n4898), 
        .QN(n3670) );
  DFFR_X1 \REGISTERS_reg[22][13]  ( .D(n2871), .CK(CLK), .RN(n1513), .Q(n4897), 
        .QN(n3645) );
  DFFR_X1 \REGISTERS_reg[22][12]  ( .D(n2870), .CK(CLK), .RN(n1513), .Q(n4896), 
        .QN(n3620) );
  DFFR_X1 \REGISTERS_reg[22][11]  ( .D(n2869), .CK(CLK), .RN(n1513), .Q(n4895), 
        .QN(n3595) );
  DFFR_X1 \REGISTERS_reg[22][10]  ( .D(n2868), .CK(CLK), .RN(n1513), .Q(n4894), 
        .QN(n3570) );
  DFFR_X1 \REGISTERS_reg[22][9]  ( .D(n2867), .CK(CLK), .RN(n1513), .Q(n4893), 
        .QN(n2489) );
  DFFR_X1 \REGISTERS_reg[22][8]  ( .D(n2866), .CK(CLK), .RN(n1513), .Q(n4892), 
        .QN(n2464) );
  DFFR_X1 \REGISTERS_reg[22][7]  ( .D(n2865), .CK(CLK), .RN(n1514), .Q(n4891), 
        .QN(n2439) );
  DFFR_X1 \REGISTERS_reg[22][6]  ( .D(n2864), .CK(CLK), .RN(n1514), .Q(n4890), 
        .QN(n2414) );
  DFFR_X1 \REGISTERS_reg[22][5]  ( .D(n2863), .CK(CLK), .RN(n1514), .Q(n4889), 
        .QN(n2389) );
  DFFR_X1 \REGISTERS_reg[22][4]  ( .D(n2862), .CK(CLK), .RN(n1514), .Q(n4888), 
        .QN(n2364) );
  DFFR_X1 \REGISTERS_reg[22][3]  ( .D(n2861), .CK(CLK), .RN(n1514), .Q(n4887), 
        .QN(n2339) );
  DFFR_X1 \REGISTERS_reg[22][2]  ( .D(n2860), .CK(CLK), .RN(n1514), .Q(n4886), 
        .QN(n2314) );
  DFFR_X1 \REGISTERS_reg[22][1]  ( .D(n2859), .CK(CLK), .RN(n1514), .Q(n4885), 
        .QN(n2289) );
  DFFR_X1 \REGISTERS_reg[22][0]  ( .D(n2858), .CK(CLK), .RN(n1514), .Q(n4884), 
        .QN(n2262) );
  DFFR_X1 \REGISTERS_reg[23][31]  ( .D(n2857), .CK(CLK), .RN(n1514), .Q(n4883)
         );
  DFFR_X1 \REGISTERS_reg[23][30]  ( .D(n2856), .CK(CLK), .RN(n1514), .Q(n4882)
         );
  DFFR_X1 \REGISTERS_reg[23][29]  ( .D(n2855), .CK(CLK), .RN(n1514), .Q(n4881)
         );
  DFFR_X1 \REGISTERS_reg[23][28]  ( .D(n2854), .CK(CLK), .RN(n1514), .Q(n4880)
         );
  DFFR_X1 \REGISTERS_reg[23][27]  ( .D(n2853), .CK(CLK), .RN(n1515), .Q(n4879)
         );
  DFFR_X1 \REGISTERS_reg[23][26]  ( .D(n2852), .CK(CLK), .RN(n1515), .Q(n4878)
         );
  DFFR_X1 \REGISTERS_reg[23][25]  ( .D(n2851), .CK(CLK), .RN(n1515), .Q(n4877)
         );
  DFFR_X1 \REGISTERS_reg[23][24]  ( .D(n2850), .CK(CLK), .RN(n1515), .Q(n4876)
         );
  DFFR_X1 \REGISTERS_reg[23][23]  ( .D(n2849), .CK(CLK), .RN(n1515), .Q(n4875)
         );
  DFFR_X1 \REGISTERS_reg[23][22]  ( .D(n2848), .CK(CLK), .RN(n1515), .Q(n4874)
         );
  DFFR_X1 \REGISTERS_reg[23][21]  ( .D(n2847), .CK(CLK), .RN(n1515), .Q(n4873)
         );
  DFFR_X1 \REGISTERS_reg[23][20]  ( .D(n2846), .CK(CLK), .RN(n1515), .Q(n4872)
         );
  DFFR_X1 \REGISTERS_reg[23][19]  ( .D(n2845), .CK(CLK), .RN(n1515), .Q(n4871)
         );
  DFFR_X1 \REGISTERS_reg[23][18]  ( .D(n2844), .CK(CLK), .RN(n1515), .Q(n4870)
         );
  DFFR_X1 \REGISTERS_reg[23][17]  ( .D(n2843), .CK(CLK), .RN(n1515), .Q(n4869)
         );
  DFFR_X1 \REGISTERS_reg[23][16]  ( .D(n2842), .CK(CLK), .RN(n1515), .Q(n4868)
         );
  DFFR_X1 \REGISTERS_reg[23][15]  ( .D(n2841), .CK(CLK), .RN(n1516), .Q(n4867)
         );
  DFFR_X1 \REGISTERS_reg[23][14]  ( .D(n2840), .CK(CLK), .RN(n1516), .Q(n4866)
         );
  DFFR_X1 \REGISTERS_reg[23][13]  ( .D(n2839), .CK(CLK), .RN(n1516), .Q(n4865)
         );
  DFFR_X1 \REGISTERS_reg[23][12]  ( .D(n2838), .CK(CLK), .RN(n1516), .Q(n4864)
         );
  DFFR_X1 \REGISTERS_reg[23][11]  ( .D(n2837), .CK(CLK), .RN(n1516), .Q(n4863)
         );
  DFFR_X1 \REGISTERS_reg[23][10]  ( .D(n2836), .CK(CLK), .RN(n1516), .Q(n4862)
         );
  DFFR_X1 \REGISTERS_reg[23][9]  ( .D(n2835), .CK(CLK), .RN(n1516), .Q(n4861)
         );
  DFFR_X1 \REGISTERS_reg[23][8]  ( .D(n2834), .CK(CLK), .RN(n1516), .Q(n4860)
         );
  DFFR_X1 \REGISTERS_reg[23][7]  ( .D(n2833), .CK(CLK), .RN(n1516), .Q(n4859)
         );
  DFFR_X1 \REGISTERS_reg[23][6]  ( .D(n2832), .CK(CLK), .RN(n1516), .Q(n4858)
         );
  DFFR_X1 \REGISTERS_reg[23][5]  ( .D(n2831), .CK(CLK), .RN(n1516), .Q(n4857)
         );
  DFFR_X1 \REGISTERS_reg[23][4]  ( .D(n2830), .CK(CLK), .RN(n1516), .Q(n4856)
         );
  DFFR_X1 \REGISTERS_reg[23][3]  ( .D(n2829), .CK(CLK), .RN(n1517), .Q(n4855)
         );
  DFFR_X1 \REGISTERS_reg[23][2]  ( .D(n2828), .CK(CLK), .RN(n1517), .Q(n4854)
         );
  DFFR_X1 \REGISTERS_reg[23][1]  ( .D(n2827), .CK(CLK), .RN(n1517), .Q(n4853)
         );
  DFFR_X1 \REGISTERS_reg[23][0]  ( .D(n2826), .CK(CLK), .RN(n1517), .Q(n4852)
         );
  DFFR_X1 \REGISTERS_reg[24][31]  ( .D(n2825), .CK(CLK), .RN(n1517), .Q(n4851), 
        .QN(n4104) );
  DFFR_X1 \REGISTERS_reg[24][30]  ( .D(n2824), .CK(CLK), .RN(n1517), .Q(n4850), 
        .QN(n4070) );
  DFFR_X1 \REGISTERS_reg[24][29]  ( .D(n2823), .CK(CLK), .RN(n1517), .Q(n4849), 
        .QN(n4044) );
  DFFR_X1 \REGISTERS_reg[24][28]  ( .D(n2822), .CK(CLK), .RN(n1517), .Q(n4848), 
        .QN(n4018) );
  DFFR_X1 \REGISTERS_reg[24][27]  ( .D(n2821), .CK(CLK), .RN(n1517), .Q(n4847), 
        .QN(n3992) );
  DFFR_X1 \REGISTERS_reg[24][26]  ( .D(n2820), .CK(CLK), .RN(n1517), .Q(n4846), 
        .QN(n3966) );
  DFFR_X1 \REGISTERS_reg[24][25]  ( .D(n2819), .CK(CLK), .RN(n1517), .Q(n4845), 
        .QN(n3940) );
  DFFR_X1 \REGISTERS_reg[24][24]  ( .D(n2818), .CK(CLK), .RN(n1517), .Q(n4844), 
        .QN(n3914) );
  DFFR_X1 \REGISTERS_reg[24][23]  ( .D(n2817), .CK(CLK), .RN(n1518), .Q(n4843), 
        .QN(n3888) );
  DFFR_X1 \REGISTERS_reg[24][22]  ( .D(n2816), .CK(CLK), .RN(n1518), .Q(n4842), 
        .QN(n3863) );
  DFFR_X1 \REGISTERS_reg[24][21]  ( .D(n2815), .CK(CLK), .RN(n1518), .Q(n4841), 
        .QN(n3838) );
  DFFR_X1 \REGISTERS_reg[24][20]  ( .D(n2814), .CK(CLK), .RN(n1518), .Q(n4840), 
        .QN(n3813) );
  DFFR_X1 \REGISTERS_reg[24][19]  ( .D(n2813), .CK(CLK), .RN(n1518), .Q(n4839), 
        .QN(n3788) );
  DFFR_X1 \REGISTERS_reg[24][18]  ( .D(n2812), .CK(CLK), .RN(n1518), .Q(n4838), 
        .QN(n3763) );
  DFFR_X1 \REGISTERS_reg[24][17]  ( .D(n2811), .CK(CLK), .RN(n1518), .Q(n4837), 
        .QN(n3738) );
  DFFR_X1 \REGISTERS_reg[24][16]  ( .D(n2810), .CK(CLK), .RN(n1518), .Q(n4836), 
        .QN(n3713) );
  DFFR_X1 \REGISTERS_reg[24][15]  ( .D(n2809), .CK(CLK), .RN(n1518), .Q(n4835), 
        .QN(n3688) );
  DFFR_X1 \REGISTERS_reg[24][14]  ( .D(n2808), .CK(CLK), .RN(n1518), .Q(n4834), 
        .QN(n3663) );
  DFFR_X1 \REGISTERS_reg[24][13]  ( .D(n2807), .CK(CLK), .RN(n1518), .Q(n4833), 
        .QN(n3638) );
  DFFR_X1 \REGISTERS_reg[24][12]  ( .D(n2806), .CK(CLK), .RN(n1518), .Q(n4832), 
        .QN(n3613) );
  DFFR_X1 \REGISTERS_reg[24][11]  ( .D(n2805), .CK(CLK), .RN(n1519), .Q(n4831), 
        .QN(n3588) );
  DFFR_X1 \REGISTERS_reg[24][10]  ( .D(n2804), .CK(CLK), .RN(n1519), .Q(n4830), 
        .QN(n3563) );
  DFFR_X1 \REGISTERS_reg[24][9]  ( .D(n2803), .CK(CLK), .RN(n1519), .Q(n4829), 
        .QN(n2482) );
  DFFR_X1 \REGISTERS_reg[24][8]  ( .D(n2802), .CK(CLK), .RN(n1519), .Q(n4828), 
        .QN(n2457) );
  DFFR_X1 \REGISTERS_reg[24][7]  ( .D(n2801), .CK(CLK), .RN(n1519), .Q(n4827), 
        .QN(n2432) );
  DFFR_X1 \REGISTERS_reg[24][6]  ( .D(n2800), .CK(CLK), .RN(n1519), .Q(n4826), 
        .QN(n2407) );
  DFFR_X1 \REGISTERS_reg[24][5]  ( .D(n2799), .CK(CLK), .RN(n1519), .Q(n4825), 
        .QN(n2382) );
  DFFR_X1 \REGISTERS_reg[24][4]  ( .D(n2798), .CK(CLK), .RN(n1519), .Q(n4824), 
        .QN(n2357) );
  DFFR_X1 \REGISTERS_reg[24][3]  ( .D(n2797), .CK(CLK), .RN(n1519), .Q(n4823), 
        .QN(n2332) );
  DFFR_X1 \REGISTERS_reg[24][2]  ( .D(n2796), .CK(CLK), .RN(n1519), .Q(n4822), 
        .QN(n2307) );
  DFFR_X1 \REGISTERS_reg[24][1]  ( .D(n2795), .CK(CLK), .RN(n1519), .Q(n4821), 
        .QN(n2282) );
  DFFR_X1 \REGISTERS_reg[24][0]  ( .D(n2794), .CK(CLK), .RN(n1519), .Q(n4820), 
        .QN(n2253) );
  DFFR_X1 \REGISTERS_reg[25][31]  ( .D(n2793), .CK(CLK), .RN(n1520), .Q(n4819)
         );
  DFFR_X1 \REGISTERS_reg[25][30]  ( .D(n2792), .CK(CLK), .RN(n1520), .Q(n4818)
         );
  DFFR_X1 \REGISTERS_reg[25][29]  ( .D(n2791), .CK(CLK), .RN(n1520), .Q(n4817)
         );
  DFFR_X1 \REGISTERS_reg[25][28]  ( .D(n2790), .CK(CLK), .RN(n1520), .Q(n4816)
         );
  DFFR_X1 \REGISTERS_reg[25][27]  ( .D(n2789), .CK(CLK), .RN(n1520), .Q(n4815)
         );
  DFFR_X1 \REGISTERS_reg[25][26]  ( .D(n2788), .CK(CLK), .RN(n1520), .Q(n4814)
         );
  DFFR_X1 \REGISTERS_reg[25][25]  ( .D(n2787), .CK(CLK), .RN(n1520), .Q(n4813)
         );
  DFFR_X1 \REGISTERS_reg[25][24]  ( .D(n2786), .CK(CLK), .RN(n1520), .Q(n4812)
         );
  DFFR_X1 \REGISTERS_reg[25][23]  ( .D(n2785), .CK(CLK), .RN(n1520), .Q(n4811)
         );
  DFFR_X1 \REGISTERS_reg[25][22]  ( .D(n2784), .CK(CLK), .RN(n1520), .Q(n4810)
         );
  DFFR_X1 \REGISTERS_reg[25][21]  ( .D(n2783), .CK(CLK), .RN(n1520), .Q(n4809)
         );
  DFFR_X1 \REGISTERS_reg[25][20]  ( .D(n2782), .CK(CLK), .RN(n1520), .Q(n4808)
         );
  DFFR_X1 \REGISTERS_reg[25][19]  ( .D(n2781), .CK(CLK), .RN(n1521), .Q(n4807)
         );
  DFFR_X1 \REGISTERS_reg[25][18]  ( .D(n2780), .CK(CLK), .RN(n1521), .Q(n4806)
         );
  DFFR_X1 \REGISTERS_reg[25][17]  ( .D(n2779), .CK(CLK), .RN(n1521), .Q(n4805)
         );
  DFFR_X1 \REGISTERS_reg[25][16]  ( .D(n2778), .CK(CLK), .RN(n1521), .Q(n4804)
         );
  DFFR_X1 \REGISTERS_reg[25][15]  ( .D(n2777), .CK(CLK), .RN(n1521), .Q(n4803)
         );
  DFFR_X1 \REGISTERS_reg[25][14]  ( .D(n2776), .CK(CLK), .RN(n1521), .Q(n4802)
         );
  DFFR_X1 \REGISTERS_reg[25][13]  ( .D(n2775), .CK(CLK), .RN(n1521), .Q(n4801)
         );
  DFFR_X1 \REGISTERS_reg[25][12]  ( .D(n2774), .CK(CLK), .RN(n1521), .Q(n4800)
         );
  DFFR_X1 \REGISTERS_reg[25][11]  ( .D(n2773), .CK(CLK), .RN(n1521), .Q(n4799)
         );
  DFFR_X1 \REGISTERS_reg[25][10]  ( .D(n2772), .CK(CLK), .RN(n1521), .Q(n4798)
         );
  DFFR_X1 \REGISTERS_reg[25][9]  ( .D(n2771), .CK(CLK), .RN(n1521), .Q(n4797)
         );
  DFFR_X1 \REGISTERS_reg[25][8]  ( .D(n2770), .CK(CLK), .RN(n1521), .Q(n4796)
         );
  DFFR_X1 \REGISTERS_reg[25][7]  ( .D(n2769), .CK(CLK), .RN(n1522), .Q(n4795)
         );
  DFFR_X1 \REGISTERS_reg[25][6]  ( .D(n2768), .CK(CLK), .RN(n1522), .Q(n4794)
         );
  DFFR_X1 \REGISTERS_reg[25][5]  ( .D(n2767), .CK(CLK), .RN(n1522), .Q(n4793)
         );
  DFFR_X1 \REGISTERS_reg[25][4]  ( .D(n2766), .CK(CLK), .RN(n1522), .Q(n4792)
         );
  DFFR_X1 \REGISTERS_reg[25][3]  ( .D(n2765), .CK(CLK), .RN(n1522), .Q(n4791)
         );
  DFFR_X1 \REGISTERS_reg[25][2]  ( .D(n2764), .CK(CLK), .RN(n1522), .Q(n4790)
         );
  DFFR_X1 \REGISTERS_reg[25][1]  ( .D(n2763), .CK(CLK), .RN(n1522), .Q(n4789)
         );
  DFFR_X1 \REGISTERS_reg[25][0]  ( .D(n2762), .CK(CLK), .RN(n1522), .Q(n4788)
         );
  DFFR_X1 \REGISTERS_reg[26][23]  ( .D(n2753), .CK(CLK), .RN(n1523), .Q(n4296), 
        .QN(n813) );
  DFFR_X1 \REGISTERS_reg[26][22]  ( .D(n2752), .CK(CLK), .RN(n1523), .Q(n4297), 
        .QN(n814) );
  DFFR_X1 \REGISTERS_reg[26][21]  ( .D(n2751), .CK(CLK), .RN(n1523), .Q(n224), 
        .QN(n815) );
  DFFR_X1 \REGISTERS_reg[26][20]  ( .D(n2750), .CK(CLK), .RN(n1523), .Q(n4298), 
        .QN(n816) );
  DFFR_X1 \REGISTERS_reg[26][19]  ( .D(n2749), .CK(CLK), .RN(n1523), .Q(n343), 
        .QN(n817) );
  DFFR_X1 \REGISTERS_reg[26][18]  ( .D(n2748), .CK(CLK), .RN(n1523), .Q(n344), 
        .QN(n818) );
  DFFR_X1 \REGISTERS_reg[26][17]  ( .D(n2747), .CK(CLK), .RN(n1523), .Q(n225), 
        .QN(n819) );
  DFFR_X1 \REGISTERS_reg[26][16]  ( .D(n2746), .CK(CLK), .RN(n1523), .Q(n4299), 
        .QN(n820) );
  DFFR_X1 \REGISTERS_reg[26][15]  ( .D(n2745), .CK(CLK), .RN(n1524), .Q(n345), 
        .QN(n821) );
  DFFR_X1 \REGISTERS_reg[26][14]  ( .D(n2744), .CK(CLK), .RN(n1524), .Q(n4300), 
        .QN(n822) );
  DFFR_X1 \REGISTERS_reg[26][13]  ( .D(n2743), .CK(CLK), .RN(n1524), .Q(n4301), 
        .QN(n823) );
  DFFR_X1 \REGISTERS_reg[26][12]  ( .D(n2742), .CK(CLK), .RN(n1524), .Q(n346), 
        .QN(n824) );
  DFFR_X1 \REGISTERS_reg[26][11]  ( .D(n2741), .CK(CLK), .RN(n1524), .Q(n4302), 
        .QN(n825) );
  DFFR_X1 \REGISTERS_reg[26][10]  ( .D(n2740), .CK(CLK), .RN(n1524), .Q(n226), 
        .QN(n826) );
  DFFR_X1 \REGISTERS_reg[26][9]  ( .D(n2739), .CK(CLK), .RN(n1524), .Q(n4303), 
        .QN(n827) );
  DFFR_X1 \REGISTERS_reg[26][8]  ( .D(n2738), .CK(CLK), .RN(n1524), .Q(n347), 
        .QN(n828) );
  DFFR_X1 \REGISTERS_reg[26][7]  ( .D(n2737), .CK(CLK), .RN(n1524), .Q(n4304), 
        .QN(n829) );
  DFFR_X1 \REGISTERS_reg[26][6]  ( .D(n2736), .CK(CLK), .RN(n1524), .Q(n4305), 
        .QN(n830) );
  DFFR_X1 \REGISTERS_reg[26][5]  ( .D(n2735), .CK(CLK), .RN(n1524), .Q(n351), 
        .QN(n831) );
  DFFR_X1 \REGISTERS_reg[26][4]  ( .D(n2734), .CK(CLK), .RN(n1524), .Q(n348), 
        .QN(n832) );
  DFFR_X1 \REGISTERS_reg[26][3]  ( .D(n2733), .CK(CLK), .RN(n1525), .Q(n349), 
        .QN(n833) );
  DFFR_X1 \REGISTERS_reg[26][2]  ( .D(n2732), .CK(CLK), .RN(n1525), .Q(n4306), 
        .QN(n834) );
  DFFR_X1 \REGISTERS_reg[26][1]  ( .D(n2731), .CK(CLK), .RN(n1525), .Q(n350), 
        .QN(n835) );
  DFFR_X1 \REGISTERS_reg[26][0]  ( .D(n2730), .CK(CLK), .RN(n1525), .Q(n4307), 
        .QN(n836) );
  DFFR_X1 \REGISTERS_reg[27][23]  ( .D(n2721), .CK(CLK), .RN(n1526), .Q(n3891), 
        .QN(n845) );
  DFFR_X1 \REGISTERS_reg[27][22]  ( .D(n2720), .CK(CLK), .RN(n1526), .Q(n3866), 
        .QN(n846) );
  DFFR_X1 \REGISTERS_reg[27][21]  ( .D(n2719), .CK(CLK), .RN(n1526), .Q(n3841), 
        .QN(n847) );
  DFFR_X1 \REGISTERS_reg[27][20]  ( .D(n2718), .CK(CLK), .RN(n1526), .Q(n3816), 
        .QN(n848) );
  DFFR_X1 \REGISTERS_reg[27][19]  ( .D(n2717), .CK(CLK), .RN(n1526), .Q(n3791), 
        .QN(n849) );
  DFFR_X1 \REGISTERS_reg[27][18]  ( .D(n2716), .CK(CLK), .RN(n1526), .Q(n3766), 
        .QN(n850) );
  DFFR_X1 \REGISTERS_reg[27][17]  ( .D(n2715), .CK(CLK), .RN(n1526), .Q(n3741), 
        .QN(n851) );
  DFFR_X1 \REGISTERS_reg[27][16]  ( .D(n2714), .CK(CLK), .RN(n1526), .Q(n3716), 
        .QN(n852) );
  DFFR_X1 \REGISTERS_reg[27][15]  ( .D(n2713), .CK(CLK), .RN(n1526), .Q(n3691), 
        .QN(n853) );
  DFFR_X1 \REGISTERS_reg[27][14]  ( .D(n2712), .CK(CLK), .RN(n1526), .Q(n3666), 
        .QN(n854) );
  DFFR_X1 \REGISTERS_reg[27][13]  ( .D(n2711), .CK(CLK), .RN(n1526), .Q(n3641), 
        .QN(n855) );
  DFFR_X1 \REGISTERS_reg[27][12]  ( .D(n2710), .CK(CLK), .RN(n1526), .Q(n3616), 
        .QN(n856) );
  DFFR_X1 \REGISTERS_reg[27][11]  ( .D(n2709), .CK(CLK), .RN(n1527), .Q(n3591), 
        .QN(n857) );
  DFFR_X1 \REGISTERS_reg[27][10]  ( .D(n2708), .CK(CLK), .RN(n1527), .Q(n3566), 
        .QN(n858) );
  DFFR_X1 \REGISTERS_reg[27][9]  ( .D(n2707), .CK(CLK), .RN(n1527), .Q(n2485), 
        .QN(n859) );
  DFFR_X1 \REGISTERS_reg[27][8]  ( .D(n2706), .CK(CLK), .RN(n1527), .Q(n2460), 
        .QN(n860) );
  DFFR_X1 \REGISTERS_reg[27][7]  ( .D(n2705), .CK(CLK), .RN(n1527), .Q(n2435), 
        .QN(n861) );
  DFFR_X1 \REGISTERS_reg[27][6]  ( .D(n2704), .CK(CLK), .RN(n1527), .Q(n2410), 
        .QN(n862) );
  DFFR_X1 \REGISTERS_reg[27][5]  ( .D(n2703), .CK(CLK), .RN(n1527), .Q(n2385), 
        .QN(n863) );
  DFFR_X1 \REGISTERS_reg[27][4]  ( .D(n2702), .CK(CLK), .RN(n1527), .Q(n2360), 
        .QN(n864) );
  DFFR_X1 \REGISTERS_reg[27][3]  ( .D(n2701), .CK(CLK), .RN(n1527), .Q(n2335), 
        .QN(n865) );
  DFFR_X1 \REGISTERS_reg[27][2]  ( .D(n2700), .CK(CLK), .RN(n1527), .Q(n2310), 
        .QN(n866) );
  DFFR_X1 \REGISTERS_reg[27][1]  ( .D(n2699), .CK(CLK), .RN(n1527), .Q(n2285), 
        .QN(n867) );
  DFFR_X1 \REGISTERS_reg[27][0]  ( .D(n2698), .CK(CLK), .RN(n1527), .Q(n2256), 
        .QN(n868) );
  DFFR_X1 \REGISTERS_reg[28][31]  ( .D(n2697), .CK(CLK), .RN(n1528), .Q(n4787), 
        .QN(n4112) );
  DFFR_X1 \REGISTERS_reg[28][30]  ( .D(n2696), .CK(CLK), .RN(n1528), .Q(n4786), 
        .QN(n4074) );
  DFFR_X1 \REGISTERS_reg[28][29]  ( .D(n2695), .CK(CLK), .RN(n1528), .Q(n4785), 
        .QN(n4048) );
  DFFR_X1 \REGISTERS_reg[28][28]  ( .D(n2694), .CK(CLK), .RN(n1528), .Q(n4784), 
        .QN(n4022) );
  DFFR_X1 \REGISTERS_reg[28][27]  ( .D(n2693), .CK(CLK), .RN(n1528), .Q(n4783), 
        .QN(n3996) );
  DFFR_X1 \REGISTERS_reg[28][26]  ( .D(n2692), .CK(CLK), .RN(n1528), .Q(n4782), 
        .QN(n3970) );
  DFFR_X1 \REGISTERS_reg[28][25]  ( .D(n2691), .CK(CLK), .RN(n1528), .Q(n4781), 
        .QN(n3944) );
  DFFR_X1 \REGISTERS_reg[28][24]  ( .D(n2690), .CK(CLK), .RN(n1528), .Q(n4780), 
        .QN(n3918) );
  DFFR_X1 \REGISTERS_reg[28][23]  ( .D(n2689), .CK(CLK), .RN(n1528), .Q(n4779), 
        .QN(n3892) );
  DFFR_X1 \REGISTERS_reg[28][22]  ( .D(n2688), .CK(CLK), .RN(n1528), .Q(n4778), 
        .QN(n3867) );
  DFFR_X1 \REGISTERS_reg[28][21]  ( .D(n2687), .CK(CLK), .RN(n1528), .Q(n4777), 
        .QN(n3842) );
  DFFR_X1 \REGISTERS_reg[28][20]  ( .D(n2686), .CK(CLK), .RN(n1528), .Q(n4776), 
        .QN(n3817) );
  DFFR_X1 \REGISTERS_reg[28][19]  ( .D(n2685), .CK(CLK), .RN(n1529), .Q(n4775), 
        .QN(n3792) );
  DFFR_X1 \REGISTERS_reg[28][18]  ( .D(n2684), .CK(CLK), .RN(n1529), .Q(n4774), 
        .QN(n3767) );
  DFFR_X1 \REGISTERS_reg[28][17]  ( .D(n2683), .CK(CLK), .RN(n1529), .Q(n4773), 
        .QN(n3742) );
  DFFR_X1 \REGISTERS_reg[28][16]  ( .D(n2682), .CK(CLK), .RN(n1529), .Q(n4772), 
        .QN(n3717) );
  DFFR_X1 \REGISTERS_reg[28][15]  ( .D(n2681), .CK(CLK), .RN(n1529), .Q(n4771), 
        .QN(n3692) );
  DFFR_X1 \REGISTERS_reg[28][14]  ( .D(n2680), .CK(CLK), .RN(n1529), .Q(n4770), 
        .QN(n3667) );
  DFFR_X1 \REGISTERS_reg[28][13]  ( .D(n2679), .CK(CLK), .RN(n1529), .Q(n4769), 
        .QN(n3642) );
  DFFR_X1 \REGISTERS_reg[28][12]  ( .D(n2678), .CK(CLK), .RN(n1529), .Q(n4768), 
        .QN(n3617) );
  DFFR_X1 \REGISTERS_reg[28][11]  ( .D(n2677), .CK(CLK), .RN(n1529), .Q(n4767), 
        .QN(n3592) );
  DFFR_X1 \REGISTERS_reg[28][10]  ( .D(n2676), .CK(CLK), .RN(n1529), .Q(n4766), 
        .QN(n3567) );
  DFFR_X1 \REGISTERS_reg[28][9]  ( .D(n2675), .CK(CLK), .RN(n1529), .Q(n4765), 
        .QN(n2486) );
  DFFR_X1 \REGISTERS_reg[28][8]  ( .D(n2674), .CK(CLK), .RN(n1529), .Q(n4764), 
        .QN(n2461) );
  DFFR_X1 \REGISTERS_reg[28][7]  ( .D(n2673), .CK(CLK), .RN(n1530), .Q(n4763), 
        .QN(n2436) );
  DFFR_X1 \REGISTERS_reg[28][6]  ( .D(n2672), .CK(CLK), .RN(n1530), .Q(n4762), 
        .QN(n2411) );
  DFFR_X1 \REGISTERS_reg[28][5]  ( .D(n2671), .CK(CLK), .RN(n1530), .Q(n4761), 
        .QN(n2386) );
  DFFR_X1 \REGISTERS_reg[28][4]  ( .D(n2670), .CK(CLK), .RN(n1530), .Q(n4760), 
        .QN(n2361) );
  DFFR_X1 \REGISTERS_reg[28][3]  ( .D(n2669), .CK(CLK), .RN(n1530), .Q(n4759), 
        .QN(n2336) );
  DFFR_X1 \REGISTERS_reg[28][2]  ( .D(n2668), .CK(CLK), .RN(n1530), .Q(n4758), 
        .QN(n2311) );
  DFFR_X1 \REGISTERS_reg[28][1]  ( .D(n2667), .CK(CLK), .RN(n1530), .Q(n4757), 
        .QN(n2286) );
  DFFR_X1 \REGISTERS_reg[28][0]  ( .D(n2666), .CK(CLK), .RN(n1530), .Q(n4756), 
        .QN(n2257) );
  DFFR_X1 \REGISTERS_reg[29][31]  ( .D(n2665), .CK(CLK), .RN(n1530), .Q(n4755), 
        .QN(n321) );
  DFFR_X1 \REGISTERS_reg[29][30]  ( .D(n2664), .CK(CLK), .RN(n1530), .Q(n4754), 
        .QN(n320) );
  DFFR_X1 \REGISTERS_reg[29][29]  ( .D(n2663), .CK(CLK), .RN(n1530), .Q(n4753), 
        .QN(n319) );
  DFFR_X1 \REGISTERS_reg[29][28]  ( .D(n2662), .CK(CLK), .RN(n1530), .Q(n4752), 
        .QN(n318) );
  DFFR_X1 \REGISTERS_reg[29][27]  ( .D(n2661), .CK(CLK), .RN(n1531), .Q(n4751), 
        .QN(n317) );
  DFFR_X1 \REGISTERS_reg[29][26]  ( .D(n2660), .CK(CLK), .RN(n1531), .Q(n4750), 
        .QN(n316) );
  DFFR_X1 \REGISTERS_reg[29][25]  ( .D(n2659), .CK(CLK), .RN(n1531), .Q(n4749), 
        .QN(n315) );
  DFFR_X1 \REGISTERS_reg[29][24]  ( .D(n2658), .CK(CLK), .RN(n1531), .Q(n4748), 
        .QN(n314) );
  DFFR_X1 \REGISTERS_reg[29][23]  ( .D(n2657), .CK(CLK), .RN(n1531), .Q(n4747), 
        .QN(n313) );
  DFFR_X1 \REGISTERS_reg[29][22]  ( .D(n2656), .CK(CLK), .RN(n1531), .Q(n4746), 
        .QN(n312) );
  DFFR_X1 \REGISTERS_reg[29][21]  ( .D(n2655), .CK(CLK), .RN(n1531), .Q(n4745), 
        .QN(n311) );
  DFFR_X1 \REGISTERS_reg[29][20]  ( .D(n2654), .CK(CLK), .RN(n1531), .Q(n4744), 
        .QN(n310) );
  DFFR_X1 \REGISTERS_reg[29][19]  ( .D(n2653), .CK(CLK), .RN(n1531), .Q(n4743), 
        .QN(n309) );
  DFFR_X1 \REGISTERS_reg[29][18]  ( .D(n2652), .CK(CLK), .RN(n1531), .Q(n4742), 
        .QN(n308) );
  DFFR_X1 \REGISTERS_reg[29][17]  ( .D(n2651), .CK(CLK), .RN(n1531), .Q(n4741), 
        .QN(n307) );
  DFFR_X1 \REGISTERS_reg[29][16]  ( .D(n2650), .CK(CLK), .RN(n1531), .Q(n4740), 
        .QN(n306) );
  DFFR_X1 \REGISTERS_reg[29][15]  ( .D(n2649), .CK(CLK), .RN(n1532), .Q(n4739), 
        .QN(n305) );
  DFFR_X1 \REGISTERS_reg[29][14]  ( .D(n2648), .CK(CLK), .RN(n1532), .Q(n4738), 
        .QN(n304) );
  DFFR_X1 \REGISTERS_reg[29][13]  ( .D(n2647), .CK(CLK), .RN(n1532), .Q(n4737), 
        .QN(n303) );
  DFFR_X1 \REGISTERS_reg[29][12]  ( .D(n2646), .CK(CLK), .RN(n1532), .Q(n4736), 
        .QN(n461) );
  DFFR_X1 \REGISTERS_reg[29][11]  ( .D(n2645), .CK(CLK), .RN(n1532), .Q(n4735), 
        .QN(n302) );
  DFFR_X1 \REGISTERS_reg[29][10]  ( .D(n2644), .CK(CLK), .RN(n1532), .Q(n4734), 
        .QN(n301) );
  DFFR_X1 \REGISTERS_reg[29][9]  ( .D(n2643), .CK(CLK), .RN(n1532), .Q(n4733), 
        .QN(n300) );
  DFFR_X1 \REGISTERS_reg[29][8]  ( .D(n2642), .CK(CLK), .RN(n1532), .Q(n4732), 
        .QN(n299) );
  DFFR_X1 \REGISTERS_reg[29][7]  ( .D(n2641), .CK(CLK), .RN(n1532), .Q(n4731), 
        .QN(n298) );
  DFFR_X1 \REGISTERS_reg[29][6]  ( .D(n2640), .CK(CLK), .RN(n1532), .Q(n4730), 
        .QN(n297) );
  DFFR_X1 \REGISTERS_reg[29][5]  ( .D(n2639), .CK(CLK), .RN(n1532), .Q(n4729), 
        .QN(n296) );
  DFFR_X1 \REGISTERS_reg[29][4]  ( .D(n2638), .CK(CLK), .RN(n1532), .Q(n4728), 
        .QN(n295) );
  DFFR_X1 \REGISTERS_reg[29][3]  ( .D(n2637), .CK(CLK), .RN(n1533), .Q(n4727), 
        .QN(n294) );
  DFFR_X1 \REGISTERS_reg[29][2]  ( .D(n2636), .CK(CLK), .RN(n1533), .Q(n4726), 
        .QN(n293) );
  DFFR_X1 \REGISTERS_reg[29][1]  ( .D(n2635), .CK(CLK), .RN(n1533), .Q(n4725), 
        .QN(n228) );
  DFFR_X1 \REGISTERS_reg[29][0]  ( .D(n2634), .CK(CLK), .RN(n1533), .Q(n4724), 
        .QN(n227) );
  DFFR_X1 \REGISTERS_reg[30][23]  ( .D(n2625), .CK(CLK), .RN(n1534), .QN(n941)
         );
  DFFR_X1 \REGISTERS_reg[30][22]  ( .D(n2624), .CK(CLK), .RN(n1534), .QN(n942)
         );
  DFFR_X1 \REGISTERS_reg[30][21]  ( .D(n2623), .CK(CLK), .RN(n1534), .QN(n943)
         );
  DFFR_X1 \REGISTERS_reg[30][20]  ( .D(n2622), .CK(CLK), .RN(n1534), .QN(n944)
         );
  DFFR_X1 \REGISTERS_reg[30][19]  ( .D(n2621), .CK(CLK), .RN(n1534), .QN(n945)
         );
  DFFR_X1 \REGISTERS_reg[30][18]  ( .D(n2620), .CK(CLK), .RN(n1534), .QN(n946)
         );
  DFFR_X1 \REGISTERS_reg[30][17]  ( .D(n2619), .CK(CLK), .RN(n1534), .QN(n947)
         );
  DFFR_X1 \REGISTERS_reg[30][16]  ( .D(n2618), .CK(CLK), .RN(n1534), .QN(n948)
         );
  DFFR_X1 \REGISTERS_reg[30][15]  ( .D(n2617), .CK(CLK), .RN(n1534), .QN(n949)
         );
  DFFR_X1 \REGISTERS_reg[30][14]  ( .D(n2616), .CK(CLK), .RN(n1534), .QN(n950)
         );
  DFFR_X1 \REGISTERS_reg[30][13]  ( .D(n2615), .CK(CLK), .RN(n1534), .QN(n951)
         );
  DFFR_X1 \REGISTERS_reg[30][12]  ( .D(n2614), .CK(CLK), .RN(n1534), .QN(n952)
         );
  DFFR_X1 \REGISTERS_reg[30][11]  ( .D(n2613), .CK(CLK), .RN(n1535), .QN(n953)
         );
  DFFR_X1 \REGISTERS_reg[30][10]  ( .D(n2612), .CK(CLK), .RN(n1535), .QN(n954)
         );
  DFFR_X1 \REGISTERS_reg[30][9]  ( .D(n2611), .CK(CLK), .RN(n1535), .QN(n955)
         );
  DFFR_X1 \REGISTERS_reg[30][8]  ( .D(n2610), .CK(CLK), .RN(n1535), .QN(n956)
         );
  DFFR_X1 \REGISTERS_reg[30][7]  ( .D(n2609), .CK(CLK), .RN(n1535), .QN(n957)
         );
  DFFR_X1 \REGISTERS_reg[30][6]  ( .D(n2608), .CK(CLK), .RN(n1535), .QN(n958)
         );
  DFFR_X1 \REGISTERS_reg[30][5]  ( .D(n2607), .CK(CLK), .RN(n1535), .QN(n959)
         );
  DFFR_X1 \REGISTERS_reg[30][4]  ( .D(n2606), .CK(CLK), .RN(n1535), .QN(n960)
         );
  DFFR_X1 \REGISTERS_reg[30][3]  ( .D(n2605), .CK(CLK), .RN(n1535), .QN(n961)
         );
  DFFR_X1 \REGISTERS_reg[30][2]  ( .D(n2604), .CK(CLK), .RN(n1535), .QN(n962)
         );
  DFFR_X1 \REGISTERS_reg[30][1]  ( .D(n2603), .CK(CLK), .RN(n1535), .QN(n963)
         );
  DFFR_X1 \REGISTERS_reg[30][0]  ( .D(n2602), .CK(CLK), .RN(n1535), .QN(n964)
         );
  DFFR_X1 \REGISTERS_reg[31][23]  ( .D(n2593), .CK(CLK), .RN(n1536), .Q(n4316)
         );
  DFFR_X1 \REGISTERS_reg[31][22]  ( .D(n2592), .CK(CLK), .RN(n1536), .Q(n4317)
         );
  DFFR_X1 \REGISTERS_reg[31][21]  ( .D(n2591), .CK(CLK), .RN(n1536), .Q(n4318)
         );
  DFFR_X1 \REGISTERS_reg[31][20]  ( .D(n2590), .CK(CLK), .RN(n1536), .Q(n4319)
         );
  DFFR_X1 \REGISTERS_reg[31][19]  ( .D(n2589), .CK(CLK), .RN(n1537), .Q(n4320)
         );
  DFFR_X1 \REGISTERS_reg[31][18]  ( .D(n2588), .CK(CLK), .RN(n1537), .Q(n4321)
         );
  DFFR_X1 \REGISTERS_reg[31][17]  ( .D(n2587), .CK(CLK), .RN(n1537), .Q(n4322)
         );
  DFFR_X1 \REGISTERS_reg[31][16]  ( .D(n2586), .CK(CLK), .RN(n1537), .Q(n4323)
         );
  DFFR_X1 \REGISTERS_reg[31][15]  ( .D(n2585), .CK(CLK), .RN(n1537), .Q(n4324)
         );
  DFFR_X1 \REGISTERS_reg[31][14]  ( .D(n2584), .CK(CLK), .RN(n1537), .Q(n4325)
         );
  DFFR_X1 \REGISTERS_reg[31][13]  ( .D(n2583), .CK(CLK), .RN(n1537), .Q(n4326)
         );
  DFFR_X1 \REGISTERS_reg[31][12]  ( .D(n2582), .CK(CLK), .RN(n1537), .Q(n4327)
         );
  DFFR_X1 \REGISTERS_reg[31][11]  ( .D(n2581), .CK(CLK), .RN(n1537), .Q(n4328)
         );
  DFFR_X1 \REGISTERS_reg[31][10]  ( .D(n2580), .CK(CLK), .RN(n1537), .Q(n4329)
         );
  DFFR_X1 \REGISTERS_reg[31][9]  ( .D(n2579), .CK(CLK), .RN(n1537), .Q(n4330)
         );
  DFFR_X1 \REGISTERS_reg[31][8]  ( .D(n2578), .CK(CLK), .RN(n1537), .Q(n4331)
         );
  DFFR_X1 \REGISTERS_reg[31][7]  ( .D(n2577), .CK(CLK), .RN(n1538), .Q(n4332)
         );
  DFFR_X1 \REGISTERS_reg[31][6]  ( .D(n2576), .CK(CLK), .RN(n1538), .Q(n4333)
         );
  DFFR_X1 \REGISTERS_reg[31][5]  ( .D(n2575), .CK(CLK), .RN(n1538), .Q(n4334)
         );
  DFFR_X1 \REGISTERS_reg[31][4]  ( .D(n2574), .CK(CLK), .RN(n1538), .Q(n4335)
         );
  DFFR_X1 \REGISTERS_reg[31][3]  ( .D(n2573), .CK(CLK), .RN(n1538), .Q(n4336)
         );
  DFFR_X1 \REGISTERS_reg[31][2]  ( .D(n2572), .CK(CLK), .RN(n1538), .Q(n4337)
         );
  DFFR_X1 \REGISTERS_reg[31][1]  ( .D(n2571), .CK(CLK), .RN(n1538), .Q(n4338)
         );
  DFFR_X1 \REGISTERS_reg[31][0]  ( .D(n2570), .CK(CLK), .RN(n1538), .Q(n4339)
         );
  DFF_X1 \OUT2_reg[31]  ( .D(n2569), .CK(CLK), .Q(OUT2[31]), .QN(n4723) );
  DFF_X1 \OUT2_reg[30]  ( .D(n2568), .CK(CLK), .Q(OUT2[30]), .QN(n4722) );
  DFF_X1 \OUT2_reg[29]  ( .D(n2567), .CK(CLK), .Q(OUT2[29]), .QN(n4721) );
  DFF_X1 \OUT2_reg[28]  ( .D(n2566), .CK(CLK), .Q(OUT2[28]), .QN(n4720) );
  DFF_X1 \OUT2_reg[27]  ( .D(n2565), .CK(CLK), .Q(OUT2[27]), .QN(n4719) );
  DFF_X1 \OUT2_reg[26]  ( .D(n2564), .CK(CLK), .Q(OUT2[26]), .QN(n4718) );
  DFF_X1 \OUT2_reg[25]  ( .D(n2563), .CK(CLK), .Q(OUT2[25]), .QN(n4717) );
  DFF_X1 \OUT2_reg[24]  ( .D(n2562), .CK(CLK), .Q(OUT2[24]), .QN(n4716) );
  DFF_X1 \OUT2_reg[23]  ( .D(n2561), .CK(CLK), .Q(OUT2[23]), .QN(n4715) );
  DFF_X1 \OUT2_reg[22]  ( .D(n2560), .CK(CLK), .Q(OUT2[22]), .QN(n4714) );
  DFF_X1 \OUT2_reg[21]  ( .D(n2559), .CK(CLK), .Q(OUT2[21]), .QN(n4713) );
  DFF_X1 \OUT2_reg[20]  ( .D(n2558), .CK(CLK), .Q(OUT2[20]), .QN(n4712) );
  DFF_X1 \OUT2_reg[19]  ( .D(n2557), .CK(CLK), .Q(OUT2[19]), .QN(n4711) );
  DFF_X1 \OUT2_reg[18]  ( .D(n2556), .CK(CLK), .Q(OUT2[18]), .QN(n4710) );
  DFF_X1 \OUT2_reg[17]  ( .D(n2555), .CK(CLK), .Q(OUT2[17]), .QN(n4709) );
  DFF_X1 \OUT2_reg[16]  ( .D(n2554), .CK(CLK), .Q(OUT2[16]), .QN(n4708) );
  DFF_X1 \OUT2_reg[15]  ( .D(n2553), .CK(CLK), .Q(OUT2[15]), .QN(n4707) );
  DFF_X1 \OUT2_reg[14]  ( .D(n2552), .CK(CLK), .Q(OUT2[14]), .QN(n4706) );
  DFF_X1 \OUT2_reg[13]  ( .D(n2551), .CK(CLK), .Q(OUT2[13]), .QN(n4705) );
  DFF_X1 \OUT2_reg[12]  ( .D(n2550), .CK(CLK), .Q(OUT2[12]), .QN(n4704) );
  DFF_X1 \OUT2_reg[11]  ( .D(n2549), .CK(CLK), .Q(OUT2[11]), .QN(n4703) );
  DFF_X1 \OUT2_reg[10]  ( .D(n2548), .CK(CLK), .Q(OUT2[10]), .QN(n4702) );
  DFF_X1 \OUT2_reg[9]  ( .D(n2547), .CK(CLK), .Q(OUT2[9]), .QN(n4701) );
  DFF_X1 \OUT2_reg[8]  ( .D(n2546), .CK(CLK), .Q(OUT2[8]), .QN(n4700) );
  DFF_X1 \OUT2_reg[7]  ( .D(n2545), .CK(CLK), .Q(OUT2[7]), .QN(n4699) );
  DFF_X1 \OUT2_reg[6]  ( .D(n2544), .CK(CLK), .Q(OUT2[6]), .QN(n4698) );
  DFF_X1 \OUT2_reg[5]  ( .D(n2543), .CK(CLK), .Q(OUT2[5]), .QN(n4697) );
  DFF_X1 \OUT2_reg[4]  ( .D(n2542), .CK(CLK), .Q(OUT2[4]), .QN(n4696) );
  DFF_X1 \OUT2_reg[3]  ( .D(n2541), .CK(CLK), .Q(OUT2[3]), .QN(n4695) );
  DFF_X1 \OUT2_reg[2]  ( .D(n2540), .CK(CLK), .Q(OUT2[2]), .QN(n4694) );
  DFF_X1 \OUT2_reg[1]  ( .D(n2539), .CK(CLK), .Q(OUT2[1]), .QN(n4693) );
  DFF_X1 \OUT2_reg[0]  ( .D(n2538), .CK(CLK), .Q(OUT2[0]), .QN(n4692) );
  DFF_X1 \OUT1_reg[31]  ( .D(n2537), .CK(CLK), .Q(OUT1[31]), .QN(n4691) );
  DFF_X1 \OUT1_reg[30]  ( .D(n2536), .CK(CLK), .Q(OUT1[30]), .QN(n4690) );
  DFF_X1 \OUT1_reg[29]  ( .D(n2535), .CK(CLK), .Q(OUT1[29]), .QN(n4689) );
  DFF_X1 \OUT1_reg[28]  ( .D(n2534), .CK(CLK), .Q(OUT1[28]), .QN(n4688) );
  DFF_X1 \OUT1_reg[27]  ( .D(n2533), .CK(CLK), .Q(OUT1[27]), .QN(n4687) );
  DFF_X1 \OUT1_reg[26]  ( .D(n2532), .CK(CLK), .Q(OUT1[26]), .QN(n4686) );
  DFF_X1 \OUT1_reg[25]  ( .D(n2531), .CK(CLK), .Q(OUT1[25]), .QN(n4685) );
  DFF_X1 \OUT1_reg[24]  ( .D(n2530), .CK(CLK), .Q(OUT1[24]), .QN(n4684) );
  DFF_X1 \OUT1_reg[23]  ( .D(n2529), .CK(CLK), .Q(OUT1[23]), .QN(n4683) );
  DFF_X1 \OUT1_reg[22]  ( .D(n2528), .CK(CLK), .Q(OUT1[22]), .QN(n4682) );
  DFF_X1 \OUT1_reg[21]  ( .D(n2527), .CK(CLK), .Q(OUT1[21]), .QN(n4681) );
  DFF_X1 \OUT1_reg[20]  ( .D(n2526), .CK(CLK), .Q(OUT1[20]), .QN(n4680) );
  DFF_X1 \OUT1_reg[19]  ( .D(n2525), .CK(CLK), .Q(OUT1[19]), .QN(n4679) );
  DFF_X1 \OUT1_reg[18]  ( .D(n2524), .CK(CLK), .Q(OUT1[18]), .QN(n4678) );
  DFF_X1 \OUT1_reg[17]  ( .D(n2523), .CK(CLK), .Q(OUT1[17]), .QN(n4677) );
  DFF_X1 \OUT1_reg[16]  ( .D(n2522), .CK(CLK), .Q(OUT1[16]), .QN(n4676) );
  DFF_X1 \OUT1_reg[15]  ( .D(n2521), .CK(CLK), .Q(OUT1[15]), .QN(n4675) );
  DFF_X1 \OUT1_reg[14]  ( .D(n2520), .CK(CLK), .Q(OUT1[14]), .QN(n4674) );
  DFF_X1 \OUT1_reg[13]  ( .D(n2519), .CK(CLK), .Q(OUT1[13]), .QN(n4673) );
  DFF_X1 \OUT1_reg[12]  ( .D(n2518), .CK(CLK), .Q(OUT1[12]), .QN(n4672) );
  DFF_X1 \OUT1_reg[11]  ( .D(n2517), .CK(CLK), .Q(OUT1[11]), .QN(n4671) );
  DFF_X1 \OUT1_reg[10]  ( .D(n2516), .CK(CLK), .Q(OUT1[10]), .QN(n4670) );
  DFF_X1 \OUT1_reg[9]  ( .D(n2515), .CK(CLK), .Q(OUT1[9]), .QN(n4669) );
  DFF_X1 \OUT1_reg[8]  ( .D(n2514), .CK(CLK), .Q(OUT1[8]), .QN(n4668) );
  DFF_X1 \OUT1_reg[7]  ( .D(n2513), .CK(CLK), .Q(OUT1[7]), .QN(n4667) );
  DFF_X1 \OUT1_reg[6]  ( .D(n2512), .CK(CLK), .Q(OUT1[6]), .QN(n4666) );
  DFF_X1 \OUT1_reg[5]  ( .D(n2511), .CK(CLK), .Q(OUT1[5]), .QN(n4665) );
  DFF_X1 \OUT1_reg[4]  ( .D(n2510), .CK(CLK), .Q(OUT1[4]), .QN(n4664) );
  DFF_X1 \OUT1_reg[3]  ( .D(n2509), .CK(CLK), .Q(OUT1[3]), .QN(n4663) );
  DFF_X1 \OUT1_reg[2]  ( .D(n2508), .CK(CLK), .Q(OUT1[2]), .QN(n4662) );
  DFF_X1 \OUT1_reg[0]  ( .D(n2506), .CK(CLK), .Q(OUT1[0]), .QN(n4660) );
  DFFR_X1 \REGISTERS_reg[8][21]  ( .D(n3327), .CK(CLK), .RN(n1475), .QN(n239)
         );
  DFFR_X1 \REGISTERS_reg[5][31]  ( .D(n3433), .CK(CLK), .RN(n1466), .Q(n4192), 
        .QN(n133) );
  DFFR_X1 \REGISTERS_reg[5][30]  ( .D(n3432), .CK(CLK), .RN(n1466), .Q(n4193), 
        .QN(n134) );
  DFFR_X1 \REGISTERS_reg[5][29]  ( .D(n3431), .CK(CLK), .RN(n1466), .Q(n4194), 
        .QN(n135) );
  DFFR_X1 \REGISTERS_reg[5][28]  ( .D(n3430), .CK(CLK), .RN(n1466), .Q(n4195), 
        .QN(n136) );
  DFFR_X1 \REGISTERS_reg[5][27]  ( .D(n3429), .CK(CLK), .RN(n1467), .Q(n4196), 
        .QN(n137) );
  DFFR_X1 \REGISTERS_reg[5][26]  ( .D(n3428), .CK(CLK), .RN(n1467), .Q(n4197), 
        .QN(n138) );
  DFFR_X1 \REGISTERS_reg[5][25]  ( .D(n3427), .CK(CLK), .RN(n1467), .Q(n4198), 
        .QN(n139) );
  DFFR_X1 \REGISTERS_reg[5][24]  ( .D(n3426), .CK(CLK), .RN(n1467), .Q(n4199), 
        .QN(n140) );
  DFFR_X1 \REGISTERS_reg[4][31]  ( .D(n3465), .CK(CLK), .RN(n1464), .Q(n4160), 
        .QN(n101) );
  DFFR_X1 \REGISTERS_reg[4][30]  ( .D(n3464), .CK(CLK), .RN(n1464), .Q(n4161), 
        .QN(n102) );
  DFFR_X1 \REGISTERS_reg[4][29]  ( .D(n3463), .CK(CLK), .RN(n1464), .Q(n4162), 
        .QN(n103) );
  DFFR_X1 \REGISTERS_reg[4][28]  ( .D(n3462), .CK(CLK), .RN(n1464), .Q(n4163), 
        .QN(n104) );
  DFFR_X1 \REGISTERS_reg[4][27]  ( .D(n3461), .CK(CLK), .RN(n1464), .Q(n4164), 
        .QN(n105) );
  DFFR_X1 \REGISTERS_reg[4][26]  ( .D(n3460), .CK(CLK), .RN(n1464), .Q(n4165), 
        .QN(n106) );
  DFFR_X1 \REGISTERS_reg[4][25]  ( .D(n3459), .CK(CLK), .RN(n1464), .Q(n4166), 
        .QN(n107) );
  DFFR_X1 \REGISTERS_reg[4][24]  ( .D(n3458), .CK(CLK), .RN(n1464), .Q(n4167), 
        .QN(n108) );
  DFFR_X1 \REGISTERS_reg[1][31]  ( .D(n3561), .CK(CLK), .RN(n1456), .Q(n4128)
         );
  DFFR_X1 \REGISTERS_reg[1][30]  ( .D(n3560), .CK(CLK), .RN(n1456), .Q(n4129)
         );
  DFFR_X1 \REGISTERS_reg[1][29]  ( .D(n3559), .CK(CLK), .RN(n1456), .Q(n4130)
         );
  DFFR_X1 \REGISTERS_reg[1][28]  ( .D(n3558), .CK(CLK), .RN(n1456), .Q(n4131)
         );
  DFFR_X1 \REGISTERS_reg[1][27]  ( .D(n3557), .CK(CLK), .RN(n1456), .Q(n4132)
         );
  DFFR_X1 \REGISTERS_reg[1][26]  ( .D(n3556), .CK(CLK), .RN(n1456), .Q(n4133)
         );
  DFFR_X1 \REGISTERS_reg[1][25]  ( .D(n3555), .CK(CLK), .RN(n1456), .Q(n4134)
         );
  DFFR_X1 \REGISTERS_reg[1][24]  ( .D(n3554), .CK(CLK), .RN(n1456), .Q(n4135)
         );
  DFFR_X1 \REGISTERS_reg[21][31]  ( .D(n2921), .CK(CLK), .RN(n1509), .Q(n4256)
         );
  DFFR_X1 \REGISTERS_reg[21][30]  ( .D(n2920), .CK(CLK), .RN(n1509), .Q(n4257)
         );
  DFFR_X1 \REGISTERS_reg[21][29]  ( .D(n2919), .CK(CLK), .RN(n1509), .Q(n4258)
         );
  DFFR_X1 \REGISTERS_reg[21][28]  ( .D(n2918), .CK(CLK), .RN(n1509), .Q(n4259)
         );
  DFFR_X1 \REGISTERS_reg[21][27]  ( .D(n2917), .CK(CLK), .RN(n1509), .Q(n4260)
         );
  DFFR_X1 \REGISTERS_reg[21][26]  ( .D(n2916), .CK(CLK), .RN(n1509), .Q(n4261)
         );
  DFFR_X1 \REGISTERS_reg[21][25]  ( .D(n2915), .CK(CLK), .RN(n1509), .Q(n4262)
         );
  DFFR_X1 \REGISTERS_reg[21][24]  ( .D(n2914), .CK(CLK), .RN(n1509), .Q(n4263)
         );
  DFFR_X1 \REGISTERS_reg[16][31]  ( .D(n3081), .CK(CLK), .RN(n1496), .Q(n4224)
         );
  DFFR_X1 \REGISTERS_reg[16][30]  ( .D(n3080), .CK(CLK), .RN(n1496), .Q(n4225)
         );
  DFFR_X1 \REGISTERS_reg[16][29]  ( .D(n3079), .CK(CLK), .RN(n1496), .Q(n4226)
         );
  DFFR_X1 \REGISTERS_reg[16][28]  ( .D(n3078), .CK(CLK), .RN(n1496), .Q(n4227)
         );
  DFFR_X1 \REGISTERS_reg[16][27]  ( .D(n3077), .CK(CLK), .RN(n1496), .Q(n4228)
         );
  DFFR_X1 \REGISTERS_reg[16][26]  ( .D(n3076), .CK(CLK), .RN(n1496), .Q(n4229)
         );
  DFFR_X1 \REGISTERS_reg[16][25]  ( .D(n3075), .CK(CLK), .RN(n1496), .Q(n4230)
         );
  DFFR_X1 \REGISTERS_reg[16][24]  ( .D(n3074), .CK(CLK), .RN(n1496), .Q(n4231)
         );
  DFFR_X1 \REGISTERS_reg[31][31]  ( .D(n2601), .CK(CLK), .RN(n1536), .Q(n4308)
         );
  DFFR_X1 \REGISTERS_reg[31][30]  ( .D(n2600), .CK(CLK), .RN(n1536), .Q(n4309)
         );
  DFFR_X1 \REGISTERS_reg[31][29]  ( .D(n2599), .CK(CLK), .RN(n1536), .Q(n4310)
         );
  DFFR_X1 \REGISTERS_reg[31][28]  ( .D(n2598), .CK(CLK), .RN(n1536), .Q(n4311)
         );
  DFFR_X1 \REGISTERS_reg[31][27]  ( .D(n2597), .CK(CLK), .RN(n1536), .Q(n4312)
         );
  DFFR_X1 \REGISTERS_reg[31][26]  ( .D(n2596), .CK(CLK), .RN(n1536), .Q(n4313)
         );
  DFFR_X1 \REGISTERS_reg[31][25]  ( .D(n2595), .CK(CLK), .RN(n1536), .Q(n4314)
         );
  DFFR_X1 \REGISTERS_reg[31][24]  ( .D(n2594), .CK(CLK), .RN(n1536), .Q(n4315)
         );
  DFFR_X1 \REGISTERS_reg[26][31]  ( .D(n2761), .CK(CLK), .RN(n1522), .Q(n4288), 
        .QN(n805) );
  DFFR_X1 \REGISTERS_reg[26][30]  ( .D(n2760), .CK(CLK), .RN(n1522), .Q(n4289), 
        .QN(n806) );
  DFFR_X1 \REGISTERS_reg[26][29]  ( .D(n2759), .CK(CLK), .RN(n1522), .Q(n4290), 
        .QN(n807) );
  DFFR_X1 \REGISTERS_reg[26][28]  ( .D(n2758), .CK(CLK), .RN(n1522), .Q(n4291), 
        .QN(n808) );
  DFFR_X1 \REGISTERS_reg[26][27]  ( .D(n2757), .CK(CLK), .RN(n1523), .Q(n4292), 
        .QN(n809) );
  DFFR_X1 \REGISTERS_reg[26][26]  ( .D(n2756), .CK(CLK), .RN(n1523), .Q(n4293), 
        .QN(n810) );
  DFFR_X1 \REGISTERS_reg[26][25]  ( .D(n2755), .CK(CLK), .RN(n1523), .Q(n4294), 
        .QN(n811) );
  DFFR_X1 \REGISTERS_reg[26][24]  ( .D(n2754), .CK(CLK), .RN(n1523), .Q(n4295), 
        .QN(n812) );
  DFFR_X1 \REGISTERS_reg[5][23]  ( .D(n3425), .CK(CLK), .RN(n1467), .Q(n4200), 
        .QN(n141) );
  DFFR_X1 \REGISTERS_reg[5][22]  ( .D(n3424), .CK(CLK), .RN(n1467), .Q(n4201), 
        .QN(n142) );
  DFFR_X1 \REGISTERS_reg[5][21]  ( .D(n3423), .CK(CLK), .RN(n1467), .Q(n4202), 
        .QN(n143) );
  DFFR_X1 \REGISTERS_reg[5][20]  ( .D(n3422), .CK(CLK), .RN(n1467), .Q(n4203), 
        .QN(n144) );
  DFFR_X1 \REGISTERS_reg[5][19]  ( .D(n3421), .CK(CLK), .RN(n1467), .Q(n4204), 
        .QN(n145) );
  DFFR_X1 \REGISTERS_reg[5][18]  ( .D(n3420), .CK(CLK), .RN(n1467), .Q(n4205), 
        .QN(n146) );
  DFFR_X1 \REGISTERS_reg[5][17]  ( .D(n3419), .CK(CLK), .RN(n1467), .Q(n4206), 
        .QN(n147) );
  DFFR_X1 \REGISTERS_reg[5][16]  ( .D(n3418), .CK(CLK), .RN(n1467), .Q(n4207), 
        .QN(n148) );
  DFFR_X1 \REGISTERS_reg[5][15]  ( .D(n3417), .CK(CLK), .RN(n1468), .Q(n4208), 
        .QN(n149) );
  DFFR_X1 \REGISTERS_reg[5][14]  ( .D(n3416), .CK(CLK), .RN(n1468), .Q(n4209), 
        .QN(n150) );
  DFFR_X1 \REGISTERS_reg[5][13]  ( .D(n3415), .CK(CLK), .RN(n1468), .Q(n4210), 
        .QN(n151) );
  DFFR_X1 \REGISTERS_reg[5][12]  ( .D(n3414), .CK(CLK), .RN(n1468), .Q(n4211), 
        .QN(n152) );
  DFFR_X1 \REGISTERS_reg[5][11]  ( .D(n3413), .CK(CLK), .RN(n1468), .Q(n4212), 
        .QN(n153) );
  DFFR_X1 \REGISTERS_reg[5][10]  ( .D(n3412), .CK(CLK), .RN(n1468), .Q(n4213), 
        .QN(n154) );
  DFFR_X1 \REGISTERS_reg[5][9]  ( .D(n3411), .CK(CLK), .RN(n1468), .Q(n4214), 
        .QN(n155) );
  DFFR_X1 \REGISTERS_reg[5][8]  ( .D(n3410), .CK(CLK), .RN(n1468), .Q(n4215), 
        .QN(n156) );
  DFFR_X1 \REGISTERS_reg[5][7]  ( .D(n3409), .CK(CLK), .RN(n1468), .Q(n4216), 
        .QN(n157) );
  DFFR_X1 \REGISTERS_reg[5][6]  ( .D(n3408), .CK(CLK), .RN(n1468), .Q(n4217), 
        .QN(n158) );
  DFFR_X1 \REGISTERS_reg[5][5]  ( .D(n3407), .CK(CLK), .RN(n1468), .Q(n4218), 
        .QN(n159) );
  DFFR_X1 \REGISTERS_reg[5][4]  ( .D(n3406), .CK(CLK), .RN(n1468), .Q(n4219), 
        .QN(n160) );
  DFFR_X1 \REGISTERS_reg[5][3]  ( .D(n3405), .CK(CLK), .RN(n1469), .Q(n4220), 
        .QN(n161) );
  DFFR_X1 \REGISTERS_reg[5][2]  ( .D(n3404), .CK(CLK), .RN(n1469), .Q(n4221), 
        .QN(n162) );
  DFFR_X1 \REGISTERS_reg[5][1]  ( .D(n3403), .CK(CLK), .RN(n1469), .Q(n4222), 
        .QN(n163) );
  DFFR_X1 \REGISTERS_reg[5][0]  ( .D(n3402), .CK(CLK), .RN(n1469), .Q(n4223), 
        .QN(n164) );
  DFFR_X1 \REGISTERS_reg[4][23]  ( .D(n3457), .CK(CLK), .RN(n1464), .Q(n4168), 
        .QN(n109) );
  DFFR_X1 \REGISTERS_reg[4][22]  ( .D(n3456), .CK(CLK), .RN(n1464), .Q(n4169), 
        .QN(n110) );
  DFFR_X1 \REGISTERS_reg[4][21]  ( .D(n3455), .CK(CLK), .RN(n1464), .Q(n4170), 
        .QN(n111) );
  DFFR_X1 \REGISTERS_reg[4][20]  ( .D(n3454), .CK(CLK), .RN(n1464), .Q(n4171), 
        .QN(n112) );
  DFFR_X1 \REGISTERS_reg[4][19]  ( .D(n3453), .CK(CLK), .RN(n1465), .Q(n4172), 
        .QN(n113) );
  DFFR_X1 \REGISTERS_reg[4][18]  ( .D(n3452), .CK(CLK), .RN(n1465), .Q(n4173), 
        .QN(n114) );
  DFFR_X1 \REGISTERS_reg[4][17]  ( .D(n3451), .CK(CLK), .RN(n1465), .Q(n4174), 
        .QN(n115) );
  DFFR_X1 \REGISTERS_reg[4][16]  ( .D(n3450), .CK(CLK), .RN(n1465), .Q(n4175), 
        .QN(n116) );
  DFFR_X1 \REGISTERS_reg[4][15]  ( .D(n3449), .CK(CLK), .RN(n1465), .Q(n4176), 
        .QN(n117) );
  DFFR_X1 \REGISTERS_reg[4][14]  ( .D(n3448), .CK(CLK), .RN(n1465), .Q(n4177), 
        .QN(n118) );
  DFFR_X1 \REGISTERS_reg[4][13]  ( .D(n3447), .CK(CLK), .RN(n1465), .Q(n4178), 
        .QN(n119) );
  DFFR_X1 \REGISTERS_reg[4][12]  ( .D(n3446), .CK(CLK), .RN(n1465), .Q(n4179), 
        .QN(n120) );
  DFFR_X1 \REGISTERS_reg[4][11]  ( .D(n3445), .CK(CLK), .RN(n1465), .Q(n4180), 
        .QN(n121) );
  DFFR_X1 \REGISTERS_reg[4][10]  ( .D(n3444), .CK(CLK), .RN(n1465), .Q(n4181), 
        .QN(n122) );
  DFFR_X1 \REGISTERS_reg[4][9]  ( .D(n3443), .CK(CLK), .RN(n1465), .Q(n4182), 
        .QN(n123) );
  DFFR_X1 \REGISTERS_reg[4][8]  ( .D(n3442), .CK(CLK), .RN(n1465), .Q(n4183), 
        .QN(n124) );
  DFFR_X1 \REGISTERS_reg[4][7]  ( .D(n3441), .CK(CLK), .RN(n1466), .Q(n4184), 
        .QN(n125) );
  DFFR_X1 \REGISTERS_reg[4][6]  ( .D(n3440), .CK(CLK), .RN(n1466), .Q(n4185), 
        .QN(n126) );
  DFFR_X1 \REGISTERS_reg[4][5]  ( .D(n3439), .CK(CLK), .RN(n1466), .Q(n4186), 
        .QN(n127) );
  DFFR_X1 \REGISTERS_reg[4][4]  ( .D(n3438), .CK(CLK), .RN(n1466), .Q(n4187), 
        .QN(n128) );
  DFFR_X1 \REGISTERS_reg[4][3]  ( .D(n3437), .CK(CLK), .RN(n1466), .Q(n4188), 
        .QN(n129) );
  DFFR_X1 \REGISTERS_reg[4][2]  ( .D(n3436), .CK(CLK), .RN(n1466), .Q(n4189), 
        .QN(n130) );
  DFFR_X1 \REGISTERS_reg[4][1]  ( .D(n3435), .CK(CLK), .RN(n1466), .Q(n4190), 
        .QN(n131) );
  DFFR_X1 \REGISTERS_reg[4][0]  ( .D(n3434), .CK(CLK), .RN(n1466), .Q(n4191), 
        .QN(n132) );
  DFFR_X1 \REGISTERS_reg[1][23]  ( .D(n3553), .CK(CLK), .RN(n1456), .Q(n4136)
         );
  DFFR_X1 \REGISTERS_reg[1][22]  ( .D(n3552), .CK(CLK), .RN(n1456), .Q(n4137)
         );
  DFFR_X1 \REGISTERS_reg[1][21]  ( .D(n3551), .CK(CLK), .RN(n1456), .Q(n4138)
         );
  DFFR_X1 \REGISTERS_reg[1][20]  ( .D(n3550), .CK(CLK), .RN(n1456), .Q(n4139)
         );
  DFFR_X1 \REGISTERS_reg[1][19]  ( .D(n3549), .CK(CLK), .RN(n1457), .Q(n4140)
         );
  DFFR_X1 \REGISTERS_reg[1][18]  ( .D(n3548), .CK(CLK), .RN(n1457), .Q(n4141)
         );
  DFFR_X1 \REGISTERS_reg[1][17]  ( .D(n3547), .CK(CLK), .RN(n1457), .Q(n4142)
         );
  DFFR_X1 \REGISTERS_reg[1][16]  ( .D(n3546), .CK(CLK), .RN(n1457), .Q(n4143)
         );
  DFFR_X1 \REGISTERS_reg[1][15]  ( .D(n3545), .CK(CLK), .RN(n1457), .Q(n4144)
         );
  DFFR_X1 \REGISTERS_reg[1][14]  ( .D(n3544), .CK(CLK), .RN(n1457), .Q(n4145)
         );
  DFFR_X1 \REGISTERS_reg[1][13]  ( .D(n3543), .CK(CLK), .RN(n1457), .Q(n4146)
         );
  DFFR_X1 \REGISTERS_reg[1][12]  ( .D(n3542), .CK(CLK), .RN(n1457), .Q(n4147)
         );
  DFFR_X1 \REGISTERS_reg[1][11]  ( .D(n3541), .CK(CLK), .RN(n1457), .Q(n4148)
         );
  DFFR_X1 \REGISTERS_reg[1][10]  ( .D(n3540), .CK(CLK), .RN(n1457), .Q(n4149)
         );
  DFFR_X1 \REGISTERS_reg[1][9]  ( .D(n3539), .CK(CLK), .RN(n1457), .Q(n4150)
         );
  DFFR_X1 \REGISTERS_reg[1][8]  ( .D(n3538), .CK(CLK), .RN(n1457), .Q(n4151)
         );
  DFFR_X1 \REGISTERS_reg[1][7]  ( .D(n3537), .CK(CLK), .RN(n1458), .Q(n4152)
         );
  DFFR_X1 \REGISTERS_reg[1][6]  ( .D(n3536), .CK(CLK), .RN(n1458), .Q(n4153)
         );
  DFFR_X1 \REGISTERS_reg[1][5]  ( .D(n3535), .CK(CLK), .RN(n1458), .Q(n4154)
         );
  DFFR_X1 \REGISTERS_reg[1][4]  ( .D(n3534), .CK(CLK), .RN(n1458), .Q(n4155)
         );
  DFFR_X1 \REGISTERS_reg[1][3]  ( .D(n3533), .CK(CLK), .RN(n1458), .Q(n4156)
         );
  DFFR_X1 \REGISTERS_reg[1][2]  ( .D(n3532), .CK(CLK), .RN(n1458), .Q(n4157)
         );
  DFFR_X1 \REGISTERS_reg[1][1]  ( .D(n3531), .CK(CLK), .RN(n1458), .Q(n4158)
         );
  DFFR_X1 \REGISTERS_reg[1][0]  ( .D(n3530), .CK(CLK), .RN(n1458), .Q(n4159)
         );
  DFFR_X1 \REGISTERS_reg[13][31]  ( .D(n3177), .CK(CLK), .RN(n1488), .Q(n2206), 
        .QN(n389) );
  DFFR_X1 \REGISTERS_reg[13][30]  ( .D(n3176), .CK(CLK), .RN(n1488), .Q(n2181), 
        .QN(n390) );
  DFFR_X1 \REGISTERS_reg[13][29]  ( .D(n3175), .CK(CLK), .RN(n1488), .Q(n2160), 
        .QN(n391) );
  DFFR_X1 \REGISTERS_reg[13][28]  ( .D(n3174), .CK(CLK), .RN(n1488), .Q(n2139), 
        .QN(n392) );
  DFFR_X1 \REGISTERS_reg[13][27]  ( .D(n3173), .CK(CLK), .RN(n1488), .Q(n2118), 
        .QN(n393) );
  DFFR_X1 \REGISTERS_reg[13][26]  ( .D(n3172), .CK(CLK), .RN(n1488), .Q(n2097), 
        .QN(n394) );
  DFFR_X1 \REGISTERS_reg[13][25]  ( .D(n3171), .CK(CLK), .RN(n1488), .Q(n2076), 
        .QN(n395) );
  DFFR_X1 \REGISTERS_reg[13][24]  ( .D(n3170), .CK(CLK), .RN(n1488), .Q(n2055), 
        .QN(n396) );
  DFFR_X1 \REGISTERS_reg[12][31]  ( .D(n3209), .CK(CLK), .RN(n1485), .Q(n2210), 
        .QN(n357) );
  DFFR_X1 \REGISTERS_reg[12][30]  ( .D(n3208), .CK(CLK), .RN(n1485), .Q(n2183), 
        .QN(n358) );
  DFFR_X1 \REGISTERS_reg[12][29]  ( .D(n3207), .CK(CLK), .RN(n1485), .Q(n2162), 
        .QN(n359) );
  DFFR_X1 \REGISTERS_reg[12][28]  ( .D(n3206), .CK(CLK), .RN(n1485), .Q(n2141), 
        .QN(n360) );
  DFFR_X1 \REGISTERS_reg[12][27]  ( .D(n3205), .CK(CLK), .RN(n1485), .Q(n2120), 
        .QN(n361) );
  DFFR_X1 \REGISTERS_reg[12][26]  ( .D(n3204), .CK(CLK), .RN(n1485), .Q(n2099), 
        .QN(n362) );
  DFFR_X1 \REGISTERS_reg[12][25]  ( .D(n3203), .CK(CLK), .RN(n1485), .Q(n2078), 
        .QN(n363) );
  DFFR_X1 \REGISTERS_reg[12][24]  ( .D(n3202), .CK(CLK), .RN(n1485), .Q(n2057), 
        .QN(n364) );
  DFFR_X1 \REGISTERS_reg[20][31]  ( .D(n2953), .CK(CLK), .RN(n1506), .QN(n613)
         );
  DFFR_X1 \REGISTERS_reg[20][30]  ( .D(n2952), .CK(CLK), .RN(n1506), .QN(n614)
         );
  DFFR_X1 \REGISTERS_reg[20][29]  ( .D(n2951), .CK(CLK), .RN(n1506), .QN(n615)
         );
  DFFR_X1 \REGISTERS_reg[20][28]  ( .D(n2950), .CK(CLK), .RN(n1506), .QN(n616)
         );
  DFFR_X1 \REGISTERS_reg[20][27]  ( .D(n2949), .CK(CLK), .RN(n1507), .QN(n617)
         );
  DFFR_X1 \REGISTERS_reg[20][26]  ( .D(n2948), .CK(CLK), .RN(n1507), .QN(n618)
         );
  DFFR_X1 \REGISTERS_reg[20][25]  ( .D(n2947), .CK(CLK), .RN(n1507), .QN(n619)
         );
  DFFR_X1 \REGISTERS_reg[20][24]  ( .D(n2946), .CK(CLK), .RN(n1507), .QN(n620)
         );
  DFFR_X1 \REGISTERS_reg[9][31]  ( .D(n3305), .CK(CLK), .RN(n1477), .Q(n4085), 
        .QN(n261) );
  DFFR_X1 \REGISTERS_reg[9][30]  ( .D(n3304), .CK(CLK), .RN(n1477), .Q(n4059), 
        .QN(n262) );
  DFFR_X1 \REGISTERS_reg[9][29]  ( .D(n3303), .CK(CLK), .RN(n1477), .Q(n4033), 
        .QN(n263) );
  DFFR_X1 \REGISTERS_reg[9][28]  ( .D(n3302), .CK(CLK), .RN(n1477), .Q(n4007), 
        .QN(n264) );
  DFFR_X1 \REGISTERS_reg[9][27]  ( .D(n3301), .CK(CLK), .RN(n1477), .Q(n3981), 
        .QN(n265) );
  DFFR_X1 \REGISTERS_reg[9][26]  ( .D(n3300), .CK(CLK), .RN(n1477), .Q(n3955), 
        .QN(n266) );
  DFFR_X1 \REGISTERS_reg[9][25]  ( .D(n3299), .CK(CLK), .RN(n1477), .Q(n3929), 
        .QN(n267) );
  DFFR_X1 \REGISTERS_reg[9][24]  ( .D(n3298), .CK(CLK), .RN(n1477), .Q(n3903), 
        .QN(n268) );
  DFFR_X1 \REGISTERS_reg[17][31]  ( .D(n3049), .CK(CLK), .RN(n1498), .Q(n4123), 
        .QN(n517) );
  DFFR_X1 \REGISTERS_reg[17][30]  ( .D(n3048), .CK(CLK), .RN(n1498), .Q(n4080), 
        .QN(n518) );
  DFFR_X1 \REGISTERS_reg[17][29]  ( .D(n3047), .CK(CLK), .RN(n1498), .Q(n4054), 
        .QN(n519) );
  DFFR_X1 \REGISTERS_reg[17][28]  ( .D(n3046), .CK(CLK), .RN(n1498), .Q(n4028), 
        .QN(n520) );
  DFFR_X1 \REGISTERS_reg[17][27]  ( .D(n3045), .CK(CLK), .RN(n1499), .Q(n4002), 
        .QN(n521) );
  DFFR_X1 \REGISTERS_reg[17][26]  ( .D(n3044), .CK(CLK), .RN(n1499), .Q(n3976), 
        .QN(n522) );
  DFFR_X1 \REGISTERS_reg[17][25]  ( .D(n3043), .CK(CLK), .RN(n1499), .Q(n3950), 
        .QN(n523) );
  DFFR_X1 \REGISTERS_reg[17][24]  ( .D(n3042), .CK(CLK), .RN(n1499), .Q(n3924), 
        .QN(n524) );
  DFFR_X1 \REGISTERS_reg[8][31]  ( .D(n3337), .CK(CLK), .RN(n1474), .QN(n229)
         );
  DFFR_X1 \REGISTERS_reg[8][30]  ( .D(n3336), .CK(CLK), .RN(n1474), .QN(n230)
         );
  DFFR_X1 \REGISTERS_reg[8][29]  ( .D(n3335), .CK(CLK), .RN(n1474), .QN(n231)
         );
  DFFR_X1 \REGISTERS_reg[8][28]  ( .D(n3334), .CK(CLK), .RN(n1474), .QN(n232)
         );
  DFFR_X1 \REGISTERS_reg[8][27]  ( .D(n3333), .CK(CLK), .RN(n1475), .QN(n233)
         );
  DFFR_X1 \REGISTERS_reg[8][26]  ( .D(n3332), .CK(CLK), .RN(n1475), .QN(n234)
         );
  DFFR_X1 \REGISTERS_reg[8][25]  ( .D(n3331), .CK(CLK), .RN(n1475), .QN(n235)
         );
  DFFR_X1 \REGISTERS_reg[8][24]  ( .D(n3330), .CK(CLK), .RN(n1475), .QN(n236)
         );
  DFFR_X1 \REGISTERS_reg[30][31]  ( .D(n2633), .CK(CLK), .RN(n1533), .QN(n933)
         );
  DFFR_X1 \REGISTERS_reg[30][30]  ( .D(n2632), .CK(CLK), .RN(n1533), .QN(n934)
         );
  DFFR_X1 \REGISTERS_reg[30][29]  ( .D(n2631), .CK(CLK), .RN(n1533), .QN(n935)
         );
  DFFR_X1 \REGISTERS_reg[30][28]  ( .D(n2630), .CK(CLK), .RN(n1533), .QN(n936)
         );
  DFFR_X1 \REGISTERS_reg[30][27]  ( .D(n2629), .CK(CLK), .RN(n1533), .QN(n937)
         );
  DFFR_X1 \REGISTERS_reg[30][26]  ( .D(n2628), .CK(CLK), .RN(n1533), .QN(n938)
         );
  DFFR_X1 \REGISTERS_reg[30][25]  ( .D(n2627), .CK(CLK), .RN(n1533), .QN(n939)
         );
  DFFR_X1 \REGISTERS_reg[30][24]  ( .D(n2626), .CK(CLK), .RN(n1533), .QN(n940)
         );
  DFFR_X1 \REGISTERS_reg[27][31]  ( .D(n2729), .CK(CLK), .RN(n1525), .Q(n4110), 
        .QN(n837) );
  DFFR_X1 \REGISTERS_reg[27][30]  ( .D(n2728), .CK(CLK), .RN(n1525), .Q(n4073), 
        .QN(n838) );
  DFFR_X1 \REGISTERS_reg[27][29]  ( .D(n2727), .CK(CLK), .RN(n1525), .Q(n4047), 
        .QN(n839) );
  DFFR_X1 \REGISTERS_reg[27][28]  ( .D(n2726), .CK(CLK), .RN(n1525), .Q(n4021), 
        .QN(n840) );
  DFFR_X1 \REGISTERS_reg[27][27]  ( .D(n2725), .CK(CLK), .RN(n1525), .Q(n3995), 
        .QN(n841) );
  DFFR_X1 \REGISTERS_reg[27][26]  ( .D(n2724), .CK(CLK), .RN(n1525), .Q(n3969), 
        .QN(n842) );
  DFFR_X1 \REGISTERS_reg[27][25]  ( .D(n2723), .CK(CLK), .RN(n1525), .Q(n3943), 
        .QN(n843) );
  DFFR_X1 \REGISTERS_reg[27][24]  ( .D(n2722), .CK(CLK), .RN(n1525), .Q(n3917), 
        .QN(n844) );
  DFFR_X2 \REGISTERS_reg[8][6]  ( .D(n3312), .CK(CLK), .RN(n1476), .QN(n254)
         );
  DFF_X2 \OUT1_reg[1]  ( .D(n2507), .CK(CLK), .Q(OUT1[1]), .QN(n4661) );
  AND2_X1 U2 ( .A1(n1030), .A2(n973), .ZN(n1) );
  AND2_X1 U3 ( .A1(n1030), .A2(n973), .ZN(n2) );
  AND2_X2 U4 ( .A1(n1030), .A2(n973), .ZN(n932) );
  AND3_X1 U5 ( .A1(ADD_RS1[0]), .A2(n706), .A3(n1560), .ZN(n1028) );
  AND2_X1 U6 ( .A1(n1182), .A2(n4256), .ZN(n3) );
  AND2_X1 U7 ( .A1(n1179), .A2(n4224), .ZN(n4) );
  NOR3_X1 U8 ( .A1(n3), .A2(n4), .A3(n2231), .ZN(n2235) );
  CLKBUF_X1 U9 ( .A(n4656), .Z(n5) );
  BUF_X2 U10 ( .A(n990), .Z(n1182) );
  BUF_X2 U11 ( .A(n992), .Z(n1179) );
  BUF_X2 U12 ( .A(n4088), .Z(n1205) );
  CLKBUF_X3 U13 ( .A(n2225), .Z(n1159) );
  CLKBUF_X3 U14 ( .A(n4091), .Z(n6) );
  BUF_X1 U15 ( .A(n4091), .Z(n1214) );
  CLKBUF_X1 U16 ( .A(n1036), .Z(n7) );
  CLKBUF_X3 U17 ( .A(n4090), .Z(n8) );
  BUF_X1 U18 ( .A(n4090), .Z(n1211) );
  CLKBUF_X3 U19 ( .A(n4099), .Z(n1230) );
  BUF_X1 U20 ( .A(n166), .Z(n55) );
  BUF_X1 U21 ( .A(n968), .Z(n9) );
  BUF_X1 U22 ( .A(n968), .Z(n1198) );
  AND2_X2 U23 ( .A1(n1554), .A2(n784), .ZN(n705) );
  OR2_X1 U24 ( .A1(n1071), .A2(n1072), .ZN(n10) );
  OR2_X1 U25 ( .A1(n1069), .A2(n1070), .ZN(n11) );
  OR2_X1 U26 ( .A1(n686), .A2(n687), .ZN(n12) );
  OR2_X1 U27 ( .A1(n602), .A2(n603), .ZN(n13) );
  OR2_X1 U28 ( .A1(n907), .A2(n906), .ZN(n14) );
  OR2_X1 U29 ( .A1(n919), .A2(n918), .ZN(n15) );
  OR2_X1 U30 ( .A1(n1042), .A2(n1041), .ZN(n16) );
  OR2_X1 U31 ( .A1(n1038), .A2(n1037), .ZN(n17) );
  OR2_X1 U32 ( .A1(n910), .A2(n911), .ZN(n18) );
  OR2_X1 U33 ( .A1(n1065), .A2(n1066), .ZN(n19) );
  OR2_X1 U34 ( .A1(n1057), .A2(n1058), .ZN(n20) );
  OR2_X1 U35 ( .A1(n765), .A2(n766), .ZN(n21) );
  OR2_X1 U36 ( .A1(n779), .A2(n780), .ZN(n22) );
  OR2_X1 U37 ( .A1(n1051), .A2(n1052), .ZN(n23) );
  OR2_X1 U38 ( .A1(n900), .A2(n901), .ZN(n24) );
  OR2_X1 U39 ( .A1(n904), .A2(n905), .ZN(n25) );
  OR2_X1 U40 ( .A1(n898), .A2(n899), .ZN(n26) );
  OR2_X1 U41 ( .A1(n777), .A2(n778), .ZN(n27) );
  OR2_X1 U42 ( .A1(n767), .A2(n768), .ZN(n28) );
  OR2_X1 U43 ( .A1(n1059), .A2(n1060), .ZN(n29) );
  OR2_X1 U44 ( .A1(n902), .A2(n903), .ZN(n30) );
  OR2_X1 U45 ( .A1(n1049), .A2(n1050), .ZN(n31) );
  OR2_X1 U46 ( .A1(n894), .A2(n895), .ZN(n32) );
  BUF_X1 U47 ( .A(n2209), .Z(n507) );
  NOR2_X1 U48 ( .A1(n2149), .A2(n21), .ZN(n2156) );
  NOR2_X1 U49 ( .A1(n2128), .A2(n31), .ZN(n2135) );
  NOR2_X1 U50 ( .A1(n2107), .A2(n28), .ZN(n2114) );
  NOR2_X1 U51 ( .A1(n1778), .A2(n26), .ZN(n1785) );
  NOR2_X1 U52 ( .A1(n1757), .A2(n30), .ZN(n1764) );
  BUF_X2 U53 ( .A(n977), .Z(n33) );
  CLKBUF_X3 U54 ( .A(n4118), .Z(n1261) );
  OR2_X1 U55 ( .A1(n385), .A2(n1214), .ZN(n34) );
  OR2_X1 U56 ( .A1(n417), .A2(n1211), .ZN(n35) );
  NAND3_X1 U57 ( .A1(n34), .A2(n35), .A3(n2323), .ZN(n2330) );
  AND2_X1 U58 ( .A1(n1181), .A2(n4274), .ZN(n36) );
  AND2_X1 U59 ( .A1(n1178), .A2(n4242), .ZN(n37) );
  NOR3_X1 U60 ( .A1(n36), .A2(n37), .A3(n1842), .ZN(n1845) );
  BUF_X2 U61 ( .A(n967), .Z(n1201) );
  AND2_X1 U62 ( .A1(n4797), .A2(n1253), .ZN(n38) );
  AND2_X1 U63 ( .A1(n1250), .A2(n4330), .ZN(n39) );
  NOR3_X1 U64 ( .A1(n38), .A2(n39), .A3(n2487), .ZN(n2495) );
  AND2_X1 U65 ( .A1(ADD_RS1[2]), .A2(n1553), .ZN(n887) );
  CLKBUF_X3 U66 ( .A(n1003), .Z(n1186) );
  CLKBUF_X3 U67 ( .A(n1003), .Z(n1187) );
  NOR2_X1 U68 ( .A1(n1694), .A2(n19), .ZN(n1701) );
  AND2_X2 U69 ( .A1(n973), .A2(n695), .ZN(n40) );
  CLKBUF_X3 U70 ( .A(n4088), .Z(n1207) );
  OR2_X1 U71 ( .A1(n1230), .A2(n186), .ZN(n41) );
  OR2_X1 U72 ( .A1(n1227), .A2(n335), .ZN(n42) );
  NAND3_X1 U73 ( .A1(n41), .A2(n42), .A3(n3909), .ZN(n3910) );
  OR2_X1 U74 ( .A1(n1228), .A2(n178), .ZN(n43) );
  OR2_X1 U75 ( .A1(n1225), .A2(n327), .ZN(n44) );
  NAND3_X1 U76 ( .A1(n43), .A2(n44), .A3(n2452), .ZN(n2453) );
  OR2_X1 U77 ( .A1(n1229), .A2(n175), .ZN(n45) );
  OR2_X1 U78 ( .A1(n1225), .A2(n324), .ZN(n46) );
  NAND3_X1 U79 ( .A1(n45), .A2(n46), .A3(n2377), .ZN(n2378) );
  OR2_X1 U80 ( .A1(n1228), .A2(n185), .ZN(n47) );
  OR2_X1 U81 ( .A1(n1226), .A2(n334), .ZN(n48) );
  NAND3_X1 U82 ( .A1(n47), .A2(n48), .A3(n3883), .ZN(n3884) );
  BUF_X1 U83 ( .A(ADD_RS1[3]), .Z(n1054) );
  NOR2_X1 U84 ( .A1(n4020), .A2(n12), .ZN(n4032) );
  BUF_X1 U85 ( .A(ADD_RS2[4]), .Z(n889) );
  NOR2_X1 U86 ( .A1(n3765), .A2(n15), .ZN(n3777) );
  OR2_X1 U87 ( .A1(n1936), .A2(n1140), .ZN(n49) );
  OR2_X1 U88 ( .A1(n114), .A2(n1137), .ZN(n50) );
  NAND3_X1 U89 ( .A1(n49), .A2(n50), .A3(n1935), .ZN(n1937) );
  BUF_X1 U90 ( .A(n494), .Z(n51) );
  BUF_X1 U91 ( .A(n494), .Z(n1121) );
  BUF_X1 U92 ( .A(n970), .Z(n52) );
  BUF_X1 U93 ( .A(n970), .Z(n1120) );
  BUF_X2 U94 ( .A(n970), .Z(n508) );
  BUF_X2 U95 ( .A(n482), .Z(n1016) );
  NOR2_X1 U96 ( .A1(n53), .A2(n2238), .ZN(n1000) );
  OR3_X1 U97 ( .A1(ADD_RS2[4]), .A2(ADD_RS2[3]), .A3(ADD_RS2[0]), .ZN(n53) );
  CLKBUF_X1 U98 ( .A(n1028), .Z(n1015) );
  BUF_X2 U99 ( .A(n166), .Z(n54) );
  BUF_X2 U100 ( .A(n965), .Z(n56) );
  BUF_X2 U101 ( .A(n965), .Z(n57) );
  AND2_X1 U102 ( .A1(n1077), .A2(n705), .ZN(n166) );
  NOR2_X1 U103 ( .A1(n3640), .A2(n16), .ZN(n3652) );
  OR2_X1 U104 ( .A1(n1874), .A2(n1140), .ZN(n58) );
  OR2_X1 U105 ( .A1(n117), .A2(n1137), .ZN(n59) );
  NAND3_X1 U106 ( .A1(n58), .A2(n59), .A3(n1873), .ZN(n1875) );
  OR2_X1 U107 ( .A1(n3959), .A2(n1127), .ZN(n60) );
  OR2_X1 U108 ( .A1(n266), .A2(n678), .ZN(n61) );
  NAND3_X1 U109 ( .A1(n60), .A2(n61), .A3(n2096), .ZN(n2104) );
  BUF_X2 U110 ( .A(n494), .Z(n512) );
  OR2_X1 U111 ( .A1(n3681), .A2(n1128), .ZN(n62) );
  OR2_X1 U112 ( .A1(n277), .A2(n1126), .ZN(n63) );
  NAND3_X1 U113 ( .A1(n1871), .A2(n63), .A3(n62), .ZN(n1877) );
  OR2_X1 U114 ( .A1(n1997), .A2(n1140), .ZN(n64) );
  OR2_X1 U115 ( .A1(n111), .A2(n1137), .ZN(n65) );
  NAND3_X1 U116 ( .A1(n64), .A2(n65), .A3(n1996), .ZN(n1998) );
  NOR2_X1 U117 ( .A1(n2086), .A2(n23), .ZN(n2093) );
  BUF_X2 U118 ( .A(n967), .Z(n66) );
  AND2_X2 U119 ( .A1(n974), .A2(n2265), .ZN(n967) );
  NOR2_X1 U120 ( .A1(n2434), .A2(n11), .ZN(n2446) );
  NOR2_X1 U121 ( .A1(n1736), .A2(n20), .ZN(n1743) );
  OR2_X1 U122 ( .A1(n1730), .A2(n1139), .ZN(n67) );
  OR2_X1 U123 ( .A1(n124), .A2(n1136), .ZN(n68) );
  NAND3_X1 U124 ( .A1(n67), .A2(n68), .A3(n1729), .ZN(n1731) );
  NOR2_X1 U125 ( .A1(n1715), .A2(n29), .ZN(n1722) );
  OR2_X1 U126 ( .A1(n1709), .A2(n1139), .ZN(n69) );
  OR2_X1 U127 ( .A1(n125), .A2(n1136), .ZN(n70) );
  NAND3_X1 U128 ( .A1(n69), .A2(n70), .A3(n1708), .ZN(n1710) );
  NOR2_X1 U129 ( .A1(n1611), .A2(n27), .ZN(n1618) );
  OR2_X1 U130 ( .A1(n1605), .A2(n1139), .ZN(n71) );
  OR2_X1 U131 ( .A1(n130), .A2(n1136), .ZN(n72) );
  NAND3_X1 U132 ( .A1(n71), .A2(n72), .A3(n1604), .ZN(n1606) );
  NOR2_X1 U133 ( .A1(n2044), .A2(n24), .ZN(n2051) );
  OR2_X1 U134 ( .A1(n2038), .A2(n1140), .ZN(n73) );
  OR2_X1 U135 ( .A1(n109), .A2(n1137), .ZN(n74) );
  NAND3_X1 U136 ( .A1(n73), .A2(n74), .A3(n2037), .ZN(n2039) );
  NOR2_X1 U137 ( .A1(n2023), .A2(n25), .ZN(n2030) );
  OR2_X1 U138 ( .A1(n2017), .A2(n1140), .ZN(n75) );
  OR2_X1 U139 ( .A1(n110), .A2(n1137), .ZN(n76) );
  NAND3_X1 U140 ( .A1(n75), .A2(n76), .A3(n2016), .ZN(n2018) );
  NOR2_X1 U141 ( .A1(n1982), .A2(n18), .ZN(n1989) );
  NOR3_X1 U142 ( .A1(n4656), .A2(n4645), .A3(n4657), .ZN(n77) );
  NOR3_X1 U143 ( .A1(n4657), .A2(n4645), .A3(n5), .ZN(n78) );
  AND2_X1 U144 ( .A1(n1268), .A2(n4278), .ZN(n79) );
  AND2_X1 U145 ( .A1(n1265), .A2(n4246), .ZN(n80) );
  NOR3_X1 U146 ( .A1(n79), .A2(n80), .A3(n2490), .ZN(n2494) );
  OR2_X1 U147 ( .A1(n635), .A2(n1262), .ZN(n81) );
  OR2_X1 U148 ( .A1(n1259), .A2(n2489), .ZN(n82) );
  OR2_X1 U149 ( .A1(n590), .A2(n2488), .ZN(n83) );
  NAND3_X1 U150 ( .A1(n81), .A2(n82), .A3(n83), .ZN(n2490) );
  BUF_X2 U151 ( .A(n986), .Z(n1268) );
  BUF_X2 U152 ( .A(n985), .Z(n1265) );
  BUF_X1 U153 ( .A(ADD_RS1[3]), .Z(n84) );
  OR2_X1 U154 ( .A1(n376), .A2(n1213), .ZN(n85) );
  OR2_X1 U155 ( .A1(n408), .A2(n8), .ZN(n86) );
  NAND3_X1 U156 ( .A1(n85), .A2(n86), .A3(n3604), .ZN(n3611) );
  CLKBUF_X1 U157 ( .A(n998), .Z(n87) );
  NOR2_X1 U158 ( .A1(n1861), .A2(n22), .ZN(n1868) );
  NOR2_X1 U159 ( .A1(n1799), .A2(n32), .ZN(n1806) );
  OR2_X1 U160 ( .A1(n1230), .A2(n187), .ZN(n88) );
  OR2_X1 U161 ( .A1(n1227), .A2(n336), .ZN(n89) );
  NAND3_X1 U162 ( .A1(n88), .A2(n89), .A3(n3935), .ZN(n3936) );
  BUF_X2 U163 ( .A(n4098), .Z(n1227) );
  NOR2_X1 U164 ( .A1(n4046), .A2(n13), .ZN(n4058) );
  OR2_X1 U165 ( .A1(n1205), .A2(n319), .ZN(n90) );
  OR2_X1 U166 ( .A1(n231), .A2(n1204), .ZN(n91) );
  NAND3_X1 U167 ( .A1(n90), .A2(n91), .A3(n4034), .ZN(n4043) );
  BUF_X2 U168 ( .A(n4087), .Z(n1204) );
  OR2_X1 U169 ( .A1(n1205), .A2(n308), .ZN(n92) );
  OR2_X1 U170 ( .A1(n242), .A2(n1203), .ZN(n93) );
  NAND3_X1 U171 ( .A1(n92), .A2(n93), .A3(n3753), .ZN(n3762) );
  OR2_X1 U172 ( .A1(n1205), .A2(n303), .ZN(n94) );
  OR2_X1 U173 ( .A1(n247), .A2(n1203), .ZN(n95) );
  NAND3_X1 U174 ( .A1(n94), .A2(n95), .A3(n3628), .ZN(n3637) );
  NOR2_X1 U175 ( .A1(n2409), .A2(n10), .ZN(n2421) );
  OR2_X1 U176 ( .A1(n1228), .A2(n176), .ZN(n96) );
  OR2_X1 U177 ( .A1(n1225), .A2(n325), .ZN(n97) );
  NAND3_X1 U178 ( .A1(n96), .A2(n97), .A3(n2402), .ZN(n2403) );
  NOR2_X1 U179 ( .A1(n3665), .A2(n17), .ZN(n3677) );
  OR2_X1 U180 ( .A1(n1230), .A2(n182), .ZN(n98) );
  OR2_X1 U181 ( .A1(n1226), .A2(n331), .ZN(n99) );
  NAND3_X1 U182 ( .A1(n98), .A2(n99), .A3(n3658), .ZN(n3659) );
  OR2_X1 U183 ( .A1(n1229), .A2(n184), .ZN(n100) );
  OR2_X1 U184 ( .A1(n1226), .A2(n333), .ZN(n165) );
  NAND3_X1 U185 ( .A1(n100), .A2(n165), .A3(n3758), .ZN(n3759) );
  AND2_X1 U186 ( .A1(n1077), .A2(n705), .ZN(n965) );
  NOR2_X1 U187 ( .A1(n3890), .A2(n14), .ZN(n3902) );
  OR2_X1 U188 ( .A1(n1205), .A2(n313), .ZN(n167) );
  OR2_X1 U189 ( .A1(n237), .A2(n1203), .ZN(n168) );
  NAND3_X1 U190 ( .A1(n167), .A2(n168), .A3(n3878), .ZN(n3887) );
  OR2_X1 U191 ( .A1(n1205), .A2(n297), .ZN(n169) );
  OR2_X1 U192 ( .A1(n254), .A2(n1202), .ZN(n170) );
  NAND3_X1 U193 ( .A1(n169), .A2(n170), .A3(n2397), .ZN(n2406) );
  CLKBUF_X3 U194 ( .A(n4087), .Z(n1202) );
  BUF_X2 U195 ( .A(n4111), .Z(n1245) );
  AND2_X1 U196 ( .A1(ADD_RS1[2]), .A2(n784), .ZN(n171) );
  AND2_X1 U197 ( .A1(ADD_RS1[0]), .A2(n1002), .ZN(n172) );
  AND2_X1 U198 ( .A1(n4004), .A2(n4003), .ZN(n222) );
  AND2_X1 U199 ( .A1(n3952), .A2(n3951), .ZN(n223) );
  NAND2_X1 U200 ( .A1(n693), .A2(n694), .ZN(n352) );
  OR2_X1 U201 ( .A1(n709), .A2(n708), .ZN(n353) );
  OR2_X1 U202 ( .A1(n1107), .A2(n1108), .ZN(n354) );
  OR2_X1 U203 ( .A1(n908), .A2(n909), .ZN(n355) );
  OR2_X1 U204 ( .A1(n1103), .A2(n1104), .ZN(n356) );
  OR2_X1 U205 ( .A1(n912), .A2(n913), .ZN(n421) );
  OR2_X1 U206 ( .A1(n920), .A2(n921), .ZN(n422) );
  OR2_X1 U207 ( .A1(n923), .A2(n924), .ZN(n423) );
  OR2_X1 U208 ( .A1(n1095), .A2(n1096), .ZN(n424) );
  OR2_X1 U209 ( .A1(n1109), .A2(n1110), .ZN(n425) );
  OR2_X1 U210 ( .A1(n914), .A2(n915), .ZN(n426) );
  OR2_X1 U211 ( .A1(n916), .A2(n917), .ZN(n427) );
  OR2_X1 U212 ( .A1(n1043), .A2(n1044), .ZN(n428) );
  OR2_X1 U213 ( .A1(n772), .A2(n771), .ZN(n429) );
  OR2_X1 U214 ( .A1(n1105), .A2(n1106), .ZN(n430) );
  OR2_X1 U215 ( .A1(n1064), .A2(n1063), .ZN(n431) );
  OR2_X1 U216 ( .A1(n897), .A2(n896), .ZN(n432) );
  OR2_X1 U217 ( .A1(n758), .A2(n757), .ZN(n433) );
  OR2_X1 U218 ( .A1(n683), .A2(n682), .ZN(n434) );
  OR2_X1 U219 ( .A1(n761), .A2(n762), .ZN(n435) );
  OR2_X1 U220 ( .A1(n774), .A2(n773), .ZN(n436) );
  OR2_X1 U221 ( .A1(n770), .A2(n769), .ZN(n437) );
  OR2_X1 U222 ( .A1(n782), .A2(n781), .ZN(n438) );
  AND2_X1 U223 ( .A1(ENABLE), .A2(n1538), .ZN(n462) );
  CLKBUF_X3 U224 ( .A(n4113), .Z(n1248) );
  AND4_X1 U225 ( .A1(n979), .A2(n2260), .A3(n1274), .A4(n926), .ZN(n463) );
  OR2_X1 U226 ( .A1(n1048), .A2(n1047), .ZN(n464) );
  BUF_X2 U227 ( .A(n988), .Z(n1281) );
  AND2_X1 U228 ( .A1(n3978), .A2(n3977), .ZN(n465) );
  AND2_X1 U229 ( .A1(n3926), .A2(n3925), .ZN(n466) );
  BUF_X2 U230 ( .A(n988), .Z(n1283) );
  BUF_X1 U231 ( .A(n972), .Z(n739) );
  BUF_X1 U232 ( .A(n1208), .Z(n892) );
  OR2_X1 U233 ( .A1(n785), .A2(n786), .ZN(n467) );
  AND2_X2 U234 ( .A1(n1554), .A2(n1553), .ZN(n468) );
  AND2_X1 U235 ( .A1(n4030), .A2(n4029), .ZN(n469) );
  AND2_X2 U236 ( .A1(n1031), .A2(n705), .ZN(n888) );
  AND3_X1 U237 ( .A1(n4648), .A2(n4646), .A3(n4647), .ZN(n470) );
  AND2_X1 U238 ( .A1(n4081), .A2(n4082), .ZN(n471) );
  AND3_X1 U239 ( .A1(n4648), .A2(n4646), .A3(n4647), .ZN(n1006) );
  AND2_X1 U240 ( .A1(n4056), .A2(n4055), .ZN(n472) );
  CLKBUF_X1 U241 ( .A(n976), .Z(n473) );
  BUF_X1 U242 ( .A(ADD_RS2[0]), .Z(n882) );
  NOR2_X1 U243 ( .A1(n474), .A2(n475), .ZN(n1968) );
  NAND3_X1 U244 ( .A1(n515), .A2(n516), .A3(n549), .ZN(n474) );
  OR2_X1 U245 ( .A1(n1067), .A2(n1068), .ZN(n475) );
  NOR2_X1 U246 ( .A1(n476), .A2(n477), .ZN(n1948) );
  NAND3_X1 U247 ( .A1(n499), .A2(n500), .A3(n501), .ZN(n476) );
  OR2_X1 U248 ( .A1(n1075), .A2(n1076), .ZN(n477) );
  NOR2_X1 U249 ( .A1(n478), .A2(n479), .ZN(n1826) );
  NAND3_X1 U250 ( .A1(n793), .A2(n794), .A3(n795), .ZN(n478) );
  OR2_X1 U251 ( .A1(n1100), .A2(n1099), .ZN(n479) );
  CLKBUF_X3 U252 ( .A(n4111), .Z(n480) );
  BUF_X1 U253 ( .A(n2208), .Z(n1132) );
  BUF_X1 U254 ( .A(n968), .Z(n1196) );
  AND2_X1 U255 ( .A1(n705), .A2(n692), .ZN(n481) );
  AND2_X1 U256 ( .A1(n705), .A2(n880), .ZN(n482) );
  AND2_X1 U257 ( .A1(n705), .A2(n880), .ZN(n877) );
  AND2_X1 U258 ( .A1(n172), .A2(n887), .ZN(n483) );
  AND2_X1 U259 ( .A1(n172), .A2(n887), .ZN(n484) );
  AND2_X1 U260 ( .A1(n172), .A2(n887), .ZN(n972) );
  BUF_X1 U261 ( .A(n2209), .Z(n1134) );
  AND2_X2 U262 ( .A1(n2260), .A2(n883), .ZN(n987) );
  AND2_X2 U263 ( .A1(n2260), .A2(n883), .ZN(n704) );
  AND2_X2 U264 ( .A1(n2260), .A2(n883), .ZN(n589) );
  NAND2_X1 U265 ( .A1(n886), .A2(n468), .ZN(n485) );
  CLKBUF_X1 U266 ( .A(n972), .Z(n486) );
  CLKBUF_X1 U267 ( .A(n972), .Z(n487) );
  INV_X1 U268 ( .A(ADD_RS2[3]), .ZN(n488) );
  BUF_X1 U269 ( .A(n702), .Z(n489) );
  BUF_X1 U270 ( .A(n702), .Z(n490) );
  BUF_X1 U271 ( .A(n702), .Z(n577) );
  NOR2_X1 U272 ( .A1(n2284), .A2(n354), .ZN(n2296) );
  OR2_X1 U273 ( .A1(n1229), .A2(n439), .ZN(n491) );
  OR2_X1 U274 ( .A1(n1225), .A2(n440), .ZN(n492) );
  NAND3_X1 U275 ( .A1(n491), .A2(n492), .A3(n2277), .ZN(n2278) );
  AND2_X1 U276 ( .A1(n1028), .A2(n171), .ZN(n493) );
  AND2_X1 U277 ( .A1(n1028), .A2(n171), .ZN(n494) );
  AND2_X1 U278 ( .A1(n1028), .A2(n171), .ZN(n970) );
  BUF_X1 U279 ( .A(n968), .Z(n495) );
  BUF_X1 U280 ( .A(n968), .Z(n496) );
  CLKBUF_X3 U281 ( .A(n4088), .Z(n1206) );
  BUF_X1 U282 ( .A(n484), .Z(n497) );
  CLKBUF_X3 U283 ( .A(n4119), .Z(n1262) );
  CLKBUF_X3 U284 ( .A(n4119), .Z(n1263) );
  CLKBUF_X3 U285 ( .A(n4119), .Z(n1264) );
  BUF_X1 U286 ( .A(n4116), .Z(n1257) );
  NAND4_X1 U287 ( .A1(n926), .A2(n878), .A3(n1274), .A4(n980), .ZN(n498) );
  BUF_X1 U288 ( .A(n1036), .Z(n878) );
  OR2_X1 U289 ( .A1(n1941), .A2(n1146), .ZN(n499) );
  OR2_X1 U290 ( .A1(n818), .A2(n1149), .ZN(n500) );
  OR2_X1 U291 ( .A1(n3763), .A2(n1143), .ZN(n501) );
  NOR2_X1 U292 ( .A1(n502), .A2(n503), .ZN(n1638) );
  NAND3_X1 U293 ( .A1(n796), .A2(n797), .A3(n798), .ZN(n502) );
  OR2_X1 U294 ( .A1(n1087), .A2(n1086), .ZN(n503) );
  BUF_X1 U295 ( .A(n702), .Z(n578) );
  NOR2_X1 U296 ( .A1(n3865), .A2(n355), .ZN(n3877) );
  OR2_X1 U297 ( .A1(n1229), .A2(n441), .ZN(n504) );
  OR2_X1 U298 ( .A1(n1226), .A2(n442), .ZN(n505) );
  NAND3_X1 U299 ( .A1(n504), .A2(n505), .A3(n3858), .ZN(n3859) );
  INV_X1 U300 ( .A(n1561), .ZN(n1014) );
  CLKBUF_X3 U301 ( .A(n2208), .Z(n506) );
  CLKBUF_X3 U302 ( .A(n4113), .Z(n509) );
  NOR2_X1 U303 ( .A1(n2309), .A2(n356), .ZN(n2321) );
  OR2_X1 U304 ( .A1(n386), .A2(n1214), .ZN(n510) );
  OR2_X1 U305 ( .A1(n418), .A2(n1211), .ZN(n511) );
  NAND3_X1 U306 ( .A1(n510), .A2(n511), .A3(n2298), .ZN(n2305) );
  CLKBUF_X3 U307 ( .A(n4091), .Z(n1213) );
  CLKBUF_X3 U308 ( .A(n4090), .Z(n1210) );
  NOR2_X1 U309 ( .A1(n4109), .A2(n435), .ZN(n4127) );
  AND2_X1 U310 ( .A1(n4791), .A2(n1253), .ZN(n513) );
  AND2_X1 U311 ( .A1(n1250), .A2(n4336), .ZN(n514) );
  NOR3_X1 U312 ( .A1(n513), .A2(n2337), .A3(n514), .ZN(n2345) );
  BUF_X2 U313 ( .A(n977), .Z(n1253) );
  BUF_X2 U314 ( .A(n989), .Z(n1250) );
  OR2_X1 U315 ( .A1(n1961), .A2(n1146), .ZN(n515) );
  OR2_X1 U316 ( .A1(n817), .A2(n1149), .ZN(n516) );
  OR2_X1 U317 ( .A1(n3788), .A2(n1143), .ZN(n549) );
  AND3_X1 U318 ( .A1(n1560), .A2(n706), .A3(n881), .ZN(n1031) );
  BUF_X1 U319 ( .A(n702), .Z(n579) );
  OR2_X1 U320 ( .A1(n161), .A2(n1117), .ZN(n550) );
  OR2_X1 U321 ( .A1(n1620), .A2(n2200), .ZN(n551) );
  NAND3_X1 U322 ( .A1(n550), .A2(n551), .A3(n1619), .ZN(n1630) );
  NOR2_X1 U323 ( .A1(n3840), .A2(n421), .ZN(n3852) );
  OR2_X1 U324 ( .A1(n1230), .A2(n443), .ZN(n552) );
  OR2_X1 U325 ( .A1(n1226), .A2(n444), .ZN(n553) );
  NAND3_X1 U326 ( .A1(n552), .A2(n553), .A3(n3833), .ZN(n3834) );
  NOR2_X1 U327 ( .A1(n3740), .A2(n422), .ZN(n3752) );
  OR2_X1 U328 ( .A1(n1228), .A2(n445), .ZN(n554) );
  OR2_X1 U329 ( .A1(n1226), .A2(n446), .ZN(n555) );
  NAND3_X1 U330 ( .A1(n554), .A2(n555), .A3(n3733), .ZN(n3734) );
  NOR2_X1 U331 ( .A1(n3715), .A2(n423), .ZN(n3727) );
  OR2_X1 U332 ( .A1(n1229), .A2(n447), .ZN(n556) );
  OR2_X1 U333 ( .A1(n1226), .A2(n448), .ZN(n557) );
  NAND3_X1 U334 ( .A1(n556), .A2(n557), .A3(n3708), .ZN(n3709) );
  NOR2_X1 U335 ( .A1(n2359), .A2(n424), .ZN(n2371) );
  OR2_X1 U336 ( .A1(n1228), .A2(n449), .ZN(n558) );
  OR2_X1 U337 ( .A1(n1225), .A2(n450), .ZN(n559) );
  NAND3_X1 U338 ( .A1(n558), .A2(n559), .A3(n2352), .ZN(n2353) );
  NOR2_X1 U339 ( .A1(n2255), .A2(n425), .ZN(n2271) );
  OR2_X1 U340 ( .A1(n1230), .A2(n451), .ZN(n560) );
  OR2_X1 U341 ( .A1(n1225), .A2(n452), .ZN(n561) );
  NAND3_X1 U342 ( .A1(n560), .A2(n561), .A3(n2248), .ZN(n2249) );
  CLKBUF_X3 U343 ( .A(n4099), .Z(n1228) );
  CLKBUF_X3 U344 ( .A(n4098), .Z(n1225) );
  NOR2_X1 U345 ( .A1(n3815), .A2(n426), .ZN(n3827) );
  OR2_X1 U346 ( .A1(n1230), .A2(n453), .ZN(n562) );
  OR2_X1 U347 ( .A1(n1226), .A2(n454), .ZN(n563) );
  NAND3_X1 U348 ( .A1(n562), .A2(n563), .A3(n3808), .ZN(n3809) );
  NOR2_X1 U349 ( .A1(n3790), .A2(n427), .ZN(n3802) );
  OR2_X1 U350 ( .A1(n1228), .A2(n455), .ZN(n564) );
  OR2_X1 U351 ( .A1(n1226), .A2(n456), .ZN(n565) );
  NAND3_X1 U352 ( .A1(n564), .A2(n565), .A3(n3783), .ZN(n3784) );
  CLKBUF_X3 U353 ( .A(n4098), .Z(n1226) );
  OR2_X1 U354 ( .A1(n3581), .A2(n1129), .ZN(n566) );
  OR2_X1 U355 ( .A1(n281), .A2(n1125), .ZN(n567) );
  NAND3_X1 U356 ( .A1(n566), .A2(n567), .A3(n1788), .ZN(n1796) );
  OR2_X1 U357 ( .A1(n2475), .A2(n1128), .ZN(n568) );
  OR2_X1 U358 ( .A1(n283), .A2(n1125), .ZN(n569) );
  NAND3_X1 U359 ( .A1(n568), .A2(n569), .A3(n1746), .ZN(n1754) );
  OR2_X1 U360 ( .A1(n3656), .A2(n1127), .ZN(n570) );
  OR2_X1 U361 ( .A1(n278), .A2(n1126), .ZN(n571) );
  NAND3_X1 U362 ( .A1(n570), .A2(n571), .A3(n1850), .ZN(n1858) );
  OR2_X1 U363 ( .A1(n3631), .A2(n1128), .ZN(n572) );
  OR2_X1 U364 ( .A1(n279), .A2(n1126), .ZN(n573) );
  NAND3_X1 U365 ( .A1(n1829), .A2(n573), .A3(n572), .ZN(n1837) );
  NOR2_X1 U366 ( .A1(n1673), .A2(n467), .ZN(n1680) );
  OR2_X1 U367 ( .A1(n831), .A2(n1148), .ZN(n574) );
  OR2_X1 U368 ( .A1(n1672), .A2(n1145), .ZN(n575) );
  OR2_X1 U369 ( .A1(n2382), .A2(n1142), .ZN(n576) );
  NAND3_X1 U370 ( .A1(n575), .A2(n574), .A3(n576), .ZN(n1673) );
  CLKBUF_X3 U371 ( .A(n2220), .Z(n1142) );
  BUF_X2 U372 ( .A(n783), .Z(n668) );
  BUF_X2 U373 ( .A(n482), .Z(n1123) );
  NOR2_X1 U374 ( .A1(n2224), .A2(n434), .ZN(n2237) );
  OR2_X1 U375 ( .A1(n805), .A2(n1150), .ZN(n580) );
  OR2_X1 U376 ( .A1(n2222), .A2(n1147), .ZN(n581) );
  OR2_X1 U377 ( .A1(n4104), .A2(n1144), .ZN(n582) );
  NAND3_X1 U378 ( .A1(n580), .A2(n581), .A3(n582), .ZN(n2224) );
  OR2_X1 U379 ( .A1(n1646), .A2(n1139), .ZN(n583) );
  OR2_X1 U380 ( .A1(n128), .A2(n1136), .ZN(n584) );
  NAND3_X1 U381 ( .A1(n583), .A2(n584), .A3(n1645), .ZN(n1647) );
  CLKBUF_X3 U382 ( .A(n4118), .Z(n1260) );
  OR2_X1 U383 ( .A1(n3606), .A2(n1129), .ZN(n585) );
  OR2_X1 U384 ( .A1(n280), .A2(n1126), .ZN(n586) );
  NAND3_X1 U385 ( .A1(n1809), .A2(n586), .A3(n585), .ZN(n1817) );
  CLKBUF_X3 U386 ( .A(n4111), .Z(n1246) );
  OR2_X1 U387 ( .A1(n1587), .A2(n1139), .ZN(n587) );
  OR2_X1 U388 ( .A1(n131), .A2(n1136), .ZN(n588) );
  NAND3_X1 U389 ( .A1(n587), .A2(n588), .A3(n1586), .ZN(n1588) );
  CLKBUF_X3 U390 ( .A(n4116), .Z(n590) );
  CLKBUF_X1 U391 ( .A(n1092), .Z(n763) );
  NOR2_X1 U392 ( .A1(n3690), .A2(n353), .ZN(n3702) );
  OR2_X1 U393 ( .A1(n821), .A2(n1238), .ZN(n591) );
  OR2_X1 U394 ( .A1(n3689), .A2(n1235), .ZN(n592) );
  OR2_X1 U395 ( .A1(n1232), .A2(n3688), .ZN(n593) );
  NAND3_X1 U396 ( .A1(n592), .A2(n591), .A3(n593), .ZN(n3690) );
  CLKBUF_X3 U397 ( .A(n4108), .Z(n1238) );
  CLKBUF_X3 U398 ( .A(n4106), .Z(n1235) );
  CLKBUF_X3 U399 ( .A(n4105), .Z(n1232) );
  AND2_X1 U400 ( .A1(n4882), .A2(n1244), .ZN(n594) );
  AND2_X1 U401 ( .A1(n1242), .A2(n4073), .ZN(n595) );
  NOR3_X1 U402 ( .A1(n4072), .A2(n595), .A3(n594), .ZN(n4084) );
  NOR2_X1 U403 ( .A1(n2065), .A2(n429), .ZN(n2072) );
  OR2_X1 U404 ( .A1(n812), .A2(n1150), .ZN(n596) );
  OR2_X1 U405 ( .A1(n2064), .A2(n1147), .ZN(n597) );
  OR2_X1 U406 ( .A1(n3914), .A2(n1144), .ZN(n598) );
  NAND3_X1 U407 ( .A1(n597), .A2(n596), .A3(n598), .ZN(n2065) );
  CLKBUF_X3 U408 ( .A(n2226), .Z(n1161) );
  CLKBUF_X3 U409 ( .A(n2226), .Z(n1160) );
  NOR2_X1 U410 ( .A1(n2170), .A2(n433), .ZN(n2177) );
  OR2_X1 U411 ( .A1(n807), .A2(n1150), .ZN(n599) );
  OR2_X1 U412 ( .A1(n2169), .A2(n1147), .ZN(n600) );
  OR2_X1 U413 ( .A1(n4044), .A2(n1144), .ZN(n601) );
  NAND3_X1 U414 ( .A1(n600), .A2(n599), .A3(n601), .ZN(n2170) );
  BUF_X2 U415 ( .A(n2223), .Z(n1150) );
  BUF_X2 U416 ( .A(n2221), .Z(n1147) );
  AND2_X1 U417 ( .A1(n4881), .A2(n1244), .ZN(n602) );
  AND2_X1 U418 ( .A1(n1242), .A2(n4047), .ZN(n603) );
  AND2_X1 U419 ( .A1(n1077), .A2(n887), .ZN(n966) );
  NOR2_X1 U420 ( .A1(n3615), .A2(n428), .ZN(n3627) );
  OR2_X1 U421 ( .A1(n1205), .A2(n461), .ZN(n604) );
  OR2_X1 U422 ( .A1(n248), .A2(n1203), .ZN(n605) );
  NAND3_X1 U423 ( .A1(n604), .A2(n605), .A3(n3603), .ZN(n3612) );
  CLKBUF_X3 U424 ( .A(n4087), .Z(n1203) );
  NOR2_X1 U425 ( .A1(n1570), .A2(n430), .ZN(n1579) );
  AND2_X1 U426 ( .A1(n1270), .A2(n4259), .ZN(n606) );
  AND2_X1 U427 ( .A1(n1267), .A2(n4227), .ZN(n607) );
  NOR3_X1 U428 ( .A1(n4026), .A2(n607), .A3(n606), .ZN(n4030) );
  OR2_X1 U429 ( .A1(n616), .A2(n1264), .ZN(n608) );
  OR2_X1 U430 ( .A1(n1261), .A2(n4025), .ZN(n609) );
  OR2_X1 U431 ( .A1(n1256), .A2(n4024), .ZN(n610) );
  NAND3_X1 U432 ( .A1(n608), .A2(n609), .A3(n610), .ZN(n4026) );
  AND2_X1 U433 ( .A1(n1270), .A2(n4260), .ZN(n611) );
  AND2_X1 U434 ( .A1(n1267), .A2(n4228), .ZN(n612) );
  NOR3_X1 U435 ( .A1(n4000), .A2(n612), .A3(n611), .ZN(n4004) );
  OR2_X1 U436 ( .A1(n617), .A2(n1264), .ZN(n645) );
  OR2_X1 U437 ( .A1(n1261), .A2(n3999), .ZN(n646) );
  OR2_X1 U438 ( .A1(n3998), .A2(n1258), .ZN(n647) );
  NAND3_X1 U439 ( .A1(n645), .A2(n646), .A3(n647), .ZN(n4000) );
  AND2_X1 U440 ( .A1(n1270), .A2(n4261), .ZN(n648) );
  AND2_X1 U441 ( .A1(n1267), .A2(n4229), .ZN(n649) );
  NOR3_X1 U442 ( .A1(n648), .A2(n649), .A3(n3974), .ZN(n3978) );
  OR2_X1 U443 ( .A1(n618), .A2(n1264), .ZN(n650) );
  OR2_X1 U444 ( .A1(n1261), .A2(n3973), .ZN(n651) );
  OR2_X1 U445 ( .A1(n3972), .A2(n1257), .ZN(n652) );
  NAND3_X1 U446 ( .A1(n650), .A2(n651), .A3(n652), .ZN(n3974) );
  AND2_X1 U447 ( .A1(n1270), .A2(n4262), .ZN(n653) );
  AND2_X1 U448 ( .A1(n1267), .A2(n4230), .ZN(n654) );
  NOR3_X1 U449 ( .A1(n653), .A2(n654), .A3(n3948), .ZN(n3952) );
  OR2_X1 U450 ( .A1(n619), .A2(n1264), .ZN(n655) );
  OR2_X1 U451 ( .A1(n1261), .A2(n3947), .ZN(n656) );
  OR2_X1 U452 ( .A1(n3946), .A2(n1257), .ZN(n657) );
  NAND3_X1 U453 ( .A1(n655), .A2(n656), .A3(n657), .ZN(n3948) );
  AND2_X1 U454 ( .A1(n1270), .A2(n4263), .ZN(n658) );
  AND2_X1 U455 ( .A1(n1267), .A2(n4231), .ZN(n659) );
  NOR3_X1 U456 ( .A1(n658), .A2(n659), .A3(n3922), .ZN(n3926) );
  OR2_X1 U457 ( .A1(n620), .A2(n1264), .ZN(n660) );
  OR2_X1 U458 ( .A1(n1261), .A2(n3921), .ZN(n661) );
  OR2_X1 U459 ( .A1(n3920), .A2(n1257), .ZN(n662) );
  NAND3_X1 U460 ( .A1(n660), .A2(n661), .A3(n662), .ZN(n3922) );
  BUF_X2 U461 ( .A(n986), .Z(n1270) );
  BUF_X2 U462 ( .A(n985), .Z(n1267) );
  AND2_X1 U463 ( .A1(n1156), .A2(n4882), .ZN(n663) );
  AND2_X1 U464 ( .A1(n1151), .A2(n4073), .ZN(n664) );
  NOR3_X1 U465 ( .A1(n2191), .A2(n664), .A3(n663), .ZN(n2198) );
  NOR2_X1 U466 ( .A1(n3968), .A2(n436), .ZN(n3980) );
  OR2_X1 U467 ( .A1(n810), .A2(n1239), .ZN(n665) );
  OR2_X1 U468 ( .A1(n3967), .A2(n1236), .ZN(n666) );
  OR2_X1 U469 ( .A1(n1233), .A2(n3966), .ZN(n667) );
  NAND3_X1 U470 ( .A1(n666), .A2(n665), .A3(n667), .ZN(n3968) );
  AND2_X1 U471 ( .A1(n1077), .A2(n887), .ZN(n702) );
  BUF_X2 U472 ( .A(n783), .Z(n669) );
  NOR2_X1 U473 ( .A1(n2459), .A2(n431), .ZN(n2471) );
  OR2_X1 U474 ( .A1(n828), .A2(n1237), .ZN(n670) );
  OR2_X1 U475 ( .A1(n2458), .A2(n1234), .ZN(n671) );
  OR2_X1 U476 ( .A1(n1231), .A2(n2457), .ZN(n672) );
  NAND3_X1 U477 ( .A1(n671), .A2(n670), .A3(n672), .ZN(n2459) );
  NOR2_X1 U478 ( .A1(n2384), .A2(n432), .ZN(n2396) );
  OR2_X1 U479 ( .A1(n831), .A2(n1237), .ZN(n673) );
  OR2_X1 U480 ( .A1(n2383), .A2(n1234), .ZN(n674) );
  OR2_X1 U481 ( .A1(n1231), .A2(n2382), .ZN(n675) );
  NAND3_X1 U482 ( .A1(n674), .A2(n673), .A3(n675), .ZN(n2384) );
  CLKBUF_X3 U483 ( .A(n4108), .Z(n1237) );
  CLKBUF_X3 U484 ( .A(n4106), .Z(n1234) );
  CLKBUF_X3 U485 ( .A(n4105), .Z(n1231) );
  NOR2_X1 U486 ( .A1(n3994), .A2(n437), .ZN(n4006) );
  OR2_X1 U487 ( .A1(n1222), .A2(n3986), .ZN(n676) );
  OR2_X1 U488 ( .A1(n1221), .A2(n3985), .ZN(n677) );
  NAND3_X1 U489 ( .A1(n676), .A2(n677), .A3(n3984), .ZN(n3989) );
  BUF_X2 U490 ( .A(n4096), .Z(n1224) );
  BUF_X2 U491 ( .A(n4094), .Z(n1221) );
  BUF_X2 U492 ( .A(n485), .Z(n678) );
  NOR2_X1 U493 ( .A1(n3916), .A2(n438), .ZN(n3928) );
  OR2_X1 U494 ( .A1(n812), .A2(n1239), .ZN(n679) );
  OR2_X1 U495 ( .A1(n3915), .A2(n1236), .ZN(n680) );
  OR2_X1 U496 ( .A1(n1233), .A2(n3914), .ZN(n681) );
  NAND3_X1 U497 ( .A1(n680), .A2(n679), .A3(n681), .ZN(n3916) );
  BUF_X2 U498 ( .A(n4108), .Z(n1239) );
  BUF_X2 U499 ( .A(n4106), .Z(n1236) );
  BUF_X2 U500 ( .A(n4105), .Z(n1233) );
  AND2_X1 U501 ( .A1(n1028), .A2(n468), .ZN(n783) );
  NOR2_X1 U502 ( .A1(n3590), .A2(n464), .ZN(n3602) );
  AND2_X1 U503 ( .A1(n1155), .A2(n4883), .ZN(n682) );
  AND2_X1 U504 ( .A1(n1151), .A2(n4110), .ZN(n683) );
  OR2_X1 U505 ( .A1(n2185), .A2(n1141), .ZN(n684) );
  OR2_X1 U506 ( .A1(n102), .A2(n1138), .ZN(n685) );
  NAND3_X1 U507 ( .A1(n684), .A2(n685), .A3(n2184), .ZN(n2186) );
  BUF_X2 U508 ( .A(n2214), .Z(n1141) );
  BUF_X2 U509 ( .A(n2213), .Z(n1138) );
  NAND3_X1 U510 ( .A1(n472), .A2(n4057), .A3(n4058), .ZN(n2567) );
  NAND3_X1 U511 ( .A1(n4032), .A2(n4031), .A3(n469), .ZN(n2566) );
  AND2_X1 U512 ( .A1(n4880), .A2(n1244), .ZN(n686) );
  AND2_X1 U513 ( .A1(n1242), .A2(n4021), .ZN(n687) );
  AND4_X1 U514 ( .A1(n978), .A2(n171), .A3(n1186), .A4(n875), .ZN(n982) );
  CLKBUF_X3 U515 ( .A(n4099), .Z(n1229) );
  BUF_X1 U516 ( .A(n968), .Z(n688) );
  AND2_X2 U517 ( .A1(n2265), .A2(n884), .ZN(n968) );
  AND2_X1 U518 ( .A1(n884), .A2(n1036), .ZN(n689) );
  AND3_X1 U519 ( .A1(n4652), .A2(n4653), .A3(n4654), .ZN(n690) );
  AND3_X1 U520 ( .A1(n4652), .A2(n4653), .A3(n4654), .ZN(n1005) );
  BUF_X1 U521 ( .A(n483), .Z(n691) );
  AND3_X1 U522 ( .A1(n1054), .A2(ADD_RS1[0]), .A3(n1560), .ZN(n692) );
  NAND2_X1 U523 ( .A1(n1151), .A2(n2360), .ZN(n693) );
  NAND2_X1 U524 ( .A1(n1156), .A2(n4856), .ZN(n694) );
  NOR3_X1 U525 ( .A1(ADD_RS2[0]), .A2(ADD_RS2[4]), .A3(ADD_RS2[3]), .ZN(n695)
         );
  INV_X1 U526 ( .A(ADD_RS2[2]), .ZN(n696) );
  BUF_X2 U527 ( .A(n967), .Z(n697) );
  NOR2_X1 U528 ( .A1(n2240), .A2(ADD_RS2[1]), .ZN(n1036) );
  CLKBUF_X3 U529 ( .A(n2225), .Z(n1157) );
  CLKBUF_X3 U530 ( .A(n2225), .Z(n1158) );
  AND2_X1 U531 ( .A1(n1166), .A2(n4791), .ZN(n698) );
  AND2_X1 U532 ( .A1(n1163), .A2(n4336), .ZN(n699) );
  NOR3_X1 U533 ( .A1(n698), .A2(n699), .A3(n1632), .ZN(n1637) );
  BUF_X2 U534 ( .A(n991), .Z(n1166) );
  BUF_X2 U535 ( .A(n996), .Z(n1163) );
  BUF_X1 U536 ( .A(n968), .Z(n1197) );
  BUF_X2 U537 ( .A(n481), .Z(n1124) );
  AND2_X1 U538 ( .A1(n4862), .A2(n1243), .ZN(n700) );
  AND2_X1 U539 ( .A1(n1240), .A2(n3566), .ZN(n701) );
  NOR3_X1 U540 ( .A1(n3565), .A2(n701), .A3(n700), .ZN(n3577) );
  CLKBUF_X2 U541 ( .A(n2220), .Z(n1143) );
  CLKBUF_X3 U542 ( .A(n2230), .Z(n1176) );
  AND2_X1 U543 ( .A1(n1036), .A2(n695), .ZN(n879) );
  BUF_X2 U544 ( .A(n2220), .Z(n1144) );
  INV_X1 U545 ( .A(n2241), .ZN(n703) );
  NAND3_X1 U546 ( .A1(n4084), .A2(n4083), .A3(n471), .ZN(n2568) );
  INV_X1 U547 ( .A(ADD_RS1[3]), .ZN(n706) );
  BUF_X1 U548 ( .A(n2226), .Z(n707) );
  AND2_X1 U549 ( .A1(n4867), .A2(n463), .ZN(n708) );
  AND2_X1 U550 ( .A1(n1241), .A2(n3691), .ZN(n709) );
  AND2_X1 U551 ( .A1(n883), .A2(n973), .ZN(n710) );
  AND2_X1 U552 ( .A1(n1181), .A2(n4266), .ZN(n711) );
  AND2_X1 U553 ( .A1(n1178), .A2(n4234), .ZN(n712) );
  NOR3_X1 U554 ( .A1(n711), .A2(n712), .A3(n2004), .ZN(n2007) );
  OR2_X1 U555 ( .A1(n623), .A2(n1176), .ZN(n713) );
  OR2_X1 U556 ( .A1(n3845), .A2(n1172), .ZN(n714) );
  OR2_X1 U557 ( .A1(n3844), .A2(n1169), .ZN(n715) );
  NAND3_X1 U558 ( .A1(n713), .A2(n714), .A3(n715), .ZN(n2004) );
  AND2_X1 U559 ( .A1(n1180), .A2(n4286), .ZN(n716) );
  AND2_X1 U560 ( .A1(n1177), .A2(n4254), .ZN(n717) );
  NOR3_X1 U561 ( .A1(n716), .A2(n717), .A3(n1594), .ZN(n1597) );
  OR2_X1 U562 ( .A1(n643), .A2(n1176), .ZN(n718) );
  OR2_X1 U563 ( .A1(n2289), .A2(n1172), .ZN(n719) );
  OR2_X1 U564 ( .A1(n2288), .A2(n1169), .ZN(n720) );
  NAND3_X1 U565 ( .A1(n718), .A2(n719), .A3(n720), .ZN(n1594) );
  AND2_X1 U566 ( .A1(n1181), .A2(n4268), .ZN(n721) );
  AND2_X1 U567 ( .A1(n1178), .A2(n4236), .ZN(n722) );
  NOR3_X1 U568 ( .A1(n721), .A2(n722), .A3(n1963), .ZN(n1966) );
  OR2_X1 U569 ( .A1(n625), .A2(n1174), .ZN(n723) );
  OR2_X1 U570 ( .A1(n3795), .A2(n1171), .ZN(n724) );
  OR2_X1 U571 ( .A1(n3794), .A2(n1170), .ZN(n725) );
  NAND3_X1 U572 ( .A1(n723), .A2(n724), .A3(n725), .ZN(n1963) );
  AND2_X1 U573 ( .A1(n1168), .A2(n4813), .ZN(n726) );
  AND2_X1 U574 ( .A1(n1165), .A2(n4314), .ZN(n727) );
  NOR3_X1 U575 ( .A1(n726), .A2(n727), .A3(n2087), .ZN(n2092) );
  BUF_X2 U576 ( .A(n991), .Z(n1168) );
  BUF_X2 U577 ( .A(n996), .Z(n1165) );
  AND2_X1 U578 ( .A1(n1181), .A2(n4269), .ZN(n728) );
  AND2_X1 U579 ( .A1(n1178), .A2(n4237), .ZN(n729) );
  NOR3_X1 U580 ( .A1(n728), .A2(n729), .A3(n1943), .ZN(n1946) );
  OR2_X1 U581 ( .A1(n626), .A2(n1174), .ZN(n730) );
  OR2_X1 U582 ( .A1(n3770), .A2(n1172), .ZN(n731) );
  OR2_X1 U583 ( .A1(n3769), .A2(n1170), .ZN(n732) );
  NAND3_X1 U584 ( .A1(n730), .A2(n731), .A3(n732), .ZN(n1943) );
  AND2_X1 U585 ( .A1(n1181), .A2(n4270), .ZN(n733) );
  AND2_X1 U586 ( .A1(n1178), .A2(n4238), .ZN(n734) );
  NOR3_X1 U587 ( .A1(n733), .A2(n734), .A3(n1923), .ZN(n1926) );
  OR2_X1 U588 ( .A1(n627), .A2(n1174), .ZN(n735) );
  OR2_X1 U589 ( .A1(n3745), .A2(n1173), .ZN(n736) );
  OR2_X1 U590 ( .A1(n3744), .A2(n1170), .ZN(n737) );
  NAND3_X1 U591 ( .A1(n735), .A2(n736), .A3(n737), .ZN(n1923) );
  BUF_X1 U592 ( .A(n483), .Z(n738) );
  AND2_X1 U593 ( .A1(n1181), .A2(n4271), .ZN(n740) );
  AND2_X1 U594 ( .A1(n1178), .A2(n4239), .ZN(n741) );
  NOR3_X1 U595 ( .A1(n740), .A2(n741), .A3(n1903), .ZN(n1906) );
  OR2_X1 U596 ( .A1(n628), .A2(n1174), .ZN(n742) );
  OR2_X1 U597 ( .A1(n3720), .A2(n1173), .ZN(n743) );
  OR2_X1 U598 ( .A1(n3719), .A2(n1169), .ZN(n744) );
  NAND3_X1 U599 ( .A1(n742), .A2(n743), .A3(n744), .ZN(n1903) );
  BUF_X2 U600 ( .A(n990), .Z(n1181) );
  BUF_X2 U601 ( .A(n992), .Z(n1178) );
  AND2_X1 U602 ( .A1(n1180), .A2(n4287), .ZN(n745) );
  AND2_X1 U603 ( .A1(n1177), .A2(n4255), .ZN(n746) );
  NOR3_X1 U604 ( .A1(n745), .A2(n746), .A3(n1573), .ZN(n1577) );
  OR2_X1 U605 ( .A1(n644), .A2(n1175), .ZN(n747) );
  OR2_X1 U606 ( .A1(n2262), .A2(n1171), .ZN(n748) );
  OR2_X1 U607 ( .A1(n2261), .A2(n1169), .ZN(n749) );
  NAND3_X1 U608 ( .A1(n747), .A2(n748), .A3(n749), .ZN(n1573) );
  BUF_X2 U609 ( .A(n990), .Z(n1180) );
  BUF_X2 U610 ( .A(n992), .Z(n1177) );
  AND2_X1 U611 ( .A1(n695), .A2(n973), .ZN(n750) );
  OR2_X1 U612 ( .A1(n4093), .A2(n1128), .ZN(n751) );
  OR2_X1 U613 ( .A1(n261), .A2(n485), .ZN(n752) );
  NAND3_X1 U614 ( .A1(n2203), .A2(n752), .A3(n751), .ZN(n2218) );
  OR2_X1 U615 ( .A1(n4063), .A2(n1127), .ZN(n753) );
  OR2_X1 U616 ( .A1(n262), .A2(n485), .ZN(n754) );
  NAND3_X1 U617 ( .A1(n2180), .A2(n754), .A3(n753), .ZN(n2188) );
  BUF_X2 U618 ( .A(n2205), .Z(n1129) );
  INV_X1 U619 ( .A(ADD_RS2[4]), .ZN(n755) );
  BUF_X2 U620 ( .A(n1000), .Z(n1217) );
  INV_X1 U621 ( .A(n84), .ZN(n756) );
  AND2_X1 U622 ( .A1(n1154), .A2(n4881), .ZN(n757) );
  AND2_X1 U623 ( .A1(n1152), .A2(n4047), .ZN(n758) );
  AND2_X2 U624 ( .A1(n880), .A2(n887), .ZN(n759) );
  AND2_X2 U625 ( .A1(n692), .A2(n887), .ZN(n760) );
  AND2_X1 U626 ( .A1(n692), .A2(n887), .ZN(n1029) );
  BUF_X2 U627 ( .A(n1000), .Z(n1218) );
  AND2_X1 U628 ( .A1(n4883), .A2(n1244), .ZN(n761) );
  AND2_X1 U629 ( .A1(n1242), .A2(n4110), .ZN(n762) );
  INV_X1 U630 ( .A(n1554), .ZN(n764) );
  BUF_X1 U631 ( .A(ADD_RS1[4]), .Z(n1092) );
  AND2_X1 U632 ( .A1(n1155), .A2(n4880), .ZN(n765) );
  AND2_X1 U633 ( .A1(n1152), .A2(n4021), .ZN(n766) );
  AND2_X1 U634 ( .A1(n1156), .A2(n4878), .ZN(n767) );
  AND2_X1 U635 ( .A1(n1153), .A2(n3969), .ZN(n768) );
  NAND3_X1 U636 ( .A1(n4006), .A2(n4005), .A3(n222), .ZN(n2565) );
  AND2_X1 U637 ( .A1(n4879), .A2(n1244), .ZN(n769) );
  AND2_X1 U638 ( .A1(n1242), .A2(n3995), .ZN(n770) );
  AND2_X1 U639 ( .A1(n1156), .A2(n4876), .ZN(n771) );
  AND2_X1 U640 ( .A1(n1153), .A2(n3917), .ZN(n772) );
  BUF_X2 U641 ( .A(n982), .Z(n1156) );
  BUF_X2 U642 ( .A(n981), .Z(n1153) );
  NAND3_X1 U643 ( .A1(n3980), .A2(n3979), .A3(n465), .ZN(n2564) );
  AND2_X1 U644 ( .A1(n4878), .A2(n1244), .ZN(n773) );
  AND2_X1 U645 ( .A1(n1242), .A2(n3969), .ZN(n774) );
  NAND3_X1 U646 ( .A1(n3954), .A2(n3953), .A3(n223), .ZN(n2563) );
  AND2_X1 U647 ( .A1(n4877), .A2(n1244), .ZN(n775) );
  AND2_X1 U648 ( .A1(n1242), .A2(n3943), .ZN(n776) );
  NOR3_X1 U649 ( .A1(n3942), .A2(n776), .A3(n775), .ZN(n3954) );
  AND2_X1 U650 ( .A1(n1156), .A2(n4854), .ZN(n777) );
  AND2_X1 U651 ( .A1(n1151), .A2(n2310), .ZN(n778) );
  AND2_X1 U652 ( .A1(n1154), .A2(n4866), .ZN(n779) );
  AND2_X1 U653 ( .A1(n1152), .A2(n3666), .ZN(n780) );
  NAND3_X1 U654 ( .A1(n3928), .A2(n3927), .A3(n466), .ZN(n2562) );
  AND2_X1 U655 ( .A1(n4876), .A2(n1244), .ZN(n781) );
  AND2_X1 U656 ( .A1(n1242), .A2(n3917), .ZN(n782) );
  BUF_X2 U657 ( .A(n984), .Z(n1244) );
  BUF_X2 U658 ( .A(n983), .Z(n1242) );
  BUF_X1 U659 ( .A(ADD_RS1[1]), .Z(n784) );
  AND2_X2 U660 ( .A1(n1028), .A2(n468), .ZN(n969) );
  AND2_X1 U661 ( .A1(n1155), .A2(n4857), .ZN(n785) );
  AND2_X1 U662 ( .A1(n1153), .A2(n2385), .ZN(n786) );
  NAND3_X1 U663 ( .A1(n787), .A2(n788), .A3(n789), .ZN(n2340) );
  OR2_X1 U664 ( .A1(n641), .A2(n1262), .ZN(n787) );
  OR2_X1 U665 ( .A1(n1260), .A2(n2339), .ZN(n788) );
  OR2_X1 U666 ( .A1(n590), .A2(n2338), .ZN(n789) );
  NOR3_X1 U667 ( .A1(n4656), .A2(n4645), .A3(n4657), .ZN(n4655) );
  AND2_X1 U668 ( .A1(n2470), .A2(n2468), .ZN(n790) );
  AND2_X1 U669 ( .A1(n2445), .A2(n2443), .ZN(n791) );
  AND2_X1 U670 ( .A1(n2395), .A2(n2393), .ZN(n792) );
  OR2_X1 U671 ( .A1(n824), .A2(n1149), .ZN(n793) );
  OR2_X1 U672 ( .A1(n1819), .A2(n1146), .ZN(n794) );
  OR2_X1 U673 ( .A1(n3613), .A2(n1143), .ZN(n795) );
  OR2_X1 U674 ( .A1(n833), .A2(n1148), .ZN(n796) );
  OR2_X1 U675 ( .A1(n1631), .A2(n1145), .ZN(n797) );
  OR2_X1 U676 ( .A1(n2332), .A2(n1142), .ZN(n798) );
  OR2_X1 U677 ( .A1(n835), .A2(n1148), .ZN(n799) );
  OR2_X1 U678 ( .A1(n1592), .A2(n1145), .ZN(n800) );
  OR2_X1 U679 ( .A1(n2282), .A2(n1142), .ZN(n801) );
  NOR2_X1 U680 ( .A1(n802), .A2(n803), .ZN(n1599) );
  NAND3_X1 U681 ( .A1(n800), .A2(n799), .A3(n801), .ZN(n802) );
  OR2_X1 U682 ( .A1(n1102), .A2(n1101), .ZN(n803) );
  AND2_X1 U683 ( .A1(n804), .A2(n922), .ZN(n2009) );
  NOR3_X1 U684 ( .A1(n1011), .A2(n1010), .A3(n1012), .ZN(n804) );
  AND2_X1 U685 ( .A1(n869), .A2(n927), .ZN(n1928) );
  NOR3_X1 U686 ( .A1(n1008), .A2(n1007), .A3(n1009), .ZN(n869) );
  NAND3_X1 U687 ( .A1(n870), .A2(n871), .A3(n872), .ZN(n1652) );
  OR2_X1 U688 ( .A1(n1651), .A2(n1145), .ZN(n870) );
  OR2_X1 U689 ( .A1(n832), .A2(n1148), .ZN(n871) );
  OR2_X1 U690 ( .A1(n2357), .A2(n1142), .ZN(n872) );
  BUF_X2 U691 ( .A(n1000), .Z(n1216) );
  BUF_X2 U692 ( .A(n967), .Z(n1199) );
  AND3_X1 U693 ( .A1(n2344), .A2(n2343), .A3(n2345), .ZN(n873) );
  NAND2_X1 U694 ( .A1(n1005), .A2(n1027), .ZN(n874) );
  NAND2_X1 U695 ( .A1(n690), .A2(n77), .ZN(n875) );
  NAND4_X1 U696 ( .A1(n1574), .A2(n705), .A3(n1187), .A4(n978), .ZN(n876) );
  NAND2_X1 U697 ( .A1(n4655), .A2(n1005), .ZN(n1574) );
  CLKBUF_X3 U698 ( .A(n2230), .Z(n1175) );
  CLKBUF_X3 U699 ( .A(n2229), .Z(n1173) );
  CLKBUF_X3 U700 ( .A(n2230), .Z(n1174) );
  AND2_X2 U701 ( .A1(n884), .A2(n1036), .ZN(n998) );
  CLKBUF_X3 U702 ( .A(n2228), .Z(n1170) );
  CLKBUF_X3 U703 ( .A(n2229), .Z(n1172) );
  AND2_X1 U704 ( .A1(n695), .A2(n1036), .ZN(n997) );
  CLKBUF_X3 U705 ( .A(n2228), .Z(n1169) );
  CLKBUF_X3 U706 ( .A(n2229), .Z(n1171) );
  AND3_X1 U707 ( .A1(n1054), .A2(ADD_RS1[0]), .A3(n1560), .ZN(n880) );
  CLKBUF_X1 U708 ( .A(n4116), .Z(n1256) );
  CLKBUF_X3 U709 ( .A(n4116), .Z(n1258) );
  INV_X1 U710 ( .A(ADD_RS1[0]), .ZN(n881) );
  AND3_X1 U711 ( .A1(n882), .A2(n1062), .A3(n2243), .ZN(n883) );
  AND3_X1 U712 ( .A1(n2243), .A2(n882), .A3(n488), .ZN(n884) );
  AND3_X1 U713 ( .A1(n882), .A2(n755), .A3(n1061), .ZN(n1030) );
  CLKBUF_X1 U714 ( .A(ADD_RS2[3]), .Z(n885) );
  AND3_X1 U715 ( .A1(ADD_RS1[0]), .A2(n1054), .A3(n1560), .ZN(n886) );
  BUF_X1 U716 ( .A(n1077), .Z(n1053) );
  CLKBUF_X1 U717 ( .A(ADD_RS1[0]), .Z(n890) );
  CLKBUF_X1 U718 ( .A(n889), .Z(n891) );
  NOR3_X1 U719 ( .A1(n4650), .A2(n4651), .A3(n4645), .ZN(n893) );
  NOR3_X1 U720 ( .A1(n4650), .A2(n4651), .A3(n4645), .ZN(n4649) );
  BUF_X2 U721 ( .A(n967), .Z(n1200) );
  BUF_X2 U722 ( .A(n997), .Z(n1209) );
  CLKBUF_X3 U723 ( .A(n4118), .Z(n1259) );
  BUF_X2 U724 ( .A(n997), .Z(n1208) );
  BUF_X2 U725 ( .A(n481), .Z(n1024) );
  AND2_X1 U726 ( .A1(n1155), .A2(n4863), .ZN(n894) );
  AND2_X1 U727 ( .A1(n1153), .A2(n3591), .ZN(n895) );
  AND2_X1 U728 ( .A1(n4857), .A2(n1243), .ZN(n896) );
  AND2_X1 U729 ( .A1(n1240), .A2(n2385), .ZN(n897) );
  BUF_X2 U730 ( .A(n984), .Z(n1243) );
  BUF_X2 U731 ( .A(n983), .Z(n1240) );
  AND2_X1 U732 ( .A1(n1154), .A2(n4862), .ZN(n898) );
  AND2_X1 U733 ( .A1(n1151), .A2(n3566), .ZN(n899) );
  AND2_X1 U734 ( .A1(n1154), .A2(n4875), .ZN(n900) );
  AND2_X1 U735 ( .A1(n1151), .A2(n3891), .ZN(n901) );
  AND2_X1 U736 ( .A1(n1155), .A2(n4861), .ZN(n902) );
  AND2_X1 U737 ( .A1(n1153), .A2(n2485), .ZN(n903) );
  BUF_X2 U738 ( .A(n981), .Z(n1151) );
  AND2_X1 U739 ( .A1(n1155), .A2(n4874), .ZN(n904) );
  AND2_X1 U740 ( .A1(n1151), .A2(n3866), .ZN(n905) );
  AND2_X1 U741 ( .A1(n4875), .A2(n463), .ZN(n906) );
  AND2_X1 U742 ( .A1(n1241), .A2(n3891), .ZN(n907) );
  AND2_X1 U743 ( .A1(n4874), .A2(n463), .ZN(n908) );
  AND2_X1 U744 ( .A1(n1241), .A2(n3866), .ZN(n909) );
  AND2_X1 U745 ( .A1(n1156), .A2(n4872), .ZN(n910) );
  AND2_X1 U746 ( .A1(n1152), .A2(n3816), .ZN(n911) );
  BUF_X2 U747 ( .A(n982), .Z(n1155) );
  BUF_X2 U748 ( .A(n981), .Z(n1152) );
  AND2_X1 U749 ( .A1(n4873), .A2(n463), .ZN(n912) );
  AND2_X1 U750 ( .A1(n1241), .A2(n3841), .ZN(n913) );
  AND2_X1 U751 ( .A1(n4872), .A2(n463), .ZN(n914) );
  AND2_X1 U752 ( .A1(n1241), .A2(n3816), .ZN(n915) );
  AND2_X1 U753 ( .A1(n4871), .A2(n463), .ZN(n916) );
  AND2_X1 U754 ( .A1(n1241), .A2(n3791), .ZN(n917) );
  BUF_X2 U755 ( .A(n983), .Z(n1241) );
  AND2_X1 U756 ( .A1(n4870), .A2(n463), .ZN(n918) );
  AND2_X1 U757 ( .A1(n1241), .A2(n3766), .ZN(n919) );
  AND2_X1 U758 ( .A1(n4869), .A2(n463), .ZN(n920) );
  AND2_X1 U759 ( .A1(n1241), .A2(n3741), .ZN(n921) );
  NOR2_X1 U760 ( .A1(n1033), .A2(n1032), .ZN(n922) );
  AND2_X1 U761 ( .A1(n4868), .A2(n463), .ZN(n923) );
  AND2_X1 U762 ( .A1(n1241), .A2(n3716), .ZN(n924) );
  NAND2_X1 U763 ( .A1(n1006), .A2(n893), .ZN(n925) );
  NAND2_X1 U764 ( .A1(n4649), .A2(n470), .ZN(n926) );
  NAND2_X1 U765 ( .A1(n1006), .A2(n4649), .ZN(n2264) );
  NOR2_X1 U766 ( .A1(n1079), .A2(n1078), .ZN(n927) );
  NOR2_X1 U767 ( .A1(n1652), .A2(n352), .ZN(n1659) );
  OR2_X1 U768 ( .A1(n1134), .A2(n3832), .ZN(n928) );
  OR2_X1 U769 ( .A1(n239), .A2(n1132), .ZN(n929) );
  NAND3_X1 U770 ( .A1(n928), .A2(n929), .A3(n1994), .ZN(n1999) );
  BUF_X2 U771 ( .A(n982), .Z(n1154) );
  CLKBUF_X1 U772 ( .A(n1004), .Z(n1276) );
  BUF_X2 U773 ( .A(n1004), .Z(n1275) );
  BUF_X1 U774 ( .A(n1539), .Z(n1538) );
  BUF_X1 U775 ( .A(n483), .Z(n1113) );
  BUF_X1 U776 ( .A(n484), .Z(n1112) );
  BUF_X1 U777 ( .A(n484), .Z(n1111) );
  BUF_X1 U778 ( .A(n1449), .Z(n1539) );
  BUF_X1 U779 ( .A(n1449), .Z(n1540) );
  BUF_X1 U780 ( .A(n1449), .Z(n1541) );
  BUF_X1 U781 ( .A(n1450), .Z(n1542) );
  BUF_X1 U782 ( .A(n1450), .Z(n1543) );
  BUF_X1 U783 ( .A(n1450), .Z(n1544) );
  BUF_X1 U784 ( .A(n1451), .Z(n1545) );
  BUF_X1 U785 ( .A(n1451), .Z(n1546) );
  BUF_X1 U786 ( .A(n1451), .Z(n1547) );
  BUF_X1 U787 ( .A(n1452), .Z(n1548) );
  BUF_X1 U788 ( .A(n1452), .Z(n1549) );
  BUF_X1 U789 ( .A(n1452), .Z(n1550) );
  BUF_X1 U790 ( .A(n1453), .Z(n1551) );
  BUF_X1 U791 ( .A(n1453), .Z(n1552) );
  BUF_X2 U792 ( .A(n4096), .Z(n1223) );
  BUF_X2 U793 ( .A(n4096), .Z(n1222) );
  BUF_X1 U794 ( .A(n985), .Z(n1266) );
  BUF_X1 U795 ( .A(n994), .Z(n1278) );
  BUF_X1 U796 ( .A(n996), .Z(n1164) );
  BUF_X1 U797 ( .A(n993), .Z(n1190) );
  BUF_X1 U798 ( .A(n993), .Z(n1191) );
  BUF_X1 U799 ( .A(n989), .Z(n1251) );
  BUF_X1 U800 ( .A(n994), .Z(n1279) );
  BUF_X1 U801 ( .A(n977), .Z(n1254) );
  BUF_X1 U802 ( .A(n988), .Z(n1282) );
  BUF_X1 U803 ( .A(n986), .Z(n1269) );
  BUF_X1 U804 ( .A(n991), .Z(n1167) );
  BUF_X1 U805 ( .A(n995), .Z(n1193) );
  BUF_X1 U806 ( .A(n995), .Z(n1194) );
  BUF_X2 U807 ( .A(n4094), .Z(n1220) );
  BUF_X2 U808 ( .A(n4094), .Z(n1219) );
  AND2_X1 U809 ( .A1(n1002), .A2(n1572), .ZN(n930) );
  BUF_X1 U810 ( .A(n4113), .Z(n1249) );
  BUF_X1 U811 ( .A(n4111), .Z(n1247) );
  BUF_X1 U812 ( .A(n989), .Z(n1252) );
  BUF_X1 U813 ( .A(n993), .Z(n1192) );
  BUF_X1 U814 ( .A(n994), .Z(n1280) );
  BUF_X1 U815 ( .A(n977), .Z(n1255) );
  BUF_X1 U816 ( .A(n2226), .Z(n1162) );
  BUF_X1 U817 ( .A(n4091), .Z(n1215) );
  BUF_X1 U818 ( .A(n4090), .Z(n1212) );
  BUF_X1 U819 ( .A(n995), .Z(n1195) );
  AND2_X1 U820 ( .A1(n973), .A2(n695), .ZN(n931) );
  AND3_X1 U821 ( .A1(n763), .A2(n1572), .A3(n756), .ZN(n971) );
  BUF_X1 U822 ( .A(n1454), .Z(n1451) );
  BUF_X1 U823 ( .A(n1454), .Z(n1452) );
  BUF_X1 U824 ( .A(n1455), .Z(n1449) );
  BUF_X1 U825 ( .A(n1455), .Z(n1450) );
  BUF_X1 U826 ( .A(n1454), .Z(n1453) );
  AND2_X2 U827 ( .A1(n696), .A2(ADD_RS2[1]), .ZN(n973) );
  BUF_X1 U828 ( .A(n4576), .Z(n1362) );
  BUF_X1 U829 ( .A(n4576), .Z(n1363) );
  BUF_X1 U830 ( .A(n4611), .Z(n1371) );
  BUF_X1 U831 ( .A(n4611), .Z(n1372) );
  BUF_X1 U832 ( .A(n4359), .Z(n1305) );
  BUF_X1 U833 ( .A(n4359), .Z(n1306) );
  BUF_X1 U834 ( .A(n4499), .Z(n1332) );
  BUF_X1 U835 ( .A(n4499), .Z(n1333) );
  BUF_X1 U836 ( .A(n4394), .Z(n1308) );
  BUF_X1 U837 ( .A(n4394), .Z(n1309) );
  BUF_X1 U838 ( .A(n4534), .Z(n1341) );
  BUF_X1 U839 ( .A(n4534), .Z(n1342) );
  BUF_X1 U840 ( .A(n4462), .Z(n1320) );
  BUF_X1 U841 ( .A(n4462), .Z(n1321) );
  BUF_X1 U842 ( .A(n4429), .Z(n1317) );
  BUF_X1 U843 ( .A(n4429), .Z(n1318) );
  BUF_X1 U844 ( .A(n4569), .Z(n1353) );
  BUF_X1 U845 ( .A(n4569), .Z(n1354) );
  BUF_X1 U846 ( .A(n4573), .Z(n1359) );
  BUF_X1 U847 ( .A(n4573), .Z(n1360) );
  BUF_X1 U848 ( .A(n4571), .Z(n1356) );
  BUF_X1 U849 ( .A(n4571), .Z(n1357) );
  BUF_X1 U850 ( .A(n4643), .Z(n1374) );
  BUF_X1 U851 ( .A(n4643), .Z(n1375) );
  BUF_X1 U852 ( .A(n4609), .Z(n1368) );
  BUF_X1 U853 ( .A(n4609), .Z(n1369) );
  BUF_X1 U854 ( .A(n4608), .Z(n1365) );
  BUF_X1 U855 ( .A(n4608), .Z(n1366) );
  BUF_X1 U856 ( .A(n4496), .Z(n1329) );
  BUF_X1 U857 ( .A(n4496), .Z(n1330) );
  BUF_X1 U858 ( .A(n4532), .Z(n1338) );
  BUF_X1 U859 ( .A(n4532), .Z(n1339) );
  BUF_X1 U860 ( .A(n4531), .Z(n1335) );
  BUF_X1 U861 ( .A(n4531), .Z(n1336) );
  BUF_X1 U862 ( .A(n4427), .Z(n1314) );
  BUF_X1 U863 ( .A(n4427), .Z(n1315) );
  BUF_X1 U864 ( .A(n4426), .Z(n1311) );
  BUF_X1 U865 ( .A(n4426), .Z(n1312) );
  BUF_X1 U866 ( .A(n4568), .Z(n1350) );
  BUF_X1 U867 ( .A(n4568), .Z(n1351) );
  BUF_X1 U868 ( .A(n4567), .Z(n1347) );
  BUF_X1 U869 ( .A(n4567), .Z(n1348) );
  BUF_X1 U870 ( .A(n4566), .Z(n1344) );
  BUF_X1 U871 ( .A(n4566), .Z(n1345) );
  BUF_X1 U872 ( .A(n4495), .Z(n1326) );
  BUF_X1 U873 ( .A(n4495), .Z(n1327) );
  BUF_X1 U874 ( .A(n4494), .Z(n1323) );
  BUF_X1 U875 ( .A(n4494), .Z(n1324) );
  BUF_X1 U876 ( .A(n4345), .Z(n1290) );
  BUF_X1 U877 ( .A(n4345), .Z(n1291) );
  BUF_X1 U878 ( .A(n4343), .Z(n1287) );
  BUF_X1 U879 ( .A(n4343), .Z(n1288) );
  BUF_X1 U880 ( .A(n4340), .Z(n1284) );
  BUF_X1 U881 ( .A(n4340), .Z(n1285) );
  BUF_X1 U882 ( .A(n4353), .Z(n1302) );
  BUF_X1 U883 ( .A(n4353), .Z(n1303) );
  BUF_X1 U884 ( .A(n4351), .Z(n1299) );
  BUF_X1 U885 ( .A(n4351), .Z(n1300) );
  BUF_X1 U886 ( .A(n4349), .Z(n1296) );
  BUF_X1 U887 ( .A(n4349), .Z(n1297) );
  BUF_X1 U888 ( .A(n4347), .Z(n1293) );
  BUF_X1 U889 ( .A(n4347), .Z(n1294) );
  BUF_X1 U890 ( .A(n1004), .Z(n1274) );
  BUF_X2 U891 ( .A(n4121), .Z(n1271) );
  BUF_X2 U892 ( .A(n2232), .Z(n1183) );
  BUF_X2 U893 ( .A(n2232), .Z(n1184) );
  BUF_X2 U894 ( .A(n4121), .Z(n1272) );
  BUF_X1 U895 ( .A(n1004), .Z(n1277) );
  BUF_X1 U896 ( .A(n1003), .Z(n1189) );
  BUF_X1 U897 ( .A(n1003), .Z(n1188) );
  AND3_X1 U898 ( .A1(ADD_RS2[3]), .A2(n755), .A3(n882), .ZN(n974) );
  AND3_X1 U899 ( .A1(ADD_RS2[3]), .A2(n2259), .A3(n2243), .ZN(n975) );
  AND2_X1 U900 ( .A1(ADD_RS2[3]), .A2(n999), .ZN(n976) );
  AND4_X1 U901 ( .A1(n703), .A2(n473), .A3(n1274), .A4(n926), .ZN(n977) );
  AND3_X1 U902 ( .A1(n763), .A2(ADD_RS1[0]), .A3(n756), .ZN(n978) );
  AND2_X1 U903 ( .A1(n999), .A2(n1062), .ZN(n979) );
  AND3_X1 U904 ( .A1(n2259), .A2(n885), .A3(n891), .ZN(n980) );
  BUF_X1 U905 ( .A(n4576), .Z(n1364) );
  BUF_X1 U906 ( .A(n4611), .Z(n1373) );
  BUF_X1 U907 ( .A(n4359), .Z(n1307) );
  BUF_X1 U908 ( .A(n4499), .Z(n1334) );
  BUF_X1 U909 ( .A(n4394), .Z(n1310) );
  BUF_X1 U910 ( .A(n4534), .Z(n1343) );
  BUF_X1 U911 ( .A(n4462), .Z(n1322) );
  BUF_X1 U912 ( .A(n4429), .Z(n1319) );
  BUF_X1 U913 ( .A(n4569), .Z(n1355) );
  BUF_X1 U914 ( .A(n4573), .Z(n1361) );
  BUF_X1 U915 ( .A(n4571), .Z(n1358) );
  BUF_X1 U916 ( .A(n4643), .Z(n1376) );
  BUF_X1 U917 ( .A(n4609), .Z(n1370) );
  BUF_X1 U918 ( .A(n4608), .Z(n1367) );
  BUF_X1 U919 ( .A(n4496), .Z(n1331) );
  BUF_X1 U920 ( .A(n4532), .Z(n1340) );
  BUF_X1 U921 ( .A(n4531), .Z(n1337) );
  BUF_X1 U922 ( .A(n4427), .Z(n1316) );
  BUF_X1 U923 ( .A(n4426), .Z(n1313) );
  BUF_X1 U924 ( .A(n4345), .Z(n1292) );
  BUF_X1 U925 ( .A(n4343), .Z(n1289) );
  BUF_X1 U926 ( .A(n4340), .Z(n1286) );
  BUF_X1 U927 ( .A(n4568), .Z(n1352) );
  BUF_X1 U928 ( .A(n4567), .Z(n1349) );
  BUF_X1 U929 ( .A(n4566), .Z(n1346) );
  BUF_X1 U930 ( .A(n4495), .Z(n1328) );
  BUF_X1 U931 ( .A(n4494), .Z(n1325) );
  BUF_X1 U932 ( .A(n4353), .Z(n1304) );
  BUF_X1 U933 ( .A(n4351), .Z(n1301) );
  BUF_X1 U934 ( .A(n4349), .Z(n1298) );
  BUF_X1 U935 ( .A(n4347), .Z(n1295) );
  AND4_X1 U936 ( .A1(n874), .A2(n172), .A3(n1186), .A4(n705), .ZN(n981) );
  AND4_X1 U937 ( .A1(n473), .A2(n973), .A3(n1274), .A4(n925), .ZN(n983) );
  AND4_X1 U938 ( .A1(n979), .A2(n2260), .A3(n1274), .A4(n926), .ZN(n984) );
  BUF_X1 U939 ( .A(n2232), .Z(n1185) );
  BUF_X1 U940 ( .A(n4121), .Z(n1273) );
  AND4_X1 U941 ( .A1(n1001), .A2(n703), .A3(n1274), .A4(n925), .ZN(n985) );
  AND4_X1 U942 ( .A1(n979), .A2(n878), .A3(n1274), .A4(n925), .ZN(n986) );
  AND4_X1 U943 ( .A1(n1001), .A2(n973), .A3(n1275), .A4(n925), .ZN(n988) );
  AND4_X1 U944 ( .A1(n473), .A2(n2260), .A3(n1274), .A4(n925), .ZN(n989) );
  AND4_X1 U945 ( .A1(n1574), .A2(n887), .A3(n1186), .A4(n978), .ZN(n990) );
  AND4_X1 U946 ( .A1(n172), .A2(n468), .A3(n1186), .A4(n875), .ZN(n991) );
  AND4_X1 U947 ( .A1(n1574), .A2(n468), .A3(n1186), .A4(n971), .ZN(n992) );
  AND4_X1 U948 ( .A1(n978), .A2(n468), .A3(n1187), .A4(n875), .ZN(n993) );
  AND4_X1 U949 ( .A1(n979), .A2(n703), .A3(n1275), .A4(n926), .ZN(n994) );
  AND4_X1 U950 ( .A1(n1574), .A2(n705), .A3(n1187), .A4(n971), .ZN(n995) );
  AND4_X1 U951 ( .A1(n172), .A2(n171), .A3(n1186), .A4(n875), .ZN(n996) );
  AND2_X1 U952 ( .A1(n889), .A2(n882), .ZN(n999) );
  AND3_X1 U953 ( .A1(n891), .A2(n2259), .A3(n1062), .ZN(n1001) );
  AND2_X1 U954 ( .A1(ADD_RS1[4]), .A2(ADD_RS1[3]), .ZN(n1002) );
  BUF_X1 U955 ( .A(RST), .Z(n1454) );
  BUF_X1 U956 ( .A(RST), .Z(n1455) );
  AND2_X1 U957 ( .A1(RD1), .A2(n462), .ZN(n1003) );
  AND2_X1 U958 ( .A1(RD2), .A2(n462), .ZN(n1004) );
  INV_X1 U959 ( .A(DATAIN[0]), .ZN(n1378) );
  INV_X1 U960 ( .A(DATAIN[1]), .ZN(n1380) );
  INV_X1 U961 ( .A(DATAIN[2]), .ZN(n1382) );
  INV_X1 U962 ( .A(DATAIN[3]), .ZN(n1384) );
  INV_X1 U963 ( .A(DATAIN[4]), .ZN(n1386) );
  INV_X1 U964 ( .A(DATAIN[5]), .ZN(n1388) );
  INV_X1 U965 ( .A(DATAIN[6]), .ZN(n1390) );
  INV_X1 U966 ( .A(DATAIN[7]), .ZN(n1392) );
  INV_X1 U967 ( .A(DATAIN[8]), .ZN(n1394) );
  INV_X1 U968 ( .A(DATAIN[12]), .ZN(n1402) );
  INV_X1 U969 ( .A(DATAIN[13]), .ZN(n1404) );
  INV_X1 U970 ( .A(DATAIN[14]), .ZN(n1406) );
  INV_X1 U971 ( .A(DATAIN[15]), .ZN(n1408) );
  INV_X1 U972 ( .A(DATAIN[16]), .ZN(n1410) );
  INV_X1 U973 ( .A(DATAIN[17]), .ZN(n1412) );
  INV_X1 U974 ( .A(DATAIN[18]), .ZN(n1414) );
  INV_X1 U975 ( .A(DATAIN[19]), .ZN(n1416) );
  INV_X1 U976 ( .A(DATAIN[21]), .ZN(n1420) );
  INV_X1 U977 ( .A(DATAIN[22]), .ZN(n1422) );
  INV_X1 U978 ( .A(DATAIN[23]), .ZN(n1424) );
  INV_X1 U979 ( .A(DATAIN[25]), .ZN(n1430) );
  INV_X1 U980 ( .A(DATAIN[26]), .ZN(n1433) );
  INV_X1 U981 ( .A(DATAIN[27]), .ZN(n1436) );
  INV_X1 U982 ( .A(DATAIN[28]), .ZN(n1439) );
  INV_X1 U983 ( .A(DATAIN[29]), .ZN(n1442) );
  INV_X1 U984 ( .A(DATAIN[30]), .ZN(n1445) );
  INV_X1 U985 ( .A(DATAIN[31]), .ZN(n1448) );
  INV_X1 U986 ( .A(DATAIN[10]), .ZN(n1398) );
  INV_X1 U987 ( .A(DATAIN[20]), .ZN(n1418) );
  INV_X1 U988 ( .A(DATAIN[24]), .ZN(n1427) );
  INV_X1 U989 ( .A(DATAIN[11]), .ZN(n1400) );
  INV_X1 U990 ( .A(DATAIN[9]), .ZN(n1396) );
  AOI221_X1 U991 ( .B1(n1268), .B2(n4280), .C1(n1265), .C2(n4248), .A(n2440), 
        .ZN(n2444) );
  AOI221_X1 U992 ( .B1(n1268), .B2(n4279), .C1(n1265), .C2(n4247), .A(n2465), 
        .ZN(n2469) );
  AOI221_X1 U993 ( .B1(n1268), .B2(n4282), .C1(n1265), .C2(n4250), .A(n2390), 
        .ZN(n2394) );
  NOR2_X1 U994 ( .A1(n819), .A2(n1149), .ZN(n1007) );
  NOR2_X1 U995 ( .A1(n1921), .A2(n1146), .ZN(n1008) );
  NOR2_X1 U996 ( .A1(n3738), .A2(n1143), .ZN(n1009) );
  NOR2_X1 U997 ( .A1(n815), .A2(n1149), .ZN(n1010) );
  NOR2_X1 U998 ( .A1(n2002), .A2(n1146), .ZN(n1011) );
  NOR2_X1 U999 ( .A1(n3838), .A2(n1143), .ZN(n1012) );
  AND3_X1 U1000 ( .A1(n3574), .A2(n3575), .A3(n3576), .ZN(n1013) );
  AND2_X1 U1001 ( .A1(n1268), .A2(n4277), .ZN(n1017) );
  AND2_X1 U1002 ( .A1(n1265), .A2(n4245), .ZN(n1018) );
  NOR3_X1 U1003 ( .A1(n1017), .A2(n1018), .A3(n3571), .ZN(n3575) );
  OR2_X1 U1004 ( .A1(n634), .A2(n1262), .ZN(n1019) );
  OR2_X1 U1005 ( .A1(n1261), .A2(n3570), .ZN(n1020) );
  OR2_X1 U1006 ( .A1(n590), .A2(n3569), .ZN(n1021) );
  NAND3_X1 U1007 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n3571) );
  NOR3_X1 U1008 ( .A1(n1092), .A2(n706), .A3(ADD_RS1[0]), .ZN(n1077) );
  AND3_X1 U1009 ( .A1(n2494), .A2(n2493), .A3(n2495), .ZN(n1022) );
  BUF_X1 U1010 ( .A(n877), .Z(n1023) );
  BUF_X1 U1011 ( .A(n877), .Z(n1122) );
  AND2_X1 U1012 ( .A1(n1268), .A2(n4284), .ZN(n1025) );
  AND2_X1 U1013 ( .A1(n1265), .A2(n4252), .ZN(n1026) );
  NOR3_X1 U1014 ( .A1(n1025), .A2(n1026), .A3(n2340), .ZN(n2344) );
  NOR3_X1 U1015 ( .A1(n4656), .A2(n4645), .A3(n4657), .ZN(n1027) );
  AND2_X1 U1016 ( .A1(n1155), .A2(n4873), .ZN(n1032) );
  AND2_X1 U1017 ( .A1(n1153), .A2(n3841), .ZN(n1033) );
  OR2_X1 U1018 ( .A1(n373), .A2(n1214), .ZN(n1034) );
  OR2_X1 U1019 ( .A1(n405), .A2(n1211), .ZN(n1035) );
  NAND3_X1 U1020 ( .A1(n1034), .A2(n1035), .A3(n3679), .ZN(n3686) );
  AND2_X1 U1021 ( .A1(n4866), .A2(n463), .ZN(n1037) );
  AND2_X1 U1022 ( .A1(n1241), .A2(n3666), .ZN(n1038) );
  OR2_X1 U1023 ( .A1(n1228), .A2(n457), .ZN(n1039) );
  OR2_X1 U1024 ( .A1(n1226), .A2(n458), .ZN(n1040) );
  NAND3_X1 U1025 ( .A1(n1039), .A2(n1040), .A3(n3633), .ZN(n3634) );
  AND2_X1 U1026 ( .A1(n4865), .A2(n463), .ZN(n1041) );
  AND2_X1 U1027 ( .A1(n1241), .A2(n3641), .ZN(n1042) );
  AND2_X1 U1028 ( .A1(n4864), .A2(n463), .ZN(n1043) );
  AND2_X1 U1029 ( .A1(n1241), .A2(n3616), .ZN(n1044) );
  OR2_X1 U1030 ( .A1(n1229), .A2(n459), .ZN(n1045) );
  OR2_X1 U1031 ( .A1(n1225), .A2(n460), .ZN(n1046) );
  NAND3_X1 U1032 ( .A1(n1045), .A2(n1046), .A3(n3583), .ZN(n3584) );
  AND2_X1 U1033 ( .A1(n4863), .A2(n1243), .ZN(n1047) );
  AND2_X1 U1034 ( .A1(n1240), .A2(n3591), .ZN(n1048) );
  NAND2_X1 U1035 ( .A1(n1013), .A2(n3577), .ZN(n2548) );
  AND2_X1 U1036 ( .A1(n1156), .A2(n4879), .ZN(n1049) );
  AND2_X1 U1037 ( .A1(n1153), .A2(n3995), .ZN(n1050) );
  AND2_X1 U1038 ( .A1(n1156), .A2(n4877), .ZN(n1051) );
  AND2_X1 U1039 ( .A1(n1151), .A2(n3943), .ZN(n1052) );
  NAND2_X1 U1040 ( .A1(n2496), .A2(n1022), .ZN(n2547) );
  AND2_X1 U1041 ( .A1(n4861), .A2(n1243), .ZN(n1055) );
  AND2_X1 U1042 ( .A1(n1240), .A2(n2485), .ZN(n1056) );
  NOR3_X1 U1043 ( .A1(n2484), .A2(n1056), .A3(n1055), .ZN(n2496) );
  AND2_X1 U1044 ( .A1(n1155), .A2(n4860), .ZN(n1057) );
  AND2_X1 U1045 ( .A1(n1152), .A2(n2460), .ZN(n1058) );
  AND2_X1 U1046 ( .A1(n1154), .A2(n4859), .ZN(n1059) );
  AND2_X1 U1047 ( .A1(n1153), .A2(n2435), .ZN(n1060) );
  INV_X1 U1048 ( .A(ADD_RS2[3]), .ZN(n1061) );
  INV_X1 U1049 ( .A(ADD_RS2[3]), .ZN(n1062) );
  NAND3_X1 U1050 ( .A1(n790), .A2(n2471), .A3(n2469), .ZN(n2546) );
  AND2_X1 U1051 ( .A1(n4860), .A2(n1243), .ZN(n1063) );
  AND2_X1 U1052 ( .A1(n1240), .A2(n2460), .ZN(n1064) );
  AND2_X1 U1053 ( .A1(n1154), .A2(n4858), .ZN(n1065) );
  AND2_X1 U1054 ( .A1(n1152), .A2(n2410), .ZN(n1066) );
  AND2_X1 U1055 ( .A1(n1154), .A2(n4871), .ZN(n1067) );
  AND2_X1 U1056 ( .A1(n1151), .A2(n3791), .ZN(n1068) );
  NAND3_X1 U1057 ( .A1(n2446), .A2(n791), .A3(n2444), .ZN(n2545) );
  AND2_X1 U1058 ( .A1(n4859), .A2(n1243), .ZN(n1069) );
  AND2_X1 U1059 ( .A1(n1240), .A2(n2435), .ZN(n1070) );
  AND2_X1 U1060 ( .A1(n4858), .A2(n1243), .ZN(n1071) );
  AND2_X1 U1061 ( .A1(n1240), .A2(n2410), .ZN(n1072) );
  OR2_X1 U1062 ( .A1(n2376), .A2(n1134), .ZN(n1073) );
  OR2_X1 U1063 ( .A1(n255), .A2(n1132), .ZN(n1074) );
  NAND3_X1 U1064 ( .A1(n1073), .A2(n1074), .A3(n1664), .ZN(n1669) );
  AND2_X1 U1065 ( .A1(n1155), .A2(n4870), .ZN(n1075) );
  AND2_X1 U1066 ( .A1(n1152), .A2(n3766), .ZN(n1076) );
  AND2_X1 U1067 ( .A1(n1154), .A2(n4869), .ZN(n1078) );
  AND2_X1 U1068 ( .A1(n1152), .A2(n3741), .ZN(n1079) );
  OR2_X1 U1069 ( .A1(n1895), .A2(n1140), .ZN(n1080) );
  OR2_X1 U1070 ( .A1(n116), .A2(n1137), .ZN(n1081) );
  NAND3_X1 U1071 ( .A1(n1894), .A2(n1081), .A3(n1080), .ZN(n1896) );
  AND2_X1 U1072 ( .A1(n1154), .A2(n4868), .ZN(n1082) );
  AND2_X1 U1073 ( .A1(n1152), .A2(n3716), .ZN(n1083) );
  NOR3_X1 U1074 ( .A1(n1901), .A2(n1083), .A3(n1082), .ZN(n1908) );
  AND2_X1 U1075 ( .A1(n1155), .A2(n4867), .ZN(n1084) );
  AND2_X1 U1076 ( .A1(n1153), .A2(n3691), .ZN(n1085) );
  NOR3_X1 U1077 ( .A1(n1880), .A2(n1085), .A3(n1084), .ZN(n1887) );
  AND2_X1 U1078 ( .A1(n1154), .A2(n4855), .ZN(n1086) );
  AND2_X1 U1079 ( .A1(n1152), .A2(n2335), .ZN(n1087) );
  OR2_X1 U1080 ( .A1(n3657), .A2(n1134), .ZN(n1088) );
  OR2_X1 U1081 ( .A1(n1132), .A2(n246), .ZN(n1089) );
  NAND3_X1 U1082 ( .A1(n1088), .A2(n1089), .A3(n1852), .ZN(n1857) );
  NAND3_X1 U1083 ( .A1(n792), .A2(n2396), .A3(n2394), .ZN(n2543) );
  AND2_X1 U1084 ( .A1(n1156), .A2(n4865), .ZN(n1090) );
  AND2_X1 U1085 ( .A1(n1151), .A2(n3641), .ZN(n1091) );
  NOR3_X1 U1086 ( .A1(n1840), .A2(n1091), .A3(n1090), .ZN(n1847) );
  OR2_X1 U1087 ( .A1(n2301), .A2(n1134), .ZN(n1093) );
  OR2_X1 U1088 ( .A1(n258), .A2(n1132), .ZN(n1094) );
  NAND3_X1 U1089 ( .A1(n1093), .A2(n1094), .A3(n1603), .ZN(n1607) );
  AND2_X1 U1090 ( .A1(n4856), .A2(n1243), .ZN(n1095) );
  AND2_X1 U1091 ( .A1(n1240), .A2(n2360), .ZN(n1096) );
  NAND2_X1 U1092 ( .A1(n2346), .A2(n873), .ZN(n2541) );
  AND2_X1 U1093 ( .A1(n4855), .A2(n1243), .ZN(n1097) );
  AND2_X1 U1094 ( .A1(n1240), .A2(n2335), .ZN(n1098) );
  NOR3_X1 U1095 ( .A1(n2334), .A2(n1098), .A3(n1097), .ZN(n2346) );
  AND2_X1 U1096 ( .A1(n1156), .A2(n4864), .ZN(n1099) );
  AND2_X1 U1097 ( .A1(n1153), .A2(n3616), .ZN(n1100) );
  AND2_X1 U1098 ( .A1(n1154), .A2(n4853), .ZN(n1101) );
  AND2_X1 U1099 ( .A1(n1153), .A2(n2285), .ZN(n1102) );
  AND2_X1 U1100 ( .A1(n4854), .A2(n1243), .ZN(n1103) );
  AND2_X1 U1101 ( .A1(n1240), .A2(n2310), .ZN(n1104) );
  AND2_X1 U1102 ( .A1(n1156), .A2(n4852), .ZN(n1105) );
  AND2_X1 U1103 ( .A1(n1151), .A2(n2256), .ZN(n1106) );
  AND2_X1 U1104 ( .A1(n4853), .A2(n1243), .ZN(n1107) );
  AND2_X1 U1105 ( .A1(n1240), .A2(n2285), .ZN(n1108) );
  AND2_X1 U1106 ( .A1(n4852), .A2(n1243), .ZN(n1109) );
  AND2_X1 U1107 ( .A1(n1240), .A2(n2256), .ZN(n1110) );
  CLKBUF_X3 U1108 ( .A(n2200), .Z(n1114) );
  CLKBUF_X3 U1109 ( .A(n2200), .Z(n1115) );
  CLKBUF_X3 U1110 ( .A(n2200), .Z(n1116) );
  CLKBUF_X3 U1111 ( .A(n2202), .Z(n1117) );
  CLKBUF_X3 U1112 ( .A(n2202), .Z(n1118) );
  CLKBUF_X3 U1113 ( .A(n2202), .Z(n1119) );
  CLKBUF_X3 U1114 ( .A(n2204), .Z(n1125) );
  CLKBUF_X3 U1115 ( .A(n2204), .Z(n1126) );
  CLKBUF_X3 U1116 ( .A(n2205), .Z(n1127) );
  CLKBUF_X3 U1117 ( .A(n2205), .Z(n1128) );
  CLKBUF_X3 U1118 ( .A(n2208), .Z(n1130) );
  CLKBUF_X3 U1119 ( .A(n2208), .Z(n1131) );
  CLKBUF_X3 U1120 ( .A(n2209), .Z(n1133) );
  CLKBUF_X3 U1121 ( .A(n2209), .Z(n1135) );
  CLKBUF_X3 U1122 ( .A(n2213), .Z(n1136) );
  CLKBUF_X3 U1123 ( .A(n2213), .Z(n1137) );
  CLKBUF_X3 U1124 ( .A(n2214), .Z(n1139) );
  CLKBUF_X3 U1125 ( .A(n2214), .Z(n1140) );
  CLKBUF_X3 U1126 ( .A(n2221), .Z(n1145) );
  CLKBUF_X3 U1127 ( .A(n2221), .Z(n1146) );
  CLKBUF_X3 U1128 ( .A(n2223), .Z(n1148) );
  CLKBUF_X3 U1129 ( .A(n2223), .Z(n1149) );
  INV_X1 U1130 ( .A(n1378), .ZN(n1377) );
  INV_X1 U1131 ( .A(n1380), .ZN(n1379) );
  INV_X1 U1132 ( .A(n1382), .ZN(n1381) );
  INV_X1 U1133 ( .A(n1384), .ZN(n1383) );
  INV_X1 U1134 ( .A(n1386), .ZN(n1385) );
  INV_X1 U1135 ( .A(n1388), .ZN(n1387) );
  INV_X1 U1136 ( .A(n1390), .ZN(n1389) );
  INV_X1 U1137 ( .A(n1392), .ZN(n1391) );
  INV_X1 U1138 ( .A(n1394), .ZN(n1393) );
  INV_X1 U1139 ( .A(n1396), .ZN(n1395) );
  INV_X1 U1140 ( .A(n1398), .ZN(n1397) );
  INV_X1 U1141 ( .A(n1400), .ZN(n1399) );
  INV_X1 U1142 ( .A(n1402), .ZN(n1401) );
  INV_X1 U1143 ( .A(n1404), .ZN(n1403) );
  INV_X1 U1144 ( .A(n1406), .ZN(n1405) );
  INV_X1 U1145 ( .A(n1408), .ZN(n1407) );
  INV_X1 U1146 ( .A(n1410), .ZN(n1409) );
  INV_X1 U1147 ( .A(n1412), .ZN(n1411) );
  INV_X1 U1148 ( .A(n1414), .ZN(n1413) );
  INV_X1 U1149 ( .A(n1416), .ZN(n1415) );
  INV_X1 U1150 ( .A(n1418), .ZN(n1417) );
  INV_X1 U1151 ( .A(n1420), .ZN(n1419) );
  INV_X1 U1152 ( .A(n1422), .ZN(n1421) );
  INV_X1 U1153 ( .A(n1424), .ZN(n1423) );
  INV_X1 U1154 ( .A(n1427), .ZN(n1425) );
  INV_X1 U1155 ( .A(n1427), .ZN(n1426) );
  INV_X1 U1156 ( .A(n1430), .ZN(n1428) );
  INV_X1 U1157 ( .A(n1430), .ZN(n1429) );
  INV_X1 U1158 ( .A(n1433), .ZN(n1431) );
  INV_X1 U1159 ( .A(n1433), .ZN(n1432) );
  INV_X1 U1160 ( .A(n1436), .ZN(n1434) );
  INV_X1 U1161 ( .A(n1436), .ZN(n1435) );
  INV_X1 U1162 ( .A(n1439), .ZN(n1437) );
  INV_X1 U1163 ( .A(n1439), .ZN(n1438) );
  INV_X1 U1164 ( .A(n1442), .ZN(n1440) );
  INV_X1 U1165 ( .A(n1442), .ZN(n1441) );
  INV_X1 U1166 ( .A(n1445), .ZN(n1443) );
  INV_X1 U1167 ( .A(n1445), .ZN(n1444) );
  INV_X1 U1168 ( .A(n1448), .ZN(n1446) );
  INV_X1 U1169 ( .A(n1448), .ZN(n1447) );
  CLKBUF_X1 U1170 ( .A(n1552), .Z(n1456) );
  CLKBUF_X1 U1171 ( .A(n1552), .Z(n1457) );
  CLKBUF_X1 U1172 ( .A(n1552), .Z(n1458) );
  CLKBUF_X1 U1173 ( .A(n1552), .Z(n1459) );
  CLKBUF_X1 U1174 ( .A(n1552), .Z(n1460) );
  CLKBUF_X1 U1175 ( .A(n1551), .Z(n1461) );
  CLKBUF_X1 U1176 ( .A(n1551), .Z(n1462) );
  CLKBUF_X1 U1177 ( .A(n1551), .Z(n1463) );
  CLKBUF_X1 U1178 ( .A(n1551), .Z(n1464) );
  CLKBUF_X1 U1179 ( .A(n1551), .Z(n1465) );
  CLKBUF_X1 U1180 ( .A(n1551), .Z(n1466) );
  CLKBUF_X1 U1181 ( .A(n1550), .Z(n1467) );
  CLKBUF_X1 U1182 ( .A(n1550), .Z(n1468) );
  CLKBUF_X1 U1183 ( .A(n1550), .Z(n1469) );
  CLKBUF_X1 U1184 ( .A(n1550), .Z(n1470) );
  CLKBUF_X1 U1185 ( .A(n1550), .Z(n1471) );
  CLKBUF_X1 U1186 ( .A(n1550), .Z(n1472) );
  CLKBUF_X1 U1187 ( .A(n1549), .Z(n1473) );
  CLKBUF_X1 U1188 ( .A(n1549), .Z(n1474) );
  CLKBUF_X1 U1189 ( .A(n1549), .Z(n1475) );
  CLKBUF_X1 U1190 ( .A(n1549), .Z(n1476) );
  CLKBUF_X1 U1191 ( .A(n1549), .Z(n1477) );
  CLKBUF_X1 U1192 ( .A(n1549), .Z(n1478) );
  CLKBUF_X1 U1193 ( .A(n1548), .Z(n1479) );
  CLKBUF_X1 U1194 ( .A(n1548), .Z(n1480) );
  CLKBUF_X1 U1195 ( .A(n1548), .Z(n1481) );
  CLKBUF_X1 U1196 ( .A(n1548), .Z(n1482) );
  CLKBUF_X1 U1197 ( .A(n1548), .Z(n1483) );
  CLKBUF_X1 U1198 ( .A(n1548), .Z(n1484) );
  CLKBUF_X1 U1199 ( .A(n1547), .Z(n1485) );
  CLKBUF_X1 U1200 ( .A(n1547), .Z(n1486) );
  CLKBUF_X1 U1201 ( .A(n1547), .Z(n1487) );
  CLKBUF_X1 U1202 ( .A(n1547), .Z(n1488) );
  CLKBUF_X1 U1203 ( .A(n1547), .Z(n1489) );
  CLKBUF_X1 U1204 ( .A(n1547), .Z(n1490) );
  CLKBUF_X1 U1205 ( .A(n1546), .Z(n1491) );
  CLKBUF_X1 U1206 ( .A(n1546), .Z(n1492) );
  CLKBUF_X1 U1207 ( .A(n1546), .Z(n1493) );
  CLKBUF_X1 U1208 ( .A(n1546), .Z(n1494) );
  CLKBUF_X1 U1209 ( .A(n1546), .Z(n1495) );
  CLKBUF_X1 U1210 ( .A(n1546), .Z(n1496) );
  CLKBUF_X1 U1211 ( .A(n1545), .Z(n1497) );
  CLKBUF_X1 U1212 ( .A(n1545), .Z(n1498) );
  CLKBUF_X1 U1213 ( .A(n1545), .Z(n1499) );
  CLKBUF_X1 U1214 ( .A(n1545), .Z(n1500) );
  CLKBUF_X1 U1215 ( .A(n1545), .Z(n1501) );
  CLKBUF_X1 U1216 ( .A(n1545), .Z(n1502) );
  CLKBUF_X1 U1217 ( .A(n1544), .Z(n1503) );
  CLKBUF_X1 U1218 ( .A(n1544), .Z(n1504) );
  CLKBUF_X1 U1219 ( .A(n1544), .Z(n1505) );
  CLKBUF_X1 U1220 ( .A(n1544), .Z(n1506) );
  CLKBUF_X1 U1221 ( .A(n1544), .Z(n1507) );
  CLKBUF_X1 U1222 ( .A(n1544), .Z(n1508) );
  CLKBUF_X1 U1223 ( .A(n1543), .Z(n1509) );
  CLKBUF_X1 U1224 ( .A(n1543), .Z(n1510) );
  CLKBUF_X1 U1225 ( .A(n1543), .Z(n1511) );
  CLKBUF_X1 U1226 ( .A(n1543), .Z(n1512) );
  CLKBUF_X1 U1227 ( .A(n1543), .Z(n1513) );
  CLKBUF_X1 U1228 ( .A(n1543), .Z(n1514) );
  CLKBUF_X1 U1229 ( .A(n1542), .Z(n1515) );
  CLKBUF_X1 U1230 ( .A(n1542), .Z(n1516) );
  CLKBUF_X1 U1231 ( .A(n1542), .Z(n1517) );
  CLKBUF_X1 U1232 ( .A(n1542), .Z(n1518) );
  CLKBUF_X1 U1233 ( .A(n1542), .Z(n1519) );
  CLKBUF_X1 U1234 ( .A(n1542), .Z(n1520) );
  CLKBUF_X1 U1235 ( .A(n1541), .Z(n1521) );
  CLKBUF_X1 U1236 ( .A(n1541), .Z(n1522) );
  CLKBUF_X1 U1237 ( .A(n1541), .Z(n1523) );
  CLKBUF_X1 U1238 ( .A(n1541), .Z(n1524) );
  CLKBUF_X1 U1239 ( .A(n1541), .Z(n1525) );
  CLKBUF_X1 U1240 ( .A(n1541), .Z(n1526) );
  CLKBUF_X1 U1241 ( .A(n1540), .Z(n1527) );
  CLKBUF_X1 U1242 ( .A(n1540), .Z(n1528) );
  CLKBUF_X1 U1243 ( .A(n1540), .Z(n1529) );
  CLKBUF_X1 U1244 ( .A(n1540), .Z(n1530) );
  CLKBUF_X1 U1245 ( .A(n1540), .Z(n1531) );
  CLKBUF_X1 U1246 ( .A(n1540), .Z(n1532) );
  CLKBUF_X1 U1247 ( .A(n1539), .Z(n1533) );
  CLKBUF_X1 U1248 ( .A(n1539), .Z(n1534) );
  CLKBUF_X1 U1249 ( .A(n1539), .Z(n1535) );
  CLKBUF_X1 U1250 ( .A(n1539), .Z(n1536) );
  CLKBUF_X1 U1251 ( .A(n1539), .Z(n1537) );
  INV_X1 U1252 ( .A(ADD_RS1[2]), .ZN(n1554) );
  INV_X1 U1253 ( .A(n890), .ZN(n1572) );
  NAND4_X1 U1254 ( .A1(n930), .A2(n705), .A3(n1186), .A4(n875), .ZN(n2223) );
  INV_X1 U1255 ( .A(ADD_RS1[4]), .ZN(n1560) );
  INV_X1 U1256 ( .A(ADD_RS1[1]), .ZN(n1553) );
  NAND2_X1 U1257 ( .A1(n1015), .A2(n887), .ZN(n2202) );
  NAND2_X1 U1258 ( .A1(n1015), .A2(n705), .ZN(n2200) );
  AOI22_X1 U1259 ( .A1(n969), .A2(n4159), .B1(n739), .B2(n4724), .ZN(n1555) );
  OAI221_X1 U1260 ( .B1(n164), .B2(n1117), .C1(n1556), .C2(n1115), .A(n1555), 
        .ZN(n1568) );
  NAND2_X1 U1261 ( .A1(n886), .A2(n171), .ZN(n2205) );
  NAND2_X1 U1262 ( .A1(n886), .A2(n468), .ZN(n2204) );
  AOI22_X1 U1263 ( .A1(n1124), .A2(n5044), .B1(n512), .B2(n5108), .ZN(n1557)
         );
  OAI221_X1 U1264 ( .B1(n2246), .B2(n1129), .C1(n292), .C2(n1125), .A(n1557), 
        .ZN(n1567) );
  NAND2_X1 U1265 ( .A1(n1053), .A2(n171), .ZN(n2209) );
  NAND2_X1 U1266 ( .A1(n1053), .A2(n468), .ZN(n2208) );
  AOI22_X1 U1267 ( .A1(n56), .A2(n5076), .B1(n760), .B2(n1558), .ZN(n1559) );
  OAI221_X1 U1268 ( .B1(n2247), .B2(n1135), .C1(n260), .C2(n1130), .A(n1559), 
        .ZN(n1566) );
  NAND2_X1 U1269 ( .A1(n1031), .A2(n171), .ZN(n2214) );
  NAND2_X1 U1270 ( .A1(n1031), .A2(n887), .ZN(n2213) );
  NAND2_X1 U1271 ( .A1(n1031), .A2(n705), .ZN(n1561) );
  INV_X1 U1272 ( .A(n1561), .ZN(n2211) );
  AOI22_X1 U1273 ( .A1(n1014), .A2(n5204), .B1(n489), .B2(n1562), .ZN(n1563)
         );
  OAI221_X1 U1274 ( .B1(n1564), .B2(n1139), .C1(n132), .C2(n1136), .A(n1563), 
        .ZN(n1565) );
  NOR4_X1 U1275 ( .A1(n1568), .A2(n1567), .A3(n1565), .A4(n1566), .ZN(n1569)
         );
  NAND2_X1 U1276 ( .A1(n1574), .A2(n1187), .ZN(n2221) );
  NAND4_X1 U1277 ( .A1(n874), .A2(n468), .A3(n1186), .A4(n930), .ZN(n2220) );
  OAI222_X1 U1278 ( .A1(n836), .A2(n1148), .B1(n1569), .B2(n1145), .C1(n2253), 
        .C2(n1142), .ZN(n1570) );
  NAND4_X1 U1279 ( .A1(n875), .A2(n887), .A3(n1186), .A4(n930), .ZN(n2226) );
  NAND4_X1 U1280 ( .A1(n874), .A2(n171), .A3(n1186), .A4(n930), .ZN(n2225) );
  OAI22_X1 U1281 ( .A1(n2257), .A2(n707), .B1(n964), .B2(n1157), .ZN(n1571) );
  AOI221_X1 U1282 ( .B1(n1166), .B2(n4788), .C1(n1163), .C2(n4339), .A(n1571), 
        .ZN(n1578) );
  NAND4_X1 U1283 ( .A1(n1574), .A2(n887), .A3(n1186), .A4(n971), .ZN(n2230) );
  NAND4_X1 U1284 ( .A1(n874), .A2(n171), .A3(n1186), .A4(n971), .ZN(n2229) );
  NAND4_X1 U1285 ( .A1(n874), .A2(n705), .A3(n1187), .A4(n978), .ZN(n2228) );
  NAND3_X1 U1286 ( .A1(n1187), .A2(n78), .A3(n690), .ZN(n2232) );
  OAI22_X1 U1287 ( .A1(n4660), .A2(n1187), .B1(n1378), .B2(n1183), .ZN(n1575)
         );
  AOI221_X1 U1288 ( .B1(n1193), .B2(n4948), .C1(n1190), .C2(n2267), .A(n1575), 
        .ZN(n1576) );
  NAND4_X1 U1289 ( .A1(n1579), .A2(n1577), .A3(n1576), .A4(n1578), .ZN(n2506)
         );
  AOI22_X1 U1290 ( .A1(n969), .A2(n4158), .B1(n486), .B2(n4725), .ZN(n1580) );
  OAI221_X1 U1291 ( .B1(n163), .B2(n1118), .C1(n1581), .C2(n1115), .A(n1580), 
        .ZN(n1591) );
  AOI22_X1 U1292 ( .A1(n1122), .A2(n5045), .B1(n493), .B2(n5109), .ZN(n1582)
         );
  OAI221_X1 U1293 ( .B1(n2275), .B2(n1127), .C1(n291), .C2(n1125), .A(n1582), 
        .ZN(n1590) );
  AOI22_X1 U1294 ( .A1(n54), .A2(n5077), .B1(n759), .B2(n1583), .ZN(n1584) );
  OAI221_X1 U1295 ( .B1(n2276), .B2(n1133), .C1(n259), .C2(n1130), .A(n1584), 
        .ZN(n1589) );
  AOI22_X1 U1296 ( .A1(n1014), .A2(n5205), .B1(n966), .B2(n1585), .ZN(n1586)
         );
  NOR4_X1 U1297 ( .A1(n1591), .A2(n1589), .A3(n1590), .A4(n1588), .ZN(n1592)
         );
  OAI22_X1 U1298 ( .A1(n2286), .A2(n1161), .B1(n963), .B2(n1157), .ZN(n1593)
         );
  AOI221_X1 U1299 ( .B1(n1166), .B2(n4789), .C1(n1163), .C2(n4338), .A(n1593), 
        .ZN(n1598) );
  OAI22_X1 U1300 ( .A1(n4661), .A2(n1189), .B1(n1380), .B2(n1183), .ZN(n1595)
         );
  AOI221_X1 U1301 ( .B1(n1193), .B2(n4949), .C1(n1190), .C2(n2292), .A(n1595), 
        .ZN(n1596) );
  NAND4_X1 U1302 ( .A1(n1599), .A2(n1597), .A3(n1596), .A4(n1598), .ZN(n2507)
         );
  AOI22_X1 U1303 ( .A1(n969), .A2(n4157), .B1(n486), .B2(n4726), .ZN(n1600) );
  OAI221_X1 U1304 ( .B1(n162), .B2(n1118), .C1(n1601), .C2(n1115), .A(n1600), 
        .ZN(n1609) );
  AOI22_X1 U1305 ( .A1(n1123), .A2(n5046), .B1(n493), .B2(n5110), .ZN(n1602)
         );
  OAI221_X1 U1306 ( .B1(n2300), .B2(n1127), .C1(n290), .C2(n1125), .A(n1602), 
        .ZN(n1608) );
  AOI22_X1 U1307 ( .A1(n56), .A2(n5078), .B1(n1029), .B2(n218), .ZN(n1603) );
  AOI22_X1 U1308 ( .A1(n888), .A2(n5206), .B1(n579), .B2(n219), .ZN(n1604) );
  NOR4_X1 U1309 ( .A1(n1609), .A2(n1608), .A3(n1606), .A4(n1607), .ZN(n1610)
         );
  OAI222_X1 U1310 ( .A1(n834), .A2(n1148), .B1(n1610), .B2(n1145), .C1(n2307), 
        .C2(n1142), .ZN(n1611) );
  OAI22_X1 U1311 ( .A1(n2311), .A2(n1160), .B1(n962), .B2(n1157), .ZN(n1612)
         );
  AOI221_X1 U1312 ( .B1(n1166), .B2(n4790), .C1(n1163), .C2(n4337), .A(n1612), 
        .ZN(n1617) );
  OAI222_X1 U1313 ( .A1(n642), .A2(n1175), .B1(n2314), .B2(n1173), .C1(n2313), 
        .C2(n1169), .ZN(n1613) );
  AOI221_X1 U1314 ( .B1(n1180), .B2(n4285), .C1(n1177), .C2(n4253), .A(n1613), 
        .ZN(n1616) );
  OAI22_X1 U1315 ( .A1(n4662), .A2(n1189), .B1(n1382), .B2(n1183), .ZN(n1614)
         );
  AOI221_X1 U1316 ( .B1(n1193), .B2(n4950), .C1(n1190), .C2(n2317), .A(n1614), 
        .ZN(n1615) );
  NAND4_X1 U1317 ( .A1(n1618), .A2(n1615), .A3(n1617), .A4(n1616), .ZN(n2508)
         );
  AOI22_X1 U1318 ( .A1(n969), .A2(n4156), .B1(n738), .B2(n4727), .ZN(n1619) );
  AOI22_X1 U1319 ( .A1(n1122), .A2(n5047), .B1(n493), .B2(n5111), .ZN(n1621)
         );
  OAI221_X1 U1320 ( .B1(n2325), .B2(n1127), .C1(n289), .C2(n1125), .A(n1621), 
        .ZN(n1629) );
  AOI22_X1 U1321 ( .A1(n56), .A2(n5079), .B1(n760), .B2(n1622), .ZN(n1623) );
  OAI221_X1 U1322 ( .B1(n507), .B2(n2326), .C1(n257), .C2(n1131), .A(n1623), 
        .ZN(n1628) );
  AOI22_X1 U1323 ( .A1(n888), .A2(n5207), .B1(n966), .B2(n1624), .ZN(n1625) );
  OAI221_X1 U1324 ( .B1(n1626), .B2(n1139), .C1(n129), .C2(n1136), .A(n1625), 
        .ZN(n1627) );
  NOR4_X1 U1325 ( .A1(n1630), .A2(n1628), .A3(n1629), .A4(n1627), .ZN(n1631)
         );
  OAI22_X1 U1326 ( .A1(n2336), .A2(n707), .B1(n961), .B2(n1157), .ZN(n1632) );
  OAI222_X1 U1327 ( .A1(n641), .A2(n1175), .B1(n2339), .B2(n1173), .C1(n2338), 
        .C2(n1169), .ZN(n1633) );
  AOI221_X1 U1328 ( .B1(n1180), .B2(n4284), .C1(n1177), .C2(n4252), .A(n1633), 
        .ZN(n1636) );
  OAI22_X1 U1329 ( .A1(n4663), .A2(n1189), .B1(n1384), .B2(n1183), .ZN(n1634)
         );
  AOI221_X1 U1330 ( .B1(n1193), .B2(n4951), .C1(n1190), .C2(n2342), .A(n1634), 
        .ZN(n1635) );
  NAND4_X1 U1331 ( .A1(n1636), .A2(n1637), .A3(n1638), .A4(n1635), .ZN(n2509)
         );
  AOI22_X1 U1332 ( .A1(n669), .A2(n4155), .B1(n1111), .B2(n4728), .ZN(n1639)
         );
  OAI221_X1 U1333 ( .B1(n160), .B2(n1118), .C1(n1640), .C2(n1114), .A(n1639), 
        .ZN(n1650) );
  AOI22_X1 U1334 ( .A1(n1122), .A2(n5048), .B1(n493), .B2(n5112), .ZN(n1641)
         );
  OAI221_X1 U1335 ( .B1(n2350), .B2(n1129), .C1(n288), .C2(n1125), .A(n1641), 
        .ZN(n1649) );
  AOI22_X1 U1336 ( .A1(n55), .A2(n5080), .B1(n759), .B2(n1642), .ZN(n1643) );
  OAI221_X1 U1337 ( .B1(n1133), .B2(n2351), .C1(n256), .C2(n1131), .A(n1643), 
        .ZN(n1648) );
  AOI22_X1 U1338 ( .A1(n1014), .A2(n5208), .B1(n966), .B2(n1644), .ZN(n1645)
         );
  NOR4_X1 U1339 ( .A1(n1650), .A2(n1648), .A3(n1649), .A4(n1647), .ZN(n1651)
         );
  OAI22_X1 U1340 ( .A1(n2361), .A2(n707), .B1(n960), .B2(n1157), .ZN(n1653) );
  AOI221_X1 U1341 ( .B1(n1166), .B2(n4792), .C1(n1163), .C2(n4335), .A(n1653), 
        .ZN(n1658) );
  OAI222_X1 U1342 ( .A1(n640), .A2(n1176), .B1(n2364), .B2(n1173), .C1(n2363), 
        .C2(n1169), .ZN(n1654) );
  AOI221_X1 U1343 ( .B1(n1180), .B2(n4283), .C1(n1177), .C2(n4251), .A(n1654), 
        .ZN(n1657) );
  OAI22_X1 U1344 ( .A1(n4664), .A2(n1189), .B1(n1386), .B2(n1183), .ZN(n1655)
         );
  AOI221_X1 U1345 ( .B1(n1193), .B2(n4952), .C1(n1190), .C2(n2367), .A(n1655), 
        .ZN(n1656) );
  NAND4_X1 U1346 ( .A1(n1657), .A2(n1659), .A3(n1656), .A4(n1658), .ZN(n2510)
         );
  AOI22_X1 U1347 ( .A1(n668), .A2(n4154), .B1(n739), .B2(n4729), .ZN(n1660) );
  OAI221_X1 U1348 ( .B1(n159), .B2(n1119), .C1(n1661), .C2(n1114), .A(n1660), 
        .ZN(n1671) );
  AOI22_X1 U1349 ( .A1(n1023), .A2(n5049), .B1(n52), .B2(n5113), .ZN(n1662) );
  OAI221_X1 U1350 ( .B1(n2375), .B2(n1128), .C1(n287), .C2(n1125), .A(n1662), 
        .ZN(n1670) );
  AOI22_X1 U1351 ( .A1(n56), .A2(n5081), .B1(n1029), .B2(n1663), .ZN(n1664) );
  AOI22_X1 U1352 ( .A1(n2211), .A2(n5209), .B1(n966), .B2(n1665), .ZN(n1666)
         );
  OAI221_X1 U1353 ( .B1(n1667), .B2(n1139), .C1(n127), .C2(n1136), .A(n1666), 
        .ZN(n1668) );
  NOR4_X1 U1354 ( .A1(n1671), .A2(n1670), .A3(n1668), .A4(n1669), .ZN(n1672)
         );
  OAI22_X1 U1355 ( .A1(n2386), .A2(n1161), .B1(n959), .B2(n1157), .ZN(n1674)
         );
  AOI221_X1 U1356 ( .B1(n1166), .B2(n4793), .C1(n1163), .C2(n4334), .A(n1674), 
        .ZN(n1679) );
  OAI222_X1 U1357 ( .A1(n639), .A2(n1175), .B1(n2389), .B2(n1173), .C1(n2388), 
        .C2(n1169), .ZN(n1675) );
  AOI221_X1 U1358 ( .B1(n1180), .B2(n4282), .C1(n1177), .C2(n4250), .A(n1675), 
        .ZN(n1678) );
  OAI22_X1 U1359 ( .A1(n4665), .A2(n1189), .B1(n1388), .B2(n1183), .ZN(n1676)
         );
  AOI221_X1 U1360 ( .B1(n1193), .B2(n4953), .C1(n1190), .C2(n2392), .A(n1676), 
        .ZN(n1677) );
  NAND4_X1 U1361 ( .A1(n1678), .A2(n1680), .A3(n1677), .A4(n1679), .ZN(n2511)
         );
  AOI22_X1 U1362 ( .A1(n969), .A2(n4153), .B1(n738), .B2(n4730), .ZN(n1681) );
  OAI221_X1 U1363 ( .B1(n158), .B2(n1117), .C1(n1682), .C2(n1114), .A(n1681), 
        .ZN(n1692) );
  AOI22_X1 U1364 ( .A1(n1024), .A2(n5050), .B1(n1120), .B2(n5114), .ZN(n1683)
         );
  OAI221_X1 U1365 ( .B1(n2400), .B2(n1129), .C1(n286), .C2(n1125), .A(n1683), 
        .ZN(n1691) );
  AOI22_X1 U1366 ( .A1(n57), .A2(n5082), .B1(n759), .B2(n1684), .ZN(n1685) );
  OAI221_X1 U1367 ( .B1(n2401), .B2(n1135), .C1(n254), .C2(n1130), .A(n1685), 
        .ZN(n1690) );
  AOI22_X1 U1368 ( .A1(n888), .A2(n5210), .B1(n966), .B2(n1686), .ZN(n1687) );
  OAI221_X1 U1369 ( .B1(n1688), .B2(n1139), .C1(n126), .C2(n1136), .A(n1687), 
        .ZN(n1689) );
  NOR4_X1 U1370 ( .A1(n1692), .A2(n1691), .A3(n1690), .A4(n1689), .ZN(n1693)
         );
  OAI222_X1 U1371 ( .A1(n830), .A2(n1148), .B1(n1693), .B2(n1145), .C1(n2407), 
        .C2(n1142), .ZN(n1694) );
  OAI22_X1 U1372 ( .A1(n2411), .A2(n1161), .B1(n958), .B2(n1157), .ZN(n1695)
         );
  AOI221_X1 U1373 ( .B1(n1166), .B2(n4794), .C1(n1163), .C2(n4333), .A(n1695), 
        .ZN(n1700) );
  OAI222_X1 U1374 ( .A1(n638), .A2(n1174), .B1(n1171), .B2(n2414), .C1(n2413), 
        .C2(n1169), .ZN(n1696) );
  AOI221_X1 U1375 ( .B1(n1180), .B2(n4281), .C1(n1177), .C2(n4249), .A(n1696), 
        .ZN(n1699) );
  OAI22_X1 U1376 ( .A1(n4666), .A2(n1189), .B1(n1390), .B2(n1183), .ZN(n1697)
         );
  AOI221_X1 U1377 ( .B1(n1193), .B2(n4954), .C1(n1190), .C2(n2417), .A(n1697), 
        .ZN(n1698) );
  NAND4_X1 U1378 ( .A1(n1699), .A2(n1701), .A3(n1700), .A4(n1698), .ZN(n2512)
         );
  AOI22_X1 U1379 ( .A1(n669), .A2(n4152), .B1(n738), .B2(n4731), .ZN(n1702) );
  OAI221_X1 U1380 ( .B1(n157), .B2(n1118), .C1(n1703), .C2(n1114), .A(n1702), 
        .ZN(n1713) );
  AOI22_X1 U1381 ( .A1(n1024), .A2(n5051), .B1(n508), .B2(n5115), .ZN(n1704)
         );
  OAI221_X1 U1382 ( .B1(n2425), .B2(n1129), .C1(n285), .C2(n1125), .A(n1704), 
        .ZN(n1712) );
  AOI22_X1 U1383 ( .A1(n54), .A2(n5083), .B1(n1029), .B2(n1705), .ZN(n1706) );
  OAI221_X1 U1384 ( .B1(n2426), .B2(n1133), .C1(n253), .C2(n506), .A(n1706), 
        .ZN(n1711) );
  AOI22_X1 U1385 ( .A1(n888), .A2(n5211), .B1(n578), .B2(n1707), .ZN(n1708) );
  NOR4_X1 U1386 ( .A1(n1713), .A2(n1712), .A3(n1710), .A4(n1711), .ZN(n1714)
         );
  OAI222_X1 U1387 ( .A1(n829), .A2(n1148), .B1(n1714), .B2(n1145), .C1(n2432), 
        .C2(n1142), .ZN(n1715) );
  OAI22_X1 U1388 ( .A1(n2436), .A2(n1162), .B1(n957), .B2(n1157), .ZN(n1716)
         );
  AOI221_X1 U1389 ( .B1(n1166), .B2(n4795), .C1(n1163), .C2(n4332), .A(n1716), 
        .ZN(n1721) );
  OAI222_X1 U1390 ( .A1(n637), .A2(n1174), .B1(n1171), .B2(n2439), .C1(n2438), 
        .C2(n1169), .ZN(n1717) );
  AOI221_X1 U1391 ( .B1(n1180), .B2(n4280), .C1(n1177), .C2(n4248), .A(n1717), 
        .ZN(n1720) );
  OAI22_X1 U1392 ( .A1(n4667), .A2(n1189), .B1(n1392), .B2(n1183), .ZN(n1718)
         );
  AOI221_X1 U1393 ( .B1(n1193), .B2(n4955), .C1(n1190), .C2(n2442), .A(n1718), 
        .ZN(n1719) );
  NAND4_X1 U1394 ( .A1(n1722), .A2(n1721), .A3(n1719), .A4(n1720), .ZN(n2513)
         );
  AOI22_X1 U1395 ( .A1(n669), .A2(n4151), .B1(n739), .B2(n4732), .ZN(n1723) );
  OAI221_X1 U1396 ( .B1(n156), .B2(n1118), .C1(n1724), .C2(n1116), .A(n1723), 
        .ZN(n1734) );
  AOI22_X1 U1397 ( .A1(n1123), .A2(n5052), .B1(n52), .B2(n5116), .ZN(n1725) );
  OAI221_X1 U1398 ( .B1(n2450), .B2(n1128), .C1(n284), .C2(n1125), .A(n1725), 
        .ZN(n1733) );
  AOI22_X1 U1399 ( .A1(n54), .A2(n5084), .B1(n760), .B2(n1726), .ZN(n1727) );
  OAI221_X1 U1400 ( .B1(n2451), .B2(n1135), .C1(n252), .C2(n1130), .A(n1727), 
        .ZN(n1732) );
  AOI22_X1 U1401 ( .A1(n1014), .A2(n5212), .B1(n577), .B2(n1728), .ZN(n1729)
         );
  NOR4_X1 U1402 ( .A1(n1734), .A2(n1733), .A3(n1731), .A4(n1732), .ZN(n1735)
         );
  OAI222_X1 U1403 ( .A1(n828), .A2(n1148), .B1(n1735), .B2(n1145), .C1(n2457), 
        .C2(n1142), .ZN(n1736) );
  OAI22_X1 U1404 ( .A1(n2461), .A2(n707), .B1(n956), .B2(n1157), .ZN(n1737) );
  AOI221_X1 U1405 ( .B1(n1166), .B2(n4796), .C1(n1163), .C2(n4331), .A(n1737), 
        .ZN(n1742) );
  OAI222_X1 U1406 ( .A1(n636), .A2(n1175), .B1(n2464), .B2(n1172), .C1(n2463), 
        .C2(n1169), .ZN(n1738) );
  AOI221_X1 U1407 ( .B1(n1180), .B2(n4279), .C1(n1177), .C2(n4247), .A(n1738), 
        .ZN(n1741) );
  OAI22_X1 U1408 ( .A1(n4668), .A2(n1189), .B1(n1394), .B2(n1183), .ZN(n1739)
         );
  AOI221_X1 U1409 ( .B1(n1193), .B2(n4956), .C1(n1190), .C2(n2467), .A(n1739), 
        .ZN(n1740) );
  NAND4_X1 U1410 ( .A1(n1743), .A2(n1742), .A3(n1740), .A4(n1741), .ZN(n2514)
         );
  AOI22_X1 U1411 ( .A1(n969), .A2(n4150), .B1(n739), .B2(n4733), .ZN(n1744) );
  OAI221_X1 U1412 ( .B1(n155), .B2(n1118), .C1(n1745), .C2(n1116), .A(n1744), 
        .ZN(n1755) );
  AOI22_X1 U1413 ( .A1(n1016), .A2(n5053), .B1(n1121), .B2(n5117), .ZN(n1746)
         );
  AOI22_X1 U1414 ( .A1(n54), .A2(n5085), .B1(n760), .B2(n1747), .ZN(n1748) );
  OAI221_X1 U1415 ( .B1(n2476), .B2(n1133), .C1(n251), .C2(n1131), .A(n1748), 
        .ZN(n1753) );
  AOI22_X1 U1416 ( .A1(n888), .A2(n5213), .B1(n578), .B2(n1749), .ZN(n1750) );
  OAI221_X1 U1417 ( .B1(n1751), .B2(n1139), .C1(n123), .C2(n1136), .A(n1750), 
        .ZN(n1752) );
  NOR4_X1 U1418 ( .A1(n1755), .A2(n1752), .A3(n1753), .A4(n1754), .ZN(n1756)
         );
  OAI222_X1 U1419 ( .A1(n827), .A2(n1148), .B1(n1756), .B2(n1145), .C1(n2482), 
        .C2(n1142), .ZN(n1757) );
  OAI22_X1 U1420 ( .A1(n2486), .A2(n1161), .B1(n955), .B2(n1157), .ZN(n1758)
         );
  AOI221_X1 U1421 ( .B1(n1166), .B2(n4797), .C1(n1163), .C2(n4330), .A(n1758), 
        .ZN(n1763) );
  OAI222_X1 U1422 ( .A1(n635), .A2(n1176), .B1(n2489), .B2(n1173), .C1(n2488), 
        .C2(n1169), .ZN(n1759) );
  AOI221_X1 U1423 ( .B1(n1180), .B2(n4278), .C1(n1177), .C2(n4246), .A(n1759), 
        .ZN(n1762) );
  OAI22_X1 U1424 ( .A1(n4669), .A2(n1189), .B1(n1396), .B2(n1183), .ZN(n1760)
         );
  AOI221_X1 U1425 ( .B1(n1193), .B2(n4957), .C1(n1190), .C2(n2492), .A(n1760), 
        .ZN(n1761) );
  NAND4_X1 U1426 ( .A1(n1762), .A2(n1761), .A3(n1763), .A4(n1764), .ZN(n2515)
         );
  AOI22_X1 U1427 ( .A1(n669), .A2(n4149), .B1(n487), .B2(n4734), .ZN(n1765) );
  OAI221_X1 U1428 ( .B1(n154), .B2(n1118), .C1(n1766), .C2(n1115), .A(n1765), 
        .ZN(n1776) );
  AOI22_X1 U1429 ( .A1(n1016), .A2(n5054), .B1(n1121), .B2(n5118), .ZN(n1767)
         );
  OAI221_X1 U1430 ( .B1(n2500), .B2(n1128), .C1(n282), .C2(n1125), .A(n1767), 
        .ZN(n1775) );
  AOI22_X1 U1431 ( .A1(n54), .A2(n5086), .B1(n759), .B2(n1768), .ZN(n1769) );
  OAI221_X1 U1432 ( .B1(n2501), .B2(n1135), .C1(n250), .C2(n1130), .A(n1769), 
        .ZN(n1774) );
  AOI22_X1 U1433 ( .A1(n888), .A2(n5214), .B1(n966), .B2(n1770), .ZN(n1771) );
  OAI221_X1 U1434 ( .B1(n1772), .B2(n1139), .C1(n122), .C2(n1136), .A(n1771), 
        .ZN(n1773) );
  NOR4_X1 U1435 ( .A1(n1776), .A2(n1775), .A3(n1774), .A4(n1773), .ZN(n1777)
         );
  OAI222_X1 U1436 ( .A1(n826), .A2(n1148), .B1(n1777), .B2(n1145), .C1(n3563), 
        .C2(n1142), .ZN(n1778) );
  OAI22_X1 U1437 ( .A1(n3567), .A2(n1161), .B1(n954), .B2(n1157), .ZN(n1779)
         );
  AOI221_X1 U1438 ( .B1(n1166), .B2(n4798), .C1(n1163), .C2(n4329), .A(n1779), 
        .ZN(n1784) );
  OAI222_X1 U1439 ( .A1(n634), .A2(n1174), .B1(n3570), .B2(n1173), .C1(n3569), 
        .C2(n1170), .ZN(n1780) );
  AOI221_X1 U1440 ( .B1(n1180), .B2(n4277), .C1(n1177), .C2(n4245), .A(n1780), 
        .ZN(n1783) );
  OAI22_X1 U1441 ( .A1(n4670), .A2(n1189), .B1(n1398), .B2(n1183), .ZN(n1781)
         );
  AOI221_X1 U1442 ( .B1(n1193), .B2(n4958), .C1(n1190), .C2(n3573), .A(n1781), 
        .ZN(n1782) );
  NAND4_X1 U1443 ( .A1(n1783), .A2(n1782), .A3(n1784), .A4(n1785), .ZN(n2516)
         );
  AOI22_X1 U1444 ( .A1(n969), .A2(n4148), .B1(n497), .B2(n4735), .ZN(n1786) );
  OAI221_X1 U1445 ( .B1(n153), .B2(n1118), .C1(n1787), .C2(n1114), .A(n1786), 
        .ZN(n1797) );
  AOI22_X1 U1446 ( .A1(n1024), .A2(n5055), .B1(n493), .B2(n5119), .ZN(n1788)
         );
  AOI22_X1 U1447 ( .A1(n55), .A2(n5087), .B1(n1029), .B2(n1789), .ZN(n1790) );
  OAI221_X1 U1448 ( .B1(n3582), .B2(n1133), .C1(n249), .C2(n1130), .A(n1790), 
        .ZN(n1795) );
  AOI22_X1 U1449 ( .A1(n1014), .A2(n5215), .B1(n579), .B2(n1791), .ZN(n1792)
         );
  OAI221_X1 U1450 ( .B1(n1793), .B2(n1139), .C1(n121), .C2(n1136), .A(n1792), 
        .ZN(n1794) );
  NOR4_X1 U1451 ( .A1(n1797), .A2(n1794), .A3(n1796), .A4(n1795), .ZN(n1798)
         );
  OAI222_X1 U1452 ( .A1(n825), .A2(n1148), .B1(n1798), .B2(n1145), .C1(n3588), 
        .C2(n1142), .ZN(n1799) );
  OAI22_X1 U1453 ( .A1(n3592), .A2(n1162), .B1(n953), .B2(n1157), .ZN(n1800)
         );
  AOI221_X1 U1454 ( .B1(n1166), .B2(n4799), .C1(n1163), .C2(n4328), .A(n1800), 
        .ZN(n1805) );
  OAI222_X1 U1455 ( .A1(n633), .A2(n1175), .B1(n3595), .B2(n1172), .C1(n3594), 
        .C2(n1170), .ZN(n1801) );
  AOI221_X1 U1456 ( .B1(n1180), .B2(n4276), .C1(n1177), .C2(n4244), .A(n1801), 
        .ZN(n1804) );
  OAI22_X1 U1457 ( .A1(n4671), .A2(n1189), .B1(n1400), .B2(n1183), .ZN(n1802)
         );
  AOI221_X1 U1458 ( .B1(n1193), .B2(n4959), .C1(n1190), .C2(n3598), .A(n1802), 
        .ZN(n1803) );
  NAND4_X1 U1459 ( .A1(n1804), .A2(n1806), .A3(n1803), .A4(n1805), .ZN(n2517)
         );
  AOI22_X1 U1460 ( .A1(n668), .A2(n4147), .B1(n691), .B2(n4736), .ZN(n1807) );
  OAI221_X1 U1461 ( .B1(n152), .B2(n1119), .C1(n1808), .C2(n1114), .A(n1807), 
        .ZN(n1818) );
  AOI22_X1 U1462 ( .A1(n1124), .A2(n5056), .B1(n493), .B2(n5120), .ZN(n1809)
         );
  AOI22_X1 U1463 ( .A1(n54), .A2(n5088), .B1(n759), .B2(n1810), .ZN(n1811) );
  OAI221_X1 U1464 ( .B1(n507), .B2(n3607), .C1(n248), .C2(n1131), .A(n1811), 
        .ZN(n1816) );
  AOI22_X1 U1465 ( .A1(n888), .A2(n5216), .B1(n966), .B2(n1812), .ZN(n1813) );
  OAI221_X1 U1466 ( .B1(n1814), .B2(n1140), .C1(n120), .C2(n1137), .A(n1813), 
        .ZN(n1815) );
  NOR4_X1 U1467 ( .A1(n1818), .A2(n1816), .A3(n1817), .A4(n1815), .ZN(n1819)
         );
  OAI22_X1 U1468 ( .A1(n3617), .A2(n707), .B1(n952), .B2(n1158), .ZN(n1820) );
  AOI221_X1 U1469 ( .B1(n1167), .B2(n4800), .C1(n1164), .C2(n4327), .A(n1820), 
        .ZN(n1825) );
  OAI222_X1 U1470 ( .A1(n632), .A2(n1176), .B1(n3620), .B2(n1171), .C1(n3619), 
        .C2(n1170), .ZN(n1821) );
  AOI221_X1 U1471 ( .B1(n1181), .B2(n4275), .C1(n1178), .C2(n4243), .A(n1821), 
        .ZN(n1824) );
  OAI22_X1 U1472 ( .A1(n4672), .A2(n1189), .B1(n1402), .B2(n1184), .ZN(n1822)
         );
  AOI221_X1 U1473 ( .B1(n1194), .B2(n4960), .C1(n1191), .C2(n3623), .A(n1822), 
        .ZN(n1823) );
  NAND4_X1 U1474 ( .A1(n1824), .A2(n1825), .A3(n1826), .A4(n1823), .ZN(n2518)
         );
  AOI22_X1 U1475 ( .A1(n969), .A2(n4146), .B1(n1111), .B2(n4737), .ZN(n1827)
         );
  OAI221_X1 U1476 ( .B1(n151), .B2(n1117), .C1(n1828), .C2(n1115), .A(n1827), 
        .ZN(n1838) );
  AOI22_X1 U1477 ( .A1(n1124), .A2(n5057), .B1(n52), .B2(n5121), .ZN(n1829) );
  AOI22_X1 U1478 ( .A1(n56), .A2(n5089), .B1(n1029), .B2(n1830), .ZN(n1831) );
  OAI221_X1 U1479 ( .B1(n3632), .B2(n1135), .C1(n247), .C2(n1130), .A(n1831), 
        .ZN(n1836) );
  AOI22_X1 U1480 ( .A1(n888), .A2(n5217), .B1(n966), .B2(n1832), .ZN(n1833) );
  OAI221_X1 U1481 ( .B1(n1834), .B2(n1140), .C1(n119), .C2(n1137), .A(n1833), 
        .ZN(n1835) );
  NOR4_X1 U1482 ( .A1(n1838), .A2(n1836), .A3(n1837), .A4(n1835), .ZN(n1839)
         );
  OAI222_X1 U1483 ( .A1(n823), .A2(n1149), .B1(n1839), .B2(n1146), .C1(n3638), 
        .C2(n1143), .ZN(n1840) );
  OAI22_X1 U1484 ( .A1(n3642), .A2(n1161), .B1(n951), .B2(n1158), .ZN(n1841)
         );
  AOI221_X1 U1485 ( .B1(n1167), .B2(n4801), .C1(n1164), .C2(n4326), .A(n1841), 
        .ZN(n1846) );
  OAI222_X1 U1486 ( .A1(n631), .A2(n1174), .B1(n3645), .B2(n1171), .C1(n3644), 
        .C2(n1170), .ZN(n1842) );
  OAI22_X1 U1487 ( .A1(n4673), .A2(n1189), .B1(n1404), .B2(n1184), .ZN(n1843)
         );
  AOI221_X1 U1488 ( .B1(n1194), .B2(n4961), .C1(n1191), .C2(n3648), .A(n1843), 
        .ZN(n1844) );
  NAND4_X1 U1489 ( .A1(n1847), .A2(n1845), .A3(n1844), .A4(n1846), .ZN(n2519)
         );
  AOI22_X1 U1490 ( .A1(n669), .A2(n4145), .B1(n1113), .B2(n4738), .ZN(n1848)
         );
  OAI221_X1 U1491 ( .B1(n150), .B2(n1119), .C1(n1849), .C2(n1116), .A(n1848), 
        .ZN(n1859) );
  AOI22_X1 U1492 ( .A1(n1024), .A2(n5058), .B1(n493), .B2(n5122), .ZN(n1850)
         );
  AOI22_X1 U1493 ( .A1(n54), .A2(n5090), .B1(n759), .B2(n1851), .ZN(n1852) );
  AOI22_X1 U1494 ( .A1(n1014), .A2(n5218), .B1(n490), .B2(n1853), .ZN(n1854)
         );
  OAI221_X1 U1495 ( .B1(n1855), .B2(n1140), .C1(n118), .C2(n1137), .A(n1854), 
        .ZN(n1856) );
  NOR4_X1 U1496 ( .A1(n1859), .A2(n1856), .A3(n1858), .A4(n1857), .ZN(n1860)
         );
  OAI222_X1 U1497 ( .A1(n822), .A2(n1149), .B1(n1860), .B2(n1146), .C1(n3663), 
        .C2(n1143), .ZN(n1861) );
  OAI22_X1 U1498 ( .A1(n3667), .A2(n1162), .B1(n950), .B2(n1158), .ZN(n1862)
         );
  AOI221_X1 U1499 ( .B1(n1167), .B2(n4802), .C1(n1164), .C2(n4325), .A(n1862), 
        .ZN(n1867) );
  OAI222_X1 U1500 ( .A1(n630), .A2(n1176), .B1(n3670), .B2(n1171), .C1(n3669), 
        .C2(n1170), .ZN(n1863) );
  AOI221_X1 U1501 ( .B1(n1181), .B2(n4273), .C1(n1178), .C2(n4241), .A(n1863), 
        .ZN(n1866) );
  OAI22_X1 U1502 ( .A1(n4674), .A2(n1188), .B1(n1406), .B2(n1184), .ZN(n1864)
         );
  AOI221_X1 U1503 ( .B1(n1194), .B2(n4962), .C1(n1191), .C2(n3673), .A(n1864), 
        .ZN(n1865) );
  NAND4_X1 U1504 ( .A1(n1866), .A2(n1868), .A3(n1867), .A4(n1865), .ZN(n2520)
         );
  AOI22_X1 U1505 ( .A1(n969), .A2(n4144), .B1(n1112), .B2(n4739), .ZN(n1869)
         );
  OAI221_X1 U1506 ( .B1(n149), .B2(n1119), .C1(n1870), .C2(n1114), .A(n1869), 
        .ZN(n1878) );
  AOI22_X1 U1507 ( .A1(n1024), .A2(n5059), .B1(n508), .B2(n5123), .ZN(n1871)
         );
  AOI22_X1 U1508 ( .A1(n54), .A2(n5091), .B1(n760), .B2(n220), .ZN(n1872) );
  OAI221_X1 U1509 ( .B1(n3682), .B2(n1135), .C1(n245), .C2(n506), .A(n1872), 
        .ZN(n1876) );
  AOI22_X1 U1510 ( .A1(n2211), .A2(n5219), .B1(n489), .B2(n221), .ZN(n1873) );
  NOR4_X1 U1511 ( .A1(n1878), .A2(n1876), .A3(n1877), .A4(n1875), .ZN(n1879)
         );
  OAI222_X1 U1512 ( .A1(n821), .A2(n1149), .B1(n1879), .B2(n1146), .C1(n3688), 
        .C2(n1143), .ZN(n1880) );
  OAI22_X1 U1513 ( .A1(n3692), .A2(n1161), .B1(n949), .B2(n1158), .ZN(n1881)
         );
  AOI221_X1 U1514 ( .B1(n1167), .B2(n4803), .C1(n1164), .C2(n4324), .A(n1881), 
        .ZN(n1886) );
  OAI222_X1 U1515 ( .A1(n629), .A2(n1176), .B1(n3695), .B2(n1171), .C1(n3694), 
        .C2(n1170), .ZN(n1882) );
  AOI221_X1 U1516 ( .B1(n1181), .B2(n4272), .C1(n1178), .C2(n4240), .A(n1882), 
        .ZN(n1885) );
  OAI22_X1 U1517 ( .A1(n4675), .A2(n1188), .B1(n1408), .B2(n1184), .ZN(n1883)
         );
  AOI221_X1 U1518 ( .B1(n1194), .B2(n4963), .C1(n1191), .C2(n3698), .A(n1883), 
        .ZN(n1884) );
  NAND4_X1 U1519 ( .A1(n1887), .A2(n1884), .A3(n1886), .A4(n1885), .ZN(n2521)
         );
  AOI22_X1 U1520 ( .A1(n669), .A2(n4143), .B1(n486), .B2(n4740), .ZN(n1888) );
  OAI221_X1 U1521 ( .B1(n148), .B2(n1117), .C1(n1889), .C2(n1115), .A(n1888), 
        .ZN(n1899) );
  AOI22_X1 U1522 ( .A1(n1123), .A2(n5060), .B1(n493), .B2(n5124), .ZN(n1890)
         );
  OAI221_X1 U1523 ( .B1(n3706), .B2(n1129), .C1(n276), .C2(n1126), .A(n1890), 
        .ZN(n1898) );
  AOI22_X1 U1524 ( .A1(n55), .A2(n5092), .B1(n1029), .B2(n1891), .ZN(n1892) );
  OAI221_X1 U1525 ( .B1(n3707), .B2(n1134), .C1(n506), .C2(n244), .A(n1892), 
        .ZN(n1897) );
  AOI22_X1 U1526 ( .A1(n2211), .A2(n5220), .B1(n489), .B2(n1893), .ZN(n1894)
         );
  NOR4_X1 U1527 ( .A1(n1899), .A2(n1898), .A3(n1897), .A4(n1896), .ZN(n1900)
         );
  OAI222_X1 U1528 ( .A1(n820), .A2(n1149), .B1(n1900), .B2(n1146), .C1(n3713), 
        .C2(n1143), .ZN(n1901) );
  OAI22_X1 U1529 ( .A1(n3717), .A2(n1162), .B1(n948), .B2(n1158), .ZN(n1902)
         );
  AOI221_X1 U1530 ( .B1(n1167), .B2(n4804), .C1(n1164), .C2(n4323), .A(n1902), 
        .ZN(n1907) );
  OAI22_X1 U1531 ( .A1(n4676), .A2(n1188), .B1(n1410), .B2(n1184), .ZN(n1904)
         );
  AOI221_X1 U1532 ( .B1(n1194), .B2(n4964), .C1(n1191), .C2(n3723), .A(n1904), 
        .ZN(n1905) );
  NAND4_X1 U1533 ( .A1(n1908), .A2(n1907), .A3(n1905), .A4(n1906), .ZN(n2522)
         );
  AOI22_X1 U1534 ( .A1(n669), .A2(n4142), .B1(n487), .B2(n4741), .ZN(n1909) );
  OAI221_X1 U1535 ( .B1(n147), .B2(n1119), .C1(n1910), .C2(n1115), .A(n1909), 
        .ZN(n1920) );
  AOI22_X1 U1536 ( .A1(n1024), .A2(n5061), .B1(n1120), .B2(n5125), .ZN(n1911)
         );
  OAI221_X1 U1537 ( .B1(n3731), .B2(n1128), .C1(n275), .C2(n1126), .A(n1911), 
        .ZN(n1919) );
  AOI22_X1 U1538 ( .A1(n57), .A2(n5093), .B1(n1029), .B2(n1912), .ZN(n1913) );
  OAI221_X1 U1539 ( .B1(n507), .B2(n3732), .C1(n243), .C2(n1131), .A(n1913), 
        .ZN(n1918) );
  AOI22_X1 U1540 ( .A1(n888), .A2(n5221), .B1(n966), .B2(n1914), .ZN(n1915) );
  OAI221_X1 U1541 ( .B1(n1916), .B2(n1140), .C1(n115), .C2(n1137), .A(n1915), 
        .ZN(n1917) );
  NOR4_X1 U1542 ( .A1(n1920), .A2(n1919), .A3(n1917), .A4(n1918), .ZN(n1921)
         );
  OAI22_X1 U1543 ( .A1(n3742), .A2(n707), .B1(n947), .B2(n1158), .ZN(n1922) );
  AOI221_X1 U1544 ( .B1(n1167), .B2(n4805), .C1(n1164), .C2(n4322), .A(n1922), 
        .ZN(n1927) );
  OAI22_X1 U1545 ( .A1(n4677), .A2(n1188), .B1(n1412), .B2(n1184), .ZN(n1924)
         );
  AOI221_X1 U1546 ( .B1(n1194), .B2(n4965), .C1(n1191), .C2(n3748), .A(n1924), 
        .ZN(n1925) );
  NAND4_X1 U1547 ( .A1(n1928), .A2(n1927), .A3(n1925), .A4(n1926), .ZN(n2523)
         );
  AOI22_X1 U1548 ( .A1(n669), .A2(n4141), .B1(n691), .B2(n4742), .ZN(n1929) );
  OAI221_X1 U1549 ( .B1(n146), .B2(n1119), .C1(n1930), .C2(n1116), .A(n1929), 
        .ZN(n1940) );
  AOI22_X1 U1550 ( .A1(n1122), .A2(n5062), .B1(n508), .B2(n5126), .ZN(n1931)
         );
  OAI221_X1 U1551 ( .B1(n3756), .B2(n1127), .C1(n274), .C2(n1126), .A(n1931), 
        .ZN(n1939) );
  AOI22_X1 U1552 ( .A1(n54), .A2(n5094), .B1(n1029), .B2(n1932), .ZN(n1933) );
  OAI221_X1 U1553 ( .B1(n3757), .B2(n1135), .C1(n242), .C2(n1131), .A(n1933), 
        .ZN(n1938) );
  AOI22_X1 U1554 ( .A1(n888), .A2(n5222), .B1(n578), .B2(n1934), .ZN(n1935) );
  NOR4_X1 U1555 ( .A1(n1940), .A2(n1939), .A3(n1938), .A4(n1937), .ZN(n1941)
         );
  OAI22_X1 U1556 ( .A1(n3767), .A2(n1161), .B1(n946), .B2(n1158), .ZN(n1942)
         );
  AOI221_X1 U1557 ( .B1(n1167), .B2(n4806), .C1(n1164), .C2(n4321), .A(n1942), 
        .ZN(n1947) );
  OAI22_X1 U1558 ( .A1(n4678), .A2(n1188), .B1(n1414), .B2(n1184), .ZN(n1944)
         );
  AOI221_X1 U1559 ( .B1(n1194), .B2(n4966), .C1(n1191), .C2(n3773), .A(n1944), 
        .ZN(n1945) );
  NAND4_X1 U1560 ( .A1(n1948), .A2(n1947), .A3(n1945), .A4(n1946), .ZN(n2524)
         );
  AOI22_X1 U1561 ( .A1(n969), .A2(n4140), .B1(n691), .B2(n4743), .ZN(n1949) );
  OAI221_X1 U1562 ( .B1(n145), .B2(n1118), .C1(n1950), .C2(n1115), .A(n1949), 
        .ZN(n1960) );
  AOI22_X1 U1563 ( .A1(n1123), .A2(n5063), .B1(n51), .B2(n5127), .ZN(n1951) );
  OAI221_X1 U1564 ( .B1(n3781), .B2(n1129), .C1(n273), .C2(n1126), .A(n1951), 
        .ZN(n1959) );
  AOI22_X1 U1565 ( .A1(n55), .A2(n5095), .B1(n759), .B2(n1952), .ZN(n1953) );
  OAI221_X1 U1566 ( .B1(n3782), .B2(n507), .C1(n241), .C2(n1131), .A(n1953), 
        .ZN(n1958) );
  AOI22_X1 U1567 ( .A1(n2211), .A2(n5223), .B1(n966), .B2(n1954), .ZN(n1955)
         );
  OAI221_X1 U1568 ( .B1(n1956), .B2(n1140), .C1(n113), .C2(n1137), .A(n1955), 
        .ZN(n1957) );
  NOR4_X1 U1569 ( .A1(n1960), .A2(n1959), .A3(n1957), .A4(n1958), .ZN(n1961)
         );
  OAI22_X1 U1570 ( .A1(n3792), .A2(n1161), .B1(n945), .B2(n1158), .ZN(n1962)
         );
  AOI221_X1 U1571 ( .B1(n1167), .B2(n4807), .C1(n1164), .C2(n4320), .A(n1962), 
        .ZN(n1967) );
  OAI22_X1 U1572 ( .A1(n4679), .A2(n1188), .B1(n1416), .B2(n1184), .ZN(n1964)
         );
  AOI221_X1 U1573 ( .B1(n1194), .B2(n4967), .C1(n1191), .C2(n3798), .A(n1964), 
        .ZN(n1965) );
  NAND4_X1 U1574 ( .A1(n1968), .A2(n1966), .A3(n1965), .A4(n1967), .ZN(n2525)
         );
  AOI22_X1 U1575 ( .A1(n669), .A2(n4139), .B1(n497), .B2(n4744), .ZN(n1969) );
  OAI221_X1 U1576 ( .B1(n144), .B2(n1119), .C1(n1970), .C2(n1116), .A(n1969), 
        .ZN(n1980) );
  AOI22_X1 U1577 ( .A1(n1023), .A2(n5064), .B1(n508), .B2(n5128), .ZN(n1971)
         );
  OAI221_X1 U1578 ( .B1(n3806), .B2(n1127), .C1(n272), .C2(n1126), .A(n1971), 
        .ZN(n1979) );
  AOI22_X1 U1579 ( .A1(n56), .A2(n5096), .B1(n1029), .B2(n1972), .ZN(n1973) );
  OAI221_X1 U1580 ( .B1(n3807), .B2(n1135), .C1(n240), .C2(n506), .A(n1973), 
        .ZN(n1978) );
  AOI22_X1 U1581 ( .A1(n1014), .A2(n5224), .B1(n578), .B2(n1974), .ZN(n1975)
         );
  OAI221_X1 U1582 ( .B1(n1976), .B2(n1140), .C1(n112), .C2(n1137), .A(n1975), 
        .ZN(n1977) );
  NOR4_X1 U1583 ( .A1(n1980), .A2(n1979), .A3(n1977), .A4(n1978), .ZN(n1981)
         );
  OAI222_X1 U1584 ( .A1(n816), .A2(n1149), .B1(n1981), .B2(n1146), .C1(n3813), 
        .C2(n1143), .ZN(n1982) );
  OAI22_X1 U1585 ( .A1(n3817), .A2(n1161), .B1(n944), .B2(n1158), .ZN(n1983)
         );
  AOI221_X1 U1586 ( .B1(n1167), .B2(n4808), .C1(n1164), .C2(n4319), .A(n1983), 
        .ZN(n1988) );
  OAI222_X1 U1587 ( .A1(n624), .A2(n1175), .B1(n3820), .B2(n1171), .C1(n3819), 
        .C2(n1170), .ZN(n1984) );
  AOI221_X1 U1588 ( .B1(n1181), .B2(n4267), .C1(n1178), .C2(n4235), .A(n1984), 
        .ZN(n1987) );
  OAI22_X1 U1589 ( .A1(n4680), .A2(n1188), .B1(n1418), .B2(n1184), .ZN(n1985)
         );
  AOI221_X1 U1590 ( .B1(n1194), .B2(n4968), .C1(n1191), .C2(n3823), .A(n1985), 
        .ZN(n1986) );
  NAND4_X1 U1591 ( .A1(n1989), .A2(n1986), .A3(n1988), .A4(n1987), .ZN(n2526)
         );
  AOI22_X1 U1592 ( .A1(n969), .A2(n4138), .B1(n1113), .B2(n4745), .ZN(n1990)
         );
  OAI221_X1 U1593 ( .B1(n143), .B2(n1118), .C1(n1991), .C2(n1116), .A(n1990), 
        .ZN(n2001) );
  AOI22_X1 U1594 ( .A1(n1124), .A2(n5065), .B1(n51), .B2(n5129), .ZN(n1992) );
  OAI221_X1 U1595 ( .B1(n3831), .B2(n1129), .C1(n271), .C2(n1126), .A(n1992), 
        .ZN(n2000) );
  AOI22_X1 U1596 ( .A1(n56), .A2(n5097), .B1(n760), .B2(n1993), .ZN(n1994) );
  AOI22_X1 U1597 ( .A1(n1014), .A2(n5225), .B1(n579), .B2(n1995), .ZN(n1996)
         );
  NOR4_X1 U1598 ( .A1(n2001), .A2(n2000), .A3(n1999), .A4(n1998), .ZN(n2002)
         );
  OAI22_X1 U1599 ( .A1(n3842), .A2(n1162), .B1(n943), .B2(n1158), .ZN(n2003)
         );
  AOI221_X1 U1600 ( .B1(n1167), .B2(n4809), .C1(n1164), .C2(n4318), .A(n2003), 
        .ZN(n2008) );
  OAI22_X1 U1601 ( .A1(n4681), .A2(n1188), .B1(n1420), .B2(n1184), .ZN(n2005)
         );
  AOI221_X1 U1602 ( .B1(n1194), .B2(n4969), .C1(n1191), .C2(n3848), .A(n2005), 
        .ZN(n2006) );
  NAND4_X1 U1603 ( .A1(n2009), .A2(n2008), .A3(n2006), .A4(n2007), .ZN(n2527)
         );
  AOI22_X1 U1604 ( .A1(n669), .A2(n4137), .B1(n738), .B2(n4746), .ZN(n2010) );
  OAI221_X1 U1605 ( .B1(n142), .B2(n1119), .C1(n2011), .C2(n1114), .A(n2010), 
        .ZN(n2021) );
  AOI22_X1 U1606 ( .A1(n1124), .A2(n5066), .B1(n493), .B2(n5130), .ZN(n2012)
         );
  OAI221_X1 U1607 ( .B1(n3856), .B2(n1128), .C1(n270), .C2(n1126), .A(n2012), 
        .ZN(n2020) );
  AOI22_X1 U1608 ( .A1(n54), .A2(n5098), .B1(n760), .B2(n2013), .ZN(n2014) );
  OAI221_X1 U1609 ( .B1(n3857), .B2(n1133), .C1(n238), .C2(n1130), .A(n2014), 
        .ZN(n2019) );
  AOI22_X1 U1610 ( .A1(n1014), .A2(n5226), .B1(n490), .B2(n2015), .ZN(n2016)
         );
  NOR4_X1 U1611 ( .A1(n2021), .A2(n2020), .A3(n2018), .A4(n2019), .ZN(n2022)
         );
  OAI222_X1 U1612 ( .A1(n814), .A2(n1149), .B1(n2022), .B2(n1146), .C1(n3863), 
        .C2(n1143), .ZN(n2023) );
  OAI22_X1 U1613 ( .A1(n3867), .A2(n1160), .B1(n942), .B2(n1158), .ZN(n2024)
         );
  AOI221_X1 U1614 ( .B1(n1167), .B2(n4810), .C1(n1164), .C2(n4317), .A(n2024), 
        .ZN(n2029) );
  OAI222_X1 U1615 ( .A1(n622), .A2(n1175), .B1(n3870), .B2(n1172), .C1(n3869), 
        .C2(n1170), .ZN(n2025) );
  AOI221_X1 U1616 ( .B1(n1181), .B2(n4265), .C1(n1178), .C2(n4233), .A(n2025), 
        .ZN(n2028) );
  OAI22_X1 U1617 ( .A1(n4682), .A2(n1188), .B1(n1422), .B2(n1184), .ZN(n2026)
         );
  AOI221_X1 U1618 ( .B1(n1194), .B2(n4970), .C1(n1191), .C2(n3873), .A(n2026), 
        .ZN(n2027) );
  NAND4_X1 U1619 ( .A1(n2030), .A2(n2029), .A3(n2027), .A4(n2028), .ZN(n2528)
         );
  AOI22_X1 U1620 ( .A1(n969), .A2(n4136), .B1(n487), .B2(n4747), .ZN(n2031) );
  OAI221_X1 U1621 ( .B1(n141), .B2(n1119), .C1(n2032), .C2(n1116), .A(n2031), 
        .ZN(n2042) );
  AOI22_X1 U1622 ( .A1(n1124), .A2(n5067), .B1(n512), .B2(n5131), .ZN(n2033)
         );
  OAI221_X1 U1623 ( .B1(n3881), .B2(n1127), .C1(n269), .C2(n1126), .A(n2033), 
        .ZN(n2041) );
  AOI22_X1 U1624 ( .A1(n54), .A2(n5099), .B1(n759), .B2(n2034), .ZN(n2035) );
  OAI221_X1 U1625 ( .B1(n3882), .B2(n1133), .C1(n237), .C2(n506), .A(n2035), 
        .ZN(n2040) );
  AOI22_X1 U1626 ( .A1(n1014), .A2(n5227), .B1(n577), .B2(n2036), .ZN(n2037)
         );
  NOR4_X1 U1627 ( .A1(n2042), .A2(n2041), .A3(n2039), .A4(n2040), .ZN(n2043)
         );
  OAI222_X1 U1628 ( .A1(n813), .A2(n1149), .B1(n2043), .B2(n1146), .C1(n3888), 
        .C2(n1143), .ZN(n2044) );
  OAI22_X1 U1629 ( .A1(n3892), .A2(n1160), .B1(n941), .B2(n1158), .ZN(n2045)
         );
  AOI221_X1 U1630 ( .B1(n1167), .B2(n4811), .C1(n1164), .C2(n4316), .A(n2045), 
        .ZN(n2050) );
  OAI222_X1 U1631 ( .A1(n621), .A2(n1176), .B1(n3895), .B2(n1172), .C1(n3894), 
        .C2(n1170), .ZN(n2046) );
  AOI221_X1 U1632 ( .B1(n1181), .B2(n4264), .C1(n1178), .C2(n4232), .A(n2046), 
        .ZN(n2049) );
  OAI22_X1 U1633 ( .A1(n4683), .A2(n1188), .B1(n1424), .B2(n1184), .ZN(n2047)
         );
  AOI221_X1 U1634 ( .B1(n1194), .B2(n4971), .C1(n1191), .C2(n3898), .A(n2047), 
        .ZN(n2048) );
  NAND4_X1 U1635 ( .A1(n2051), .A2(n2050), .A3(n2048), .A4(n2049), .ZN(n2529)
         );
  AOI22_X1 U1636 ( .A1(n969), .A2(n4135), .B1(n1113), .B2(n4748), .ZN(n2052)
         );
  OAI221_X1 U1637 ( .B1(n140), .B2(n1119), .C1(n2053), .C2(n1114), .A(n2052), 
        .ZN(n2063) );
  AOI22_X1 U1638 ( .A1(n1016), .A2(n5068), .B1(n512), .B2(n5132), .ZN(n2054)
         );
  OAI221_X1 U1639 ( .B1(n3907), .B2(n1129), .C1(n268), .C2(n678), .A(n2054), 
        .ZN(n2062) );
  AOI22_X1 U1640 ( .A1(n56), .A2(n5100), .B1(n760), .B2(n2055), .ZN(n2056) );
  OAI221_X1 U1641 ( .B1(n3908), .B2(n1133), .C1(n236), .C2(n1131), .A(n2056), 
        .ZN(n2061) );
  AOI22_X1 U1642 ( .A1(n888), .A2(n5228), .B1(n490), .B2(n2057), .ZN(n2058) );
  OAI221_X1 U1643 ( .B1(n2059), .B2(n1141), .C1(n108), .C2(n1138), .A(n2058), 
        .ZN(n2060) );
  NOR4_X1 U1644 ( .A1(n2063), .A2(n2062), .A3(n2060), .A4(n2061), .ZN(n2064)
         );
  OAI22_X1 U1645 ( .A1(n3918), .A2(n1160), .B1(n940), .B2(n1159), .ZN(n2066)
         );
  AOI221_X1 U1646 ( .B1(n1168), .B2(n4812), .C1(n1165), .C2(n4315), .A(n2066), 
        .ZN(n2071) );
  OAI222_X1 U1647 ( .A1(n620), .A2(n1175), .B1(n3921), .B2(n1172), .C1(n3920), 
        .C2(n876), .ZN(n2067) );
  AOI221_X1 U1648 ( .B1(n1182), .B2(n4263), .C1(n1179), .C2(n4231), .A(n2067), 
        .ZN(n2070) );
  OAI22_X1 U1649 ( .A1(n4684), .A2(n1188), .B1(n1427), .B2(n1185), .ZN(n2068)
         );
  AOI221_X1 U1650 ( .B1(n1195), .B2(n4972), .C1(n1192), .C2(n3924), .A(n2068), 
        .ZN(n2069) );
  NAND4_X1 U1651 ( .A1(n2072), .A2(n2071), .A3(n2069), .A4(n2070), .ZN(n2530)
         );
  AOI22_X1 U1652 ( .A1(n669), .A2(n4134), .B1(n1112), .B2(n4749), .ZN(n2073)
         );
  OAI221_X1 U1653 ( .B1(n139), .B2(n1119), .C1(n2074), .C2(n1116), .A(n2073), 
        .ZN(n2084) );
  AOI22_X1 U1654 ( .A1(n1123), .A2(n5069), .B1(n52), .B2(n5133), .ZN(n2075) );
  OAI221_X1 U1655 ( .B1(n3933), .B2(n1127), .C1(n267), .C2(n678), .A(n2075), 
        .ZN(n2083) );
  AOI22_X1 U1656 ( .A1(n56), .A2(n5101), .B1(n760), .B2(n2076), .ZN(n2077) );
  OAI221_X1 U1657 ( .B1(n3934), .B2(n1133), .C1(n235), .C2(n1130), .A(n2077), 
        .ZN(n2082) );
  AOI22_X1 U1658 ( .A1(n1014), .A2(n5229), .B1(n490), .B2(n2078), .ZN(n2079)
         );
  OAI221_X1 U1659 ( .B1(n2080), .B2(n1141), .C1(n107), .C2(n1138), .A(n2079), 
        .ZN(n2081) );
  NOR4_X1 U1660 ( .A1(n2084), .A2(n2083), .A3(n2081), .A4(n2082), .ZN(n2085)
         );
  OAI222_X1 U1661 ( .A1(n811), .A2(n1150), .B1(n2085), .B2(n1147), .C1(n3940), 
        .C2(n1144), .ZN(n2086) );
  OAI22_X1 U1662 ( .A1(n3944), .A2(n1162), .B1(n939), .B2(n1159), .ZN(n2087)
         );
  OAI222_X1 U1663 ( .A1(n619), .A2(n1176), .B1(n3947), .B2(n1172), .C1(n3946), 
        .C2(n876), .ZN(n2088) );
  AOI221_X1 U1664 ( .B1(n1182), .B2(n4262), .C1(n1179), .C2(n4230), .A(n2088), 
        .ZN(n2091) );
  OAI22_X1 U1665 ( .A1(n4685), .A2(n1187), .B1(n1430), .B2(n1185), .ZN(n2089)
         );
  AOI221_X1 U1666 ( .B1(n1195), .B2(n4973), .C1(n1192), .C2(n3950), .A(n2089), 
        .ZN(n2090) );
  NAND4_X1 U1667 ( .A1(n2093), .A2(n2092), .A3(n2090), .A4(n2091), .ZN(n2531)
         );
  AOI22_X1 U1668 ( .A1(n668), .A2(n4133), .B1(n1113), .B2(n4750), .ZN(n2094)
         );
  OAI221_X1 U1669 ( .B1(n138), .B2(n1119), .C1(n2095), .C2(n1114), .A(n2094), 
        .ZN(n2105) );
  AOI22_X1 U1670 ( .A1(n1016), .A2(n5070), .B1(n1120), .B2(n5134), .ZN(n2096)
         );
  AOI22_X1 U1671 ( .A1(n57), .A2(n5102), .B1(n1029), .B2(n2097), .ZN(n2098) );
  OAI221_X1 U1672 ( .B1(n3960), .B2(n1135), .C1(n234), .C2(n506), .A(n2098), 
        .ZN(n2103) );
  AOI22_X1 U1673 ( .A1(n888), .A2(n5230), .B1(n577), .B2(n2099), .ZN(n2100) );
  OAI221_X1 U1674 ( .B1(n2101), .B2(n1141), .C1(n106), .C2(n1138), .A(n2100), 
        .ZN(n2102) );
  NOR4_X1 U1675 ( .A1(n2105), .A2(n2102), .A3(n2103), .A4(n2104), .ZN(n2106)
         );
  OAI222_X1 U1676 ( .A1(n810), .A2(n1150), .B1(n2106), .B2(n1147), .C1(n3966), 
        .C2(n1144), .ZN(n2107) );
  OAI22_X1 U1677 ( .A1(n3970), .A2(n1160), .B1(n938), .B2(n1159), .ZN(n2108)
         );
  AOI221_X1 U1678 ( .B1(n1168), .B2(n4814), .C1(n1165), .C2(n4313), .A(n2108), 
        .ZN(n2113) );
  OAI222_X1 U1679 ( .A1(n618), .A2(n1176), .B1(n3973), .B2(n1173), .C1(n3972), 
        .C2(n876), .ZN(n2109) );
  AOI221_X1 U1680 ( .B1(n1182), .B2(n4261), .C1(n1179), .C2(n4229), .A(n2109), 
        .ZN(n2112) );
  OAI22_X1 U1681 ( .A1(n4686), .A2(n1187), .B1(n1433), .B2(n1185), .ZN(n2110)
         );
  AOI221_X1 U1682 ( .B1(n1195), .B2(n4974), .C1(n1192), .C2(n3976), .A(n2110), 
        .ZN(n2111) );
  NAND4_X1 U1683 ( .A1(n2112), .A2(n2113), .A3(n2111), .A4(n2114), .ZN(n2532)
         );
  AOI22_X1 U1684 ( .A1(n969), .A2(n4132), .B1(n497), .B2(n4751), .ZN(n2115) );
  OAI221_X1 U1685 ( .B1(n137), .B2(n1118), .C1(n2116), .C2(n1115), .A(n2115), 
        .ZN(n2126) );
  AOI22_X1 U1686 ( .A1(n1023), .A2(n5071), .B1(n493), .B2(n5135), .ZN(n2117)
         );
  OAI221_X1 U1687 ( .B1(n3985), .B2(n1128), .C1(n265), .C2(n678), .A(n2117), 
        .ZN(n2125) );
  AOI22_X1 U1688 ( .A1(n57), .A2(n5103), .B1(n759), .B2(n2118), .ZN(n2119) );
  OAI221_X1 U1689 ( .B1(n3986), .B2(n1133), .C1(n233), .C2(n506), .A(n2119), 
        .ZN(n2124) );
  AOI22_X1 U1690 ( .A1(n888), .A2(n5231), .B1(n966), .B2(n2120), .ZN(n2121) );
  OAI221_X1 U1691 ( .B1(n2122), .B2(n1141), .C1(n105), .C2(n1138), .A(n2121), 
        .ZN(n2123) );
  NOR4_X1 U1692 ( .A1(n2126), .A2(n2125), .A3(n2124), .A4(n2123), .ZN(n2127)
         );
  OAI222_X1 U1693 ( .A1(n809), .A2(n1150), .B1(n2127), .B2(n1147), .C1(n3992), 
        .C2(n1144), .ZN(n2128) );
  OAI22_X1 U1694 ( .A1(n3996), .A2(n1160), .B1(n937), .B2(n1159), .ZN(n2129)
         );
  AOI221_X1 U1695 ( .B1(n1168), .B2(n4815), .C1(n1165), .C2(n4312), .A(n2129), 
        .ZN(n2134) );
  OAI222_X1 U1696 ( .A1(n617), .A2(n1174), .B1(n1173), .B2(n3999), .C1(n3998), 
        .C2(n876), .ZN(n2130) );
  AOI221_X1 U1697 ( .B1(n1182), .B2(n4260), .C1(n1179), .C2(n4228), .A(n2130), 
        .ZN(n2133) );
  OAI22_X1 U1698 ( .A1(n4687), .A2(n1187), .B1(n1436), .B2(n1185), .ZN(n2131)
         );
  AOI221_X1 U1699 ( .B1(n1195), .B2(n4975), .C1(n1192), .C2(n4002), .A(n2131), 
        .ZN(n2132) );
  NAND4_X1 U1700 ( .A1(n2133), .A2(n2132), .A3(n2135), .A4(n2134), .ZN(n2533)
         );
  AOI22_X1 U1701 ( .A1(n969), .A2(n4131), .B1(n1111), .B2(n4752), .ZN(n2136)
         );
  OAI221_X1 U1702 ( .B1(n136), .B2(n1118), .C1(n2137), .C2(n1116), .A(n2136), 
        .ZN(n2147) );
  AOI22_X1 U1703 ( .A1(n1023), .A2(n5072), .B1(n1121), .B2(n5136), .ZN(n2138)
         );
  OAI221_X1 U1704 ( .B1(n4011), .B2(n1129), .C1(n264), .C2(n678), .A(n2138), 
        .ZN(n2146) );
  AOI22_X1 U1705 ( .A1(n57), .A2(n5104), .B1(n759), .B2(n2139), .ZN(n2140) );
  OAI221_X1 U1706 ( .B1(n4012), .B2(n1133), .C1(n232), .C2(n506), .A(n2140), 
        .ZN(n2145) );
  AOI22_X1 U1707 ( .A1(n888), .A2(n5232), .B1(n966), .B2(n2141), .ZN(n2142) );
  OAI221_X1 U1708 ( .B1(n2143), .B2(n1141), .C1(n104), .C2(n1138), .A(n2142), 
        .ZN(n2144) );
  NOR4_X1 U1709 ( .A1(n2147), .A2(n2146), .A3(n2145), .A4(n2144), .ZN(n2148)
         );
  OAI222_X1 U1710 ( .A1(n808), .A2(n1150), .B1(n2148), .B2(n1147), .C1(n4018), 
        .C2(n1144), .ZN(n2149) );
  OAI22_X1 U1711 ( .A1(n4022), .A2(n1160), .B1(n936), .B2(n1159), .ZN(n2150)
         );
  AOI221_X1 U1712 ( .B1(n1168), .B2(n4816), .C1(n1165), .C2(n4311), .A(n2150), 
        .ZN(n2155) );
  OAI222_X1 U1713 ( .A1(n616), .A2(n1175), .B1(n4025), .B2(n1172), .C1(n4024), 
        .C2(n876), .ZN(n2151) );
  AOI221_X1 U1714 ( .B1(n1182), .B2(n4259), .C1(n1179), .C2(n4227), .A(n2151), 
        .ZN(n2154) );
  OAI22_X1 U1715 ( .A1(n4688), .A2(n1187), .B1(n1439), .B2(n1185), .ZN(n2152)
         );
  AOI221_X1 U1716 ( .B1(n1195), .B2(n4976), .C1(n1192), .C2(n4028), .A(n2152), 
        .ZN(n2153) );
  NAND4_X1 U1717 ( .A1(n2154), .A2(n2155), .A3(n2153), .A4(n2156), .ZN(n2534)
         );
  AOI22_X1 U1718 ( .A1(n668), .A2(n4130), .B1(n1112), .B2(n4753), .ZN(n2157)
         );
  OAI221_X1 U1719 ( .B1(n135), .B2(n1118), .C1(n2158), .C2(n1116), .A(n2157), 
        .ZN(n2168) );
  AOI22_X1 U1720 ( .A1(n1123), .A2(n5073), .B1(n51), .B2(n5137), .ZN(n2159) );
  OAI221_X1 U1721 ( .B1(n4037), .B2(n1128), .C1(n263), .C2(n678), .A(n2159), 
        .ZN(n2167) );
  AOI22_X1 U1722 ( .A1(n56), .A2(n5105), .B1(n1029), .B2(n2160), .ZN(n2161) );
  OAI221_X1 U1723 ( .B1(n4038), .B2(n507), .C1(n231), .C2(n506), .A(n2161), 
        .ZN(n2166) );
  AOI22_X1 U1724 ( .A1(n2211), .A2(n5233), .B1(n577), .B2(n2162), .ZN(n2163)
         );
  OAI221_X1 U1725 ( .B1(n2164), .B2(n1141), .C1(n103), .C2(n1138), .A(n2163), 
        .ZN(n2165) );
  NOR4_X1 U1726 ( .A1(n2168), .A2(n2167), .A3(n2165), .A4(n2166), .ZN(n2169)
         );
  OAI22_X1 U1727 ( .A1(n4048), .A2(n1160), .B1(n935), .B2(n1159), .ZN(n2171)
         );
  AOI221_X1 U1728 ( .B1(n1168), .B2(n4817), .C1(n1165), .C2(n4310), .A(n2171), 
        .ZN(n2176) );
  OAI222_X1 U1729 ( .A1(n615), .A2(n1174), .B1(n1171), .B2(n4051), .C1(n4050), 
        .C2(n876), .ZN(n2172) );
  AOI221_X1 U1730 ( .B1(n1182), .B2(n4258), .C1(n1179), .C2(n4226), .A(n2172), 
        .ZN(n2175) );
  OAI22_X1 U1731 ( .A1(n4689), .A2(n1187), .B1(n1442), .B2(n1185), .ZN(n2173)
         );
  AOI221_X1 U1732 ( .B1(n1195), .B2(n4977), .C1(n1192), .C2(n4054), .A(n2173), 
        .ZN(n2174) );
  NAND4_X1 U1733 ( .A1(n2177), .A2(n2176), .A3(n2174), .A4(n2175), .ZN(n2535)
         );
  AOI22_X1 U1734 ( .A1(n969), .A2(n4129), .B1(n1111), .B2(n4754), .ZN(n2178)
         );
  OAI221_X1 U1735 ( .B1(n134), .B2(n1117), .C1(n2179), .C2(n1115), .A(n2178), 
        .ZN(n2189) );
  AOI22_X1 U1736 ( .A1(n1016), .A2(n5074), .B1(n512), .B2(n5138), .ZN(n2180)
         );
  AOI22_X1 U1737 ( .A1(n57), .A2(n5106), .B1(n759), .B2(n2181), .ZN(n2182) );
  OAI221_X1 U1738 ( .B1(n4064), .B2(n1135), .C1(n230), .C2(n506), .A(n2182), 
        .ZN(n2187) );
  AOI22_X1 U1739 ( .A1(n2211), .A2(n5234), .B1(n966), .B2(n2183), .ZN(n2184)
         );
  NOR4_X1 U1740 ( .A1(n2189), .A2(n2187), .A3(n2188), .A4(n2186), .ZN(n2190)
         );
  OAI222_X1 U1741 ( .A1(n806), .A2(n1150), .B1(n2190), .B2(n1147), .C1(n4070), 
        .C2(n1144), .ZN(n2191) );
  OAI22_X1 U1742 ( .A1(n4074), .A2(n1160), .B1(n934), .B2(n1159), .ZN(n2192)
         );
  AOI221_X1 U1743 ( .B1(n1168), .B2(n4818), .C1(n1165), .C2(n4309), .A(n2192), 
        .ZN(n2197) );
  OAI222_X1 U1744 ( .A1(n614), .A2(n1174), .B1(n1171), .B2(n4077), .C1(n4076), 
        .C2(n876), .ZN(n2193) );
  AOI221_X1 U1745 ( .B1(n1182), .B2(n4257), .C1(n1179), .C2(n4225), .A(n2193), 
        .ZN(n2196) );
  OAI22_X1 U1746 ( .A1(n4690), .A2(n1187), .B1(n1445), .B2(n1185), .ZN(n2194)
         );
  AOI221_X1 U1747 ( .B1(n1195), .B2(n4978), .C1(n1192), .C2(n4080), .A(n2194), 
        .ZN(n2195) );
  NAND4_X1 U1748 ( .A1(n2198), .A2(n2197), .A3(n2195), .A4(n2196), .ZN(n2536)
         );
  AOI22_X1 U1749 ( .A1(n668), .A2(n4128), .B1(n497), .B2(n4755), .ZN(n2199) );
  OAI221_X1 U1750 ( .B1(n133), .B2(n1119), .C1(n2201), .C2(n1115), .A(n2199), 
        .ZN(n2219) );
  AOI22_X1 U1751 ( .A1(n1023), .A2(n5075), .B1(n508), .B2(n5139), .ZN(n2203)
         );
  AOI22_X1 U1752 ( .A1(n55), .A2(n5107), .B1(n760), .B2(n2206), .ZN(n2207) );
  OAI221_X1 U1753 ( .B1(n4095), .B2(n1135), .C1(n229), .C2(n1130), .A(n2207), 
        .ZN(n2217) );
  AOI22_X1 U1754 ( .A1(n2211), .A2(n5235), .B1(n579), .B2(n2210), .ZN(n2212)
         );
  OAI221_X1 U1755 ( .B1(n2215), .B2(n1141), .C1(n101), .C2(n1138), .A(n2212), 
        .ZN(n2216) );
  NOR4_X1 U1756 ( .A1(n2219), .A2(n2218), .A3(n2216), .A4(n2217), .ZN(n2222)
         );
  OAI22_X1 U1757 ( .A1(n4112), .A2(n1160), .B1(n933), .B2(n1159), .ZN(n2227)
         );
  AOI221_X1 U1758 ( .B1(n1168), .B2(n4819), .C1(n1165), .C2(n4308), .A(n2227), 
        .ZN(n2236) );
  OAI222_X1 U1759 ( .A1(n613), .A2(n1176), .B1(n4117), .B2(n1173), .C1(n4115), 
        .C2(n876), .ZN(n2231) );
  OAI22_X1 U1760 ( .A1(n4691), .A2(n1188), .B1(n1448), .B2(n1185), .ZN(n2233)
         );
  AOI221_X1 U1761 ( .B1(n1195), .B2(n4979), .C1(n1192), .C2(n4123), .A(n2233), 
        .ZN(n2234) );
  NAND4_X1 U1762 ( .A1(n2237), .A2(n2236), .A3(n2234), .A4(n2235), .ZN(n2537)
         );
  NAND2_X1 U1763 ( .A1(ADD_RS2[1]), .A2(ADD_RS2[2]), .ZN(n2238) );
  INV_X1 U1764 ( .A(n2238), .ZN(n2260) );
  INV_X1 U1765 ( .A(ADD_RS2[2]), .ZN(n2240) );
  INV_X1 U1766 ( .A(ADD_RS2[0]), .ZN(n2259) );
  NAND4_X1 U1767 ( .A1(n980), .A2(n973), .A3(n1274), .A4(n926), .ZN(n4108) );
  INV_X1 U1768 ( .A(ADD_RS2[1]), .ZN(n2239) );
  NAND2_X1 U1769 ( .A1(n976), .A2(n878), .ZN(n4088) );
  NAND2_X1 U1770 ( .A1(n2239), .A2(n2240), .ZN(n2241) );
  INV_X1 U1771 ( .A(n2241), .ZN(n2265) );
  INV_X1 U1772 ( .A(ADD_RS2[4]), .ZN(n2243) );
  NAND2_X1 U1773 ( .A1(n975), .A2(n2265), .ZN(n4087) );
  AOI22_X1 U1774 ( .A1(n1200), .A2(n194), .B1(n1198), .B2(n4159), .ZN(n2242)
         );
  OAI221_X1 U1775 ( .B1(n1207), .B2(n227), .C1(n260), .C2(n1202), .A(n2242), 
        .ZN(n2252) );
  NAND2_X1 U1776 ( .A1(n975), .A2(n1036), .ZN(n4091) );
  NAND2_X1 U1777 ( .A1(n7), .A2(n974), .ZN(n4090) );
  AOI22_X1 U1778 ( .A1(n689), .A2(n4223), .B1(n879), .B2(n4191), .ZN(n2244) );
  OAI221_X1 U1779 ( .B1(n388), .B2(n6), .C1(n420), .C2(n1210), .A(n2244), .ZN(
        n2251) );
  NAND2_X1 U1780 ( .A1(n975), .A2(n2260), .ZN(n4096) );
  NAND2_X1 U1781 ( .A1(n2260), .A2(n974), .ZN(n4094) );
  AOI22_X1 U1782 ( .A1(n5108), .A2(n704), .B1(n5140), .B2(n1216), .ZN(n2245)
         );
  OAI221_X1 U1783 ( .B1(n1223), .B2(n2247), .C1(n1219), .C2(n2246), .A(n2245), 
        .ZN(n2250) );
  NAND2_X1 U1784 ( .A1(n975), .A2(n973), .ZN(n4099) );
  NAND2_X1 U1785 ( .A1(n974), .A2(n973), .ZN(n4098) );
  AOI22_X1 U1786 ( .A1(n5172), .A2(n932), .B1(n5204), .B2(n750), .ZN(n2248) );
  NOR4_X1 U1787 ( .A1(n2252), .A2(n2251), .A3(n2250), .A4(n2249), .ZN(n2254)
         );
  NAND2_X1 U1788 ( .A1(n1275), .A2(n926), .ZN(n4106) );
  NAND4_X1 U1789 ( .A1(n980), .A2(n703), .A3(n1274), .A4(n925), .ZN(n4105) );
  OAI222_X1 U1790 ( .A1(n836), .A2(n1237), .B1(n2254), .B2(n1234), .C1(n1231), 
        .C2(n2253), .ZN(n2255) );
  NAND4_X1 U1791 ( .A1(n980), .A2(n878), .A3(n1274), .A4(n926), .ZN(n4113) );
  NAND4_X1 U1792 ( .A1(n925), .A2(n2260), .A3(n1274), .A4(n980), .ZN(n4111) );
  OAI22_X1 U1793 ( .A1(n509), .A2(n2257), .B1(n964), .B2(n480), .ZN(n2258) );
  AOI221_X1 U1794 ( .B1(n4788), .B2(n1255), .C1(n1250), .C2(n4339), .A(n2258), 
        .ZN(n2270) );
  NAND4_X1 U1795 ( .A1(n2264), .A2(n878), .A3(n1274), .A4(n1001), .ZN(n4119)
         );
  NAND4_X1 U1796 ( .A1(n2264), .A2(n2260), .A3(n1274), .A4(n1001), .ZN(n4118)
         );
  NAND4_X1 U1797 ( .A1(n2264), .A2(n973), .A3(n1275), .A4(n979), .ZN(n4116) );
  OAI222_X1 U1798 ( .A1(n644), .A2(n1262), .B1(n1259), .B2(n2262), .C1(n1258), 
        .C2(n2261), .ZN(n2263) );
  AOI221_X1 U1799 ( .B1(n1268), .B2(n4287), .C1(n1265), .C2(n4255), .A(n2263), 
        .ZN(n2269) );
  NAND3_X1 U1800 ( .A1(n1275), .A2(n893), .A3(n470), .ZN(n4121) );
  OAI22_X1 U1801 ( .A1(n4692), .A2(n1275), .B1(n1378), .B2(n1271), .ZN(n2266)
         );
  AOI221_X1 U1802 ( .B1(n4948), .B2(n1281), .C1(n1278), .C2(n2267), .A(n2266), 
        .ZN(n2268) );
  NAND4_X1 U1803 ( .A1(n2271), .A2(n2270), .A3(n2269), .A4(n2268), .ZN(n2538)
         );
  AOI22_X1 U1804 ( .A1(n1201), .A2(n195), .B1(n495), .B2(n4158), .ZN(n2272) );
  OAI221_X1 U1805 ( .B1(n1206), .B2(n228), .C1(n259), .C2(n1202), .A(n2272), 
        .ZN(n2281) );
  AOI22_X1 U1806 ( .A1(n689), .A2(n4222), .B1(n879), .B2(n4190), .ZN(n2273) );
  OAI221_X1 U1807 ( .B1(n387), .B2(n1213), .C1(n419), .C2(n1212), .A(n2273), 
        .ZN(n2280) );
  AOI22_X1 U1808 ( .A1(n5109), .A2(n589), .B1(n5141), .B2(n1216), .ZN(n2274)
         );
  OAI221_X1 U1809 ( .B1(n1222), .B2(n2276), .C1(n1219), .C2(n2275), .A(n2274), 
        .ZN(n2279) );
  AOI22_X1 U1810 ( .A1(n5173), .A2(n2), .B1(n5205), .B2(n931), .ZN(n2277) );
  NOR4_X1 U1811 ( .A1(n2281), .A2(n2280), .A3(n2279), .A4(n2278), .ZN(n2283)
         );
  OAI222_X1 U1812 ( .A1(n835), .A2(n1237), .B1(n2283), .B2(n1234), .C1(n1231), 
        .C2(n2282), .ZN(n2284) );
  OAI22_X1 U1813 ( .A1(n1249), .A2(n2286), .B1(n963), .B2(n1246), .ZN(n2287)
         );
  AOI221_X1 U1814 ( .B1(n4789), .B2(n33), .C1(n1250), .C2(n4338), .A(n2287), 
        .ZN(n2295) );
  OAI222_X1 U1815 ( .A1(n643), .A2(n1262), .B1(n1259), .B2(n2289), .C1(n1256), 
        .C2(n2288), .ZN(n2290) );
  AOI221_X1 U1816 ( .B1(n1268), .B2(n4286), .C1(n1265), .C2(n4254), .A(n2290), 
        .ZN(n2294) );
  OAI22_X1 U1817 ( .A1(n4693), .A2(n1277), .B1(n1380), .B2(n1271), .ZN(n2291)
         );
  AOI221_X1 U1818 ( .B1(n4949), .B2(n1281), .C1(n1278), .C2(n2292), .A(n2291), 
        .ZN(n2293) );
  NAND4_X1 U1819 ( .A1(n2296), .A2(n2295), .A3(n2294), .A4(n2293), .ZN(n2539)
         );
  AOI22_X1 U1820 ( .A1(n1200), .A2(n196), .B1(n1196), .B2(n4157), .ZN(n2297)
         );
  OAI221_X1 U1821 ( .B1(n1207), .B2(n293), .C1(n258), .C2(n1202), .A(n2297), 
        .ZN(n2306) );
  AOI22_X1 U1822 ( .A1(n998), .A2(n4221), .B1(n879), .B2(n4189), .ZN(n2298) );
  AOI22_X1 U1823 ( .A1(n5110), .A2(n704), .B1(n5142), .B2(n1216), .ZN(n2299)
         );
  OAI221_X1 U1824 ( .B1(n1224), .B2(n2301), .C1(n1219), .C2(n2300), .A(n2299), 
        .ZN(n2304) );
  AOI22_X1 U1825 ( .A1(n5174), .A2(n932), .B1(n5206), .B2(n931), .ZN(n2302) );
  OAI221_X1 U1826 ( .B1(n1230), .B2(n173), .C1(n1225), .C2(n322), .A(n2302), 
        .ZN(n2303) );
  NOR4_X1 U1827 ( .A1(n2306), .A2(n2303), .A3(n2305), .A4(n2304), .ZN(n2308)
         );
  OAI222_X1 U1828 ( .A1(n834), .A2(n1237), .B1(n2308), .B2(n1234), .C1(n1231), 
        .C2(n2307), .ZN(n2309) );
  OAI22_X1 U1829 ( .A1(n1248), .A2(n2311), .B1(n962), .B2(n1246), .ZN(n2312)
         );
  AOI221_X1 U1830 ( .B1(n4790), .B2(n33), .C1(n1250), .C2(n4337), .A(n2312), 
        .ZN(n2320) );
  OAI222_X1 U1831 ( .A1(n642), .A2(n1262), .B1(n1260), .B2(n2314), .C1(n1256), 
        .C2(n2313), .ZN(n2315) );
  AOI221_X1 U1832 ( .B1(n1268), .B2(n4285), .C1(n1265), .C2(n4253), .A(n2315), 
        .ZN(n2319) );
  OAI22_X1 U1833 ( .A1(n4694), .A2(n1277), .B1(n1382), .B2(n1271), .ZN(n2316)
         );
  AOI221_X1 U1834 ( .B1(n4950), .B2(n1281), .C1(n1278), .C2(n2317), .A(n2316), 
        .ZN(n2318) );
  NAND4_X1 U1835 ( .A1(n2321), .A2(n2320), .A3(n2319), .A4(n2318), .ZN(n2540)
         );
  AOI22_X1 U1836 ( .A1(n66), .A2(n197), .B1(n1196), .B2(n4156), .ZN(n2322) );
  OAI221_X1 U1837 ( .B1(n1206), .B2(n294), .C1(n257), .C2(n1202), .A(n2322), 
        .ZN(n2331) );
  AOI22_X1 U1838 ( .A1(n998), .A2(n4220), .B1(n879), .B2(n4188), .ZN(n2323) );
  AOI22_X1 U1839 ( .A1(n5111), .A2(n987), .B1(n5143), .B2(n1216), .ZN(n2324)
         );
  OAI221_X1 U1840 ( .B1(n1222), .B2(n2326), .C1(n1219), .C2(n2325), .A(n2324), 
        .ZN(n2329) );
  AOI22_X1 U1841 ( .A1(n5175), .A2(n1), .B1(n5207), .B2(n40), .ZN(n2327) );
  OAI221_X1 U1842 ( .B1(n1230), .B2(n174), .C1(n1225), .C2(n323), .A(n2327), 
        .ZN(n2328) );
  NOR4_X1 U1843 ( .A1(n2331), .A2(n2328), .A3(n2330), .A4(n2329), .ZN(n2333)
         );
  OAI222_X1 U1844 ( .A1(n833), .A2(n1237), .B1(n2333), .B2(n1234), .C1(n1231), 
        .C2(n2332), .ZN(n2334) );
  OAI22_X1 U1845 ( .A1(n509), .A2(n2336), .B1(n961), .B2(n1247), .ZN(n2337) );
  OAI22_X1 U1846 ( .A1(n4695), .A2(n1277), .B1(n1384), .B2(n1271), .ZN(n2341)
         );
  AOI221_X1 U1847 ( .B1(n4951), .B2(n1281), .C1(n1278), .C2(n2342), .A(n2341), 
        .ZN(n2343) );
  AOI22_X1 U1848 ( .A1(n697), .A2(n198), .B1(n9), .B2(n4155), .ZN(n2347) );
  OAI221_X1 U1849 ( .B1(n1207), .B2(n295), .C1(n256), .C2(n1202), .A(n2347), 
        .ZN(n2356) );
  AOI22_X1 U1850 ( .A1(n998), .A2(n4219), .B1(n879), .B2(n4187), .ZN(n2348) );
  OAI221_X1 U1851 ( .B1(n384), .B2(n1215), .C1(n416), .C2(n8), .A(n2348), .ZN(
        n2355) );
  AOI22_X1 U1852 ( .A1(n5112), .A2(n987), .B1(n5144), .B2(n1216), .ZN(n2349)
         );
  OAI221_X1 U1853 ( .B1(n1224), .B2(n2351), .C1(n1219), .C2(n2350), .A(n2349), 
        .ZN(n2354) );
  AOI22_X1 U1854 ( .A1(n5176), .A2(n1), .B1(n5208), .B2(n750), .ZN(n2352) );
  NOR4_X1 U1855 ( .A1(n2356), .A2(n2355), .A3(n2354), .A4(n2353), .ZN(n2358)
         );
  OAI222_X1 U1856 ( .A1(n832), .A2(n1237), .B1(n2358), .B2(n1234), .C1(n1231), 
        .C2(n2357), .ZN(n2359) );
  OAI22_X1 U1857 ( .A1(n509), .A2(n2361), .B1(n960), .B2(n1246), .ZN(n2362) );
  AOI221_X1 U1858 ( .B1(n4792), .B2(n1254), .C1(n1250), .C2(n4335), .A(n2362), 
        .ZN(n2370) );
  OAI222_X1 U1859 ( .A1(n640), .A2(n1262), .B1(n1259), .B2(n2364), .C1(n590), 
        .C2(n2363), .ZN(n2365) );
  AOI221_X1 U1860 ( .B1(n1268), .B2(n4283), .C1(n1265), .C2(n4251), .A(n2365), 
        .ZN(n2369) );
  OAI22_X1 U1861 ( .A1(n4696), .A2(n1277), .B1(n1386), .B2(n1271), .ZN(n2366)
         );
  AOI221_X1 U1862 ( .B1(n4952), .B2(n1281), .C1(n1278), .C2(n2367), .A(n2366), 
        .ZN(n2368) );
  NAND4_X1 U1863 ( .A1(n2371), .A2(n2370), .A3(n2369), .A4(n2368), .ZN(n2542)
         );
  AOI22_X1 U1864 ( .A1(n1200), .A2(n199), .B1(n495), .B2(n4154), .ZN(n2372) );
  OAI221_X1 U1865 ( .B1(n1207), .B2(n296), .C1(n255), .C2(n1202), .A(n2372), 
        .ZN(n2381) );
  AOI22_X1 U1866 ( .A1(n998), .A2(n4218), .B1(n879), .B2(n4186), .ZN(n2373) );
  OAI221_X1 U1867 ( .B1(n383), .B2(n6), .C1(n415), .C2(n1212), .A(n2373), .ZN(
        n2380) );
  AOI22_X1 U1868 ( .A1(n5113), .A2(n704), .B1(n5145), .B2(n1216), .ZN(n2374)
         );
  OAI221_X1 U1869 ( .B1(n1223), .B2(n2376), .C1(n1219), .C2(n2375), .A(n2374), 
        .ZN(n2379) );
  AOI22_X1 U1870 ( .A1(n5177), .A2(n2), .B1(n5209), .B2(n750), .ZN(n2377) );
  NOR4_X1 U1871 ( .A1(n2381), .A2(n2380), .A3(n2379), .A4(n2378), .ZN(n2383)
         );
  OAI22_X1 U1872 ( .A1(n498), .A2(n2386), .B1(n959), .B2(n1245), .ZN(n2387) );
  AOI221_X1 U1873 ( .B1(n4793), .B2(n1253), .C1(n1250), .C2(n4334), .A(n2387), 
        .ZN(n2395) );
  OAI222_X1 U1874 ( .A1(n639), .A2(n1262), .B1(n1260), .B2(n2389), .C1(n590), 
        .C2(n2388), .ZN(n2390) );
  OAI22_X1 U1875 ( .A1(n4697), .A2(n1277), .B1(n1388), .B2(n1271), .ZN(n2391)
         );
  AOI221_X1 U1876 ( .B1(n4953), .B2(n1281), .C1(n1278), .C2(n2392), .A(n2391), 
        .ZN(n2393) );
  AOI22_X1 U1877 ( .A1(n1200), .A2(n200), .B1(n9), .B2(n4153), .ZN(n2397) );
  AOI22_X1 U1878 ( .A1(n998), .A2(n4217), .B1(n879), .B2(n4185), .ZN(n2398) );
  OAI221_X1 U1879 ( .B1(n382), .B2(n1213), .C1(n414), .C2(n8), .A(n2398), .ZN(
        n2405) );
  AOI22_X1 U1880 ( .A1(n5114), .A2(n704), .B1(n5146), .B2(n1216), .ZN(n2399)
         );
  OAI221_X1 U1881 ( .B1(n1223), .B2(n2401), .C1(n1219), .C2(n2400), .A(n2399), 
        .ZN(n2404) );
  AOI22_X1 U1882 ( .A1(n5178), .A2(n932), .B1(n5210), .B2(n931), .ZN(n2402) );
  NOR4_X1 U1883 ( .A1(n2406), .A2(n2405), .A3(n2403), .A4(n2404), .ZN(n2408)
         );
  OAI222_X1 U1884 ( .A1(n830), .A2(n1237), .B1(n2408), .B2(n1234), .C1(n1231), 
        .C2(n2407), .ZN(n2409) );
  OAI22_X1 U1885 ( .A1(n1248), .A2(n2411), .B1(n958), .B2(n480), .ZN(n2412) );
  AOI221_X1 U1886 ( .B1(n4794), .B2(n1255), .C1(n1250), .C2(n4333), .A(n2412), 
        .ZN(n2420) );
  OAI222_X1 U1887 ( .A1(n638), .A2(n1262), .B1(n1260), .B2(n2414), .C1(n590), 
        .C2(n2413), .ZN(n2415) );
  AOI221_X1 U1888 ( .B1(n1268), .B2(n4281), .C1(n1265), .C2(n4249), .A(n2415), 
        .ZN(n2419) );
  OAI22_X1 U1889 ( .A1(n4698), .A2(n1277), .B1(n1390), .B2(n1271), .ZN(n2416)
         );
  AOI221_X1 U1890 ( .B1(n4954), .B2(n1281), .C1(n1278), .C2(n2417), .A(n2416), 
        .ZN(n2418) );
  NAND4_X1 U1891 ( .A1(n2421), .A2(n2418), .A3(n2419), .A4(n2420), .ZN(n2544)
         );
  AOI22_X1 U1892 ( .A1(n66), .A2(n201), .B1(n496), .B2(n4152), .ZN(n2422) );
  OAI221_X1 U1893 ( .B1(n1206), .B2(n298), .C1(n253), .C2(n1202), .A(n2422), 
        .ZN(n2431) );
  AOI22_X1 U1894 ( .A1(n998), .A2(n4216), .B1(n879), .B2(n4184), .ZN(n2423) );
  OAI221_X1 U1895 ( .B1(n381), .B2(n1215), .C1(n413), .C2(n1212), .A(n2423), 
        .ZN(n2430) );
  AOI22_X1 U1896 ( .A1(n5115), .A2(n589), .B1(n5147), .B2(n1216), .ZN(n2424)
         );
  OAI221_X1 U1897 ( .B1(n1222), .B2(n2426), .C1(n1219), .C2(n2425), .A(n2424), 
        .ZN(n2429) );
  AOI22_X1 U1898 ( .A1(n5179), .A2(n932), .B1(n5211), .B2(n931), .ZN(n2427) );
  OAI221_X1 U1899 ( .B1(n1230), .B2(n177), .C1(n1225), .C2(n326), .A(n2427), 
        .ZN(n2428) );
  NOR4_X1 U1900 ( .A1(n2431), .A2(n2430), .A3(n2428), .A4(n2429), .ZN(n2433)
         );
  OAI222_X1 U1901 ( .A1(n829), .A2(n1237), .B1(n2433), .B2(n1234), .C1(n1231), 
        .C2(n2432), .ZN(n2434) );
  OAI22_X1 U1902 ( .A1(n498), .A2(n2436), .B1(n957), .B2(n1245), .ZN(n2437) );
  AOI221_X1 U1903 ( .B1(n4795), .B2(n1253), .C1(n1250), .C2(n4332), .A(n2437), 
        .ZN(n2445) );
  OAI222_X1 U1904 ( .A1(n637), .A2(n1262), .B1(n1259), .B2(n2439), .C1(n1258), 
        .C2(n2438), .ZN(n2440) );
  OAI22_X1 U1905 ( .A1(n4699), .A2(n1277), .B1(n1392), .B2(n1271), .ZN(n2441)
         );
  AOI221_X1 U1906 ( .B1(n4955), .B2(n1281), .C1(n1278), .C2(n2442), .A(n2441), 
        .ZN(n2443) );
  AOI22_X1 U1907 ( .A1(n1201), .A2(n202), .B1(n496), .B2(n4151), .ZN(n2447) );
  OAI221_X1 U1908 ( .B1(n1207), .B2(n299), .C1(n252), .C2(n1202), .A(n2447), 
        .ZN(n2456) );
  AOI22_X1 U1909 ( .A1(n998), .A2(n4215), .B1(n879), .B2(n4183), .ZN(n2448) );
  OAI221_X1 U1910 ( .B1(n380), .B2(n1213), .C1(n412), .C2(n1210), .A(n2448), 
        .ZN(n2455) );
  AOI22_X1 U1911 ( .A1(n5116), .A2(n987), .B1(n5148), .B2(n1216), .ZN(n2449)
         );
  OAI221_X1 U1912 ( .B1(n1223), .B2(n2451), .C1(n1219), .C2(n2450), .A(n2449), 
        .ZN(n2454) );
  AOI22_X1 U1913 ( .A1(n5180), .A2(n932), .B1(n5212), .B2(n750), .ZN(n2452) );
  NOR4_X1 U1914 ( .A1(n2456), .A2(n2455), .A3(n2453), .A4(n2454), .ZN(n2458)
         );
  OAI22_X1 U1915 ( .A1(n498), .A2(n2461), .B1(n956), .B2(n1245), .ZN(n2462) );
  AOI221_X1 U1916 ( .B1(n4796), .B2(n1253), .C1(n1250), .C2(n4331), .A(n2462), 
        .ZN(n2470) );
  OAI222_X1 U1917 ( .A1(n636), .A2(n1262), .B1(n1259), .B2(n2464), .C1(n1258), 
        .C2(n2463), .ZN(n2465) );
  OAI22_X1 U1918 ( .A1(n4700), .A2(n1277), .B1(n1394), .B2(n1271), .ZN(n2466)
         );
  AOI221_X1 U1919 ( .B1(n4956), .B2(n1281), .C1(n1278), .C2(n2467), .A(n2466), 
        .ZN(n2468) );
  AOI22_X1 U1920 ( .A1(n66), .A2(n213), .B1(n9), .B2(n4150), .ZN(n2472) );
  OAI221_X1 U1921 ( .B1(n1206), .B2(n300), .C1(n251), .C2(n1202), .A(n2472), 
        .ZN(n2481) );
  AOI22_X1 U1922 ( .A1(n689), .A2(n4214), .B1(n879), .B2(n4182), .ZN(n2473) );
  OAI221_X1 U1923 ( .B1(n379), .B2(n6), .C1(n411), .C2(n8), .A(n2473), .ZN(
        n2480) );
  AOI22_X1 U1924 ( .A1(n5117), .A2(n589), .B1(n5149), .B2(n1216), .ZN(n2474)
         );
  OAI221_X1 U1925 ( .B1(n1222), .B2(n2476), .C1(n1219), .C2(n2475), .A(n2474), 
        .ZN(n2479) );
  AOI22_X1 U1926 ( .A1(n5181), .A2(n932), .B1(n5213), .B2(n40), .ZN(n2477) );
  OAI221_X1 U1927 ( .B1(n1228), .B2(n179), .C1(n1225), .C2(n328), .A(n2477), 
        .ZN(n2478) );
  NOR4_X1 U1928 ( .A1(n2481), .A2(n2478), .A3(n2479), .A4(n2480), .ZN(n2483)
         );
  OAI222_X1 U1929 ( .A1(n827), .A2(n1237), .B1(n2483), .B2(n1234), .C1(n1231), 
        .C2(n2482), .ZN(n2484) );
  OAI22_X1 U1930 ( .A1(n498), .A2(n2486), .B1(n955), .B2(n1245), .ZN(n2487) );
  OAI22_X1 U1931 ( .A1(n4701), .A2(n1277), .B1(n1396), .B2(n1271), .ZN(n2491)
         );
  AOI221_X1 U1932 ( .B1(n4957), .B2(n1281), .C1(n1278), .C2(n2492), .A(n2491), 
        .ZN(n2493) );
  AOI22_X1 U1933 ( .A1(n1200), .A2(n203), .B1(n1198), .B2(n4149), .ZN(n2497)
         );
  OAI221_X1 U1934 ( .B1(n1206), .B2(n301), .C1(n250), .C2(n1202), .A(n2497), 
        .ZN(n3562) );
  AOI22_X1 U1935 ( .A1(n689), .A2(n4213), .B1(n879), .B2(n4181), .ZN(n2498) );
  OAI221_X1 U1936 ( .B1(n378), .B2(n1213), .C1(n410), .C2(n1210), .A(n2498), 
        .ZN(n2505) );
  AOI22_X1 U1937 ( .A1(n5118), .A2(n589), .B1(n5150), .B2(n1216), .ZN(n2499)
         );
  OAI221_X1 U1938 ( .B1(n1223), .B2(n2501), .C1(n1219), .C2(n2500), .A(n2499), 
        .ZN(n2504) );
  AOI22_X1 U1939 ( .A1(n5182), .A2(n2), .B1(n5214), .B2(n750), .ZN(n2502) );
  OAI221_X1 U1940 ( .B1(n1228), .B2(n180), .C1(n1225), .C2(n329), .A(n2502), 
        .ZN(n2503) );
  NOR4_X1 U1941 ( .A1(n3562), .A2(n2503), .A3(n2505), .A4(n2504), .ZN(n3564)
         );
  OAI222_X1 U1942 ( .A1(n826), .A2(n1237), .B1(n3564), .B2(n1234), .C1(n1231), 
        .C2(n3563), .ZN(n3565) );
  OAI22_X1 U1943 ( .A1(n498), .A2(n3567), .B1(n954), .B2(n1245), .ZN(n3568) );
  AOI221_X1 U1944 ( .B1(n4798), .B2(n1253), .C1(n1250), .C2(n4329), .A(n3568), 
        .ZN(n3576) );
  OAI22_X1 U1945 ( .A1(n4702), .A2(n1277), .B1(n1398), .B2(n1271), .ZN(n3572)
         );
  AOI221_X1 U1946 ( .B1(n4958), .B2(n1281), .C1(n1278), .C2(n3573), .A(n3572), 
        .ZN(n3574) );
  AOI22_X1 U1947 ( .A1(n697), .A2(n214), .B1(n688), .B2(n4148), .ZN(n3578) );
  OAI221_X1 U1948 ( .B1(n1206), .B2(n302), .C1(n249), .C2(n1202), .A(n3578), 
        .ZN(n3587) );
  AOI22_X1 U1949 ( .A1(n689), .A2(n4212), .B1(n879), .B2(n4180), .ZN(n3579) );
  OAI221_X1 U1950 ( .B1(n377), .B2(n1213), .C1(n409), .C2(n1210), .A(n3579), 
        .ZN(n3586) );
  AOI22_X1 U1951 ( .A1(n987), .A2(n5119), .B1(n5151), .B2(n1216), .ZN(n3580)
         );
  OAI221_X1 U1952 ( .B1(n1223), .B2(n3582), .C1(n1219), .C2(n3581), .A(n3580), 
        .ZN(n3585) );
  AOI22_X1 U1953 ( .A1(n5183), .A2(n1), .B1(n5215), .B2(n750), .ZN(n3583) );
  NOR4_X1 U1954 ( .A1(n3587), .A2(n3586), .A3(n3585), .A4(n3584), .ZN(n3589)
         );
  OAI222_X1 U1955 ( .A1(n825), .A2(n1237), .B1(n3589), .B2(n1234), .C1(n1231), 
        .C2(n3588), .ZN(n3590) );
  OAI22_X1 U1956 ( .A1(n509), .A2(n3592), .B1(n953), .B2(n480), .ZN(n3593) );
  AOI221_X1 U1957 ( .B1(n4799), .B2(n33), .C1(n1250), .C2(n4328), .A(n3593), 
        .ZN(n3601) );
  OAI222_X1 U1958 ( .A1(n633), .A2(n1262), .B1(n1260), .B2(n3595), .C1(n1258), 
        .C2(n3594), .ZN(n3596) );
  AOI221_X1 U1959 ( .B1(n1268), .B2(n4276), .C1(n1265), .C2(n4244), .A(n3596), 
        .ZN(n3600) );
  OAI22_X1 U1960 ( .A1(n4703), .A2(n1277), .B1(n1400), .B2(n1271), .ZN(n3597)
         );
  AOI221_X1 U1961 ( .B1(n4959), .B2(n1281), .C1(n1278), .C2(n3598), .A(n3597), 
        .ZN(n3599) );
  NAND4_X1 U1962 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n2549)
         );
  AOI22_X1 U1963 ( .A1(n1199), .A2(n215), .B1(n1197), .B2(n4147), .ZN(n3603)
         );
  AOI22_X1 U1964 ( .A1(n87), .A2(n4211), .B1(n892), .B2(n4179), .ZN(n3604) );
  AOI22_X1 U1965 ( .A1(n5120), .A2(n589), .B1(n5152), .B2(n1217), .ZN(n3605)
         );
  OAI221_X1 U1966 ( .B1(n1224), .B2(n3607), .C1(n1220), .C2(n3606), .A(n3605), 
        .ZN(n3610) );
  AOI22_X1 U1967 ( .A1(n2), .A2(n5184), .B1(n5216), .B2(n931), .ZN(n3608) );
  OAI221_X1 U1968 ( .B1(n1230), .B2(n181), .C1(n1226), .C2(n330), .A(n3608), 
        .ZN(n3609) );
  NOR4_X1 U1969 ( .A1(n3611), .A2(n3612), .A3(n3609), .A4(n3610), .ZN(n3614)
         );
  OAI222_X1 U1970 ( .A1(n824), .A2(n1238), .B1(n3614), .B2(n1235), .C1(n1232), 
        .C2(n3613), .ZN(n3615) );
  OAI22_X1 U1971 ( .A1(n1249), .A2(n3617), .B1(n952), .B2(n1246), .ZN(n3618)
         );
  AOI221_X1 U1972 ( .B1(n4800), .B2(n1255), .C1(n1251), .C2(n4327), .A(n3618), 
        .ZN(n3626) );
  OAI222_X1 U1973 ( .A1(n632), .A2(n1263), .B1(n1259), .B2(n3620), .C1(n590), 
        .C2(n3619), .ZN(n3621) );
  AOI221_X1 U1974 ( .B1(n1269), .B2(n4275), .C1(n1266), .C2(n4243), .A(n3621), 
        .ZN(n3625) );
  OAI22_X1 U1975 ( .A1(n4704), .A2(n1277), .B1(n1402), .B2(n1272), .ZN(n3622)
         );
  AOI221_X1 U1976 ( .B1(n4960), .B2(n1282), .C1(n1279), .C2(n3623), .A(n3622), 
        .ZN(n3624) );
  NAND4_X1 U1977 ( .A1(n3627), .A2(n3626), .A3(n3625), .A4(n3624), .ZN(n2550)
         );
  AOI22_X1 U1978 ( .A1(n697), .A2(n216), .B1(n688), .B2(n4146), .ZN(n3628) );
  AOI22_X1 U1979 ( .A1(n998), .A2(n4210), .B1(n1208), .B2(n4178), .ZN(n3629)
         );
  OAI221_X1 U1980 ( .B1(n375), .B2(n1215), .C1(n407), .C2(n1210), .A(n3629), 
        .ZN(n3636) );
  AOI22_X1 U1981 ( .A1(n5121), .A2(n704), .B1(n5153), .B2(n1217), .ZN(n3630)
         );
  OAI221_X1 U1982 ( .B1(n1222), .B2(n3632), .C1(n1220), .C2(n3631), .A(n3630), 
        .ZN(n3635) );
  AOI22_X1 U1983 ( .A1(n5185), .A2(n1), .B1(n5217), .B2(n750), .ZN(n3633) );
  NOR4_X1 U1984 ( .A1(n3637), .A2(n3636), .A3(n3634), .A4(n3635), .ZN(n3639)
         );
  OAI222_X1 U1985 ( .A1(n823), .A2(n1238), .B1(n3639), .B2(n1235), .C1(n1232), 
        .C2(n3638), .ZN(n3640) );
  OAI22_X1 U1986 ( .A1(n1248), .A2(n3642), .B1(n951), .B2(n480), .ZN(n3643) );
  AOI221_X1 U1987 ( .B1(n4801), .B2(n33), .C1(n1251), .C2(n4326), .A(n3643), 
        .ZN(n3651) );
  OAI222_X1 U1988 ( .A1(n631), .A2(n1263), .B1(n1259), .B2(n3645), .C1(n590), 
        .C2(n3644), .ZN(n3646) );
  AOI221_X1 U1989 ( .B1(n1269), .B2(n4274), .C1(n1266), .C2(n4242), .A(n3646), 
        .ZN(n3650) );
  OAI22_X1 U1990 ( .A1(n4705), .A2(n1277), .B1(n1404), .B2(n1272), .ZN(n3647)
         );
  AOI221_X1 U1991 ( .B1(n4961), .B2(n1282), .C1(n1279), .C2(n3648), .A(n3647), 
        .ZN(n3649) );
  NAND4_X1 U1992 ( .A1(n3652), .A2(n3649), .A3(n3650), .A4(n3651), .ZN(n2551)
         );
  AOI22_X1 U1993 ( .A1(n697), .A2(n217), .B1(n496), .B2(n4145), .ZN(n3653) );
  OAI221_X1 U1994 ( .B1(n1206), .B2(n304), .C1(n246), .C2(n1203), .A(n3653), 
        .ZN(n3662) );
  AOI22_X1 U1995 ( .A1(n689), .A2(n4209), .B1(n1209), .B2(n4177), .ZN(n3654)
         );
  OAI221_X1 U1996 ( .B1(n374), .B2(n6), .C1(n406), .C2(n8), .A(n3654), .ZN(
        n3661) );
  AOI22_X1 U1997 ( .A1(n5122), .A2(n987), .B1(n5154), .B2(n1217), .ZN(n3655)
         );
  OAI221_X1 U1998 ( .B1(n1223), .B2(n3657), .C1(n1220), .C2(n3656), .A(n3655), 
        .ZN(n3660) );
  AOI22_X1 U1999 ( .A1(n5186), .A2(n932), .B1(n5218), .B2(n40), .ZN(n3658) );
  NOR4_X1 U2000 ( .A1(n3662), .A2(n3661), .A3(n3659), .A4(n3660), .ZN(n3664)
         );
  OAI222_X1 U2001 ( .A1(n822), .A2(n1238), .B1(n3664), .B2(n1235), .C1(n1232), 
        .C2(n3663), .ZN(n3665) );
  OAI22_X1 U2002 ( .A1(n509), .A2(n3667), .B1(n950), .B2(n1247), .ZN(n3668) );
  AOI221_X1 U2003 ( .B1(n4802), .B2(n1254), .C1(n1251), .C2(n4325), .A(n3668), 
        .ZN(n3676) );
  OAI222_X1 U2004 ( .A1(n630), .A2(n1263), .B1(n1260), .B2(n3670), .C1(n1258), 
        .C2(n3669), .ZN(n3671) );
  AOI221_X1 U2005 ( .B1(n1269), .B2(n4273), .C1(n1266), .C2(n4241), .A(n3671), 
        .ZN(n3675) );
  OAI22_X1 U2006 ( .A1(n4706), .A2(n1276), .B1(n1406), .B2(n1272), .ZN(n3672)
         );
  AOI221_X1 U2007 ( .B1(n4962), .B2(n1282), .C1(n1279), .C2(n3673), .A(n3672), 
        .ZN(n3674) );
  NAND4_X1 U2008 ( .A1(n3677), .A2(n3676), .A3(n3675), .A4(n3674), .ZN(n2552)
         );
  AOI22_X1 U2009 ( .A1(n1199), .A2(n204), .B1(n1198), .B2(n4144), .ZN(n3678)
         );
  OAI221_X1 U2010 ( .B1(n1207), .B2(n305), .C1(n245), .C2(n1203), .A(n3678), 
        .ZN(n3687) );
  AOI22_X1 U2011 ( .A1(n998), .A2(n4208), .B1(n1208), .B2(n4176), .ZN(n3679)
         );
  AOI22_X1 U2012 ( .A1(n5123), .A2(n704), .B1(n5155), .B2(n1217), .ZN(n3680)
         );
  OAI221_X1 U2013 ( .B1(n1224), .B2(n3682), .C1(n1220), .C2(n3681), .A(n3680), 
        .ZN(n3685) );
  AOI22_X1 U2014 ( .A1(n5187), .A2(n710), .B1(n5219), .B2(n40), .ZN(n3683) );
  OAI221_X1 U2015 ( .B1(n1229), .B2(n183), .C1(n1226), .C2(n332), .A(n3683), 
        .ZN(n3684) );
  NOR4_X1 U2016 ( .A1(n3687), .A2(n3685), .A3(n3686), .A4(n3684), .ZN(n3689)
         );
  OAI22_X1 U2017 ( .A1(n1249), .A2(n3692), .B1(n949), .B2(n1246), .ZN(n3693)
         );
  AOI221_X1 U2018 ( .B1(n4803), .B2(n1255), .C1(n1251), .C2(n4324), .A(n3693), 
        .ZN(n3701) );
  OAI222_X1 U2019 ( .A1(n629), .A2(n1263), .B1(n1260), .B2(n3695), .C1(n1258), 
        .C2(n3694), .ZN(n3696) );
  AOI221_X1 U2020 ( .B1(n1269), .B2(n4272), .C1(n1266), .C2(n4240), .A(n3696), 
        .ZN(n3700) );
  OAI22_X1 U2021 ( .A1(n4707), .A2(n1276), .B1(n1408), .B2(n1272), .ZN(n3697)
         );
  AOI221_X1 U2022 ( .B1(n4963), .B2(n1282), .C1(n1279), .C2(n3698), .A(n3697), 
        .ZN(n3699) );
  NAND4_X1 U2023 ( .A1(n3702), .A2(n3699), .A3(n3700), .A4(n3701), .ZN(n2553)
         );
  AOI22_X1 U2024 ( .A1(n1200), .A2(n205), .B1(n495), .B2(n4143), .ZN(n3703) );
  OAI221_X1 U2025 ( .B1(n1207), .B2(n306), .C1(n244), .C2(n1203), .A(n3703), 
        .ZN(n3712) );
  AOI22_X1 U2026 ( .A1(n998), .A2(n4207), .B1(n1208), .B2(n4175), .ZN(n3704)
         );
  OAI221_X1 U2027 ( .B1(n372), .B2(n1213), .C1(n404), .C2(n8), .A(n3704), .ZN(
        n3711) );
  AOI22_X1 U2028 ( .A1(n5124), .A2(n704), .B1(n5156), .B2(n1217), .ZN(n3705)
         );
  OAI221_X1 U2029 ( .B1(n1224), .B2(n3707), .C1(n1220), .C2(n3706), .A(n3705), 
        .ZN(n3710) );
  AOI22_X1 U2030 ( .A1(n5188), .A2(n1), .B1(n5220), .B2(n931), .ZN(n3708) );
  NOR4_X1 U2031 ( .A1(n3712), .A2(n3711), .A3(n3710), .A4(n3709), .ZN(n3714)
         );
  OAI222_X1 U2032 ( .A1(n820), .A2(n1238), .B1(n3714), .B2(n1235), .C1(n1232), 
        .C2(n3713), .ZN(n3715) );
  OAI22_X1 U2033 ( .A1(n509), .A2(n3717), .B1(n948), .B2(n1247), .ZN(n3718) );
  AOI221_X1 U2034 ( .B1(n4804), .B2(n33), .C1(n1251), .C2(n4323), .A(n3718), 
        .ZN(n3726) );
  OAI222_X1 U2035 ( .A1(n628), .A2(n1263), .B1(n1259), .B2(n3720), .C1(n1256), 
        .C2(n3719), .ZN(n3721) );
  AOI221_X1 U2036 ( .B1(n1269), .B2(n4271), .C1(n1266), .C2(n4239), .A(n3721), 
        .ZN(n3725) );
  OAI22_X1 U2037 ( .A1(n4708), .A2(n1276), .B1(n1410), .B2(n1272), .ZN(n3722)
         );
  AOI221_X1 U2038 ( .B1(n4964), .B2(n1282), .C1(n1279), .C2(n3723), .A(n3722), 
        .ZN(n3724) );
  NAND4_X1 U2039 ( .A1(n3727), .A2(n3726), .A3(n3725), .A4(n3724), .ZN(n2554)
         );
  AOI22_X1 U2040 ( .A1(n697), .A2(n206), .B1(n495), .B2(n4142), .ZN(n3728) );
  OAI221_X1 U2041 ( .B1(n1206), .B2(n307), .C1(n243), .C2(n1203), .A(n3728), 
        .ZN(n3737) );
  AOI22_X1 U2042 ( .A1(n998), .A2(n4206), .B1(n1209), .B2(n4174), .ZN(n3729)
         );
  OAI221_X1 U2043 ( .B1(n371), .B2(n6), .C1(n403), .C2(n1210), .A(n3729), .ZN(
        n3736) );
  AOI22_X1 U2044 ( .A1(n5125), .A2(n987), .B1(n5157), .B2(n1217), .ZN(n3730)
         );
  OAI221_X1 U2045 ( .B1(n1222), .B2(n3732), .C1(n1220), .C2(n3731), .A(n3730), 
        .ZN(n3735) );
  AOI22_X1 U2046 ( .A1(n5189), .A2(n2), .B1(n5221), .B2(n40), .ZN(n3733) );
  NOR4_X1 U2047 ( .A1(n3737), .A2(n3736), .A3(n3735), .A4(n3734), .ZN(n3739)
         );
  OAI222_X1 U2048 ( .A1(n819), .A2(n1238), .B1(n3739), .B2(n1235), .C1(n1232), 
        .C2(n3738), .ZN(n3740) );
  OAI22_X1 U2049 ( .A1(n509), .A2(n3742), .B1(n947), .B2(n1246), .ZN(n3743) );
  AOI221_X1 U2050 ( .B1(n4805), .B2(n33), .C1(n1251), .C2(n4322), .A(n3743), 
        .ZN(n3751) );
  OAI222_X1 U2051 ( .A1(n627), .A2(n1263), .B1(n1260), .B2(n3745), .C1(n1258), 
        .C2(n3744), .ZN(n3746) );
  AOI221_X1 U2052 ( .B1(n1269), .B2(n4270), .C1(n1266), .C2(n4238), .A(n3746), 
        .ZN(n3750) );
  OAI22_X1 U2053 ( .A1(n4709), .A2(n1276), .B1(n1412), .B2(n1272), .ZN(n3747)
         );
  AOI221_X1 U2054 ( .B1(n4965), .B2(n1282), .C1(n1279), .C2(n3748), .A(n3747), 
        .ZN(n3749) );
  NAND4_X1 U2055 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(n2555)
         );
  AOI22_X1 U2056 ( .A1(n66), .A2(n207), .B1(n495), .B2(n4141), .ZN(n3753) );
  AOI22_X1 U2057 ( .A1(n998), .A2(n4205), .B1(n1208), .B2(n4173), .ZN(n3754)
         );
  OAI221_X1 U2058 ( .B1(n370), .B2(n6), .C1(n402), .C2(n1212), .A(n3754), .ZN(
        n3761) );
  AOI22_X1 U2059 ( .A1(n589), .A2(n5126), .B1(n5158), .B2(n1217), .ZN(n3755)
         );
  OAI221_X1 U2060 ( .B1(n1224), .B2(n3757), .C1(n1220), .C2(n3756), .A(n3755), 
        .ZN(n3760) );
  AOI22_X1 U2061 ( .A1(n5190), .A2(n932), .B1(n5222), .B2(n750), .ZN(n3758) );
  NOR4_X1 U2062 ( .A1(n3762), .A2(n3761), .A3(n3759), .A4(n3760), .ZN(n3764)
         );
  OAI222_X1 U2063 ( .A1(n818), .A2(n1238), .B1(n3764), .B2(n1235), .C1(n1232), 
        .C2(n3763), .ZN(n3765) );
  OAI22_X1 U2064 ( .A1(n1248), .A2(n3767), .B1(n946), .B2(n1246), .ZN(n3768)
         );
  AOI221_X1 U2065 ( .B1(n4806), .B2(n1254), .C1(n1251), .C2(n4321), .A(n3768), 
        .ZN(n3776) );
  OAI222_X1 U2066 ( .A1(n626), .A2(n1263), .B1(n1259), .B2(n3770), .C1(n1258), 
        .C2(n3769), .ZN(n3771) );
  AOI221_X1 U2067 ( .B1(n1269), .B2(n4269), .C1(n1266), .C2(n4237), .A(n3771), 
        .ZN(n3775) );
  OAI22_X1 U2068 ( .A1(n4710), .A2(n1276), .B1(n1414), .B2(n1272), .ZN(n3772)
         );
  AOI221_X1 U2069 ( .B1(n4966), .B2(n1282), .C1(n1279), .C2(n3773), .A(n3772), 
        .ZN(n3774) );
  NAND4_X1 U2070 ( .A1(n3777), .A2(n3774), .A3(n3775), .A4(n3776), .ZN(n2556)
         );
  AOI22_X1 U2071 ( .A1(n1201), .A2(n208), .B1(n688), .B2(n4140), .ZN(n3778) );
  OAI221_X1 U2072 ( .B1(n1206), .B2(n309), .C1(n241), .C2(n1203), .A(n3778), 
        .ZN(n3787) );
  AOI22_X1 U2073 ( .A1(n689), .A2(n4204), .B1(n1208), .B2(n4172), .ZN(n3779)
         );
  OAI221_X1 U2074 ( .B1(n369), .B2(n1213), .C1(n401), .C2(n8), .A(n3779), .ZN(
        n3786) );
  AOI22_X1 U2075 ( .A1(n5127), .A2(n987), .B1(n5159), .B2(n1217), .ZN(n3780)
         );
  OAI221_X1 U2076 ( .B1(n1223), .B2(n3782), .C1(n1220), .C2(n3781), .A(n3780), 
        .ZN(n3785) );
  AOI22_X1 U2077 ( .A1(n5191), .A2(n2), .B1(n5223), .B2(n750), .ZN(n3783) );
  NOR4_X1 U2078 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3789)
         );
  OAI222_X1 U2079 ( .A1(n817), .A2(n1238), .B1(n3789), .B2(n1235), .C1(n1232), 
        .C2(n3788), .ZN(n3790) );
  OAI22_X1 U2080 ( .A1(n509), .A2(n3792), .B1(n945), .B2(n480), .ZN(n3793) );
  AOI221_X1 U2081 ( .B1(n4807), .B2(n1255), .C1(n1251), .C2(n4320), .A(n3793), 
        .ZN(n3801) );
  OAI222_X1 U2082 ( .A1(n625), .A2(n1263), .B1(n1259), .B2(n3795), .C1(n590), 
        .C2(n3794), .ZN(n3796) );
  AOI221_X1 U2083 ( .B1(n1269), .B2(n4268), .C1(n1266), .C2(n4236), .A(n3796), 
        .ZN(n3800) );
  OAI22_X1 U2084 ( .A1(n4711), .A2(n1276), .B1(n1416), .B2(n1272), .ZN(n3797)
         );
  AOI221_X1 U2085 ( .B1(n4967), .B2(n1282), .C1(n1279), .C2(n3798), .A(n3797), 
        .ZN(n3799) );
  NAND4_X1 U2086 ( .A1(n3802), .A2(n3801), .A3(n3800), .A4(n3799), .ZN(n2557)
         );
  AOI22_X1 U2087 ( .A1(n1200), .A2(n209), .B1(n1196), .B2(n4139), .ZN(n3803)
         );
  OAI221_X1 U2088 ( .B1(n1206), .B2(n310), .C1(n240), .C2(n1203), .A(n3803), 
        .ZN(n3812) );
  AOI22_X1 U2089 ( .A1(n689), .A2(n4203), .B1(n1209), .B2(n4171), .ZN(n3804)
         );
  OAI221_X1 U2090 ( .B1(n368), .B2(n1215), .C1(n400), .C2(n1212), .A(n3804), 
        .ZN(n3811) );
  AOI22_X1 U2091 ( .A1(n5128), .A2(n589), .B1(n5160), .B2(n1217), .ZN(n3805)
         );
  OAI221_X1 U2092 ( .B1(n1224), .B2(n3807), .C1(n1220), .C2(n3806), .A(n3805), 
        .ZN(n3810) );
  AOI22_X1 U2093 ( .A1(n5192), .A2(n1), .B1(n5224), .B2(n750), .ZN(n3808) );
  NOR4_X1 U2094 ( .A1(n3812), .A2(n3811), .A3(n3810), .A4(n3809), .ZN(n3814)
         );
  OAI222_X1 U2095 ( .A1(n816), .A2(n1238), .B1(n3814), .B2(n1235), .C1(n1232), 
        .C2(n3813), .ZN(n3815) );
  OAI22_X1 U2096 ( .A1(n1249), .A2(n3817), .B1(n944), .B2(n480), .ZN(n3818) );
  AOI221_X1 U2097 ( .B1(n4808), .B2(n33), .C1(n1251), .C2(n4319), .A(n3818), 
        .ZN(n3826) );
  OAI222_X1 U2098 ( .A1(n624), .A2(n1263), .B1(n1259), .B2(n3820), .C1(n590), 
        .C2(n3819), .ZN(n3821) );
  AOI221_X1 U2099 ( .B1(n1269), .B2(n4267), .C1(n1266), .C2(n4235), .A(n3821), 
        .ZN(n3825) );
  OAI22_X1 U2100 ( .A1(n4712), .A2(n1276), .B1(n1418), .B2(n1272), .ZN(n3822)
         );
  AOI221_X1 U2101 ( .B1(n4968), .B2(n1282), .C1(n1279), .C2(n3823), .A(n3822), 
        .ZN(n3824) );
  NAND4_X1 U2102 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n2558)
         );
  AOI22_X1 U2103 ( .A1(n66), .A2(n210), .B1(n688), .B2(n4138), .ZN(n3828) );
  OAI221_X1 U2104 ( .B1(n1207), .B2(n311), .C1(n239), .C2(n1203), .A(n3828), 
        .ZN(n3837) );
  AOI22_X1 U2105 ( .A1(n998), .A2(n4202), .B1(n1208), .B2(n4170), .ZN(n3829)
         );
  OAI221_X1 U2106 ( .B1(n367), .B2(n6), .C1(n399), .C2(n1210), .A(n3829), .ZN(
        n3836) );
  AOI22_X1 U2107 ( .A1(n5129), .A2(n589), .B1(n5161), .B2(n1217), .ZN(n3830)
         );
  OAI221_X1 U2108 ( .B1(n1222), .B2(n3832), .C1(n1220), .C2(n3831), .A(n3830), 
        .ZN(n3835) );
  AOI22_X1 U2109 ( .A1(n5193), .A2(n932), .B1(n5225), .B2(n40), .ZN(n3833) );
  NOR4_X1 U2110 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n3839)
         );
  OAI222_X1 U2111 ( .A1(n815), .A2(n1238), .B1(n3839), .B2(n1235), .C1(n1232), 
        .C2(n3838), .ZN(n3840) );
  OAI22_X1 U2112 ( .A1(n1248), .A2(n3842), .B1(n943), .B2(n480), .ZN(n3843) );
  AOI221_X1 U2113 ( .B1(n4809), .B2(n33), .C1(n1251), .C2(n4318), .A(n3843), 
        .ZN(n3851) );
  OAI222_X1 U2114 ( .A1(n623), .A2(n1263), .B1(n1260), .B2(n3845), .C1(n1258), 
        .C2(n3844), .ZN(n3846) );
  AOI221_X1 U2115 ( .B1(n1269), .B2(n4266), .C1(n1266), .C2(n4234), .A(n3846), 
        .ZN(n3850) );
  OAI22_X1 U2116 ( .A1(n4713), .A2(n1276), .B1(n1420), .B2(n1272), .ZN(n3847)
         );
  AOI221_X1 U2117 ( .B1(n4969), .B2(n1282), .C1(n1279), .C2(n3848), .A(n3847), 
        .ZN(n3849) );
  NAND4_X1 U2118 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n2559)
         );
  AOI22_X1 U2119 ( .A1(n66), .A2(n211), .B1(n496), .B2(n4137), .ZN(n3853) );
  OAI221_X1 U2120 ( .B1(n1207), .B2(n312), .C1(n238), .C2(n1203), .A(n3853), 
        .ZN(n3862) );
  AOI22_X1 U2121 ( .A1(n998), .A2(n4201), .B1(n1209), .B2(n4169), .ZN(n3854)
         );
  OAI221_X1 U2122 ( .B1(n366), .B2(n1215), .C1(n398), .C2(n8), .A(n3854), .ZN(
        n3861) );
  AOI22_X1 U2123 ( .A1(n5130), .A2(n704), .B1(n5162), .B2(n1217), .ZN(n3855)
         );
  OAI221_X1 U2124 ( .B1(n1223), .B2(n3857), .C1(n1220), .C2(n3856), .A(n3855), 
        .ZN(n3860) );
  AOI22_X1 U2125 ( .A1(n5194), .A2(n932), .B1(n5226), .B2(n931), .ZN(n3858) );
  NOR4_X1 U2126 ( .A1(n3862), .A2(n3861), .A3(n3860), .A4(n3859), .ZN(n3864)
         );
  OAI222_X1 U2127 ( .A1(n814), .A2(n1238), .B1(n3864), .B2(n1235), .C1(n1232), 
        .C2(n3863), .ZN(n3865) );
  OAI22_X1 U2128 ( .A1(n509), .A2(n3867), .B1(n942), .B2(n1246), .ZN(n3868) );
  AOI221_X1 U2129 ( .B1(n4810), .B2(n33), .C1(n1251), .C2(n4317), .A(n3868), 
        .ZN(n3876) );
  OAI222_X1 U2130 ( .A1(n622), .A2(n1263), .B1(n1260), .B2(n3870), .C1(n1258), 
        .C2(n3869), .ZN(n3871) );
  AOI221_X1 U2131 ( .B1(n1269), .B2(n4265), .C1(n1266), .C2(n4233), .A(n3871), 
        .ZN(n3875) );
  OAI22_X1 U2132 ( .A1(n4714), .A2(n1276), .B1(n1422), .B2(n1272), .ZN(n3872)
         );
  AOI221_X1 U2133 ( .B1(n4970), .B2(n1282), .C1(n1279), .C2(n3873), .A(n3872), 
        .ZN(n3874) );
  NAND4_X1 U2134 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n3874), .ZN(n2560)
         );
  AOI22_X1 U2135 ( .A1(n697), .A2(n212), .B1(n496), .B2(n4136), .ZN(n3878) );
  AOI22_X1 U2136 ( .A1(n998), .A2(n4200), .B1(n1209), .B2(n4168), .ZN(n3879)
         );
  OAI221_X1 U2137 ( .B1(n365), .B2(n1213), .C1(n397), .C2(n1210), .A(n3879), 
        .ZN(n3886) );
  AOI22_X1 U2138 ( .A1(n5131), .A2(n589), .B1(n5163), .B2(n1217), .ZN(n3880)
         );
  OAI221_X1 U2139 ( .B1(n1222), .B2(n3882), .C1(n1220), .C2(n3881), .A(n3880), 
        .ZN(n3885) );
  AOI22_X1 U2140 ( .A1(n5195), .A2(n932), .B1(n5227), .B2(n40), .ZN(n3883) );
  NOR4_X1 U2141 ( .A1(n3887), .A2(n3886), .A3(n3884), .A4(n3885), .ZN(n3889)
         );
  OAI222_X1 U2142 ( .A1(n813), .A2(n1238), .B1(n3889), .B2(n1235), .C1(n1232), 
        .C2(n3888), .ZN(n3890) );
  OAI22_X1 U2143 ( .A1(n1248), .A2(n3892), .B1(n941), .B2(n1246), .ZN(n3893)
         );
  AOI221_X1 U2144 ( .B1(n4811), .B2(n33), .C1(n1251), .C2(n4316), .A(n3893), 
        .ZN(n3901) );
  OAI222_X1 U2145 ( .A1(n621), .A2(n1263), .B1(n1260), .B2(n3895), .C1(n1256), 
        .C2(n3894), .ZN(n3896) );
  AOI221_X1 U2146 ( .B1(n1269), .B2(n4264), .C1(n1266), .C2(n4232), .A(n3896), 
        .ZN(n3900) );
  OAI22_X1 U2147 ( .A1(n4715), .A2(n1276), .B1(n1424), .B2(n1272), .ZN(n3897)
         );
  AOI221_X1 U2148 ( .B1(n4971), .B2(n1282), .C1(n1279), .C2(n3898), .A(n3897), 
        .ZN(n3899) );
  NAND4_X1 U2149 ( .A1(n3902), .A2(n3899), .A3(n3900), .A4(n3901), .ZN(n2561)
         );
  AOI22_X1 U2150 ( .A1(n66), .A2(n3903), .B1(n9), .B2(n4135), .ZN(n3904) );
  OAI221_X1 U2151 ( .B1(n1207), .B2(n314), .C1(n236), .C2(n1204), .A(n3904), 
        .ZN(n3913) );
  AOI22_X1 U2152 ( .A1(n998), .A2(n4199), .B1(n1209), .B2(n4167), .ZN(n3905)
         );
  OAI221_X1 U2153 ( .B1(n364), .B2(n6), .C1(n396), .C2(n8), .A(n3905), .ZN(
        n3912) );
  AOI22_X1 U2154 ( .A1(n5132), .A2(n704), .B1(n5164), .B2(n1218), .ZN(n3906)
         );
  OAI221_X1 U2155 ( .B1(n1224), .B2(n3908), .C1(n1221), .C2(n3907), .A(n3906), 
        .ZN(n3911) );
  AOI22_X1 U2156 ( .A1(n5196), .A2(n2), .B1(n5228), .B2(n931), .ZN(n3909) );
  NOR4_X1 U2157 ( .A1(n3913), .A2(n3912), .A3(n3910), .A4(n3911), .ZN(n3915)
         );
  OAI22_X1 U2158 ( .A1(n509), .A2(n3918), .B1(n940), .B2(n1247), .ZN(n3919) );
  AOI221_X1 U2159 ( .B1(n4812), .B2(n1254), .C1(n1252), .C2(n4315), .A(n3919), 
        .ZN(n3927) );
  OAI22_X1 U2160 ( .A1(n4716), .A2(n1276), .B1(n1427), .B2(n1273), .ZN(n3923)
         );
  AOI221_X1 U2161 ( .B1(n4972), .B2(n1283), .C1(n1280), .C2(n3924), .A(n3923), 
        .ZN(n3925) );
  AOI22_X1 U2162 ( .A1(n1199), .A2(n3929), .B1(n1197), .B2(n4134), .ZN(n3930)
         );
  OAI221_X1 U2163 ( .B1(n1207), .B2(n315), .C1(n235), .C2(n1204), .A(n3930), 
        .ZN(n3939) );
  AOI22_X1 U2164 ( .A1(n998), .A2(n4198), .B1(n1209), .B2(n4166), .ZN(n3931)
         );
  OAI221_X1 U2165 ( .B1(n363), .B2(n6), .C1(n395), .C2(n1210), .A(n3931), .ZN(
        n3938) );
  AOI22_X1 U2166 ( .A1(n987), .A2(n5133), .B1(n5165), .B2(n1218), .ZN(n3932)
         );
  OAI221_X1 U2167 ( .B1(n1223), .B2(n3934), .C1(n1221), .C2(n3933), .A(n3932), 
        .ZN(n3937) );
  AOI22_X1 U2168 ( .A1(n5197), .A2(n1), .B1(n5229), .B2(n40), .ZN(n3935) );
  NOR4_X1 U2169 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3941)
         );
  OAI222_X1 U2170 ( .A1(n811), .A2(n1239), .B1(n3941), .B2(n1236), .C1(n1233), 
        .C2(n3940), .ZN(n3942) );
  OAI22_X1 U2171 ( .A1(n1249), .A2(n3944), .B1(n939), .B2(n1247), .ZN(n3945)
         );
  AOI221_X1 U2172 ( .B1(n4813), .B2(n1255), .C1(n1252), .C2(n4314), .A(n3945), 
        .ZN(n3953) );
  OAI22_X1 U2173 ( .A1(n4717), .A2(n1275), .B1(n1430), .B2(n1273), .ZN(n3949)
         );
  AOI221_X1 U2174 ( .B1(n4973), .B2(n1283), .C1(n1280), .C2(n3950), .A(n3949), 
        .ZN(n3951) );
  AOI22_X1 U2175 ( .A1(n697), .A2(n3955), .B1(n688), .B2(n4133), .ZN(n3956) );
  OAI221_X1 U2176 ( .B1(n1206), .B2(n316), .C1(n234), .C2(n1204), .A(n3956), 
        .ZN(n3965) );
  AOI22_X1 U2177 ( .A1(n689), .A2(n4197), .B1(n1208), .B2(n4165), .ZN(n3957)
         );
  OAI221_X1 U2178 ( .B1(n362), .B2(n1213), .C1(n394), .C2(n8), .A(n3957), .ZN(
        n3964) );
  AOI22_X1 U2179 ( .A1(n5134), .A2(n987), .B1(n5166), .B2(n1218), .ZN(n3958)
         );
  OAI221_X1 U2180 ( .B1(n1224), .B2(n3960), .C1(n1221), .C2(n3959), .A(n3958), 
        .ZN(n3963) );
  AOI22_X1 U2181 ( .A1(n5198), .A2(n2), .B1(n5230), .B2(n750), .ZN(n3961) );
  OAI221_X1 U2182 ( .B1(n1228), .B2(n188), .C1(n1227), .C2(n337), .A(n3961), 
        .ZN(n3962) );
  NOR4_X1 U2183 ( .A1(n3965), .A2(n3962), .A3(n3964), .A4(n3963), .ZN(n3967)
         );
  OAI22_X1 U2184 ( .A1(n1248), .A2(n3970), .B1(n938), .B2(n1246), .ZN(n3971)
         );
  AOI221_X1 U2185 ( .B1(n4814), .B2(n33), .C1(n1252), .C2(n4313), .A(n3971), 
        .ZN(n3979) );
  OAI22_X1 U2186 ( .A1(n4718), .A2(n1275), .B1(n1433), .B2(n1273), .ZN(n3975)
         );
  AOI221_X1 U2187 ( .B1(n4974), .B2(n1283), .C1(n1280), .C2(n3976), .A(n3975), 
        .ZN(n3977) );
  AOI22_X1 U2188 ( .A1(n1201), .A2(n3981), .B1(n9), .B2(n4132), .ZN(n3982) );
  OAI221_X1 U2189 ( .B1(n1207), .B2(n317), .C1(n233), .C2(n1204), .A(n3982), 
        .ZN(n3991) );
  AOI22_X1 U2190 ( .A1(n998), .A2(n4196), .B1(n1209), .B2(n4164), .ZN(n3983)
         );
  OAI221_X1 U2191 ( .B1(n361), .B2(n1213), .C1(n393), .C2(n1212), .A(n3983), 
        .ZN(n3990) );
  AOI22_X1 U2192 ( .A1(n5135), .A2(n987), .B1(n5167), .B2(n1218), .ZN(n3984)
         );
  AOI22_X1 U2193 ( .A1(n5199), .A2(n932), .B1(n5231), .B2(n40), .ZN(n3987) );
  OAI221_X1 U2194 ( .B1(n1229), .B2(n189), .C1(n1227), .C2(n338), .A(n3987), 
        .ZN(n3988) );
  NOR4_X1 U2195 ( .A1(n3991), .A2(n3990), .A3(n3988), .A4(n3989), .ZN(n3993)
         );
  OAI222_X1 U2196 ( .A1(n809), .A2(n1239), .B1(n3993), .B2(n1236), .C1(n1233), 
        .C2(n3992), .ZN(n3994) );
  OAI22_X1 U2197 ( .A1(n509), .A2(n3996), .B1(n937), .B2(n480), .ZN(n3997) );
  AOI221_X1 U2198 ( .B1(n4815), .B2(n1254), .C1(n1252), .C2(n4312), .A(n3997), 
        .ZN(n4005) );
  OAI22_X1 U2199 ( .A1(n4719), .A2(n1275), .B1(n1436), .B2(n1273), .ZN(n4001)
         );
  AOI221_X1 U2200 ( .B1(n4975), .B2(n1283), .C1(n1280), .C2(n4002), .A(n4001), 
        .ZN(n4003) );
  AOI22_X1 U2201 ( .A1(n1199), .A2(n4007), .B1(n1196), .B2(n4131), .ZN(n4008)
         );
  OAI221_X1 U2202 ( .B1(n1207), .B2(n318), .C1(n232), .C2(n1204), .A(n4008), 
        .ZN(n4017) );
  AOI22_X1 U2203 ( .A1(n998), .A2(n4195), .B1(n1208), .B2(n4163), .ZN(n4009)
         );
  OAI221_X1 U2204 ( .B1(n360), .B2(n1215), .C1(n392), .C2(n8), .A(n4009), .ZN(
        n4016) );
  AOI22_X1 U2205 ( .A1(n5136), .A2(n589), .B1(n5168), .B2(n1218), .ZN(n4010)
         );
  OAI221_X1 U2206 ( .B1(n1224), .B2(n4012), .C1(n1221), .C2(n4011), .A(n4010), 
        .ZN(n4015) );
  AOI22_X1 U2207 ( .A1(n5200), .A2(n710), .B1(n5232), .B2(n931), .ZN(n4013) );
  OAI221_X1 U2208 ( .B1(n1228), .B2(n190), .C1(n1227), .C2(n339), .A(n4013), 
        .ZN(n4014) );
  NOR4_X1 U2209 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4019)
         );
  OAI222_X1 U2210 ( .A1(n808), .A2(n1239), .B1(n4019), .B2(n1236), .C1(n1233), 
        .C2(n4018), .ZN(n4020) );
  OAI22_X1 U2211 ( .A1(n1248), .A2(n4022), .B1(n936), .B2(n1247), .ZN(n4023)
         );
  AOI221_X1 U2212 ( .B1(n4816), .B2(n1255), .C1(n1252), .C2(n4311), .A(n4023), 
        .ZN(n4031) );
  OAI22_X1 U2213 ( .A1(n4720), .A2(n1275), .B1(n1439), .B2(n1273), .ZN(n4027)
         );
  AOI221_X1 U2214 ( .B1(n4976), .B2(n1283), .C1(n1280), .C2(n4028), .A(n4027), 
        .ZN(n4029) );
  AOI22_X1 U2215 ( .A1(n1201), .A2(n4033), .B1(n1196), .B2(n4130), .ZN(n4034)
         );
  AOI22_X1 U2216 ( .A1(n689), .A2(n4194), .B1(n1208), .B2(n4162), .ZN(n4035)
         );
  OAI221_X1 U2217 ( .B1(n359), .B2(n6), .C1(n391), .C2(n1210), .A(n4035), .ZN(
        n4042) );
  AOI22_X1 U2218 ( .A1(n5137), .A2(n987), .B1(n5169), .B2(n1218), .ZN(n4036)
         );
  OAI221_X1 U2219 ( .B1(n1222), .B2(n4038), .C1(n1221), .C2(n4037), .A(n4036), 
        .ZN(n4041) );
  AOI22_X1 U2220 ( .A1(n5201), .A2(n710), .B1(n5233), .B2(n40), .ZN(n4039) );
  OAI221_X1 U2221 ( .B1(n1229), .B2(n191), .C1(n1227), .C2(n340), .A(n4039), 
        .ZN(n4040) );
  NOR4_X1 U2222 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4045)
         );
  OAI222_X1 U2223 ( .A1(n807), .A2(n1239), .B1(n4045), .B2(n1236), .C1(n1233), 
        .C2(n4044), .ZN(n4046) );
  OAI22_X1 U2224 ( .A1(n1249), .A2(n4048), .B1(n935), .B2(n1246), .ZN(n4049)
         );
  AOI221_X1 U2225 ( .B1(n4817), .B2(n33), .C1(n1252), .C2(n4310), .A(n4049), 
        .ZN(n4057) );
  OAI222_X1 U2226 ( .A1(n615), .A2(n1264), .B1(n1261), .B2(n4051), .C1(n1257), 
        .C2(n4050), .ZN(n4052) );
  AOI221_X1 U2227 ( .B1(n1270), .B2(n4258), .C1(n1267), .C2(n4226), .A(n4052), 
        .ZN(n4056) );
  OAI22_X1 U2228 ( .A1(n4721), .A2(n1275), .B1(n1442), .B2(n1273), .ZN(n4053)
         );
  AOI221_X1 U2229 ( .B1(n4977), .B2(n1283), .C1(n1280), .C2(n4054), .A(n4053), 
        .ZN(n4055) );
  AOI22_X1 U2230 ( .A1(n1199), .A2(n4059), .B1(n1197), .B2(n4129), .ZN(n4060)
         );
  OAI221_X1 U2231 ( .B1(n1206), .B2(n320), .C1(n230), .C2(n1204), .A(n4060), 
        .ZN(n4069) );
  AOI22_X1 U2232 ( .A1(n689), .A2(n4193), .B1(n1209), .B2(n4161), .ZN(n4061)
         );
  OAI221_X1 U2233 ( .B1(n358), .B2(n6), .C1(n390), .C2(n1210), .A(n4061), .ZN(
        n4068) );
  AOI22_X1 U2234 ( .A1(n704), .A2(n5138), .B1(n5170), .B2(n1218), .ZN(n4062)
         );
  OAI221_X1 U2235 ( .B1(n1222), .B2(n4064), .C1(n1221), .C2(n4063), .A(n4062), 
        .ZN(n4067) );
  AOI22_X1 U2236 ( .A1(n5202), .A2(n710), .B1(n5234), .B2(n40), .ZN(n4065) );
  OAI221_X1 U2237 ( .B1(n1229), .B2(n192), .C1(n1227), .C2(n341), .A(n4065), 
        .ZN(n4066) );
  NOR4_X1 U2238 ( .A1(n4069), .A2(n4068), .A3(n4067), .A4(n4066), .ZN(n4071)
         );
  OAI222_X1 U2239 ( .A1(n806), .A2(n1239), .B1(n4071), .B2(n1236), .C1(n1233), 
        .C2(n4070), .ZN(n4072) );
  OAI22_X1 U2240 ( .A1(n1248), .A2(n4074), .B1(n934), .B2(n480), .ZN(n4075) );
  AOI221_X1 U2241 ( .B1(n4818), .B2(n1254), .C1(n1252), .C2(n4309), .A(n4075), 
        .ZN(n4083) );
  OAI222_X1 U2242 ( .A1(n614), .A2(n1264), .B1(n1261), .B2(n4077), .C1(n1257), 
        .C2(n4076), .ZN(n4078) );
  AOI221_X1 U2243 ( .B1(n1270), .B2(n4257), .C1(n1267), .C2(n4225), .A(n4078), 
        .ZN(n4082) );
  OAI22_X1 U2244 ( .A1(n4722), .A2(n1275), .B1(n1445), .B2(n1273), .ZN(n4079)
         );
  AOI221_X1 U2245 ( .B1(n4978), .B2(n1283), .C1(n1280), .C2(n4080), .A(n4079), 
        .ZN(n4081) );
  AOI22_X1 U2246 ( .A1(n1201), .A2(n4085), .B1(n1198), .B2(n4128), .ZN(n4086)
         );
  OAI221_X1 U2247 ( .B1(n1206), .B2(n321), .C1(n229), .C2(n1204), .A(n4086), 
        .ZN(n4103) );
  AOI22_X1 U2248 ( .A1(n689), .A2(n4192), .B1(n1209), .B2(n4160), .ZN(n4089)
         );
  OAI221_X1 U2249 ( .B1(n357), .B2(n1214), .C1(n389), .C2(n1211), .A(n4089), 
        .ZN(n4102) );
  AOI22_X1 U2250 ( .A1(n589), .A2(n5139), .B1(n5171), .B2(n1218), .ZN(n4092)
         );
  OAI221_X1 U2251 ( .B1(n1224), .B2(n4095), .C1(n1221), .C2(n4093), .A(n4092), 
        .ZN(n4101) );
  AOI22_X1 U2252 ( .A1(n5203), .A2(n2), .B1(n5235), .B2(n931), .ZN(n4097) );
  OAI221_X1 U2253 ( .B1(n1229), .B2(n193), .C1(n1227), .C2(n342), .A(n4097), 
        .ZN(n4100) );
  NOR4_X1 U2254 ( .A1(n4103), .A2(n4100), .A3(n4102), .A4(n4101), .ZN(n4107)
         );
  OAI222_X1 U2255 ( .A1(n805), .A2(n1239), .B1(n4107), .B2(n1236), .C1(n1233), 
        .C2(n4104), .ZN(n4109) );
  OAI22_X1 U2256 ( .A1(n1248), .A2(n4112), .B1(n933), .B2(n480), .ZN(n4114) );
  AOI221_X1 U2257 ( .B1(n4819), .B2(n1254), .C1(n1252), .C2(n4308), .A(n4114), 
        .ZN(n4126) );
  OAI222_X1 U2258 ( .A1(n613), .A2(n1264), .B1(n1260), .B2(n4117), .C1(n590), 
        .C2(n4115), .ZN(n4120) );
  AOI221_X1 U2259 ( .B1(n1270), .B2(n4256), .C1(n1267), .C2(n4224), .A(n4120), 
        .ZN(n4125) );
  OAI22_X1 U2260 ( .A1(n4723), .A2(n1276), .B1(n1448), .B2(n1273), .ZN(n4122)
         );
  AOI221_X1 U2261 ( .B1(n4979), .B2(n1283), .C1(n1280), .C2(n4123), .A(n4122), 
        .ZN(n4124) );
  NAND4_X1 U2262 ( .A1(n4127), .A2(n4124), .A3(n4125), .A4(n4126), .ZN(n2569)
         );
  MUX2_X1 U2263 ( .A(n4128), .B(n1446), .S(n1286), .Z(n3561) );
  MUX2_X1 U2264 ( .A(n4129), .B(n1443), .S(n1286), .Z(n3560) );
  MUX2_X1 U2265 ( .A(n4130), .B(n1440), .S(n1286), .Z(n3559) );
  MUX2_X1 U2266 ( .A(n4131), .B(n1437), .S(n1286), .Z(n3558) );
  MUX2_X1 U2267 ( .A(n4132), .B(n1434), .S(n1286), .Z(n3557) );
  MUX2_X1 U2268 ( .A(n4133), .B(n1431), .S(n1286), .Z(n3556) );
  MUX2_X1 U2269 ( .A(n4134), .B(n1428), .S(n1286), .Z(n3555) );
  MUX2_X1 U2270 ( .A(n4135), .B(n1425), .S(n1286), .Z(n3554) );
  MUX2_X1 U2271 ( .A(n4136), .B(n1423), .S(n1285), .Z(n3553) );
  MUX2_X1 U2272 ( .A(n4137), .B(n1421), .S(n1285), .Z(n3552) );
  MUX2_X1 U2273 ( .A(n4138), .B(n1419), .S(n1285), .Z(n3551) );
  MUX2_X1 U2274 ( .A(n4139), .B(n1417), .S(n1285), .Z(n3550) );
  MUX2_X1 U2275 ( .A(n4140), .B(n1415), .S(n1285), .Z(n3549) );
  MUX2_X1 U2276 ( .A(n4141), .B(n1413), .S(n1285), .Z(n3548) );
  MUX2_X1 U2277 ( .A(n4142), .B(n1411), .S(n1285), .Z(n3547) );
  MUX2_X1 U2278 ( .A(n4143), .B(n1409), .S(n1285), .Z(n3546) );
  MUX2_X1 U2279 ( .A(n4144), .B(n1407), .S(n1285), .Z(n3545) );
  MUX2_X1 U2280 ( .A(n4145), .B(n1405), .S(n1285), .Z(n3544) );
  MUX2_X1 U2281 ( .A(n4146), .B(n1403), .S(n1285), .Z(n3543) );
  MUX2_X1 U2282 ( .A(n4147), .B(n1401), .S(n1285), .Z(n3542) );
  MUX2_X1 U2283 ( .A(n4148), .B(n1399), .S(n1284), .Z(n3541) );
  MUX2_X1 U2284 ( .A(n4149), .B(n1397), .S(n1284), .Z(n3540) );
  MUX2_X1 U2285 ( .A(n4150), .B(n1395), .S(n1284), .Z(n3539) );
  MUX2_X1 U2286 ( .A(n4151), .B(n1393), .S(n1284), .Z(n3538) );
  MUX2_X1 U2287 ( .A(n4152), .B(n1391), .S(n1284), .Z(n3537) );
  MUX2_X1 U2288 ( .A(n4153), .B(n1389), .S(n1284), .Z(n3536) );
  MUX2_X1 U2289 ( .A(n4154), .B(n1387), .S(n1284), .Z(n3535) );
  MUX2_X1 U2290 ( .A(n4155), .B(n1385), .S(n1284), .Z(n3534) );
  MUX2_X1 U2291 ( .A(n4156), .B(n1383), .S(n1284), .Z(n3533) );
  MUX2_X1 U2292 ( .A(n4157), .B(n1381), .S(n1284), .Z(n3532) );
  MUX2_X1 U2293 ( .A(n4158), .B(n1379), .S(n1284), .Z(n3531) );
  MUX2_X1 U2294 ( .A(n4159), .B(n1377), .S(n1284), .Z(n3530) );
  AND2_X1 U2295 ( .A1(n4341), .A2(n4342), .ZN(n4340) );
  MUX2_X1 U2296 ( .A(n5235), .B(n1446), .S(n1289), .Z(n3529) );
  MUX2_X1 U2297 ( .A(n5234), .B(n1443), .S(n1289), .Z(n3528) );
  MUX2_X1 U2298 ( .A(n5233), .B(n1440), .S(n1289), .Z(n3527) );
  MUX2_X1 U2299 ( .A(n5232), .B(n1437), .S(n1289), .Z(n3526) );
  MUX2_X1 U2300 ( .A(n5231), .B(n1434), .S(n1289), .Z(n3525) );
  MUX2_X1 U2301 ( .A(n5230), .B(n1431), .S(n1289), .Z(n3524) );
  MUX2_X1 U2302 ( .A(n5229), .B(n1428), .S(n1289), .Z(n3523) );
  MUX2_X1 U2303 ( .A(n5228), .B(n1425), .S(n1289), .Z(n3522) );
  MUX2_X1 U2304 ( .A(n5227), .B(n1423), .S(n1288), .Z(n3521) );
  MUX2_X1 U2305 ( .A(n5226), .B(n1421), .S(n1288), .Z(n3520) );
  MUX2_X1 U2306 ( .A(n5225), .B(n1419), .S(n1288), .Z(n3519) );
  MUX2_X1 U2307 ( .A(n5224), .B(n1417), .S(n1288), .Z(n3518) );
  MUX2_X1 U2308 ( .A(n5223), .B(n1415), .S(n1288), .Z(n3517) );
  MUX2_X1 U2309 ( .A(n5222), .B(n1413), .S(n1288), .Z(n3516) );
  MUX2_X1 U2310 ( .A(n5221), .B(n1411), .S(n1288), .Z(n3515) );
  MUX2_X1 U2311 ( .A(n5220), .B(n1409), .S(n1288), .Z(n3514) );
  MUX2_X1 U2312 ( .A(n5219), .B(n1407), .S(n1288), .Z(n3513) );
  MUX2_X1 U2313 ( .A(n5218), .B(n1405), .S(n1288), .Z(n3512) );
  MUX2_X1 U2314 ( .A(n5217), .B(n1403), .S(n1288), .Z(n3511) );
  MUX2_X1 U2315 ( .A(n5216), .B(n1401), .S(n1288), .Z(n3510) );
  MUX2_X1 U2316 ( .A(n5215), .B(n1399), .S(n1287), .Z(n3509) );
  MUX2_X1 U2317 ( .A(n5214), .B(n1397), .S(n1287), .Z(n3508) );
  MUX2_X1 U2318 ( .A(n5213), .B(n1395), .S(n1287), .Z(n3507) );
  MUX2_X1 U2319 ( .A(n5212), .B(n1393), .S(n1287), .Z(n3506) );
  MUX2_X1 U2320 ( .A(n5211), .B(n1391), .S(n1287), .Z(n3505) );
  MUX2_X1 U2321 ( .A(n5210), .B(n1389), .S(n1287), .Z(n3504) );
  MUX2_X1 U2322 ( .A(n5209), .B(n1387), .S(n1287), .Z(n3503) );
  MUX2_X1 U2323 ( .A(n5208), .B(n1385), .S(n1287), .Z(n3502) );
  MUX2_X1 U2324 ( .A(n5207), .B(n1383), .S(n1287), .Z(n3501) );
  MUX2_X1 U2325 ( .A(n5206), .B(n1381), .S(n1287), .Z(n3500) );
  MUX2_X1 U2326 ( .A(n5205), .B(n1379), .S(n1287), .Z(n3499) );
  MUX2_X1 U2327 ( .A(n5204), .B(n1377), .S(n1287), .Z(n3498) );
  AND2_X1 U2328 ( .A1(n4344), .A2(n4342), .ZN(n4343) );
  MUX2_X1 U2329 ( .A(n5203), .B(n1446), .S(n1292), .Z(n3497) );
  MUX2_X1 U2330 ( .A(n5202), .B(n1443), .S(n1292), .Z(n3496) );
  MUX2_X1 U2331 ( .A(n5201), .B(n1440), .S(n1292), .Z(n3495) );
  MUX2_X1 U2332 ( .A(n5200), .B(n1437), .S(n1292), .Z(n3494) );
  MUX2_X1 U2333 ( .A(n5199), .B(n1434), .S(n1292), .Z(n3493) );
  MUX2_X1 U2334 ( .A(n5198), .B(n1431), .S(n1292), .Z(n3492) );
  MUX2_X1 U2335 ( .A(n5197), .B(n1428), .S(n1292), .Z(n3491) );
  MUX2_X1 U2336 ( .A(n5196), .B(n1425), .S(n1292), .Z(n3490) );
  MUX2_X1 U2337 ( .A(n5195), .B(n1423), .S(n1291), .Z(n3489) );
  MUX2_X1 U2338 ( .A(n5194), .B(n1421), .S(n1291), .Z(n3488) );
  MUX2_X1 U2339 ( .A(n5193), .B(n1419), .S(n1291), .Z(n3487) );
  MUX2_X1 U2340 ( .A(n5192), .B(n1417), .S(n1291), .Z(n3486) );
  MUX2_X1 U2341 ( .A(n5191), .B(n1415), .S(n1291), .Z(n3485) );
  MUX2_X1 U2342 ( .A(n5190), .B(n1413), .S(n1291), .Z(n3484) );
  MUX2_X1 U2343 ( .A(n5189), .B(n1411), .S(n1291), .Z(n3483) );
  MUX2_X1 U2344 ( .A(n5188), .B(n1409), .S(n1291), .Z(n3482) );
  MUX2_X1 U2345 ( .A(n5187), .B(n1407), .S(n1291), .Z(n3481) );
  MUX2_X1 U2346 ( .A(n5186), .B(n1405), .S(n1291), .Z(n3480) );
  MUX2_X1 U2347 ( .A(n5185), .B(n1403), .S(n1291), .Z(n3479) );
  MUX2_X1 U2348 ( .A(n5184), .B(n1401), .S(n1291), .Z(n3478) );
  MUX2_X1 U2349 ( .A(n5183), .B(n1399), .S(n1290), .Z(n3477) );
  MUX2_X1 U2350 ( .A(n5182), .B(n1397), .S(n1290), .Z(n3476) );
  MUX2_X1 U2351 ( .A(n5181), .B(n1395), .S(n1290), .Z(n3475) );
  MUX2_X1 U2352 ( .A(n5180), .B(n1393), .S(n1290), .Z(n3474) );
  MUX2_X1 U2353 ( .A(n5179), .B(n1391), .S(n1290), .Z(n3473) );
  MUX2_X1 U2354 ( .A(n5178), .B(n1389), .S(n1290), .Z(n3472) );
  MUX2_X1 U2355 ( .A(n5177), .B(n1387), .S(n1290), .Z(n3471) );
  MUX2_X1 U2356 ( .A(n5176), .B(n1385), .S(n1290), .Z(n3470) );
  MUX2_X1 U2357 ( .A(n5175), .B(n1383), .S(n1290), .Z(n3469) );
  MUX2_X1 U2358 ( .A(n5174), .B(n1381), .S(n1290), .Z(n3468) );
  MUX2_X1 U2359 ( .A(n5173), .B(n1379), .S(n1290), .Z(n3467) );
  MUX2_X1 U2360 ( .A(n5172), .B(n1377), .S(n1290), .Z(n3466) );
  AND2_X1 U2361 ( .A1(n4346), .A2(n4342), .ZN(n4345) );
  MUX2_X1 U2362 ( .A(n4160), .B(n1446), .S(n1295), .Z(n3465) );
  MUX2_X1 U2363 ( .A(n4161), .B(n1443), .S(n1295), .Z(n3464) );
  MUX2_X1 U2364 ( .A(n4162), .B(n1440), .S(n1295), .Z(n3463) );
  MUX2_X1 U2365 ( .A(n4163), .B(n1437), .S(n1295), .Z(n3462) );
  MUX2_X1 U2366 ( .A(n4164), .B(n1434), .S(n1295), .Z(n3461) );
  MUX2_X1 U2367 ( .A(n4165), .B(n1431), .S(n1295), .Z(n3460) );
  MUX2_X1 U2368 ( .A(n4166), .B(n1428), .S(n1295), .Z(n3459) );
  MUX2_X1 U2369 ( .A(n4167), .B(n1425), .S(n1295), .Z(n3458) );
  MUX2_X1 U2370 ( .A(n4168), .B(n1423), .S(n1294), .Z(n3457) );
  MUX2_X1 U2371 ( .A(n4169), .B(n1421), .S(n1294), .Z(n3456) );
  MUX2_X1 U2372 ( .A(n4170), .B(n1419), .S(n1294), .Z(n3455) );
  MUX2_X1 U2373 ( .A(n4171), .B(n1417), .S(n1294), .Z(n3454) );
  MUX2_X1 U2374 ( .A(n4172), .B(n1415), .S(n1294), .Z(n3453) );
  MUX2_X1 U2375 ( .A(n4173), .B(n1413), .S(n1294), .Z(n3452) );
  MUX2_X1 U2376 ( .A(n4174), .B(n1411), .S(n1294), .Z(n3451) );
  MUX2_X1 U2377 ( .A(n4175), .B(n1409), .S(n1294), .Z(n3450) );
  MUX2_X1 U2378 ( .A(n4176), .B(n1407), .S(n1294), .Z(n3449) );
  MUX2_X1 U2379 ( .A(n4177), .B(n1405), .S(n1294), .Z(n3448) );
  MUX2_X1 U2380 ( .A(n4178), .B(n1403), .S(n1294), .Z(n3447) );
  MUX2_X1 U2381 ( .A(n4179), .B(n1401), .S(n1294), .Z(n3446) );
  MUX2_X1 U2382 ( .A(n4180), .B(n1399), .S(n1293), .Z(n3445) );
  MUX2_X1 U2383 ( .A(n4181), .B(n1397), .S(n1293), .Z(n3444) );
  MUX2_X1 U2384 ( .A(n4182), .B(n1395), .S(n1293), .Z(n3443) );
  MUX2_X1 U2385 ( .A(n4183), .B(n1393), .S(n1293), .Z(n3442) );
  MUX2_X1 U2386 ( .A(n4184), .B(n1391), .S(n1293), .Z(n3441) );
  MUX2_X1 U2387 ( .A(n4185), .B(n1389), .S(n1293), .Z(n3440) );
  MUX2_X1 U2388 ( .A(n4186), .B(n1387), .S(n1293), .Z(n3439) );
  MUX2_X1 U2389 ( .A(n4187), .B(n1385), .S(n1293), .Z(n3438) );
  MUX2_X1 U2390 ( .A(n4188), .B(n1383), .S(n1293), .Z(n3437) );
  MUX2_X1 U2391 ( .A(n4189), .B(n1381), .S(n1293), .Z(n3436) );
  MUX2_X1 U2392 ( .A(n4190), .B(n1379), .S(n1293), .Z(n3435) );
  MUX2_X1 U2393 ( .A(n4191), .B(n1377), .S(n1293), .Z(n3434) );
  AND2_X1 U2394 ( .A1(n4348), .A2(n4342), .ZN(n4347) );
  MUX2_X1 U2395 ( .A(n4192), .B(n1446), .S(n1298), .Z(n3433) );
  MUX2_X1 U2396 ( .A(n4193), .B(n1443), .S(n1298), .Z(n3432) );
  MUX2_X1 U2397 ( .A(n4194), .B(n1440), .S(n1298), .Z(n3431) );
  MUX2_X1 U2398 ( .A(n4195), .B(n1437), .S(n1298), .Z(n3430) );
  MUX2_X1 U2399 ( .A(n4196), .B(n1434), .S(n1298), .Z(n3429) );
  MUX2_X1 U2400 ( .A(n4197), .B(n1431), .S(n1298), .Z(n3428) );
  MUX2_X1 U2401 ( .A(n4198), .B(n1428), .S(n1298), .Z(n3427) );
  MUX2_X1 U2402 ( .A(n4199), .B(n1425), .S(n1298), .Z(n3426) );
  MUX2_X1 U2403 ( .A(n4200), .B(n1423), .S(n1297), .Z(n3425) );
  MUX2_X1 U2404 ( .A(n4201), .B(n1421), .S(n1297), .Z(n3424) );
  MUX2_X1 U2405 ( .A(n4202), .B(n1419), .S(n1297), .Z(n3423) );
  MUX2_X1 U2406 ( .A(n4203), .B(n1417), .S(n1297), .Z(n3422) );
  MUX2_X1 U2407 ( .A(n4204), .B(n1415), .S(n1297), .Z(n3421) );
  MUX2_X1 U2408 ( .A(n4205), .B(n1413), .S(n1297), .Z(n3420) );
  MUX2_X1 U2409 ( .A(n4206), .B(n1411), .S(n1297), .Z(n3419) );
  MUX2_X1 U2410 ( .A(n4207), .B(n1409), .S(n1297), .Z(n3418) );
  MUX2_X1 U2411 ( .A(n4208), .B(n1407), .S(n1297), .Z(n3417) );
  MUX2_X1 U2412 ( .A(n4209), .B(n1405), .S(n1297), .Z(n3416) );
  MUX2_X1 U2413 ( .A(n4210), .B(n1403), .S(n1297), .Z(n3415) );
  MUX2_X1 U2414 ( .A(n4211), .B(n1401), .S(n1297), .Z(n3414) );
  MUX2_X1 U2415 ( .A(n4212), .B(n1399), .S(n1296), .Z(n3413) );
  MUX2_X1 U2416 ( .A(n4213), .B(n1397), .S(n1296), .Z(n3412) );
  MUX2_X1 U2417 ( .A(n4214), .B(n1395), .S(n1296), .Z(n3411) );
  MUX2_X1 U2418 ( .A(n4215), .B(n1393), .S(n1296), .Z(n3410) );
  MUX2_X1 U2419 ( .A(n4216), .B(n1391), .S(n1296), .Z(n3409) );
  MUX2_X1 U2420 ( .A(n4217), .B(n1389), .S(n1296), .Z(n3408) );
  MUX2_X1 U2421 ( .A(n4218), .B(n1387), .S(n1296), .Z(n3407) );
  MUX2_X1 U2422 ( .A(n4219), .B(n1385), .S(n1296), .Z(n3406) );
  MUX2_X1 U2423 ( .A(n4220), .B(n1383), .S(n1296), .Z(n3405) );
  MUX2_X1 U2424 ( .A(n4221), .B(n1381), .S(n1296), .Z(n3404) );
  MUX2_X1 U2425 ( .A(n4222), .B(n1379), .S(n1296), .Z(n3403) );
  MUX2_X1 U2426 ( .A(n4223), .B(n1377), .S(n1296), .Z(n3402) );
  AND2_X1 U2427 ( .A1(n4350), .A2(n4342), .ZN(n4349) );
  MUX2_X1 U2428 ( .A(n5171), .B(n1446), .S(n1301), .Z(n3401) );
  MUX2_X1 U2429 ( .A(n5170), .B(n1443), .S(n1301), .Z(n3400) );
  MUX2_X1 U2430 ( .A(n5169), .B(n1440), .S(n1301), .Z(n3399) );
  MUX2_X1 U2431 ( .A(n5168), .B(n1437), .S(n1301), .Z(n3398) );
  MUX2_X1 U2432 ( .A(n5167), .B(n1434), .S(n1301), .Z(n3397) );
  MUX2_X1 U2433 ( .A(n5166), .B(n1431), .S(n1301), .Z(n3396) );
  MUX2_X1 U2434 ( .A(n5165), .B(n1428), .S(n1301), .Z(n3395) );
  MUX2_X1 U2435 ( .A(n5164), .B(n1425), .S(n1301), .Z(n3394) );
  MUX2_X1 U2436 ( .A(n5163), .B(n1423), .S(n1300), .Z(n3393) );
  MUX2_X1 U2437 ( .A(n5162), .B(n1421), .S(n1300), .Z(n3392) );
  MUX2_X1 U2438 ( .A(n5161), .B(n1419), .S(n1300), .Z(n3391) );
  MUX2_X1 U2439 ( .A(n5160), .B(n1417), .S(n1300), .Z(n3390) );
  MUX2_X1 U2440 ( .A(n5159), .B(n1415), .S(n1300), .Z(n3389) );
  MUX2_X1 U2441 ( .A(n5158), .B(n1413), .S(n1300), .Z(n3388) );
  MUX2_X1 U2442 ( .A(n5157), .B(n1411), .S(n1300), .Z(n3387) );
  MUX2_X1 U2443 ( .A(n5156), .B(n1409), .S(n1300), .Z(n3386) );
  MUX2_X1 U2444 ( .A(n5155), .B(n1407), .S(n1300), .Z(n3385) );
  MUX2_X1 U2445 ( .A(n5154), .B(n1405), .S(n1300), .Z(n3384) );
  MUX2_X1 U2446 ( .A(n5153), .B(n1403), .S(n1300), .Z(n3383) );
  MUX2_X1 U2447 ( .A(n5152), .B(n1401), .S(n1300), .Z(n3382) );
  MUX2_X1 U2448 ( .A(n5151), .B(n1399), .S(n1299), .Z(n3381) );
  MUX2_X1 U2449 ( .A(n5150), .B(n1397), .S(n1299), .Z(n3380) );
  MUX2_X1 U2450 ( .A(n5149), .B(n1395), .S(n1299), .Z(n3379) );
  MUX2_X1 U2451 ( .A(n5148), .B(n1393), .S(n1299), .Z(n3378) );
  MUX2_X1 U2452 ( .A(n5147), .B(n1391), .S(n1299), .Z(n3377) );
  MUX2_X1 U2453 ( .A(n5146), .B(n1389), .S(n1299), .Z(n3376) );
  MUX2_X1 U2454 ( .A(n5145), .B(n1387), .S(n1299), .Z(n3375) );
  MUX2_X1 U2455 ( .A(n5144), .B(n1385), .S(n1299), .Z(n3374) );
  MUX2_X1 U2456 ( .A(n5143), .B(n1383), .S(n1299), .Z(n3373) );
  MUX2_X1 U2457 ( .A(n5142), .B(n1381), .S(n1299), .Z(n3372) );
  MUX2_X1 U2458 ( .A(n5141), .B(n1379), .S(n1299), .Z(n3371) );
  MUX2_X1 U2459 ( .A(n5140), .B(n1377), .S(n1299), .Z(n3370) );
  AND2_X1 U2460 ( .A1(n4352), .A2(n4342), .ZN(n4351) );
  MUX2_X1 U2461 ( .A(n5139), .B(n1446), .S(n1304), .Z(n3369) );
  MUX2_X1 U2462 ( .A(n5138), .B(n1443), .S(n1304), .Z(n3368) );
  MUX2_X1 U2463 ( .A(n5137), .B(n1440), .S(n1304), .Z(n3367) );
  MUX2_X1 U2464 ( .A(n5136), .B(n1437), .S(n1304), .Z(n3366) );
  MUX2_X1 U2465 ( .A(n5135), .B(n1434), .S(n1304), .Z(n3365) );
  MUX2_X1 U2466 ( .A(n5134), .B(n1431), .S(n1304), .Z(n3364) );
  MUX2_X1 U2467 ( .A(n5133), .B(n1428), .S(n1304), .Z(n3363) );
  MUX2_X1 U2468 ( .A(n5132), .B(n1425), .S(n1304), .Z(n3362) );
  MUX2_X1 U2469 ( .A(n5131), .B(n1423), .S(n1303), .Z(n3361) );
  MUX2_X1 U2470 ( .A(n5130), .B(n1421), .S(n1303), .Z(n3360) );
  MUX2_X1 U2471 ( .A(n5129), .B(n1419), .S(n1303), .Z(n3359) );
  MUX2_X1 U2472 ( .A(n5128), .B(n1417), .S(n1303), .Z(n3358) );
  MUX2_X1 U2473 ( .A(n5127), .B(n1415), .S(n1303), .Z(n3357) );
  MUX2_X1 U2474 ( .A(n5126), .B(n1413), .S(n1303), .Z(n3356) );
  MUX2_X1 U2475 ( .A(n5125), .B(n1411), .S(n1303), .Z(n3355) );
  MUX2_X1 U2476 ( .A(n5124), .B(n1409), .S(n1303), .Z(n3354) );
  MUX2_X1 U2477 ( .A(n5123), .B(n1407), .S(n1303), .Z(n3353) );
  MUX2_X1 U2478 ( .A(n5122), .B(n1405), .S(n1303), .Z(n3352) );
  MUX2_X1 U2479 ( .A(n5121), .B(n1403), .S(n1303), .Z(n3351) );
  MUX2_X1 U2480 ( .A(n5120), .B(n1401), .S(n1303), .Z(n3350) );
  MUX2_X1 U2481 ( .A(n5119), .B(n1399), .S(n1302), .Z(n3349) );
  MUX2_X1 U2482 ( .A(n5118), .B(n1397), .S(n1302), .Z(n3348) );
  MUX2_X1 U2483 ( .A(n5117), .B(n1395), .S(n1302), .Z(n3347) );
  MUX2_X1 U2484 ( .A(n5116), .B(n1393), .S(n1302), .Z(n3346) );
  MUX2_X1 U2485 ( .A(n5115), .B(n1391), .S(n1302), .Z(n3345) );
  MUX2_X1 U2486 ( .A(n5114), .B(n1389), .S(n1302), .Z(n3344) );
  MUX2_X1 U2487 ( .A(n5113), .B(n1387), .S(n1302), .Z(n3343) );
  MUX2_X1 U2488 ( .A(n5112), .B(n1385), .S(n1302), .Z(n3342) );
  MUX2_X1 U2489 ( .A(n5111), .B(n1383), .S(n1302), .Z(n3341) );
  MUX2_X1 U2490 ( .A(n5110), .B(n1381), .S(n1302), .Z(n3340) );
  MUX2_X1 U2491 ( .A(n5109), .B(n1379), .S(n1302), .Z(n3339) );
  MUX2_X1 U2492 ( .A(n5108), .B(n1377), .S(n1302), .Z(n3338) );
  AND2_X1 U2493 ( .A1(n4354), .A2(n4342), .ZN(n4353) );
  AND3_X1 U2494 ( .A1(n4355), .A2(n4356), .A3(n4357), .ZN(n4342) );
  INV_X1 U2495 ( .A(n4358), .ZN(n3337) );
  MUX2_X1 U2496 ( .A(n229), .B(n1448), .S(n1307), .Z(n4358) );
  INV_X1 U2497 ( .A(n4360), .ZN(n3336) );
  MUX2_X1 U2498 ( .A(n230), .B(n1445), .S(n1307), .Z(n4360) );
  INV_X1 U2499 ( .A(n4361), .ZN(n3335) );
  MUX2_X1 U2500 ( .A(n231), .B(n1442), .S(n1307), .Z(n4361) );
  INV_X1 U2501 ( .A(n4362), .ZN(n3334) );
  MUX2_X1 U2502 ( .A(n232), .B(n1439), .S(n1307), .Z(n4362) );
  INV_X1 U2503 ( .A(n4363), .ZN(n3333) );
  MUX2_X1 U2504 ( .A(n233), .B(n1436), .S(n1307), .Z(n4363) );
  INV_X1 U2505 ( .A(n4364), .ZN(n3332) );
  MUX2_X1 U2506 ( .A(n234), .B(n1433), .S(n1307), .Z(n4364) );
  INV_X1 U2507 ( .A(n4365), .ZN(n3331) );
  MUX2_X1 U2508 ( .A(n235), .B(n1430), .S(n1307), .Z(n4365) );
  INV_X1 U2509 ( .A(n4366), .ZN(n3330) );
  MUX2_X1 U2510 ( .A(n236), .B(n1427), .S(n1307), .Z(n4366) );
  INV_X1 U2511 ( .A(n4367), .ZN(n3329) );
  MUX2_X1 U2512 ( .A(n237), .B(n1424), .S(n1306), .Z(n4367) );
  INV_X1 U2513 ( .A(n4368), .ZN(n3328) );
  MUX2_X1 U2514 ( .A(n238), .B(n1422), .S(n1306), .Z(n4368) );
  INV_X1 U2515 ( .A(n4369), .ZN(n3327) );
  MUX2_X1 U2516 ( .A(n239), .B(n1420), .S(n1306), .Z(n4369) );
  INV_X1 U2517 ( .A(n4370), .ZN(n3326) );
  MUX2_X1 U2518 ( .A(n240), .B(n1418), .S(n1306), .Z(n4370) );
  INV_X1 U2519 ( .A(n4371), .ZN(n3325) );
  MUX2_X1 U2520 ( .A(n241), .B(n1416), .S(n1306), .Z(n4371) );
  INV_X1 U2521 ( .A(n4372), .ZN(n3324) );
  MUX2_X1 U2522 ( .A(n242), .B(n1414), .S(n1306), .Z(n4372) );
  INV_X1 U2523 ( .A(n4373), .ZN(n3323) );
  MUX2_X1 U2524 ( .A(n243), .B(n1412), .S(n1306), .Z(n4373) );
  INV_X1 U2525 ( .A(n4374), .ZN(n3322) );
  MUX2_X1 U2526 ( .A(n244), .B(n1410), .S(n1306), .Z(n4374) );
  INV_X1 U2527 ( .A(n4375), .ZN(n3321) );
  MUX2_X1 U2528 ( .A(n245), .B(n1408), .S(n1306), .Z(n4375) );
  INV_X1 U2529 ( .A(n4376), .ZN(n3320) );
  MUX2_X1 U2530 ( .A(n246), .B(n1406), .S(n1306), .Z(n4376) );
  INV_X1 U2531 ( .A(n4377), .ZN(n3319) );
  MUX2_X1 U2532 ( .A(n247), .B(n1404), .S(n1306), .Z(n4377) );
  INV_X1 U2533 ( .A(n4378), .ZN(n3318) );
  MUX2_X1 U2534 ( .A(n248), .B(n1402), .S(n1306), .Z(n4378) );
  INV_X1 U2535 ( .A(n4379), .ZN(n3317) );
  MUX2_X1 U2536 ( .A(n249), .B(n1400), .S(n1305), .Z(n4379) );
  INV_X1 U2537 ( .A(n4380), .ZN(n3316) );
  MUX2_X1 U2538 ( .A(n250), .B(n1398), .S(n1305), .Z(n4380) );
  INV_X1 U2539 ( .A(n4381), .ZN(n3315) );
  MUX2_X1 U2540 ( .A(n251), .B(n1396), .S(n1305), .Z(n4381) );
  INV_X1 U2541 ( .A(n4382), .ZN(n3314) );
  MUX2_X1 U2542 ( .A(n252), .B(n1394), .S(n1305), .Z(n4382) );
  INV_X1 U2543 ( .A(n4383), .ZN(n3313) );
  MUX2_X1 U2544 ( .A(n253), .B(n1392), .S(n1305), .Z(n4383) );
  INV_X1 U2545 ( .A(n4384), .ZN(n3312) );
  MUX2_X1 U2546 ( .A(n254), .B(n1390), .S(n1305), .Z(n4384) );
  INV_X1 U2547 ( .A(n4385), .ZN(n3311) );
  MUX2_X1 U2548 ( .A(n255), .B(n1388), .S(n1305), .Z(n4385) );
  INV_X1 U2549 ( .A(n4386), .ZN(n3310) );
  MUX2_X1 U2550 ( .A(n256), .B(n1386), .S(n1305), .Z(n4386) );
  INV_X1 U2551 ( .A(n4387), .ZN(n3309) );
  MUX2_X1 U2552 ( .A(n257), .B(n1384), .S(n1305), .Z(n4387) );
  INV_X1 U2553 ( .A(n4388), .ZN(n3308) );
  MUX2_X1 U2554 ( .A(n258), .B(n1382), .S(n1305), .Z(n4388) );
  INV_X1 U2555 ( .A(n4389), .ZN(n3307) );
  MUX2_X1 U2556 ( .A(n259), .B(n1380), .S(n1305), .Z(n4389) );
  INV_X1 U2557 ( .A(n4390), .ZN(n3306) );
  MUX2_X1 U2558 ( .A(n260), .B(n1378), .S(n1305), .Z(n4390) );
  AND2_X1 U2559 ( .A1(n4391), .A2(n4392), .ZN(n4359) );
  INV_X1 U2560 ( .A(n4393), .ZN(n3305) );
  MUX2_X1 U2561 ( .A(n261), .B(n1448), .S(n1310), .Z(n4393) );
  INV_X1 U2562 ( .A(n4395), .ZN(n3304) );
  MUX2_X1 U2563 ( .A(n262), .B(n1445), .S(n1310), .Z(n4395) );
  INV_X1 U2564 ( .A(n4396), .ZN(n3303) );
  MUX2_X1 U2565 ( .A(n263), .B(n1442), .S(n1310), .Z(n4396) );
  INV_X1 U2566 ( .A(n4397), .ZN(n3302) );
  MUX2_X1 U2567 ( .A(n264), .B(n1439), .S(n1310), .Z(n4397) );
  INV_X1 U2568 ( .A(n4398), .ZN(n3301) );
  MUX2_X1 U2569 ( .A(n265), .B(n1436), .S(n1310), .Z(n4398) );
  INV_X1 U2570 ( .A(n4399), .ZN(n3300) );
  MUX2_X1 U2571 ( .A(n266), .B(n1433), .S(n1310), .Z(n4399) );
  INV_X1 U2572 ( .A(n4400), .ZN(n3299) );
  MUX2_X1 U2573 ( .A(n267), .B(n1430), .S(n1310), .Z(n4400) );
  INV_X1 U2574 ( .A(n4401), .ZN(n3298) );
  MUX2_X1 U2575 ( .A(n268), .B(n1427), .S(n1310), .Z(n4401) );
  INV_X1 U2576 ( .A(n4402), .ZN(n3297) );
  MUX2_X1 U2577 ( .A(n269), .B(n1424), .S(n1309), .Z(n4402) );
  INV_X1 U2578 ( .A(n4403), .ZN(n3296) );
  MUX2_X1 U2579 ( .A(n270), .B(n1422), .S(n1309), .Z(n4403) );
  INV_X1 U2580 ( .A(n4404), .ZN(n3295) );
  MUX2_X1 U2581 ( .A(n271), .B(n1420), .S(n1309), .Z(n4404) );
  INV_X1 U2582 ( .A(n4405), .ZN(n3294) );
  MUX2_X1 U2583 ( .A(n272), .B(n1418), .S(n1309), .Z(n4405) );
  INV_X1 U2584 ( .A(n4406), .ZN(n3293) );
  MUX2_X1 U2585 ( .A(n273), .B(n1416), .S(n1309), .Z(n4406) );
  INV_X1 U2586 ( .A(n4407), .ZN(n3292) );
  MUX2_X1 U2587 ( .A(n274), .B(n1414), .S(n1309), .Z(n4407) );
  INV_X1 U2588 ( .A(n4408), .ZN(n3291) );
  MUX2_X1 U2589 ( .A(n275), .B(n1412), .S(n1309), .Z(n4408) );
  INV_X1 U2590 ( .A(n4409), .ZN(n3290) );
  MUX2_X1 U2591 ( .A(n276), .B(n1410), .S(n1309), .Z(n4409) );
  INV_X1 U2592 ( .A(n4410), .ZN(n3289) );
  MUX2_X1 U2593 ( .A(n277), .B(n1408), .S(n1309), .Z(n4410) );
  INV_X1 U2594 ( .A(n4411), .ZN(n3288) );
  MUX2_X1 U2595 ( .A(n278), .B(n1406), .S(n1309), .Z(n4411) );
  INV_X1 U2596 ( .A(n4412), .ZN(n3287) );
  MUX2_X1 U2597 ( .A(n279), .B(n1404), .S(n1309), .Z(n4412) );
  INV_X1 U2598 ( .A(n4413), .ZN(n3286) );
  MUX2_X1 U2599 ( .A(n280), .B(n1402), .S(n1309), .Z(n4413) );
  INV_X1 U2600 ( .A(n4414), .ZN(n3285) );
  MUX2_X1 U2601 ( .A(n281), .B(n1400), .S(n1308), .Z(n4414) );
  INV_X1 U2602 ( .A(n4415), .ZN(n3284) );
  MUX2_X1 U2603 ( .A(n282), .B(n1398), .S(n1308), .Z(n4415) );
  INV_X1 U2604 ( .A(n4416), .ZN(n3283) );
  MUX2_X1 U2605 ( .A(n283), .B(n1396), .S(n1308), .Z(n4416) );
  INV_X1 U2606 ( .A(n4417), .ZN(n3282) );
  MUX2_X1 U2607 ( .A(n284), .B(n1394), .S(n1308), .Z(n4417) );
  INV_X1 U2608 ( .A(n4418), .ZN(n3281) );
  MUX2_X1 U2609 ( .A(n285), .B(n1392), .S(n1308), .Z(n4418) );
  INV_X1 U2610 ( .A(n4419), .ZN(n3280) );
  MUX2_X1 U2611 ( .A(n286), .B(n1390), .S(n1308), .Z(n4419) );
  INV_X1 U2612 ( .A(n4420), .ZN(n3279) );
  MUX2_X1 U2613 ( .A(n287), .B(n1388), .S(n1308), .Z(n4420) );
  INV_X1 U2614 ( .A(n4421), .ZN(n3278) );
  MUX2_X1 U2615 ( .A(n288), .B(n1386), .S(n1308), .Z(n4421) );
  INV_X1 U2616 ( .A(n4422), .ZN(n3277) );
  MUX2_X1 U2617 ( .A(n289), .B(n1384), .S(n1308), .Z(n4422) );
  INV_X1 U2618 ( .A(n4423), .ZN(n3276) );
  MUX2_X1 U2619 ( .A(n290), .B(n1382), .S(n1308), .Z(n4423) );
  INV_X1 U2620 ( .A(n4424), .ZN(n3275) );
  MUX2_X1 U2621 ( .A(n291), .B(n1380), .S(n1308), .Z(n4424) );
  INV_X1 U2622 ( .A(n4425), .ZN(n3274) );
  MUX2_X1 U2623 ( .A(n292), .B(n1378), .S(n1308), .Z(n4425) );
  AND2_X1 U2624 ( .A1(n4391), .A2(n4341), .ZN(n4394) );
  MUX2_X1 U2625 ( .A(n5107), .B(n1446), .S(n1313), .Z(n3273) );
  MUX2_X1 U2626 ( .A(n5106), .B(n1443), .S(n1313), .Z(n3272) );
  MUX2_X1 U2627 ( .A(n5105), .B(n1440), .S(n1313), .Z(n3271) );
  MUX2_X1 U2628 ( .A(n5104), .B(n1437), .S(n1313), .Z(n3270) );
  MUX2_X1 U2629 ( .A(n5103), .B(n1434), .S(n1313), .Z(n3269) );
  MUX2_X1 U2630 ( .A(n5102), .B(n1431), .S(n1313), .Z(n3268) );
  MUX2_X1 U2631 ( .A(n5101), .B(n1428), .S(n1313), .Z(n3267) );
  MUX2_X1 U2632 ( .A(n5100), .B(n1425), .S(n1313), .Z(n3266) );
  MUX2_X1 U2633 ( .A(n5099), .B(n1423), .S(n1312), .Z(n3265) );
  MUX2_X1 U2634 ( .A(n5098), .B(n1421), .S(n1312), .Z(n3264) );
  MUX2_X1 U2635 ( .A(n5097), .B(n1419), .S(n1312), .Z(n3263) );
  MUX2_X1 U2636 ( .A(n5096), .B(n1417), .S(n1312), .Z(n3262) );
  MUX2_X1 U2637 ( .A(n5095), .B(n1415), .S(n1312), .Z(n3261) );
  MUX2_X1 U2638 ( .A(n5094), .B(n1413), .S(n1312), .Z(n3260) );
  MUX2_X1 U2639 ( .A(n5093), .B(n1411), .S(n1312), .Z(n3259) );
  MUX2_X1 U2640 ( .A(n5092), .B(n1409), .S(n1312), .Z(n3258) );
  MUX2_X1 U2641 ( .A(n5091), .B(n1407), .S(n1312), .Z(n3257) );
  MUX2_X1 U2642 ( .A(n5090), .B(n1405), .S(n1312), .Z(n3256) );
  MUX2_X1 U2643 ( .A(n5089), .B(n1403), .S(n1312), .Z(n3255) );
  MUX2_X1 U2644 ( .A(n5088), .B(n1401), .S(n1312), .Z(n3254) );
  MUX2_X1 U2645 ( .A(n5087), .B(n1399), .S(n1311), .Z(n3253) );
  MUX2_X1 U2646 ( .A(n5086), .B(n1397), .S(n1311), .Z(n3252) );
  MUX2_X1 U2647 ( .A(n5085), .B(n1395), .S(n1311), .Z(n3251) );
  MUX2_X1 U2648 ( .A(n5084), .B(n1393), .S(n1311), .Z(n3250) );
  MUX2_X1 U2649 ( .A(n5083), .B(n1391), .S(n1311), .Z(n3249) );
  MUX2_X1 U2650 ( .A(n5082), .B(n1389), .S(n1311), .Z(n3248) );
  MUX2_X1 U2651 ( .A(n5081), .B(n1387), .S(n1311), .Z(n3247) );
  MUX2_X1 U2652 ( .A(n5080), .B(n1385), .S(n1311), .Z(n3246) );
  MUX2_X1 U2653 ( .A(n5079), .B(n1383), .S(n1311), .Z(n3245) );
  MUX2_X1 U2654 ( .A(n5078), .B(n1381), .S(n1311), .Z(n3244) );
  MUX2_X1 U2655 ( .A(n5077), .B(n1379), .S(n1311), .Z(n3243) );
  MUX2_X1 U2656 ( .A(n5076), .B(n1377), .S(n1311), .Z(n3242) );
  AND2_X1 U2657 ( .A1(n4391), .A2(n4344), .ZN(n4426) );
  MUX2_X1 U2658 ( .A(n5075), .B(n1446), .S(n1316), .Z(n3241) );
  MUX2_X1 U2659 ( .A(n5074), .B(n1443), .S(n1316), .Z(n3240) );
  MUX2_X1 U2660 ( .A(n5073), .B(n1440), .S(n1316), .Z(n3239) );
  MUX2_X1 U2661 ( .A(n5072), .B(n1437), .S(n1316), .Z(n3238) );
  MUX2_X1 U2662 ( .A(n5071), .B(n1434), .S(n1316), .Z(n3237) );
  MUX2_X1 U2663 ( .A(n5070), .B(n1431), .S(n1316), .Z(n3236) );
  MUX2_X1 U2664 ( .A(n5069), .B(n1428), .S(n1316), .Z(n3235) );
  MUX2_X1 U2665 ( .A(n5068), .B(n1425), .S(n1316), .Z(n3234) );
  MUX2_X1 U2666 ( .A(n5067), .B(n1423), .S(n1315), .Z(n3233) );
  MUX2_X1 U2667 ( .A(n5066), .B(n1421), .S(n1315), .Z(n3232) );
  MUX2_X1 U2668 ( .A(n5065), .B(n1419), .S(n1315), .Z(n3231) );
  MUX2_X1 U2669 ( .A(n5064), .B(n1417), .S(n1315), .Z(n3230) );
  MUX2_X1 U2670 ( .A(n5063), .B(n1415), .S(n1315), .Z(n3229) );
  MUX2_X1 U2671 ( .A(n5062), .B(n1413), .S(n1315), .Z(n3228) );
  MUX2_X1 U2672 ( .A(n5061), .B(n1411), .S(n1315), .Z(n3227) );
  MUX2_X1 U2673 ( .A(n5060), .B(n1409), .S(n1315), .Z(n3226) );
  MUX2_X1 U2674 ( .A(n5059), .B(n1407), .S(n1315), .Z(n3225) );
  MUX2_X1 U2675 ( .A(n5058), .B(n1405), .S(n1315), .Z(n3224) );
  MUX2_X1 U2676 ( .A(n5057), .B(n1403), .S(n1315), .Z(n3223) );
  MUX2_X1 U2677 ( .A(n5056), .B(n1401), .S(n1315), .Z(n3222) );
  MUX2_X1 U2678 ( .A(n5055), .B(n1399), .S(n1314), .Z(n3221) );
  MUX2_X1 U2679 ( .A(n5054), .B(n1397), .S(n1314), .Z(n3220) );
  MUX2_X1 U2680 ( .A(n5053), .B(n1395), .S(n1314), .Z(n3219) );
  MUX2_X1 U2681 ( .A(n5052), .B(n1393), .S(n1314), .Z(n3218) );
  MUX2_X1 U2682 ( .A(n5051), .B(n1391), .S(n1314), .Z(n3217) );
  MUX2_X1 U2683 ( .A(n5050), .B(n1389), .S(n1314), .Z(n3216) );
  MUX2_X1 U2684 ( .A(n5049), .B(n1387), .S(n1314), .Z(n3215) );
  MUX2_X1 U2685 ( .A(n5048), .B(n1385), .S(n1314), .Z(n3214) );
  MUX2_X1 U2686 ( .A(n5047), .B(n1383), .S(n1314), .Z(n3213) );
  MUX2_X1 U2687 ( .A(n5046), .B(n1381), .S(n1314), .Z(n3212) );
  MUX2_X1 U2688 ( .A(n5045), .B(n1379), .S(n1314), .Z(n3211) );
  MUX2_X1 U2689 ( .A(n5044), .B(n1377), .S(n1314), .Z(n3210) );
  AND2_X1 U2690 ( .A1(n4391), .A2(n4346), .ZN(n4427) );
  INV_X1 U2691 ( .A(n4428), .ZN(n3209) );
  MUX2_X1 U2692 ( .A(n357), .B(n1448), .S(n1319), .Z(n4428) );
  INV_X1 U2693 ( .A(n4430), .ZN(n3208) );
  MUX2_X1 U2694 ( .A(n358), .B(n1445), .S(n1319), .Z(n4430) );
  INV_X1 U2695 ( .A(n4431), .ZN(n3207) );
  MUX2_X1 U2696 ( .A(n359), .B(n1442), .S(n1319), .Z(n4431) );
  INV_X1 U2697 ( .A(n4432), .ZN(n3206) );
  MUX2_X1 U2698 ( .A(n360), .B(n1439), .S(n1319), .Z(n4432) );
  INV_X1 U2699 ( .A(n4433), .ZN(n3205) );
  MUX2_X1 U2700 ( .A(n361), .B(n1436), .S(n1319), .Z(n4433) );
  INV_X1 U2701 ( .A(n4434), .ZN(n3204) );
  MUX2_X1 U2702 ( .A(n362), .B(n1433), .S(n1319), .Z(n4434) );
  INV_X1 U2703 ( .A(n4435), .ZN(n3203) );
  MUX2_X1 U2704 ( .A(n363), .B(n1430), .S(n1319), .Z(n4435) );
  INV_X1 U2705 ( .A(n4436), .ZN(n3202) );
  MUX2_X1 U2706 ( .A(n364), .B(n1427), .S(n1319), .Z(n4436) );
  INV_X1 U2707 ( .A(n4437), .ZN(n3201) );
  MUX2_X1 U2708 ( .A(n365), .B(n1424), .S(n1318), .Z(n4437) );
  INV_X1 U2709 ( .A(n4438), .ZN(n3200) );
  MUX2_X1 U2710 ( .A(n366), .B(n1422), .S(n1318), .Z(n4438) );
  INV_X1 U2711 ( .A(n4439), .ZN(n3199) );
  MUX2_X1 U2712 ( .A(n367), .B(n1420), .S(n1318), .Z(n4439) );
  INV_X1 U2713 ( .A(n4440), .ZN(n3198) );
  MUX2_X1 U2714 ( .A(n368), .B(n1418), .S(n1318), .Z(n4440) );
  INV_X1 U2715 ( .A(n4441), .ZN(n3197) );
  MUX2_X1 U2716 ( .A(n369), .B(n1416), .S(n1318), .Z(n4441) );
  INV_X1 U2717 ( .A(n4442), .ZN(n3196) );
  MUX2_X1 U2718 ( .A(n370), .B(n1414), .S(n1318), .Z(n4442) );
  INV_X1 U2719 ( .A(n4443), .ZN(n3195) );
  MUX2_X1 U2720 ( .A(n371), .B(n1412), .S(n1318), .Z(n4443) );
  INV_X1 U2721 ( .A(n4444), .ZN(n3194) );
  MUX2_X1 U2722 ( .A(n372), .B(n1410), .S(n1318), .Z(n4444) );
  INV_X1 U2723 ( .A(n4445), .ZN(n3193) );
  MUX2_X1 U2724 ( .A(n373), .B(n1408), .S(n1318), .Z(n4445) );
  INV_X1 U2725 ( .A(n4446), .ZN(n3192) );
  MUX2_X1 U2726 ( .A(n374), .B(n1406), .S(n1318), .Z(n4446) );
  INV_X1 U2727 ( .A(n4447), .ZN(n3191) );
  MUX2_X1 U2728 ( .A(n375), .B(n1404), .S(n1318), .Z(n4447) );
  INV_X1 U2729 ( .A(n4448), .ZN(n3190) );
  MUX2_X1 U2730 ( .A(n376), .B(n1402), .S(n1318), .Z(n4448) );
  INV_X1 U2731 ( .A(n4449), .ZN(n3189) );
  MUX2_X1 U2732 ( .A(n377), .B(n1400), .S(n1317), .Z(n4449) );
  INV_X1 U2733 ( .A(n4450), .ZN(n3188) );
  MUX2_X1 U2734 ( .A(n378), .B(n1398), .S(n1317), .Z(n4450) );
  INV_X1 U2735 ( .A(n4451), .ZN(n3187) );
  MUX2_X1 U2736 ( .A(n379), .B(n1396), .S(n1317), .Z(n4451) );
  INV_X1 U2737 ( .A(n4452), .ZN(n3186) );
  MUX2_X1 U2738 ( .A(n380), .B(n1394), .S(n1317), .Z(n4452) );
  INV_X1 U2739 ( .A(n4453), .ZN(n3185) );
  MUX2_X1 U2740 ( .A(n381), .B(n1392), .S(n1317), .Z(n4453) );
  INV_X1 U2741 ( .A(n4454), .ZN(n3184) );
  MUX2_X1 U2742 ( .A(n382), .B(n1390), .S(n1317), .Z(n4454) );
  INV_X1 U2743 ( .A(n4455), .ZN(n3183) );
  MUX2_X1 U2744 ( .A(n383), .B(n1388), .S(n1317), .Z(n4455) );
  INV_X1 U2745 ( .A(n4456), .ZN(n3182) );
  MUX2_X1 U2746 ( .A(n384), .B(n1386), .S(n1317), .Z(n4456) );
  INV_X1 U2747 ( .A(n4457), .ZN(n3181) );
  MUX2_X1 U2748 ( .A(n385), .B(n1384), .S(n1317), .Z(n4457) );
  INV_X1 U2749 ( .A(n4458), .ZN(n3180) );
  MUX2_X1 U2750 ( .A(n386), .B(n1382), .S(n1317), .Z(n4458) );
  INV_X1 U2751 ( .A(n4459), .ZN(n3179) );
  MUX2_X1 U2752 ( .A(n387), .B(n1380), .S(n1317), .Z(n4459) );
  INV_X1 U2753 ( .A(n4460), .ZN(n3178) );
  MUX2_X1 U2754 ( .A(n388), .B(n1378), .S(n1317), .Z(n4460) );
  AND2_X1 U2755 ( .A1(n4391), .A2(n4348), .ZN(n4429) );
  INV_X1 U2756 ( .A(n4461), .ZN(n3177) );
  MUX2_X1 U2757 ( .A(n389), .B(n1448), .S(n1322), .Z(n4461) );
  INV_X1 U2758 ( .A(n4463), .ZN(n3176) );
  MUX2_X1 U2759 ( .A(n390), .B(n1445), .S(n1322), .Z(n4463) );
  INV_X1 U2760 ( .A(n4464), .ZN(n3175) );
  MUX2_X1 U2761 ( .A(n391), .B(n1442), .S(n1322), .Z(n4464) );
  INV_X1 U2762 ( .A(n4465), .ZN(n3174) );
  MUX2_X1 U2763 ( .A(n392), .B(n1439), .S(n1322), .Z(n4465) );
  INV_X1 U2764 ( .A(n4466), .ZN(n3173) );
  MUX2_X1 U2765 ( .A(n393), .B(n1436), .S(n1322), .Z(n4466) );
  INV_X1 U2766 ( .A(n4467), .ZN(n3172) );
  MUX2_X1 U2767 ( .A(n394), .B(n1433), .S(n1322), .Z(n4467) );
  INV_X1 U2768 ( .A(n4468), .ZN(n3171) );
  MUX2_X1 U2769 ( .A(n395), .B(n1430), .S(n1322), .Z(n4468) );
  INV_X1 U2770 ( .A(n4469), .ZN(n3170) );
  MUX2_X1 U2771 ( .A(n396), .B(n1427), .S(n1322), .Z(n4469) );
  INV_X1 U2772 ( .A(n4470), .ZN(n3169) );
  MUX2_X1 U2773 ( .A(n397), .B(n1424), .S(n1321), .Z(n4470) );
  INV_X1 U2774 ( .A(n4471), .ZN(n3168) );
  MUX2_X1 U2775 ( .A(n398), .B(n1422), .S(n1321), .Z(n4471) );
  INV_X1 U2776 ( .A(n4472), .ZN(n3167) );
  MUX2_X1 U2777 ( .A(n399), .B(n1420), .S(n1321), .Z(n4472) );
  INV_X1 U2778 ( .A(n4473), .ZN(n3166) );
  MUX2_X1 U2779 ( .A(n400), .B(n1418), .S(n1321), .Z(n4473) );
  INV_X1 U2780 ( .A(n4474), .ZN(n3165) );
  MUX2_X1 U2781 ( .A(n401), .B(n1416), .S(n1321), .Z(n4474) );
  INV_X1 U2782 ( .A(n4475), .ZN(n3164) );
  MUX2_X1 U2783 ( .A(n402), .B(n1414), .S(n1321), .Z(n4475) );
  INV_X1 U2784 ( .A(n4476), .ZN(n3163) );
  MUX2_X1 U2785 ( .A(n403), .B(n1412), .S(n1321), .Z(n4476) );
  INV_X1 U2786 ( .A(n4477), .ZN(n3162) );
  MUX2_X1 U2787 ( .A(n404), .B(n1410), .S(n1321), .Z(n4477) );
  INV_X1 U2788 ( .A(n4478), .ZN(n3161) );
  MUX2_X1 U2789 ( .A(n405), .B(n1408), .S(n1321), .Z(n4478) );
  INV_X1 U2790 ( .A(n4479), .ZN(n3160) );
  MUX2_X1 U2791 ( .A(n406), .B(n1406), .S(n1321), .Z(n4479) );
  INV_X1 U2792 ( .A(n4480), .ZN(n3159) );
  MUX2_X1 U2793 ( .A(n407), .B(n1404), .S(n1321), .Z(n4480) );
  INV_X1 U2794 ( .A(n4481), .ZN(n3158) );
  MUX2_X1 U2795 ( .A(n408), .B(n1402), .S(n1321), .Z(n4481) );
  INV_X1 U2796 ( .A(n4482), .ZN(n3157) );
  MUX2_X1 U2797 ( .A(n409), .B(n1400), .S(n1320), .Z(n4482) );
  INV_X1 U2798 ( .A(n4483), .ZN(n3156) );
  MUX2_X1 U2799 ( .A(n410), .B(n1398), .S(n1320), .Z(n4483) );
  INV_X1 U2800 ( .A(n4484), .ZN(n3155) );
  MUX2_X1 U2801 ( .A(n411), .B(n1396), .S(n1320), .Z(n4484) );
  INV_X1 U2802 ( .A(n4485), .ZN(n3154) );
  MUX2_X1 U2803 ( .A(n412), .B(n1394), .S(n1320), .Z(n4485) );
  INV_X1 U2804 ( .A(n4486), .ZN(n3153) );
  MUX2_X1 U2805 ( .A(n413), .B(n1392), .S(n1320), .Z(n4486) );
  INV_X1 U2806 ( .A(n4487), .ZN(n3152) );
  MUX2_X1 U2807 ( .A(n414), .B(n1390), .S(n1320), .Z(n4487) );
  INV_X1 U2808 ( .A(n4488), .ZN(n3151) );
  MUX2_X1 U2809 ( .A(n415), .B(n1388), .S(n1320), .Z(n4488) );
  INV_X1 U2810 ( .A(n4489), .ZN(n3150) );
  MUX2_X1 U2811 ( .A(n416), .B(n1386), .S(n1320), .Z(n4489) );
  INV_X1 U2812 ( .A(n4490), .ZN(n3149) );
  MUX2_X1 U2813 ( .A(n417), .B(n1384), .S(n1320), .Z(n4490) );
  INV_X1 U2814 ( .A(n4491), .ZN(n3148) );
  MUX2_X1 U2815 ( .A(n418), .B(n1382), .S(n1320), .Z(n4491) );
  INV_X1 U2816 ( .A(n4492), .ZN(n3147) );
  MUX2_X1 U2817 ( .A(n419), .B(n1380), .S(n1320), .Z(n4492) );
  INV_X1 U2818 ( .A(n4493), .ZN(n3146) );
  MUX2_X1 U2819 ( .A(n420), .B(n1378), .S(n1320), .Z(n4493) );
  AND2_X1 U2820 ( .A1(n4391), .A2(n4350), .ZN(n4462) );
  MUX2_X1 U2821 ( .A(n5043), .B(n1446), .S(n1325), .Z(n3145) );
  MUX2_X1 U2822 ( .A(n5042), .B(n1443), .S(n1325), .Z(n3144) );
  MUX2_X1 U2823 ( .A(n5041), .B(n1440), .S(n1325), .Z(n3143) );
  MUX2_X1 U2824 ( .A(n5040), .B(n1437), .S(n1325), .Z(n3142) );
  MUX2_X1 U2825 ( .A(n5039), .B(n1434), .S(n1325), .Z(n3141) );
  MUX2_X1 U2826 ( .A(n5038), .B(n1431), .S(n1325), .Z(n3140) );
  MUX2_X1 U2827 ( .A(n5037), .B(n1428), .S(n1325), .Z(n3139) );
  MUX2_X1 U2828 ( .A(n5036), .B(n1425), .S(n1325), .Z(n3138) );
  MUX2_X1 U2829 ( .A(n5035), .B(n1423), .S(n1324), .Z(n3137) );
  MUX2_X1 U2830 ( .A(n5034), .B(n1421), .S(n1324), .Z(n3136) );
  MUX2_X1 U2831 ( .A(n5033), .B(n1419), .S(n1324), .Z(n3135) );
  MUX2_X1 U2832 ( .A(n5032), .B(n1417), .S(n1324), .Z(n3134) );
  MUX2_X1 U2833 ( .A(n5031), .B(n1415), .S(n1324), .Z(n3133) );
  MUX2_X1 U2834 ( .A(n5030), .B(n1413), .S(n1324), .Z(n3132) );
  MUX2_X1 U2835 ( .A(n5029), .B(n1411), .S(n1324), .Z(n3131) );
  MUX2_X1 U2836 ( .A(n5028), .B(n1409), .S(n1324), .Z(n3130) );
  MUX2_X1 U2837 ( .A(n5027), .B(n1407), .S(n1324), .Z(n3129) );
  MUX2_X1 U2838 ( .A(n5026), .B(n1405), .S(n1324), .Z(n3128) );
  MUX2_X1 U2839 ( .A(n5025), .B(n1403), .S(n1324), .Z(n3127) );
  MUX2_X1 U2840 ( .A(n5024), .B(n1401), .S(n1324), .Z(n3126) );
  MUX2_X1 U2841 ( .A(n5023), .B(n1399), .S(n1323), .Z(n3125) );
  MUX2_X1 U2842 ( .A(n5022), .B(n1397), .S(n1323), .Z(n3124) );
  MUX2_X1 U2843 ( .A(n5021), .B(n1395), .S(n1323), .Z(n3123) );
  MUX2_X1 U2844 ( .A(n5020), .B(n1393), .S(n1323), .Z(n3122) );
  MUX2_X1 U2845 ( .A(n5019), .B(n1391), .S(n1323), .Z(n3121) );
  MUX2_X1 U2846 ( .A(n5018), .B(n1389), .S(n1323), .Z(n3120) );
  MUX2_X1 U2847 ( .A(n5017), .B(n1387), .S(n1323), .Z(n3119) );
  MUX2_X1 U2848 ( .A(n5016), .B(n1385), .S(n1323), .Z(n3118) );
  MUX2_X1 U2849 ( .A(n5015), .B(n1383), .S(n1323), .Z(n3117) );
  MUX2_X1 U2850 ( .A(n5014), .B(n1381), .S(n1323), .Z(n3116) );
  MUX2_X1 U2851 ( .A(n5013), .B(n1379), .S(n1323), .Z(n3115) );
  MUX2_X1 U2852 ( .A(n5012), .B(n1377), .S(n1323), .Z(n3114) );
  AND2_X1 U2853 ( .A1(n4391), .A2(n4352), .ZN(n4494) );
  MUX2_X1 U2854 ( .A(n5011), .B(n1446), .S(n1328), .Z(n3113) );
  MUX2_X1 U2855 ( .A(n5010), .B(n1443), .S(n1328), .Z(n3112) );
  MUX2_X1 U2856 ( .A(n5009), .B(n1440), .S(n1328), .Z(n3111) );
  MUX2_X1 U2857 ( .A(n5008), .B(n1437), .S(n1328), .Z(n3110) );
  MUX2_X1 U2858 ( .A(n5007), .B(n1434), .S(n1328), .Z(n3109) );
  MUX2_X1 U2859 ( .A(n5006), .B(n1431), .S(n1328), .Z(n3108) );
  MUX2_X1 U2860 ( .A(n5005), .B(n1428), .S(n1328), .Z(n3107) );
  MUX2_X1 U2861 ( .A(n5004), .B(n1425), .S(n1328), .Z(n3106) );
  MUX2_X1 U2862 ( .A(n5003), .B(n1423), .S(n1327), .Z(n3105) );
  MUX2_X1 U2863 ( .A(n5002), .B(n1421), .S(n1327), .Z(n3104) );
  MUX2_X1 U2864 ( .A(n5001), .B(n1419), .S(n1327), .Z(n3103) );
  MUX2_X1 U2865 ( .A(n5000), .B(n1417), .S(n1327), .Z(n3102) );
  MUX2_X1 U2866 ( .A(n4999), .B(n1415), .S(n1327), .Z(n3101) );
  MUX2_X1 U2867 ( .A(n4998), .B(n1413), .S(n1327), .Z(n3100) );
  MUX2_X1 U2868 ( .A(n4997), .B(n1411), .S(n1327), .Z(n3099) );
  MUX2_X1 U2869 ( .A(n4996), .B(n1409), .S(n1327), .Z(n3098) );
  MUX2_X1 U2870 ( .A(n4995), .B(n1407), .S(n1327), .Z(n3097) );
  MUX2_X1 U2871 ( .A(n4994), .B(n1405), .S(n1327), .Z(n3096) );
  MUX2_X1 U2872 ( .A(n4993), .B(n1403), .S(n1327), .Z(n3095) );
  MUX2_X1 U2873 ( .A(n4992), .B(n1401), .S(n1327), .Z(n3094) );
  MUX2_X1 U2874 ( .A(n4991), .B(n1399), .S(n1326), .Z(n3093) );
  MUX2_X1 U2875 ( .A(n4990), .B(n1397), .S(n1326), .Z(n3092) );
  MUX2_X1 U2876 ( .A(n4989), .B(n1395), .S(n1326), .Z(n3091) );
  MUX2_X1 U2877 ( .A(n4988), .B(n1393), .S(n1326), .Z(n3090) );
  MUX2_X1 U2878 ( .A(n4987), .B(n1391), .S(n1326), .Z(n3089) );
  MUX2_X1 U2879 ( .A(n4986), .B(n1389), .S(n1326), .Z(n3088) );
  MUX2_X1 U2880 ( .A(n4985), .B(n1387), .S(n1326), .Z(n3087) );
  MUX2_X1 U2881 ( .A(n4984), .B(n1385), .S(n1326), .Z(n3086) );
  MUX2_X1 U2882 ( .A(n4983), .B(n1383), .S(n1326), .Z(n3085) );
  MUX2_X1 U2883 ( .A(n4982), .B(n1381), .S(n1326), .Z(n3084) );
  MUX2_X1 U2884 ( .A(n4981), .B(n1379), .S(n1326), .Z(n3083) );
  MUX2_X1 U2885 ( .A(n4980), .B(n1377), .S(n1326), .Z(n3082) );
  AND2_X1 U2886 ( .A1(n4391), .A2(n4354), .ZN(n4495) );
  AND3_X1 U2887 ( .A1(n4357), .A2(n4356), .A3(ADD_WR[3]), .ZN(n4391) );
  MUX2_X1 U2888 ( .A(n4224), .B(n1447), .S(n1331), .Z(n3081) );
  MUX2_X1 U2889 ( .A(n4225), .B(n1444), .S(n1331), .Z(n3080) );
  MUX2_X1 U2890 ( .A(n4226), .B(n1441), .S(n1331), .Z(n3079) );
  MUX2_X1 U2891 ( .A(n4227), .B(n1438), .S(n1331), .Z(n3078) );
  MUX2_X1 U2892 ( .A(n4228), .B(n1435), .S(n1331), .Z(n3077) );
  MUX2_X1 U2893 ( .A(n4229), .B(n1432), .S(n1331), .Z(n3076) );
  MUX2_X1 U2894 ( .A(n4230), .B(n1429), .S(n1331), .Z(n3075) );
  MUX2_X1 U2895 ( .A(n4231), .B(n1426), .S(n1331), .Z(n3074) );
  MUX2_X1 U2896 ( .A(n4232), .B(n1423), .S(n1330), .Z(n3073) );
  MUX2_X1 U2897 ( .A(n4233), .B(n1421), .S(n1330), .Z(n3072) );
  MUX2_X1 U2898 ( .A(n4234), .B(n1419), .S(n1330), .Z(n3071) );
  MUX2_X1 U2899 ( .A(n4235), .B(n1417), .S(n1330), .Z(n3070) );
  MUX2_X1 U2900 ( .A(n4236), .B(n1415), .S(n1330), .Z(n3069) );
  MUX2_X1 U2901 ( .A(n4237), .B(n1413), .S(n1330), .Z(n3068) );
  MUX2_X1 U2902 ( .A(n4238), .B(n1411), .S(n1330), .Z(n3067) );
  MUX2_X1 U2903 ( .A(n4239), .B(n1409), .S(n1330), .Z(n3066) );
  MUX2_X1 U2904 ( .A(n4240), .B(n1407), .S(n1330), .Z(n3065) );
  MUX2_X1 U2905 ( .A(n4241), .B(n1405), .S(n1330), .Z(n3064) );
  MUX2_X1 U2906 ( .A(n4242), .B(n1403), .S(n1330), .Z(n3063) );
  MUX2_X1 U2907 ( .A(n4243), .B(n1401), .S(n1330), .Z(n3062) );
  MUX2_X1 U2908 ( .A(n4244), .B(n1399), .S(n1329), .Z(n3061) );
  MUX2_X1 U2909 ( .A(n4245), .B(n1397), .S(n1329), .Z(n3060) );
  MUX2_X1 U2910 ( .A(n4246), .B(n1395), .S(n1329), .Z(n3059) );
  MUX2_X1 U2911 ( .A(n4247), .B(n1393), .S(n1329), .Z(n3058) );
  MUX2_X1 U2912 ( .A(n4248), .B(n1391), .S(n1329), .Z(n3057) );
  MUX2_X1 U2913 ( .A(n4249), .B(n1389), .S(n1329), .Z(n3056) );
  MUX2_X1 U2914 ( .A(n4250), .B(n1387), .S(n1329), .Z(n3055) );
  MUX2_X1 U2915 ( .A(n4251), .B(n1385), .S(n1329), .Z(n3054) );
  MUX2_X1 U2916 ( .A(n4252), .B(n1383), .S(n1329), .Z(n3053) );
  MUX2_X1 U2917 ( .A(n4253), .B(n1381), .S(n1329), .Z(n3052) );
  MUX2_X1 U2918 ( .A(n4254), .B(n1379), .S(n1329), .Z(n3051) );
  MUX2_X1 U2919 ( .A(n4255), .B(n1377), .S(n1329), .Z(n3050) );
  AND2_X1 U2920 ( .A1(n4497), .A2(n4392), .ZN(n4496) );
  INV_X1 U2921 ( .A(n4498), .ZN(n3049) );
  MUX2_X1 U2922 ( .A(n517), .B(n1448), .S(n1334), .Z(n4498) );
  INV_X1 U2923 ( .A(n4500), .ZN(n3048) );
  MUX2_X1 U2924 ( .A(n518), .B(n1445), .S(n1334), .Z(n4500) );
  INV_X1 U2925 ( .A(n4501), .ZN(n3047) );
  MUX2_X1 U2926 ( .A(n519), .B(n1442), .S(n1334), .Z(n4501) );
  INV_X1 U2927 ( .A(n4502), .ZN(n3046) );
  MUX2_X1 U2928 ( .A(n520), .B(n1439), .S(n1334), .Z(n4502) );
  INV_X1 U2929 ( .A(n4503), .ZN(n3045) );
  MUX2_X1 U2930 ( .A(n521), .B(n1436), .S(n1334), .Z(n4503) );
  INV_X1 U2931 ( .A(n4504), .ZN(n3044) );
  MUX2_X1 U2932 ( .A(n522), .B(n1433), .S(n1334), .Z(n4504) );
  INV_X1 U2933 ( .A(n4505), .ZN(n3043) );
  MUX2_X1 U2934 ( .A(n523), .B(n1430), .S(n1334), .Z(n4505) );
  INV_X1 U2935 ( .A(n4506), .ZN(n3042) );
  MUX2_X1 U2936 ( .A(n524), .B(n1427), .S(n1334), .Z(n4506) );
  INV_X1 U2937 ( .A(n4507), .ZN(n3041) );
  MUX2_X1 U2938 ( .A(n525), .B(n1424), .S(n1333), .Z(n4507) );
  INV_X1 U2939 ( .A(n4508), .ZN(n3040) );
  MUX2_X1 U2940 ( .A(n526), .B(n1422), .S(n1333), .Z(n4508) );
  INV_X1 U2941 ( .A(n4509), .ZN(n3039) );
  MUX2_X1 U2942 ( .A(n527), .B(n1420), .S(n1333), .Z(n4509) );
  INV_X1 U2943 ( .A(n4510), .ZN(n3038) );
  MUX2_X1 U2944 ( .A(n528), .B(n1418), .S(n1333), .Z(n4510) );
  INV_X1 U2945 ( .A(n4511), .ZN(n3037) );
  MUX2_X1 U2946 ( .A(n529), .B(n1416), .S(n1333), .Z(n4511) );
  INV_X1 U2947 ( .A(n4512), .ZN(n3036) );
  MUX2_X1 U2948 ( .A(n530), .B(n1414), .S(n1333), .Z(n4512) );
  INV_X1 U2949 ( .A(n4513), .ZN(n3035) );
  MUX2_X1 U2950 ( .A(n531), .B(n1412), .S(n1333), .Z(n4513) );
  INV_X1 U2951 ( .A(n4514), .ZN(n3034) );
  MUX2_X1 U2952 ( .A(n532), .B(n1410), .S(n1333), .Z(n4514) );
  INV_X1 U2953 ( .A(n4515), .ZN(n3033) );
  MUX2_X1 U2954 ( .A(n533), .B(n1408), .S(n1333), .Z(n4515) );
  INV_X1 U2955 ( .A(n4516), .ZN(n3032) );
  MUX2_X1 U2956 ( .A(n534), .B(n1406), .S(n1333), .Z(n4516) );
  INV_X1 U2957 ( .A(n4517), .ZN(n3031) );
  MUX2_X1 U2958 ( .A(n535), .B(n1404), .S(n1333), .Z(n4517) );
  INV_X1 U2959 ( .A(n4518), .ZN(n3030) );
  MUX2_X1 U2960 ( .A(n536), .B(n1402), .S(n1333), .Z(n4518) );
  INV_X1 U2961 ( .A(n4519), .ZN(n3029) );
  MUX2_X1 U2962 ( .A(n537), .B(n1400), .S(n1332), .Z(n4519) );
  INV_X1 U2963 ( .A(n4520), .ZN(n3028) );
  MUX2_X1 U2964 ( .A(n538), .B(n1398), .S(n1332), .Z(n4520) );
  INV_X1 U2965 ( .A(n4521), .ZN(n3027) );
  MUX2_X1 U2966 ( .A(n539), .B(n1396), .S(n1332), .Z(n4521) );
  INV_X1 U2967 ( .A(n4522), .ZN(n3026) );
  MUX2_X1 U2968 ( .A(n540), .B(n1394), .S(n1332), .Z(n4522) );
  INV_X1 U2969 ( .A(n4523), .ZN(n3025) );
  MUX2_X1 U2970 ( .A(n541), .B(n1392), .S(n1332), .Z(n4523) );
  INV_X1 U2971 ( .A(n4524), .ZN(n3024) );
  MUX2_X1 U2972 ( .A(n542), .B(n1390), .S(n1332), .Z(n4524) );
  INV_X1 U2973 ( .A(n4525), .ZN(n3023) );
  MUX2_X1 U2974 ( .A(n543), .B(n1388), .S(n1332), .Z(n4525) );
  INV_X1 U2975 ( .A(n4526), .ZN(n3022) );
  MUX2_X1 U2976 ( .A(n544), .B(n1386), .S(n1332), .Z(n4526) );
  INV_X1 U2977 ( .A(n4527), .ZN(n3021) );
  MUX2_X1 U2978 ( .A(n545), .B(n1384), .S(n1332), .Z(n4527) );
  INV_X1 U2979 ( .A(n4528), .ZN(n3020) );
  MUX2_X1 U2980 ( .A(n546), .B(n1382), .S(n1332), .Z(n4528) );
  INV_X1 U2981 ( .A(n4529), .ZN(n3019) );
  MUX2_X1 U2982 ( .A(n547), .B(n1380), .S(n1332), .Z(n4529) );
  INV_X1 U2983 ( .A(n4530), .ZN(n3018) );
  MUX2_X1 U2984 ( .A(n548), .B(n1378), .S(n1332), .Z(n4530) );
  AND2_X1 U2985 ( .A1(n4497), .A2(n4341), .ZN(n4499) );
  MUX2_X1 U2986 ( .A(n4979), .B(n1447), .S(n1337), .Z(n3017) );
  MUX2_X1 U2987 ( .A(n4978), .B(n1444), .S(n1337), .Z(n3016) );
  MUX2_X1 U2988 ( .A(n4977), .B(n1441), .S(n1337), .Z(n3015) );
  MUX2_X1 U2989 ( .A(n4976), .B(n1438), .S(n1337), .Z(n3014) );
  MUX2_X1 U2990 ( .A(n4975), .B(n1435), .S(n1337), .Z(n3013) );
  MUX2_X1 U2991 ( .A(n4974), .B(n1432), .S(n1337), .Z(n3012) );
  MUX2_X1 U2992 ( .A(n4973), .B(n1429), .S(n1337), .Z(n3011) );
  MUX2_X1 U2993 ( .A(n4972), .B(n1426), .S(n1337), .Z(n3010) );
  MUX2_X1 U2994 ( .A(n4971), .B(n1423), .S(n1336), .Z(n3009) );
  MUX2_X1 U2995 ( .A(n4970), .B(n1421), .S(n1336), .Z(n3008) );
  MUX2_X1 U2996 ( .A(n4969), .B(n1419), .S(n1336), .Z(n3007) );
  MUX2_X1 U2997 ( .A(n4968), .B(n1417), .S(n1336), .Z(n3006) );
  MUX2_X1 U2998 ( .A(n4967), .B(n1415), .S(n1336), .Z(n3005) );
  MUX2_X1 U2999 ( .A(n4966), .B(n1413), .S(n1336), .Z(n3004) );
  MUX2_X1 U3000 ( .A(n4965), .B(n1411), .S(n1336), .Z(n3003) );
  MUX2_X1 U3001 ( .A(n4964), .B(n1409), .S(n1336), .Z(n3002) );
  MUX2_X1 U3002 ( .A(n4963), .B(n1407), .S(n1336), .Z(n3001) );
  MUX2_X1 U3003 ( .A(n4962), .B(n1405), .S(n1336), .Z(n3000) );
  MUX2_X1 U3004 ( .A(n4961), .B(n1403), .S(n1336), .Z(n2999) );
  MUX2_X1 U3005 ( .A(n4960), .B(n1401), .S(n1336), .Z(n2998) );
  MUX2_X1 U3006 ( .A(n4959), .B(n1399), .S(n1335), .Z(n2997) );
  MUX2_X1 U3007 ( .A(n4958), .B(n1397), .S(n1335), .Z(n2996) );
  MUX2_X1 U3008 ( .A(n4957), .B(n1395), .S(n1335), .Z(n2995) );
  MUX2_X1 U3009 ( .A(n4956), .B(n1393), .S(n1335), .Z(n2994) );
  MUX2_X1 U3010 ( .A(n4955), .B(n1391), .S(n1335), .Z(n2993) );
  MUX2_X1 U3011 ( .A(n4954), .B(n1389), .S(n1335), .Z(n2992) );
  MUX2_X1 U3012 ( .A(n4953), .B(n1387), .S(n1335), .Z(n2991) );
  MUX2_X1 U3013 ( .A(n4952), .B(n1385), .S(n1335), .Z(n2990) );
  MUX2_X1 U3014 ( .A(n4951), .B(n1383), .S(n1335), .Z(n2989) );
  MUX2_X1 U3015 ( .A(n4950), .B(n1381), .S(n1335), .Z(n2988) );
  MUX2_X1 U3016 ( .A(n4949), .B(n1379), .S(n1335), .Z(n2987) );
  MUX2_X1 U3017 ( .A(n4948), .B(n1377), .S(n1335), .Z(n2986) );
  AND2_X1 U3018 ( .A1(n4497), .A2(n4344), .ZN(n4531) );
  MUX2_X1 U3019 ( .A(n4947), .B(n1447), .S(n1340), .Z(n2985) );
  MUX2_X1 U3020 ( .A(n4946), .B(n1444), .S(n1340), .Z(n2984) );
  MUX2_X1 U3021 ( .A(n4945), .B(n1441), .S(n1340), .Z(n2983) );
  MUX2_X1 U3022 ( .A(n4944), .B(n1438), .S(n1340), .Z(n2982) );
  MUX2_X1 U3023 ( .A(n4943), .B(n1435), .S(n1340), .Z(n2981) );
  MUX2_X1 U3024 ( .A(n4942), .B(n1432), .S(n1340), .Z(n2980) );
  MUX2_X1 U3025 ( .A(n4941), .B(n1429), .S(n1340), .Z(n2979) );
  MUX2_X1 U3026 ( .A(n4940), .B(n1426), .S(n1340), .Z(n2978) );
  MUX2_X1 U3027 ( .A(n4939), .B(n1423), .S(n1339), .Z(n2977) );
  MUX2_X1 U3028 ( .A(n4938), .B(n1421), .S(n1339), .Z(n2976) );
  MUX2_X1 U3029 ( .A(n4937), .B(n1419), .S(n1339), .Z(n2975) );
  MUX2_X1 U3030 ( .A(n4936), .B(n1417), .S(n1339), .Z(n2974) );
  MUX2_X1 U3031 ( .A(n4935), .B(n1415), .S(n1339), .Z(n2973) );
  MUX2_X1 U3032 ( .A(n4934), .B(n1413), .S(n1339), .Z(n2972) );
  MUX2_X1 U3033 ( .A(n4933), .B(n1411), .S(n1339), .Z(n2971) );
  MUX2_X1 U3034 ( .A(n4932), .B(n1409), .S(n1339), .Z(n2970) );
  MUX2_X1 U3035 ( .A(n4931), .B(n1407), .S(n1339), .Z(n2969) );
  MUX2_X1 U3036 ( .A(n4930), .B(n1405), .S(n1339), .Z(n2968) );
  MUX2_X1 U3037 ( .A(n4929), .B(n1403), .S(n1339), .Z(n2967) );
  MUX2_X1 U3038 ( .A(n4928), .B(n1401), .S(n1339), .Z(n2966) );
  MUX2_X1 U3039 ( .A(n4927), .B(n1399), .S(n1338), .Z(n2965) );
  MUX2_X1 U3040 ( .A(n4926), .B(n1397), .S(n1338), .Z(n2964) );
  MUX2_X1 U3041 ( .A(n4925), .B(n1395), .S(n1338), .Z(n2963) );
  MUX2_X1 U3042 ( .A(n4924), .B(n1393), .S(n1338), .Z(n2962) );
  MUX2_X1 U3043 ( .A(n4923), .B(n1391), .S(n1338), .Z(n2961) );
  MUX2_X1 U3044 ( .A(n4922), .B(n1389), .S(n1338), .Z(n2960) );
  MUX2_X1 U3045 ( .A(n4921), .B(n1387), .S(n1338), .Z(n2959) );
  MUX2_X1 U3046 ( .A(n4920), .B(n1385), .S(n1338), .Z(n2958) );
  MUX2_X1 U3047 ( .A(n4919), .B(n1383), .S(n1338), .Z(n2957) );
  MUX2_X1 U3048 ( .A(n4918), .B(n1381), .S(n1338), .Z(n2956) );
  MUX2_X1 U3049 ( .A(n4917), .B(n1379), .S(n1338), .Z(n2955) );
  MUX2_X1 U3050 ( .A(n4916), .B(n1377), .S(n1338), .Z(n2954) );
  AND2_X1 U3051 ( .A1(n4497), .A2(n4346), .ZN(n4532) );
  INV_X1 U3052 ( .A(n4533), .ZN(n2953) );
  MUX2_X1 U3053 ( .A(n613), .B(n1448), .S(n1343), .Z(n4533) );
  INV_X1 U3054 ( .A(n4535), .ZN(n2952) );
  MUX2_X1 U3055 ( .A(n614), .B(n1445), .S(n1343), .Z(n4535) );
  INV_X1 U3056 ( .A(n4536), .ZN(n2951) );
  MUX2_X1 U3057 ( .A(n615), .B(n1442), .S(n1343), .Z(n4536) );
  INV_X1 U3058 ( .A(n4537), .ZN(n2950) );
  MUX2_X1 U3059 ( .A(n616), .B(n1439), .S(n1343), .Z(n4537) );
  INV_X1 U3060 ( .A(n4538), .ZN(n2949) );
  MUX2_X1 U3061 ( .A(n617), .B(n1436), .S(n1343), .Z(n4538) );
  INV_X1 U3062 ( .A(n4539), .ZN(n2948) );
  MUX2_X1 U3063 ( .A(n618), .B(n1433), .S(n1343), .Z(n4539) );
  INV_X1 U3064 ( .A(n4540), .ZN(n2947) );
  MUX2_X1 U3065 ( .A(n619), .B(n1430), .S(n1343), .Z(n4540) );
  INV_X1 U3066 ( .A(n4541), .ZN(n2946) );
  MUX2_X1 U3067 ( .A(n620), .B(n1427), .S(n1343), .Z(n4541) );
  INV_X1 U3068 ( .A(n4542), .ZN(n2945) );
  MUX2_X1 U3069 ( .A(n621), .B(n1424), .S(n1342), .Z(n4542) );
  INV_X1 U3070 ( .A(n4543), .ZN(n2944) );
  MUX2_X1 U3071 ( .A(n622), .B(n1422), .S(n1342), .Z(n4543) );
  INV_X1 U3072 ( .A(n4544), .ZN(n2943) );
  MUX2_X1 U3073 ( .A(n623), .B(n1420), .S(n1342), .Z(n4544) );
  INV_X1 U3074 ( .A(n4545), .ZN(n2942) );
  MUX2_X1 U3075 ( .A(n624), .B(n1418), .S(n1342), .Z(n4545) );
  INV_X1 U3076 ( .A(n4546), .ZN(n2941) );
  MUX2_X1 U3077 ( .A(n625), .B(n1416), .S(n1342), .Z(n4546) );
  INV_X1 U3078 ( .A(n4547), .ZN(n2940) );
  MUX2_X1 U3079 ( .A(n626), .B(n1414), .S(n1342), .Z(n4547) );
  INV_X1 U3080 ( .A(n4548), .ZN(n2939) );
  MUX2_X1 U3081 ( .A(n627), .B(n1412), .S(n1342), .Z(n4548) );
  INV_X1 U3082 ( .A(n4549), .ZN(n2938) );
  MUX2_X1 U3083 ( .A(n628), .B(n1410), .S(n1342), .Z(n4549) );
  INV_X1 U3084 ( .A(n4550), .ZN(n2937) );
  MUX2_X1 U3085 ( .A(n629), .B(n1408), .S(n1342), .Z(n4550) );
  INV_X1 U3086 ( .A(n4551), .ZN(n2936) );
  MUX2_X1 U3087 ( .A(n630), .B(n1406), .S(n1342), .Z(n4551) );
  INV_X1 U3088 ( .A(n4552), .ZN(n2935) );
  MUX2_X1 U3089 ( .A(n631), .B(n1404), .S(n1342), .Z(n4552) );
  INV_X1 U3090 ( .A(n4553), .ZN(n2934) );
  MUX2_X1 U3091 ( .A(n632), .B(n1402), .S(n1342), .Z(n4553) );
  INV_X1 U3092 ( .A(n4554), .ZN(n2933) );
  MUX2_X1 U3093 ( .A(n633), .B(n1400), .S(n1341), .Z(n4554) );
  INV_X1 U3094 ( .A(n4555), .ZN(n2932) );
  MUX2_X1 U3095 ( .A(n634), .B(n1398), .S(n1341), .Z(n4555) );
  INV_X1 U3096 ( .A(n4556), .ZN(n2931) );
  MUX2_X1 U3097 ( .A(n635), .B(n1396), .S(n1341), .Z(n4556) );
  INV_X1 U3098 ( .A(n4557), .ZN(n2930) );
  MUX2_X1 U3099 ( .A(n636), .B(n1394), .S(n1341), .Z(n4557) );
  INV_X1 U3100 ( .A(n4558), .ZN(n2929) );
  MUX2_X1 U3101 ( .A(n637), .B(n1392), .S(n1341), .Z(n4558) );
  INV_X1 U3102 ( .A(n4559), .ZN(n2928) );
  MUX2_X1 U3103 ( .A(n638), .B(n1390), .S(n1341), .Z(n4559) );
  INV_X1 U3104 ( .A(n4560), .ZN(n2927) );
  MUX2_X1 U3105 ( .A(n639), .B(n1388), .S(n1341), .Z(n4560) );
  INV_X1 U3106 ( .A(n4561), .ZN(n2926) );
  MUX2_X1 U3107 ( .A(n640), .B(n1386), .S(n1341), .Z(n4561) );
  INV_X1 U3108 ( .A(n4562), .ZN(n2925) );
  MUX2_X1 U3109 ( .A(n641), .B(n1384), .S(n1341), .Z(n4562) );
  INV_X1 U3110 ( .A(n4563), .ZN(n2924) );
  MUX2_X1 U3111 ( .A(n642), .B(n1382), .S(n1341), .Z(n4563) );
  INV_X1 U3112 ( .A(n4564), .ZN(n2923) );
  MUX2_X1 U3113 ( .A(n643), .B(n1380), .S(n1341), .Z(n4564) );
  INV_X1 U3114 ( .A(n4565), .ZN(n2922) );
  MUX2_X1 U3115 ( .A(n644), .B(n1378), .S(n1341), .Z(n4565) );
  AND2_X1 U3116 ( .A1(n4497), .A2(n4348), .ZN(n4534) );
  MUX2_X1 U3117 ( .A(n4256), .B(n1447), .S(n1346), .Z(n2921) );
  MUX2_X1 U3118 ( .A(n4257), .B(n1444), .S(n1346), .Z(n2920) );
  MUX2_X1 U3119 ( .A(n4258), .B(n1441), .S(n1346), .Z(n2919) );
  MUX2_X1 U3120 ( .A(n4259), .B(n1438), .S(n1346), .Z(n2918) );
  MUX2_X1 U3121 ( .A(n4260), .B(n1435), .S(n1346), .Z(n2917) );
  MUX2_X1 U3122 ( .A(n4261), .B(n1432), .S(n1346), .Z(n2916) );
  MUX2_X1 U3123 ( .A(n4262), .B(n1429), .S(n1346), .Z(n2915) );
  MUX2_X1 U3124 ( .A(n4263), .B(n1426), .S(n1346), .Z(n2914) );
  MUX2_X1 U3125 ( .A(n4264), .B(n1423), .S(n1345), .Z(n2913) );
  MUX2_X1 U3126 ( .A(n4265), .B(n1421), .S(n1345), .Z(n2912) );
  MUX2_X1 U3127 ( .A(n4266), .B(n1419), .S(n1345), .Z(n2911) );
  MUX2_X1 U3128 ( .A(n4267), .B(n1417), .S(n1345), .Z(n2910) );
  MUX2_X1 U3129 ( .A(n4268), .B(n1415), .S(n1345), .Z(n2909) );
  MUX2_X1 U3130 ( .A(n4269), .B(n1413), .S(n1345), .Z(n2908) );
  MUX2_X1 U3131 ( .A(n4270), .B(n1411), .S(n1345), .Z(n2907) );
  MUX2_X1 U3132 ( .A(n4271), .B(n1409), .S(n1345), .Z(n2906) );
  MUX2_X1 U3133 ( .A(n4272), .B(n1407), .S(n1345), .Z(n2905) );
  MUX2_X1 U3134 ( .A(n4273), .B(n1405), .S(n1345), .Z(n2904) );
  MUX2_X1 U3135 ( .A(n4274), .B(n1403), .S(n1345), .Z(n2903) );
  MUX2_X1 U3136 ( .A(n4275), .B(n1401), .S(n1345), .Z(n2902) );
  MUX2_X1 U3137 ( .A(n4276), .B(n1399), .S(n1344), .Z(n2901) );
  MUX2_X1 U3138 ( .A(n4277), .B(n1397), .S(n1344), .Z(n2900) );
  MUX2_X1 U3139 ( .A(n4278), .B(n1395), .S(n1344), .Z(n2899) );
  MUX2_X1 U3140 ( .A(n4279), .B(n1393), .S(n1344), .Z(n2898) );
  MUX2_X1 U3141 ( .A(n4280), .B(n1391), .S(n1344), .Z(n2897) );
  MUX2_X1 U3142 ( .A(n4281), .B(n1389), .S(n1344), .Z(n2896) );
  MUX2_X1 U3143 ( .A(n4282), .B(n1387), .S(n1344), .Z(n2895) );
  MUX2_X1 U3144 ( .A(n4283), .B(n1385), .S(n1344), .Z(n2894) );
  MUX2_X1 U3145 ( .A(n4284), .B(n1383), .S(n1344), .Z(n2893) );
  MUX2_X1 U3146 ( .A(n4285), .B(n1381), .S(n1344), .Z(n2892) );
  MUX2_X1 U3147 ( .A(n4286), .B(n1379), .S(n1344), .Z(n2891) );
  MUX2_X1 U3148 ( .A(n4287), .B(n1377), .S(n1344), .Z(n2890) );
  AND2_X1 U3149 ( .A1(n4497), .A2(n4350), .ZN(n4566) );
  MUX2_X1 U3150 ( .A(n4915), .B(n1447), .S(n1349), .Z(n2889) );
  MUX2_X1 U3151 ( .A(n4914), .B(n1444), .S(n1349), .Z(n2888) );
  MUX2_X1 U3152 ( .A(n4913), .B(n1441), .S(n1349), .Z(n2887) );
  MUX2_X1 U3153 ( .A(n4912), .B(n1438), .S(n1349), .Z(n2886) );
  MUX2_X1 U3154 ( .A(n4911), .B(n1435), .S(n1349), .Z(n2885) );
  MUX2_X1 U3155 ( .A(n4910), .B(n1432), .S(n1349), .Z(n2884) );
  MUX2_X1 U3156 ( .A(n4909), .B(n1429), .S(n1349), .Z(n2883) );
  MUX2_X1 U3157 ( .A(n4908), .B(n1426), .S(n1349), .Z(n2882) );
  MUX2_X1 U3158 ( .A(n4907), .B(n1423), .S(n1348), .Z(n2881) );
  MUX2_X1 U3159 ( .A(n4906), .B(n1421), .S(n1348), .Z(n2880) );
  MUX2_X1 U3160 ( .A(n4905), .B(n1419), .S(n1348), .Z(n2879) );
  MUX2_X1 U3161 ( .A(n4904), .B(n1417), .S(n1348), .Z(n2878) );
  MUX2_X1 U3162 ( .A(n4903), .B(n1415), .S(n1348), .Z(n2877) );
  MUX2_X1 U3163 ( .A(n4902), .B(n1413), .S(n1348), .Z(n2876) );
  MUX2_X1 U3164 ( .A(n4901), .B(n1411), .S(n1348), .Z(n2875) );
  MUX2_X1 U3165 ( .A(n4900), .B(n1409), .S(n1348), .Z(n2874) );
  MUX2_X1 U3166 ( .A(n4899), .B(n1407), .S(n1348), .Z(n2873) );
  MUX2_X1 U3167 ( .A(n4898), .B(n1405), .S(n1348), .Z(n2872) );
  MUX2_X1 U3168 ( .A(n4897), .B(n1403), .S(n1348), .Z(n2871) );
  MUX2_X1 U3169 ( .A(n4896), .B(n1401), .S(n1348), .Z(n2870) );
  MUX2_X1 U3170 ( .A(n4895), .B(n1399), .S(n1347), .Z(n2869) );
  MUX2_X1 U3171 ( .A(n4894), .B(n1397), .S(n1347), .Z(n2868) );
  MUX2_X1 U3172 ( .A(n4893), .B(n1395), .S(n1347), .Z(n2867) );
  MUX2_X1 U3173 ( .A(n4892), .B(n1393), .S(n1347), .Z(n2866) );
  MUX2_X1 U3174 ( .A(n4891), .B(n1391), .S(n1347), .Z(n2865) );
  MUX2_X1 U3175 ( .A(n4890), .B(n1389), .S(n1347), .Z(n2864) );
  MUX2_X1 U3176 ( .A(n4889), .B(n1387), .S(n1347), .Z(n2863) );
  MUX2_X1 U3177 ( .A(n4888), .B(n1385), .S(n1347), .Z(n2862) );
  MUX2_X1 U3178 ( .A(n4887), .B(n1383), .S(n1347), .Z(n2861) );
  MUX2_X1 U3179 ( .A(n4886), .B(n1381), .S(n1347), .Z(n2860) );
  MUX2_X1 U3180 ( .A(n4885), .B(n1379), .S(n1347), .Z(n2859) );
  MUX2_X1 U3181 ( .A(n4884), .B(n1377), .S(n1347), .Z(n2858) );
  AND2_X1 U3182 ( .A1(n4497), .A2(n4352), .ZN(n4567) );
  MUX2_X1 U3183 ( .A(n4883), .B(n1447), .S(n1352), .Z(n2857) );
  MUX2_X1 U3184 ( .A(n4882), .B(n1444), .S(n1352), .Z(n2856) );
  MUX2_X1 U3185 ( .A(n4881), .B(n1441), .S(n1352), .Z(n2855) );
  MUX2_X1 U3186 ( .A(n4880), .B(n1438), .S(n1352), .Z(n2854) );
  MUX2_X1 U3187 ( .A(n4879), .B(n1435), .S(n1352), .Z(n2853) );
  MUX2_X1 U3188 ( .A(n4878), .B(n1432), .S(n1352), .Z(n2852) );
  MUX2_X1 U3189 ( .A(n4877), .B(n1429), .S(n1352), .Z(n2851) );
  MUX2_X1 U3190 ( .A(n4876), .B(n1426), .S(n1352), .Z(n2850) );
  MUX2_X1 U3191 ( .A(n4875), .B(n1423), .S(n1351), .Z(n2849) );
  MUX2_X1 U3192 ( .A(n4874), .B(n1421), .S(n1351), .Z(n2848) );
  MUX2_X1 U3193 ( .A(n4873), .B(n1419), .S(n1351), .Z(n2847) );
  MUX2_X1 U3194 ( .A(n4872), .B(n1417), .S(n1351), .Z(n2846) );
  MUX2_X1 U3195 ( .A(n4871), .B(n1415), .S(n1351), .Z(n2845) );
  MUX2_X1 U3196 ( .A(n4870), .B(n1413), .S(n1351), .Z(n2844) );
  MUX2_X1 U3197 ( .A(n4869), .B(n1411), .S(n1351), .Z(n2843) );
  MUX2_X1 U3198 ( .A(n4868), .B(n1409), .S(n1351), .Z(n2842) );
  MUX2_X1 U3199 ( .A(n4867), .B(n1407), .S(n1351), .Z(n2841) );
  MUX2_X1 U3200 ( .A(n4866), .B(n1405), .S(n1351), .Z(n2840) );
  MUX2_X1 U3201 ( .A(n4865), .B(n1403), .S(n1351), .Z(n2839) );
  MUX2_X1 U3202 ( .A(n4864), .B(n1401), .S(n1351), .Z(n2838) );
  MUX2_X1 U3203 ( .A(n4863), .B(n1399), .S(n1350), .Z(n2837) );
  MUX2_X1 U3204 ( .A(n4862), .B(n1397), .S(n1350), .Z(n2836) );
  MUX2_X1 U3205 ( .A(n4861), .B(n1395), .S(n1350), .Z(n2835) );
  MUX2_X1 U3206 ( .A(n4860), .B(n1393), .S(n1350), .Z(n2834) );
  MUX2_X1 U3207 ( .A(n4859), .B(n1391), .S(n1350), .Z(n2833) );
  MUX2_X1 U3208 ( .A(n4858), .B(n1389), .S(n1350), .Z(n2832) );
  MUX2_X1 U3209 ( .A(n4857), .B(n1387), .S(n1350), .Z(n2831) );
  MUX2_X1 U3210 ( .A(n4856), .B(n1385), .S(n1350), .Z(n2830) );
  MUX2_X1 U3211 ( .A(n4855), .B(n1383), .S(n1350), .Z(n2829) );
  MUX2_X1 U3212 ( .A(n4854), .B(n1381), .S(n1350), .Z(n2828) );
  MUX2_X1 U3213 ( .A(n4853), .B(n1379), .S(n1350), .Z(n2827) );
  MUX2_X1 U3214 ( .A(n4852), .B(n1377), .S(n1350), .Z(n2826) );
  AND2_X1 U3215 ( .A1(n4497), .A2(n4354), .ZN(n4568) );
  AND3_X1 U3216 ( .A1(n4357), .A2(n4355), .A3(ADD_WR[4]), .ZN(n4497) );
  MUX2_X1 U3217 ( .A(n4851), .B(n1447), .S(n1355), .Z(n2825) );
  MUX2_X1 U3218 ( .A(n4850), .B(n1444), .S(n1355), .Z(n2824) );
  MUX2_X1 U3219 ( .A(n4849), .B(n1441), .S(n1355), .Z(n2823) );
  MUX2_X1 U3220 ( .A(n4848), .B(n1438), .S(n1355), .Z(n2822) );
  MUX2_X1 U3221 ( .A(n4847), .B(n1435), .S(n1355), .Z(n2821) );
  MUX2_X1 U3222 ( .A(n4846), .B(n1432), .S(n1355), .Z(n2820) );
  MUX2_X1 U3223 ( .A(n4845), .B(n1429), .S(n1355), .Z(n2819) );
  MUX2_X1 U3224 ( .A(n4844), .B(n1426), .S(n1355), .Z(n2818) );
  MUX2_X1 U3225 ( .A(n4843), .B(n1423), .S(n1354), .Z(n2817) );
  MUX2_X1 U3226 ( .A(n4842), .B(n1421), .S(n1354), .Z(n2816) );
  MUX2_X1 U3227 ( .A(n4841), .B(n1419), .S(n1354), .Z(n2815) );
  MUX2_X1 U3228 ( .A(n4840), .B(n1417), .S(n1354), .Z(n2814) );
  MUX2_X1 U3229 ( .A(n4839), .B(n1415), .S(n1354), .Z(n2813) );
  MUX2_X1 U3230 ( .A(n4838), .B(n1413), .S(n1354), .Z(n2812) );
  MUX2_X1 U3231 ( .A(n4837), .B(n1411), .S(n1354), .Z(n2811) );
  MUX2_X1 U3232 ( .A(n4836), .B(n1409), .S(n1354), .Z(n2810) );
  MUX2_X1 U3233 ( .A(n4835), .B(n1407), .S(n1354), .Z(n2809) );
  MUX2_X1 U3234 ( .A(n4834), .B(n1405), .S(n1354), .Z(n2808) );
  MUX2_X1 U3235 ( .A(n4833), .B(n1403), .S(n1354), .Z(n2807) );
  MUX2_X1 U3236 ( .A(n4832), .B(n1401), .S(n1354), .Z(n2806) );
  MUX2_X1 U3237 ( .A(n4831), .B(n1399), .S(n1353), .Z(n2805) );
  MUX2_X1 U3238 ( .A(n4830), .B(n1397), .S(n1353), .Z(n2804) );
  MUX2_X1 U3239 ( .A(n4829), .B(n1395), .S(n1353), .Z(n2803) );
  MUX2_X1 U3240 ( .A(n4828), .B(n1393), .S(n1353), .Z(n2802) );
  MUX2_X1 U3241 ( .A(n4827), .B(n1391), .S(n1353), .Z(n2801) );
  MUX2_X1 U3242 ( .A(n4826), .B(n1389), .S(n1353), .Z(n2800) );
  MUX2_X1 U3243 ( .A(n4825), .B(n1387), .S(n1353), .Z(n2799) );
  MUX2_X1 U3244 ( .A(n4824), .B(n1385), .S(n1353), .Z(n2798) );
  MUX2_X1 U3245 ( .A(n4823), .B(n1383), .S(n1353), .Z(n2797) );
  MUX2_X1 U3246 ( .A(n4822), .B(n1381), .S(n1353), .Z(n2796) );
  MUX2_X1 U3247 ( .A(n4821), .B(n1379), .S(n1353), .Z(n2795) );
  MUX2_X1 U3248 ( .A(n4820), .B(n1377), .S(n1353), .Z(n2794) );
  AND2_X1 U3249 ( .A1(n4570), .A2(n4392), .ZN(n4569) );
  MUX2_X1 U3250 ( .A(n4819), .B(n1447), .S(n1358), .Z(n2793) );
  MUX2_X1 U3251 ( .A(n4818), .B(n1444), .S(n1358), .Z(n2792) );
  MUX2_X1 U3252 ( .A(n4817), .B(n1441), .S(n1358), .Z(n2791) );
  MUX2_X1 U3253 ( .A(n4816), .B(n1438), .S(n1358), .Z(n2790) );
  MUX2_X1 U3254 ( .A(n4815), .B(n1435), .S(n1358), .Z(n2789) );
  MUX2_X1 U3255 ( .A(n4814), .B(n1432), .S(n1358), .Z(n2788) );
  MUX2_X1 U3256 ( .A(n4813), .B(n1429), .S(n1358), .Z(n2787) );
  MUX2_X1 U3257 ( .A(n4812), .B(n1426), .S(n1358), .Z(n2786) );
  MUX2_X1 U3258 ( .A(n4811), .B(n1423), .S(n1357), .Z(n2785) );
  MUX2_X1 U3259 ( .A(n4810), .B(n1421), .S(n1357), .Z(n2784) );
  MUX2_X1 U3260 ( .A(n4809), .B(n1419), .S(n1357), .Z(n2783) );
  MUX2_X1 U3261 ( .A(n4808), .B(n1417), .S(n1357), .Z(n2782) );
  MUX2_X1 U3262 ( .A(n4807), .B(n1415), .S(n1357), .Z(n2781) );
  MUX2_X1 U3263 ( .A(n4806), .B(n1413), .S(n1357), .Z(n2780) );
  MUX2_X1 U3264 ( .A(n4805), .B(n1411), .S(n1357), .Z(n2779) );
  MUX2_X1 U3265 ( .A(n4804), .B(n1409), .S(n1357), .Z(n2778) );
  MUX2_X1 U3266 ( .A(n4803), .B(n1407), .S(n1357), .Z(n2777) );
  MUX2_X1 U3267 ( .A(n4802), .B(n1405), .S(n1357), .Z(n2776) );
  MUX2_X1 U3268 ( .A(n4801), .B(n1403), .S(n1357), .Z(n2775) );
  MUX2_X1 U3269 ( .A(n4800), .B(n1401), .S(n1357), .Z(n2774) );
  MUX2_X1 U3270 ( .A(n4799), .B(n1399), .S(n1356), .Z(n2773) );
  MUX2_X1 U3271 ( .A(n4798), .B(n1397), .S(n1356), .Z(n2772) );
  MUX2_X1 U3272 ( .A(n4797), .B(n1395), .S(n1356), .Z(n2771) );
  MUX2_X1 U3273 ( .A(n4796), .B(n1393), .S(n1356), .Z(n2770) );
  MUX2_X1 U3274 ( .A(n4795), .B(n1391), .S(n1356), .Z(n2769) );
  MUX2_X1 U3275 ( .A(n4794), .B(n1389), .S(n1356), .Z(n2768) );
  MUX2_X1 U3276 ( .A(n4793), .B(n1387), .S(n1356), .Z(n2767) );
  MUX2_X1 U3277 ( .A(n4792), .B(n1385), .S(n1356), .Z(n2766) );
  MUX2_X1 U3278 ( .A(n4791), .B(n1383), .S(n1356), .Z(n2765) );
  MUX2_X1 U3279 ( .A(n4790), .B(n1381), .S(n1356), .Z(n2764) );
  MUX2_X1 U3280 ( .A(n4789), .B(n1379), .S(n1356), .Z(n2763) );
  MUX2_X1 U3281 ( .A(n4788), .B(n1377), .S(n1356), .Z(n2762) );
  AND2_X1 U3282 ( .A1(n4570), .A2(n4341), .ZN(n4571) );
  NOR3_X1 U3283 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(n4572), .ZN(n4341) );
  MUX2_X1 U3284 ( .A(n4288), .B(n1447), .S(n1361), .Z(n2761) );
  MUX2_X1 U3285 ( .A(n4289), .B(n1444), .S(n1361), .Z(n2760) );
  MUX2_X1 U3286 ( .A(n4290), .B(n1441), .S(n1361), .Z(n2759) );
  MUX2_X1 U3287 ( .A(n4291), .B(n1438), .S(n1361), .Z(n2758) );
  MUX2_X1 U3288 ( .A(n4292), .B(n1435), .S(n1361), .Z(n2757) );
  MUX2_X1 U3289 ( .A(n4293), .B(n1432), .S(n1361), .Z(n2756) );
  MUX2_X1 U3290 ( .A(n4294), .B(n1429), .S(n1361), .Z(n2755) );
  MUX2_X1 U3291 ( .A(n4295), .B(n1426), .S(n1361), .Z(n2754) );
  MUX2_X1 U3292 ( .A(n4296), .B(n1423), .S(n1360), .Z(n2753) );
  MUX2_X1 U3293 ( .A(n4297), .B(n1421), .S(n1360), .Z(n2752) );
  MUX2_X1 U3294 ( .A(n224), .B(n1419), .S(n1360), .Z(n2751) );
  MUX2_X1 U3295 ( .A(n4298), .B(n1417), .S(n1360), .Z(n2750) );
  MUX2_X1 U3296 ( .A(n343), .B(n1415), .S(n1360), .Z(n2749) );
  MUX2_X1 U3297 ( .A(n344), .B(n1413), .S(n1360), .Z(n2748) );
  MUX2_X1 U3298 ( .A(n225), .B(n1411), .S(n1360), .Z(n2747) );
  MUX2_X1 U3299 ( .A(n4299), .B(n1409), .S(n1360), .Z(n2746) );
  MUX2_X1 U3300 ( .A(n345), .B(n1407), .S(n1360), .Z(n2745) );
  MUX2_X1 U3301 ( .A(n4300), .B(n1405), .S(n1360), .Z(n2744) );
  MUX2_X1 U3302 ( .A(n4301), .B(n1403), .S(n1360), .Z(n2743) );
  MUX2_X1 U3303 ( .A(n346), .B(n1401), .S(n1360), .Z(n2742) );
  MUX2_X1 U3304 ( .A(n4302), .B(n1399), .S(n1359), .Z(n2741) );
  MUX2_X1 U3305 ( .A(n226), .B(n1397), .S(n1359), .Z(n2740) );
  MUX2_X1 U3306 ( .A(n4303), .B(n1395), .S(n1359), .Z(n2739) );
  MUX2_X1 U3307 ( .A(n347), .B(n1393), .S(n1359), .Z(n2738) );
  MUX2_X1 U3308 ( .A(n4304), .B(n1391), .S(n1359), .Z(n2737) );
  MUX2_X1 U3309 ( .A(n4305), .B(n1389), .S(n1359), .Z(n2736) );
  MUX2_X1 U3310 ( .A(n351), .B(n1387), .S(n1359), .Z(n2735) );
  MUX2_X1 U3311 ( .A(n348), .B(n1385), .S(n1359), .Z(n2734) );
  MUX2_X1 U3312 ( .A(n349), .B(n1383), .S(n1359), .Z(n2733) );
  MUX2_X1 U3313 ( .A(n4306), .B(n1381), .S(n1359), .Z(n2732) );
  MUX2_X1 U3314 ( .A(n350), .B(n1379), .S(n1359), .Z(n2731) );
  MUX2_X1 U3315 ( .A(n4307), .B(n1377), .S(n1359), .Z(n2730) );
  AND2_X1 U3316 ( .A1(n4570), .A2(n4344), .ZN(n4573) );
  NOR3_X1 U3317 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(n4574), .ZN(n4344) );
  INV_X1 U3318 ( .A(n4575), .ZN(n2729) );
  MUX2_X1 U3319 ( .A(n837), .B(n1448), .S(n1364), .Z(n4575) );
  INV_X1 U3320 ( .A(n4577), .ZN(n2728) );
  MUX2_X1 U3321 ( .A(n838), .B(n1445), .S(n1364), .Z(n4577) );
  INV_X1 U3322 ( .A(n4578), .ZN(n2727) );
  MUX2_X1 U3323 ( .A(n839), .B(n1442), .S(n1364), .Z(n4578) );
  INV_X1 U3324 ( .A(n4579), .ZN(n2726) );
  MUX2_X1 U3325 ( .A(n840), .B(n1439), .S(n1364), .Z(n4579) );
  INV_X1 U3326 ( .A(n4580), .ZN(n2725) );
  MUX2_X1 U3327 ( .A(n841), .B(n1436), .S(n1364), .Z(n4580) );
  INV_X1 U3328 ( .A(n4581), .ZN(n2724) );
  MUX2_X1 U3329 ( .A(n842), .B(n1433), .S(n1364), .Z(n4581) );
  INV_X1 U3330 ( .A(n4582), .ZN(n2723) );
  MUX2_X1 U3331 ( .A(n843), .B(n1430), .S(n1364), .Z(n4582) );
  INV_X1 U3332 ( .A(n4583), .ZN(n2722) );
  MUX2_X1 U3333 ( .A(n844), .B(n1427), .S(n1364), .Z(n4583) );
  INV_X1 U3334 ( .A(n4584), .ZN(n2721) );
  MUX2_X1 U3335 ( .A(n845), .B(n1424), .S(n1363), .Z(n4584) );
  INV_X1 U3336 ( .A(n4585), .ZN(n2720) );
  MUX2_X1 U3337 ( .A(n846), .B(n1422), .S(n1363), .Z(n4585) );
  INV_X1 U3338 ( .A(n4586), .ZN(n2719) );
  MUX2_X1 U3339 ( .A(n847), .B(n1420), .S(n1363), .Z(n4586) );
  INV_X1 U3340 ( .A(n4587), .ZN(n2718) );
  MUX2_X1 U3341 ( .A(n848), .B(n1418), .S(n1363), .Z(n4587) );
  INV_X1 U3342 ( .A(n4588), .ZN(n2717) );
  MUX2_X1 U3343 ( .A(n849), .B(n1416), .S(n1363), .Z(n4588) );
  INV_X1 U3344 ( .A(n4589), .ZN(n2716) );
  MUX2_X1 U3345 ( .A(n850), .B(n1414), .S(n1363), .Z(n4589) );
  INV_X1 U3346 ( .A(n4590), .ZN(n2715) );
  MUX2_X1 U3347 ( .A(n851), .B(n1412), .S(n1363), .Z(n4590) );
  INV_X1 U3348 ( .A(n4591), .ZN(n2714) );
  MUX2_X1 U3349 ( .A(n852), .B(n1410), .S(n1363), .Z(n4591) );
  INV_X1 U3350 ( .A(n4592), .ZN(n2713) );
  MUX2_X1 U3351 ( .A(n853), .B(n1408), .S(n1363), .Z(n4592) );
  INV_X1 U3352 ( .A(n4593), .ZN(n2712) );
  MUX2_X1 U3353 ( .A(n854), .B(n1406), .S(n1363), .Z(n4593) );
  INV_X1 U3354 ( .A(n4594), .ZN(n2711) );
  MUX2_X1 U3355 ( .A(n855), .B(n1404), .S(n1363), .Z(n4594) );
  INV_X1 U3356 ( .A(n4595), .ZN(n2710) );
  MUX2_X1 U3357 ( .A(n856), .B(n1402), .S(n1363), .Z(n4595) );
  INV_X1 U3358 ( .A(n4596), .ZN(n2709) );
  MUX2_X1 U3359 ( .A(n857), .B(n1400), .S(n1362), .Z(n4596) );
  INV_X1 U3360 ( .A(n4597), .ZN(n2708) );
  MUX2_X1 U3361 ( .A(n858), .B(n1398), .S(n1362), .Z(n4597) );
  INV_X1 U3362 ( .A(n4598), .ZN(n2707) );
  MUX2_X1 U3363 ( .A(n859), .B(n1396), .S(n1362), .Z(n4598) );
  INV_X1 U3364 ( .A(n4599), .ZN(n2706) );
  MUX2_X1 U3365 ( .A(n860), .B(n1394), .S(n1362), .Z(n4599) );
  INV_X1 U3366 ( .A(n4600), .ZN(n2705) );
  MUX2_X1 U3367 ( .A(n861), .B(n1392), .S(n1362), .Z(n4600) );
  INV_X1 U3368 ( .A(n4601), .ZN(n2704) );
  MUX2_X1 U3369 ( .A(n862), .B(n1390), .S(n1362), .Z(n4601) );
  INV_X1 U3370 ( .A(n4602), .ZN(n2703) );
  MUX2_X1 U3371 ( .A(n863), .B(n1388), .S(n1362), .Z(n4602) );
  INV_X1 U3372 ( .A(n4603), .ZN(n2702) );
  MUX2_X1 U3373 ( .A(n864), .B(n1386), .S(n1362), .Z(n4603) );
  INV_X1 U3374 ( .A(n4604), .ZN(n2701) );
  MUX2_X1 U3375 ( .A(n865), .B(n1384), .S(n1362), .Z(n4604) );
  INV_X1 U3376 ( .A(n4605), .ZN(n2700) );
  MUX2_X1 U3377 ( .A(n866), .B(n1382), .S(n1362), .Z(n4605) );
  INV_X1 U3378 ( .A(n4606), .ZN(n2699) );
  MUX2_X1 U3379 ( .A(n867), .B(n1380), .S(n1362), .Z(n4606) );
  INV_X1 U3380 ( .A(n4607), .ZN(n2698) );
  MUX2_X1 U3381 ( .A(n868), .B(n1378), .S(n1362), .Z(n4607) );
  AND2_X1 U3382 ( .A1(n4570), .A2(n4346), .ZN(n4576) );
  NOR3_X1 U3383 ( .A1(n4572), .A2(ADD_WR[2]), .A3(n4574), .ZN(n4346) );
  MUX2_X1 U3384 ( .A(n4787), .B(n1447), .S(n1367), .Z(n2697) );
  MUX2_X1 U3385 ( .A(n4786), .B(n1444), .S(n1367), .Z(n2696) );
  MUX2_X1 U3386 ( .A(n4785), .B(n1441), .S(n1367), .Z(n2695) );
  MUX2_X1 U3387 ( .A(n4784), .B(n1438), .S(n1367), .Z(n2694) );
  MUX2_X1 U3388 ( .A(n4783), .B(n1435), .S(n1367), .Z(n2693) );
  MUX2_X1 U3389 ( .A(n4782), .B(n1432), .S(n1367), .Z(n2692) );
  MUX2_X1 U3390 ( .A(n4781), .B(n1429), .S(n1367), .Z(n2691) );
  MUX2_X1 U3391 ( .A(n4780), .B(n1426), .S(n1367), .Z(n2690) );
  MUX2_X1 U3392 ( .A(n4779), .B(n1423), .S(n1366), .Z(n2689) );
  MUX2_X1 U3393 ( .A(n4778), .B(n1421), .S(n1366), .Z(n2688) );
  MUX2_X1 U3394 ( .A(n4777), .B(n1419), .S(n1366), .Z(n2687) );
  MUX2_X1 U3395 ( .A(n4776), .B(n1417), .S(n1366), .Z(n2686) );
  MUX2_X1 U3396 ( .A(n4775), .B(n1415), .S(n1366), .Z(n2685) );
  MUX2_X1 U3397 ( .A(n4774), .B(n1413), .S(n1366), .Z(n2684) );
  MUX2_X1 U3398 ( .A(n4773), .B(n1411), .S(n1366), .Z(n2683) );
  MUX2_X1 U3399 ( .A(n4772), .B(n1409), .S(n1366), .Z(n2682) );
  MUX2_X1 U3400 ( .A(n4771), .B(n1407), .S(n1366), .Z(n2681) );
  MUX2_X1 U3401 ( .A(n4770), .B(n1405), .S(n1366), .Z(n2680) );
  MUX2_X1 U3402 ( .A(n4769), .B(n1403), .S(n1366), .Z(n2679) );
  MUX2_X1 U3403 ( .A(n4768), .B(n1401), .S(n1366), .Z(n2678) );
  MUX2_X1 U3404 ( .A(n4767), .B(n1399), .S(n1365), .Z(n2677) );
  MUX2_X1 U3405 ( .A(n4766), .B(n1397), .S(n1365), .Z(n2676) );
  MUX2_X1 U3406 ( .A(n4765), .B(n1395), .S(n1365), .Z(n2675) );
  MUX2_X1 U3407 ( .A(n4764), .B(n1393), .S(n1365), .Z(n2674) );
  MUX2_X1 U3408 ( .A(n4763), .B(n1391), .S(n1365), .Z(n2673) );
  MUX2_X1 U3409 ( .A(n4762), .B(n1389), .S(n1365), .Z(n2672) );
  MUX2_X1 U3410 ( .A(n4761), .B(n1387), .S(n1365), .Z(n2671) );
  MUX2_X1 U3411 ( .A(n4760), .B(n1385), .S(n1365), .Z(n2670) );
  MUX2_X1 U3412 ( .A(n4759), .B(n1383), .S(n1365), .Z(n2669) );
  MUX2_X1 U3413 ( .A(n4758), .B(n1381), .S(n1365), .Z(n2668) );
  MUX2_X1 U3414 ( .A(n4757), .B(n1379), .S(n1365), .Z(n2667) );
  MUX2_X1 U3415 ( .A(n4756), .B(n1377), .S(n1365), .Z(n2666) );
  AND2_X1 U3416 ( .A1(n4570), .A2(n4348), .ZN(n4608) );
  AND3_X1 U3417 ( .A1(n4572), .A2(n4574), .A3(ADD_WR[2]), .ZN(n4348) );
  MUX2_X1 U3418 ( .A(n4755), .B(n1447), .S(n1370), .Z(n2665) );
  MUX2_X1 U3419 ( .A(n4754), .B(n1444), .S(n1370), .Z(n2664) );
  MUX2_X1 U3420 ( .A(n4753), .B(n1441), .S(n1370), .Z(n2663) );
  MUX2_X1 U3421 ( .A(n4752), .B(n1438), .S(n1370), .Z(n2662) );
  MUX2_X1 U3422 ( .A(n4751), .B(n1435), .S(n1370), .Z(n2661) );
  MUX2_X1 U3423 ( .A(n4750), .B(n1432), .S(n1370), .Z(n2660) );
  MUX2_X1 U3424 ( .A(n4749), .B(n1429), .S(n1370), .Z(n2659) );
  MUX2_X1 U3425 ( .A(n4748), .B(n1426), .S(n1370), .Z(n2658) );
  MUX2_X1 U3426 ( .A(n4747), .B(n1423), .S(n1369), .Z(n2657) );
  MUX2_X1 U3427 ( .A(n4746), .B(n1421), .S(n1369), .Z(n2656) );
  MUX2_X1 U3428 ( .A(n4745), .B(n1419), .S(n1369), .Z(n2655) );
  MUX2_X1 U3429 ( .A(n4744), .B(n1417), .S(n1369), .Z(n2654) );
  MUX2_X1 U3430 ( .A(n4743), .B(n1415), .S(n1369), .Z(n2653) );
  MUX2_X1 U3431 ( .A(n4742), .B(n1413), .S(n1369), .Z(n2652) );
  MUX2_X1 U3432 ( .A(n4741), .B(n1411), .S(n1369), .Z(n2651) );
  MUX2_X1 U3433 ( .A(n4740), .B(n1409), .S(n1369), .Z(n2650) );
  MUX2_X1 U3434 ( .A(n4739), .B(n1407), .S(n1369), .Z(n2649) );
  MUX2_X1 U3435 ( .A(n4738), .B(n1405), .S(n1369), .Z(n2648) );
  MUX2_X1 U3436 ( .A(n4737), .B(n1403), .S(n1369), .Z(n2647) );
  MUX2_X1 U3437 ( .A(n4736), .B(n1401), .S(n1369), .Z(n2646) );
  MUX2_X1 U3438 ( .A(n4735), .B(n1399), .S(n1368), .Z(n2645) );
  MUX2_X1 U3439 ( .A(n4734), .B(n1397), .S(n1368), .Z(n2644) );
  MUX2_X1 U3440 ( .A(n4733), .B(n1395), .S(n1368), .Z(n2643) );
  MUX2_X1 U3441 ( .A(n4732), .B(n1393), .S(n1368), .Z(n2642) );
  MUX2_X1 U3442 ( .A(n4731), .B(n1391), .S(n1368), .Z(n2641) );
  MUX2_X1 U3443 ( .A(n4730), .B(n1389), .S(n1368), .Z(n2640) );
  MUX2_X1 U3444 ( .A(n4729), .B(n1387), .S(n1368), .Z(n2639) );
  MUX2_X1 U3445 ( .A(n4728), .B(n1385), .S(n1368), .Z(n2638) );
  MUX2_X1 U3446 ( .A(n4727), .B(n1383), .S(n1368), .Z(n2637) );
  MUX2_X1 U3447 ( .A(n4726), .B(n1381), .S(n1368), .Z(n2636) );
  MUX2_X1 U3448 ( .A(n4725), .B(n1379), .S(n1368), .Z(n2635) );
  MUX2_X1 U3449 ( .A(n4724), .B(n1377), .S(n1368), .Z(n2634) );
  AND2_X1 U3450 ( .A1(n4570), .A2(n4350), .ZN(n4609) );
  AND3_X1 U3451 ( .A1(ADD_WR[0]), .A2(n4574), .A3(ADD_WR[2]), .ZN(n4350) );
  INV_X1 U3452 ( .A(n4610), .ZN(n2633) );
  MUX2_X1 U3453 ( .A(n933), .B(n1448), .S(n1373), .Z(n4610) );
  INV_X1 U3454 ( .A(n4612), .ZN(n2632) );
  MUX2_X1 U3455 ( .A(n934), .B(n1445), .S(n1373), .Z(n4612) );
  INV_X1 U3456 ( .A(n4613), .ZN(n2631) );
  MUX2_X1 U3457 ( .A(n935), .B(n1442), .S(n1373), .Z(n4613) );
  INV_X1 U3458 ( .A(n4614), .ZN(n2630) );
  MUX2_X1 U3459 ( .A(n936), .B(n1439), .S(n1373), .Z(n4614) );
  INV_X1 U3460 ( .A(n4615), .ZN(n2629) );
  MUX2_X1 U3461 ( .A(n937), .B(n1436), .S(n1373), .Z(n4615) );
  INV_X1 U3462 ( .A(n4616), .ZN(n2628) );
  MUX2_X1 U3463 ( .A(n938), .B(n1433), .S(n1373), .Z(n4616) );
  INV_X1 U3464 ( .A(n4617), .ZN(n2627) );
  MUX2_X1 U3465 ( .A(n939), .B(n1430), .S(n1373), .Z(n4617) );
  INV_X1 U3466 ( .A(n4618), .ZN(n2626) );
  MUX2_X1 U3467 ( .A(n940), .B(n1427), .S(n1373), .Z(n4618) );
  INV_X1 U3468 ( .A(n4619), .ZN(n2625) );
  MUX2_X1 U3469 ( .A(n941), .B(n1424), .S(n1372), .Z(n4619) );
  INV_X1 U3470 ( .A(n4620), .ZN(n2624) );
  MUX2_X1 U3471 ( .A(n942), .B(n1422), .S(n1372), .Z(n4620) );
  INV_X1 U3472 ( .A(n4621), .ZN(n2623) );
  MUX2_X1 U3473 ( .A(n943), .B(n1420), .S(n1372), .Z(n4621) );
  INV_X1 U3474 ( .A(n4622), .ZN(n2622) );
  MUX2_X1 U3475 ( .A(n944), .B(n1418), .S(n1372), .Z(n4622) );
  INV_X1 U3476 ( .A(n4623), .ZN(n2621) );
  MUX2_X1 U3477 ( .A(n945), .B(n1416), .S(n1372), .Z(n4623) );
  INV_X1 U3478 ( .A(n4624), .ZN(n2620) );
  MUX2_X1 U3479 ( .A(n946), .B(n1414), .S(n1372), .Z(n4624) );
  INV_X1 U3480 ( .A(n4625), .ZN(n2619) );
  MUX2_X1 U3481 ( .A(n947), .B(n1412), .S(n1372), .Z(n4625) );
  INV_X1 U3482 ( .A(n4626), .ZN(n2618) );
  MUX2_X1 U3483 ( .A(n948), .B(n1410), .S(n1372), .Z(n4626) );
  INV_X1 U3484 ( .A(n4627), .ZN(n2617) );
  MUX2_X1 U3485 ( .A(n949), .B(n1408), .S(n1372), .Z(n4627) );
  INV_X1 U3486 ( .A(n4628), .ZN(n2616) );
  MUX2_X1 U3487 ( .A(n950), .B(n1406), .S(n1372), .Z(n4628) );
  INV_X1 U3488 ( .A(n4629), .ZN(n2615) );
  MUX2_X1 U3489 ( .A(n951), .B(n1404), .S(n1372), .Z(n4629) );
  INV_X1 U3490 ( .A(n4630), .ZN(n2614) );
  MUX2_X1 U3491 ( .A(n952), .B(n1402), .S(n1372), .Z(n4630) );
  INV_X1 U3492 ( .A(n4631), .ZN(n2613) );
  MUX2_X1 U3493 ( .A(n953), .B(n1400), .S(n1371), .Z(n4631) );
  INV_X1 U3494 ( .A(n4632), .ZN(n2612) );
  MUX2_X1 U3495 ( .A(n954), .B(n1398), .S(n1371), .Z(n4632) );
  INV_X1 U3496 ( .A(n4633), .ZN(n2611) );
  MUX2_X1 U3497 ( .A(n955), .B(n1396), .S(n1371), .Z(n4633) );
  INV_X1 U3498 ( .A(n4634), .ZN(n2610) );
  MUX2_X1 U3499 ( .A(n956), .B(n1394), .S(n1371), .Z(n4634) );
  INV_X1 U3500 ( .A(n4635), .ZN(n2609) );
  MUX2_X1 U3501 ( .A(n957), .B(n1392), .S(n1371), .Z(n4635) );
  INV_X1 U3502 ( .A(n4636), .ZN(n2608) );
  MUX2_X1 U3503 ( .A(n958), .B(n1390), .S(n1371), .Z(n4636) );
  INV_X1 U3504 ( .A(n4637), .ZN(n2607) );
  MUX2_X1 U3505 ( .A(n959), .B(n1388), .S(n1371), .Z(n4637) );
  INV_X1 U3506 ( .A(n4638), .ZN(n2606) );
  MUX2_X1 U3507 ( .A(n960), .B(n1386), .S(n1371), .Z(n4638) );
  INV_X1 U3508 ( .A(n4639), .ZN(n2605) );
  MUX2_X1 U3509 ( .A(n961), .B(n1384), .S(n1371), .Z(n4639) );
  INV_X1 U3510 ( .A(n4640), .ZN(n2604) );
  MUX2_X1 U3511 ( .A(n962), .B(n1382), .S(n1371), .Z(n4640) );
  INV_X1 U3512 ( .A(n4641), .ZN(n2603) );
  MUX2_X1 U3513 ( .A(n963), .B(n1380), .S(n1371), .Z(n4641) );
  INV_X1 U3514 ( .A(n4642), .ZN(n2602) );
  MUX2_X1 U3515 ( .A(n964), .B(n1378), .S(n1371), .Z(n4642) );
  AND2_X1 U3516 ( .A1(n4570), .A2(n4352), .ZN(n4611) );
  AND3_X1 U3517 ( .A1(ADD_WR[1]), .A2(n4572), .A3(ADD_WR[2]), .ZN(n4352) );
  MUX2_X1 U3518 ( .A(n4308), .B(n1446), .S(n1376), .Z(n2601) );
  MUX2_X1 U3519 ( .A(n4309), .B(n1443), .S(n1376), .Z(n2600) );
  MUX2_X1 U3520 ( .A(n4310), .B(n1440), .S(n1376), .Z(n2599) );
  MUX2_X1 U3521 ( .A(n4311), .B(n1437), .S(n1376), .Z(n2598) );
  MUX2_X1 U3522 ( .A(n4312), .B(n1434), .S(n1376), .Z(n2597) );
  MUX2_X1 U3523 ( .A(n4313), .B(n1431), .S(n1376), .Z(n2596) );
  MUX2_X1 U3524 ( .A(n4314), .B(n1428), .S(n1376), .Z(n2595) );
  MUX2_X1 U3525 ( .A(n4315), .B(n1425), .S(n1376), .Z(n2594) );
  MUX2_X1 U3526 ( .A(n4316), .B(n1423), .S(n1375), .Z(n2593) );
  MUX2_X1 U3527 ( .A(n4317), .B(n1421), .S(n1375), .Z(n2592) );
  MUX2_X1 U3528 ( .A(n4318), .B(n1419), .S(n1375), .Z(n2591) );
  MUX2_X1 U3529 ( .A(n4319), .B(n1417), .S(n1375), .Z(n2590) );
  MUX2_X1 U3530 ( .A(n4320), .B(n1415), .S(n1375), .Z(n2589) );
  MUX2_X1 U3531 ( .A(n4321), .B(n1413), .S(n1375), .Z(n2588) );
  MUX2_X1 U3532 ( .A(n4322), .B(n1411), .S(n1375), .Z(n2587) );
  MUX2_X1 U3533 ( .A(n4323), .B(n1409), .S(n1375), .Z(n2586) );
  MUX2_X1 U3534 ( .A(n4324), .B(n1407), .S(n1375), .Z(n2585) );
  MUX2_X1 U3535 ( .A(n4325), .B(n1405), .S(n1375), .Z(n2584) );
  MUX2_X1 U3536 ( .A(n4326), .B(n1403), .S(n1375), .Z(n2583) );
  MUX2_X1 U3537 ( .A(n4327), .B(n1401), .S(n1375), .Z(n2582) );
  MUX2_X1 U3538 ( .A(n4328), .B(n1399), .S(n1374), .Z(n2581) );
  MUX2_X1 U3539 ( .A(n4329), .B(n1397), .S(n1374), .Z(n2580) );
  MUX2_X1 U3540 ( .A(n4330), .B(n1395), .S(n1374), .Z(n2579) );
  MUX2_X1 U3541 ( .A(n4331), .B(n1393), .S(n1374), .Z(n2578) );
  MUX2_X1 U3542 ( .A(n4332), .B(n1391), .S(n1374), .Z(n2577) );
  MUX2_X1 U3543 ( .A(n4333), .B(n1389), .S(n1374), .Z(n2576) );
  MUX2_X1 U3544 ( .A(n4334), .B(n1387), .S(n1374), .Z(n2575) );
  MUX2_X1 U3545 ( .A(n4335), .B(n1385), .S(n1374), .Z(n2574) );
  MUX2_X1 U3546 ( .A(n4336), .B(n1383), .S(n1374), .Z(n2573) );
  MUX2_X1 U3547 ( .A(n4337), .B(n1381), .S(n1374), .Z(n2572) );
  MUX2_X1 U3548 ( .A(n4338), .B(n1379), .S(n1374), .Z(n2571) );
  MUX2_X1 U3549 ( .A(n4339), .B(n1377), .S(n1374), .Z(n2570) );
  AND2_X1 U3550 ( .A1(n4570), .A2(n4354), .ZN(n4643) );
  AND3_X1 U3551 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(ADD_WR[2]), .ZN(n4354)
         );
  AND3_X1 U3552 ( .A1(ADD_WR[3]), .A2(n4357), .A3(ADD_WR[4]), .ZN(n4570) );
  NOR2_X1 U3553 ( .A1(n4644), .A2(n4645), .ZN(n4357) );
  INV_X1 U3554 ( .A(ENABLE), .ZN(n4644) );
  XNOR2_X1 U3555 ( .A(ADD_RS2[1]), .B(n4574), .ZN(n4651) );
  XNOR2_X1 U3556 ( .A(ADD_RS2[0]), .B(n4572), .ZN(n4650) );
  XNOR2_X1 U3557 ( .A(ADD_RS2[3]), .B(ADD_WR[3]), .ZN(n4648) );
  XNOR2_X1 U3558 ( .A(ADD_RS2[4]), .B(ADD_WR[4]), .ZN(n4647) );
  XNOR2_X1 U3559 ( .A(ADD_RS2[2]), .B(ADD_WR[2]), .ZN(n4646) );
  XNOR2_X1 U3560 ( .A(n4574), .B(n784), .ZN(n4657) );
  INV_X1 U3561 ( .A(ADD_WR[1]), .ZN(n4574) );
  OAI21_X1 U3562 ( .B1(n4658), .B2(n4659), .A(WR), .ZN(n4645) );
  NAND2_X1 U3563 ( .A1(n4355), .A2(n4356), .ZN(n4659) );
  INV_X1 U3564 ( .A(ADD_WR[4]), .ZN(n4356) );
  INV_X1 U3565 ( .A(ADD_WR[3]), .ZN(n4355) );
  INV_X1 U3566 ( .A(n4392), .ZN(n4658) );
  NOR3_X1 U3567 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(ADD_WR[0]), .ZN(n4392)
         );
  XNOR2_X1 U3568 ( .A(ADD_RS1[0]), .B(n4572), .ZN(n4656) );
  INV_X1 U3569 ( .A(ADD_WR[0]), .ZN(n4572) );
  XNOR2_X1 U3570 ( .A(n84), .B(ADD_WR[3]), .ZN(n4654) );
  XNOR2_X1 U3571 ( .A(n1092), .B(ADD_WR[4]), .ZN(n4653) );
  XNOR2_X1 U3572 ( .A(n764), .B(ADD_WR[2]), .ZN(n4652) );
endmodule


module Decode ( CLK, RST, Bubble, RF_WE, ZERO_FLAG, PC_IN, INS_IN, ADD_WR, 
        DATA_WR_IN, PC_OUT, A_OUT, B_OUT, IMM_OUT, ADD_RS1_HDU, ADD_RS2_HDU, 
        ADD_WR_OUT, ADD_RS1_OUT, ADD_RS2_OUT );
  input [31:0] PC_IN;
  input [31:0] INS_IN;
  input [4:0] ADD_WR;
  input [31:0] DATA_WR_IN;
  output [31:0] PC_OUT;
  output [31:0] A_OUT;
  output [31:0] B_OUT;
  output [31:0] IMM_OUT;
  output [4:0] ADD_RS1_HDU;
  output [4:0] ADD_RS2_HDU;
  output [4:0] ADD_WR_OUT;
  output [4:0] ADD_RS1_OUT;
  output [4:0] ADD_RS2_OUT;
  input CLK, RST, Bubble, RF_WE, ZERO_FLAG;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, sig_RST, sig_Rtype,
         sig_Itype, sig_Jtype, RD1, RD2, n1, n3, n4, n6, n10, n11, n12, n18,
         n19, n20;
  wire   [4:0] sig_ADD_WR;
  wire   [31:0] sig_IMM;
  wire   [4:0] sig_ADD_WRHAZ;
  wire   [4:0] sig_ADD_RS1HAZ;
  wire   [4:0] sig_ADD_RS2HAZ;

  NOR2_X2 U3 ( .A1(ZERO_FLAG), .A2(n20), .ZN(sig_RST) );
  instruction_type ins_type ( .INST_IN(INS_IN), .Rtype(sig_Rtype), .Itype(
        sig_Itype), .Jtype(sig_Jtype) );
  instruction_decomposition ins_dec ( .INST_IN({INS_IN[31:28], n12, n11, 
        INS_IN[25:0]}), .Rtype(sig_Rtype), .Itype(sig_Itype), .Jtype(sig_Jtype), .ADD_RS1({n21, n22, n23, n24, n25}), .ADD_RS2({n26, n27, n28, n29, n30}), 
        .ADD_WR(sig_ADD_WR), .IMM(sig_IMM), .RD1(RD1), .RD2(RD2) );
  regn_N32_7 regPC ( .DIN(PC_IN), .CLK(CLK), .EN(1'b1), .RST(sig_RST), .DOUT(
        PC_OUT) );
  regn_N32_6 regIMM ( .DIN(sig_IMM), .CLK(CLK), .EN(1'b1), .RST(sig_RST), 
        .DOUT(IMM_OUT) );
  regn_N5_0 regWR ( .DIN(sig_ADD_WRHAZ), .CLK(CLK), .EN(1'b1), .RST(sig_RST), 
        .DOUT(ADD_WR_OUT) );
  regn_N5_4 regRS1 ( .DIN(sig_ADD_RS1HAZ), .CLK(CLK), .EN(1'b1), .RST(sig_RST), 
        .DOUT(ADD_RS1_OUT) );
  regn_N5_3 regRS2 ( .DIN(sig_ADD_RS2HAZ), .CLK(CLK), .EN(1'b1), .RST(sig_RST), 
        .DOUT(ADD_RS2_OUT) );
  mux21_NBIT5_0 muxRS1 ( .A({ADD_RS1_HDU[4:3], n10, ADD_RS1_HDU[1], n4}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(Bubble), .Z(sig_ADD_RS1HAZ) );
  mux21_NBIT5_2 muxRS2 ( .A({n3, n1, n6, n29, ADD_RS2_HDU[0]}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .S(Bubble), .Z(sig_ADD_RS2HAZ) );
  mux21_NBIT5_1 muxWR ( .A(sig_ADD_WR), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .S(Bubble), .Z(sig_ADD_WRHAZ) );
  register_file_NBIT_ADD5_NBIT_DATA32 rf ( .CLK(CLK), .RST(RST), .ENABLE(1'b1), 
        .RD1(RD1), .RD2(RD2), .WR(RF_WE), .ADD_WR(ADD_WR), .ADD_RS1({n21, n22, 
        n23, n24, n25}), .ADD_RS2({n19, n18, n28, n29, n30}), .DATAIN(
        DATA_WR_IN), .OUT1(A_OUT), .OUT2(B_OUT) );
  CLKBUF_X1 U4 ( .A(n30), .Z(ADD_RS2_HDU[0]) );
  BUF_X1 U5 ( .A(n22), .Z(ADD_RS1_HDU[3]) );
  CLKBUF_X1 U6 ( .A(INS_IN[27]), .Z(n12) );
  CLKBUF_X1 U7 ( .A(n18), .Z(n1) );
  CLKBUF_X1 U8 ( .A(n24), .Z(ADD_RS1_HDU[1]) );
  CLKBUF_X1 U9 ( .A(n19), .Z(n3) );
  BUF_X2 U10 ( .A(n26), .Z(n19) );
  CLKBUF_X1 U11 ( .A(n25), .Z(n4) );
  CLKBUF_X1 U12 ( .A(n4), .Z(ADD_RS1_HDU[0]) );
  CLKBUF_X1 U13 ( .A(n28), .Z(n6) );
  CLKBUF_X1 U14 ( .A(n29), .Z(ADD_RS2_HDU[1]) );
  CLKBUF_X1 U15 ( .A(n1), .Z(ADD_RS2_HDU[3]) );
  CLKBUF_X1 U16 ( .A(n3), .Z(ADD_RS2_HDU[4]) );
  CLKBUF_X1 U17 ( .A(n21), .Z(ADD_RS1_HDU[4]) );
  CLKBUF_X3 U18 ( .A(n27), .Z(n18) );
  CLKBUF_X1 U19 ( .A(n23), .Z(n10) );
  CLKBUF_X1 U20 ( .A(INS_IN[26]), .Z(n11) );
  CLKBUF_X1 U21 ( .A(n10), .Z(ADD_RS1_HDU[2]) );
  CLKBUF_X1 U22 ( .A(n6), .Z(ADD_RS2_HDU[2]) );
  INV_X1 U23 ( .A(RST), .ZN(n20) );
endmodule


module Branch_Cond_Unit_NBIT32 ( RST, A, .ALU_OPC({\ALU_OPC[4] , \ALU_OPC[3] , 
        \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), JUMP_TYPE, PC_SEL, ZERO );
  input [31:0] A;
  input [1:0] JUMP_TYPE;
  output [1:0] PC_SEL;
  input RST, \ALU_OPC[4] , \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] ,
         \ALU_OPC[0] ;
  output ZERO;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n1, n2;
  wire   [4:0] ALU_OPC;

  NAND3_X1 U24 ( .A1(ALU_OPC[2]), .A2(n7), .A3(ALU_OPC[3]), .ZN(n9) );
  NAND3_X1 U25 ( .A1(ALU_OPC[3]), .A2(ALU_OPC[2]), .A3(n20), .ZN(n7) );
  NOR4_X1 U3 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n15) );
  NOR4_X1 U4 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n19) );
  NOR4_X1 U5 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n14) );
  NOR4_X1 U6 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n18) );
  NOR4_X1 U7 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n13) );
  NOR4_X1 U8 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n17) );
  NOR4_X1 U9 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n12) );
  NOR2_X1 U10 ( .A1(n10), .A2(n11), .ZN(n8) );
  NAND4_X1 U11 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .ZN(n10) );
  NAND4_X1 U12 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .ZN(n11) );
  NOR4_X1 U13 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n16) );
  NOR3_X1 U14 ( .A1(ALU_OPC[0]), .A2(ALU_OPC[4]), .A3(ALU_OPC[1]), .ZN(n20) );
  OAI211_X1 U15 ( .C1(n5), .C2(n6), .A(JUMP_TYPE[0]), .B(RST), .ZN(n4) );
  NOR2_X1 U16 ( .A1(n7), .A2(n1), .ZN(n6) );
  NOR4_X1 U17 ( .A1(n9), .A2(n8), .A3(ALU_OPC[4]), .A4(ALU_OPC[1]), .ZN(n5) );
  INV_X1 U18 ( .A(n8), .ZN(n1) );
  NAND2_X1 U19 ( .A1(JUMP_TYPE[1]), .A2(RST), .ZN(n3) );
  NAND2_X1 U20 ( .A1(n3), .A2(n4), .ZN(ZERO) );
  OAI22_X1 U21 ( .A1(JUMP_TYPE[0]), .A2(n3), .B1(JUMP_TYPE[1]), .B2(n4), .ZN(
        PC_SEL[0]) );
  NOR2_X1 U22 ( .A1(n2), .A2(n3), .ZN(PC_SEL[1]) );
  INV_X1 U23 ( .A(JUMP_TYPE[0]), .ZN(n2) );
endmodule


module ff_1 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n4, n5, n6;

  DFFR_X1 Q_reg ( .D(n4), .CK(CLK), .RN(RST), .Q(Q), .QN(n5) );
  OAI21_X1 U2 ( .B1(n5), .B2(EN), .A(n6), .ZN(n4) );
  NAND2_X1 U3 ( .A1(EN), .A2(D), .ZN(n6) );
endmodule


module regn_N2 ( DIN, CLK, EN, RST, DOUT );
  input [1:0] DIN;
  output [1:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n4, n5, n6;

  DFFR_X1 \DOUT_reg[1]  ( .D(n6), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n4) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n5), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n3) );
  OAI21_X1 U2 ( .B1(n3), .B2(EN), .A(n1), .ZN(n5) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n1) );
  OAI21_X1 U4 ( .B1(n4), .B2(EN), .A(n2), .ZN(n6) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n2) );
endmodule


module FWD_Unit ( RST, ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB, RF_WE_MEM, 
        RF_WE_WB, FWDA, FWDB );
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [4:0] ADD_WR_MEM;
  input [4:0] ADD_WR_WB;
  output [1:0] FWDA;
  output [1:0] FWDB;
  input RST, RF_WE_MEM, RF_WE_WB;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42;

  NOR2_X1 U3 ( .A1(n1), .A2(n2), .ZN(FWDB[1]) );
  AOI21_X1 U4 ( .B1(n3), .B2(n4), .A(n5), .ZN(n1) );
  INV_X1 U5 ( .A(n6), .ZN(n3) );
  NOR2_X1 U6 ( .A1(n2), .A2(n7), .ZN(FWDB[0]) );
  MUX2_X1 U7 ( .A(n6), .B(n8), .S(n5), .Z(n7) );
  AND4_X1 U8 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n5) );
  NOR2_X1 U9 ( .A1(n13), .A2(n14), .ZN(n12) );
  XOR2_X1 U10 ( .A(ADD_WR_MEM[4]), .B(ADD_RS2[4]), .Z(n14) );
  XOR2_X1 U11 ( .A(ADD_WR_MEM[3]), .B(ADD_RS2[3]), .Z(n13) );
  XNOR2_X1 U12 ( .A(ADD_RS2[1]), .B(ADD_WR_MEM[1]), .ZN(n11) );
  XNOR2_X1 U13 ( .A(ADD_RS2[2]), .B(ADD_WR_MEM[2]), .ZN(n10) );
  XNOR2_X1 U14 ( .A(ADD_RS2[0]), .B(ADD_WR_MEM[0]), .ZN(n9) );
  NAND4_X1 U15 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(n6) );
  NOR2_X1 U16 ( .A1(n19), .A2(n20), .ZN(n18) );
  XOR2_X1 U17 ( .A(ADD_WR_WB[3]), .B(ADD_RS2[3]), .Z(n20) );
  XOR2_X1 U18 ( .A(ADD_WR_WB[2]), .B(ADD_RS2[2]), .Z(n19) );
  XNOR2_X1 U19 ( .A(ADD_RS2[4]), .B(ADD_WR_WB[4]), .ZN(n17) );
  XNOR2_X1 U20 ( .A(ADD_RS2[1]), .B(ADD_WR_WB[1]), .ZN(n16) );
  XNOR2_X1 U21 ( .A(ADD_RS2[0]), .B(ADD_WR_WB[0]), .ZN(n15) );
  NOR2_X1 U22 ( .A1(n21), .A2(n2), .ZN(FWDA[1]) );
  AOI21_X1 U23 ( .B1(n22), .B2(n4), .A(n23), .ZN(n21) );
  OAI21_X1 U24 ( .B1(n24), .B2(n25), .A(RF_WE_WB), .ZN(n4) );
  OR2_X1 U25 ( .A1(ADD_WR_WB[0]), .A2(ADD_WR_WB[1]), .ZN(n25) );
  OR3_X1 U26 ( .A1(ADD_WR_WB[3]), .A2(ADD_WR_WB[4]), .A3(ADD_WR_WB[2]), .ZN(
        n24) );
  INV_X1 U27 ( .A(n26), .ZN(n22) );
  NOR2_X1 U28 ( .A1(n2), .A2(n27), .ZN(FWDA[0]) );
  MUX2_X1 U29 ( .A(n26), .B(n8), .S(n23), .Z(n27) );
  AND4_X1 U30 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n23) );
  NOR2_X1 U31 ( .A1(n32), .A2(n33), .ZN(n31) );
  XOR2_X1 U32 ( .A(ADD_WR_MEM[4]), .B(ADD_RS1[4]), .Z(n33) );
  XOR2_X1 U33 ( .A(ADD_WR_MEM[3]), .B(ADD_RS1[3]), .Z(n32) );
  XNOR2_X1 U34 ( .A(ADD_RS1[1]), .B(ADD_WR_MEM[1]), .ZN(n30) );
  XNOR2_X1 U35 ( .A(ADD_RS1[2]), .B(ADD_WR_MEM[2]), .ZN(n29) );
  XNOR2_X1 U36 ( .A(ADD_RS1[0]), .B(ADD_WR_MEM[0]), .ZN(n28) );
  INV_X1 U37 ( .A(n34), .ZN(n8) );
  OAI21_X1 U38 ( .B1(n35), .B2(n36), .A(RF_WE_MEM), .ZN(n34) );
  OR2_X1 U39 ( .A1(ADD_WR_MEM[0]), .A2(ADD_WR_MEM[1]), .ZN(n36) );
  OR3_X1 U40 ( .A1(ADD_WR_MEM[3]), .A2(ADD_WR_MEM[4]), .A3(ADD_WR_MEM[2]), 
        .ZN(n35) );
  NAND4_X1 U41 ( .A1(n37), .A2(n38), .A3(n39), .A4(n40), .ZN(n26) );
  NOR2_X1 U42 ( .A1(n41), .A2(n42), .ZN(n40) );
  XOR2_X1 U43 ( .A(ADD_WR_WB[3]), .B(ADD_RS1[3]), .Z(n42) );
  XOR2_X1 U44 ( .A(ADD_WR_WB[2]), .B(ADD_RS1[2]), .Z(n41) );
  XNOR2_X1 U45 ( .A(ADD_RS1[4]), .B(ADD_WR_WB[4]), .ZN(n39) );
  XNOR2_X1 U46 ( .A(ADD_RS1[1]), .B(ADD_WR_WB[1]), .ZN(n38) );
  XNOR2_X1 U47 ( .A(ADD_RS1[0]), .B(ADD_WR_WB[0]), .ZN(n37) );
  INV_X1 U48 ( .A(RST), .ZN(n2) );
endmodule


module mux41_NBIT32_0 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n1, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  BUF_X1 U1 ( .A(n6), .Z(n72) );
  BUF_X1 U2 ( .A(n6), .Z(n73) );
  BUF_X1 U3 ( .A(n4), .Z(n78) );
  BUF_X1 U4 ( .A(n4), .Z(n79) );
  BUF_X1 U5 ( .A(n7), .Z(n1) );
  BUF_X1 U6 ( .A(n7), .Z(n70) );
  BUF_X1 U7 ( .A(n5), .Z(n75) );
  BUF_X1 U8 ( .A(n5), .Z(n76) );
  BUF_X1 U9 ( .A(n6), .Z(n74) );
  BUF_X1 U10 ( .A(n4), .Z(n80) );
  BUF_X1 U11 ( .A(n7), .Z(n71) );
  BUF_X1 U12 ( .A(n5), .Z(n77) );
  NOR2_X1 U13 ( .A1(n81), .A2(S[1]), .ZN(n6) );
  NOR2_X1 U14 ( .A1(S[0]), .A2(S[1]), .ZN(n7) );
  AND2_X1 U15 ( .A1(S[1]), .A2(S[0]), .ZN(n4) );
  AND2_X1 U16 ( .A1(S[1]), .A2(n81), .ZN(n5) );
  INV_X1 U17 ( .A(S[0]), .ZN(n81) );
  NAND2_X1 U18 ( .A1(n68), .A2(n69), .ZN(Z[0]) );
  AOI22_X1 U19 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n68) );
  AOI22_X1 U20 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n69) );
  NAND2_X1 U21 ( .A1(n44), .A2(n45), .ZN(Z[20]) );
  NAND2_X1 U22 ( .A1(n36), .A2(n37), .ZN(Z[24]) );
  NAND2_X1 U23 ( .A1(n52), .A2(n53), .ZN(Z[17]) );
  AOI22_X1 U24 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n52) );
  AOI22_X1 U25 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n53) );
  NAND2_X1 U26 ( .A1(n60), .A2(n61), .ZN(Z[13]) );
  AOI22_X1 U27 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n60) );
  AOI22_X1 U28 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n61) );
  NAND2_X1 U29 ( .A1(n12), .A2(n13), .ZN(Z[6]) );
  AOI22_X1 U30 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n12) );
  AOI22_X1 U31 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n20), .A2(n21), .ZN(Z[31]) );
  AOI22_X1 U33 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n20) );
  AOI22_X1 U34 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n21) );
  NAND2_X1 U35 ( .A1(n28), .A2(n29), .ZN(Z[28]) );
  AOI22_X1 U36 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n28) );
  AOI22_X1 U37 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n29) );
  NAND2_X1 U38 ( .A1(n66), .A2(n67), .ZN(Z[10]) );
  NAND2_X1 U39 ( .A1(n42), .A2(n43), .ZN(Z[21]) );
  AOI22_X1 U40 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n42) );
  AOI22_X1 U41 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n43) );
  NAND2_X1 U42 ( .A1(n50), .A2(n51), .ZN(Z[18]) );
  AOI22_X1 U43 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n50) );
  AOI22_X1 U44 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n51) );
  NAND2_X1 U45 ( .A1(n58), .A2(n59), .ZN(Z[14]) );
  AOI22_X1 U46 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n58) );
  AOI22_X1 U47 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n59) );
  NAND2_X1 U48 ( .A1(n10), .A2(n11), .ZN(Z[7]) );
  AOI22_X1 U49 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n10) );
  AOI22_X1 U50 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n11) );
  NAND2_X1 U51 ( .A1(n18), .A2(n19), .ZN(Z[3]) );
  AOI22_X1 U52 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n18) );
  AOI22_X1 U53 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n19) );
  NAND2_X1 U54 ( .A1(n26), .A2(n27), .ZN(Z[29]) );
  AOI22_X1 U55 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n26) );
  AOI22_X1 U56 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n27) );
  NAND2_X1 U57 ( .A1(n34), .A2(n35), .ZN(Z[25]) );
  AOI22_X1 U58 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n34) );
  AOI22_X1 U59 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n35) );
  NAND2_X1 U60 ( .A1(n2), .A2(n3), .ZN(Z[9]) );
  NAND2_X1 U61 ( .A1(n64), .A2(n65), .ZN(Z[11]) );
  NAND2_X1 U62 ( .A1(n40), .A2(n41), .ZN(Z[22]) );
  AOI22_X1 U63 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n40) );
  AOI22_X1 U64 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n41) );
  NAND2_X1 U65 ( .A1(n48), .A2(n49), .ZN(Z[19]) );
  AOI22_X1 U66 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n48) );
  AOI22_X1 U67 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n49) );
  NAND2_X1 U68 ( .A1(n56), .A2(n57), .ZN(Z[15]) );
  AOI22_X1 U69 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n56) );
  AOI22_X1 U70 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n57) );
  NAND2_X1 U71 ( .A1(n8), .A2(n9), .ZN(Z[8]) );
  AOI22_X1 U72 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n8) );
  AOI22_X1 U73 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n9) );
  NAND2_X1 U74 ( .A1(n16), .A2(n17), .ZN(Z[4]) );
  AOI22_X1 U75 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n16) );
  AOI22_X1 U76 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n17) );
  NAND2_X1 U77 ( .A1(n24), .A2(n25), .ZN(Z[2]) );
  AOI22_X1 U78 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n24) );
  AOI22_X1 U79 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n25) );
  NAND2_X1 U80 ( .A1(n32), .A2(n33), .ZN(Z[26]) );
  AOI22_X1 U81 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n32) );
  AOI22_X1 U82 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n33) );
  NAND2_X1 U83 ( .A1(n38), .A2(n39), .ZN(Z[23]) );
  AOI22_X1 U84 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n38) );
  AOI22_X1 U85 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n39) );
  NAND2_X1 U86 ( .A1(n46), .A2(n47), .ZN(Z[1]) );
  AOI22_X1 U87 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n46) );
  AOI22_X1 U88 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n47) );
  NAND2_X1 U89 ( .A1(n54), .A2(n55), .ZN(Z[16]) );
  AOI22_X1 U90 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n54) );
  AOI22_X1 U91 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n55) );
  NAND2_X1 U92 ( .A1(n62), .A2(n63), .ZN(Z[12]) );
  AOI22_X1 U93 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n62) );
  AOI22_X1 U94 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n63) );
  NAND2_X1 U95 ( .A1(n14), .A2(n15), .ZN(Z[5]) );
  AOI22_X1 U96 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n14) );
  AOI22_X1 U97 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n15) );
  NAND2_X1 U98 ( .A1(n22), .A2(n23), .ZN(Z[30]) );
  AOI22_X1 U99 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n22) );
  AOI22_X1 U100 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n23) );
  NAND2_X1 U101 ( .A1(n30), .A2(n31), .ZN(Z[27]) );
  AOI22_X1 U102 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n30) );
  AOI22_X1 U103 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n31) );
  AOI22_X1 U104 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n64) );
  AOI22_X1 U105 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n65) );
  AOI22_X1 U106 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n66) );
  AOI22_X1 U107 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n67) );
  AOI22_X1 U108 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n44) );
  AOI22_X1 U109 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n45) );
  AOI22_X1 U110 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n36) );
  AOI22_X1 U111 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n37) );
  AOI22_X1 U112 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n2) );
  AOI22_X1 U113 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n3) );
endmodule


module mux41_NBIT32_4 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149;

  BUF_X1 U1 ( .A(n145), .Z(n73) );
  BUF_X1 U2 ( .A(n147), .Z(n79) );
  BUF_X1 U3 ( .A(n144), .Z(n70) );
  BUF_X1 U4 ( .A(n146), .Z(n76) );
  BUF_X1 U5 ( .A(n145), .Z(n72) );
  BUF_X1 U6 ( .A(n147), .Z(n78) );
  BUF_X1 U7 ( .A(n144), .Z(n1) );
  BUF_X1 U8 ( .A(n146), .Z(n75) );
  BUF_X1 U9 ( .A(n145), .Z(n74) );
  BUF_X1 U10 ( .A(n147), .Z(n80) );
  BUF_X1 U11 ( .A(n144), .Z(n71) );
  BUF_X1 U12 ( .A(n146), .Z(n77) );
  NOR2_X1 U13 ( .A1(n81), .A2(S[1]), .ZN(n145) );
  NOR2_X1 U14 ( .A1(S[0]), .A2(S[1]), .ZN(n144) );
  AND2_X1 U15 ( .A1(S[1]), .A2(S[0]), .ZN(n147) );
  AND2_X1 U16 ( .A1(S[1]), .A2(n81), .ZN(n146) );
  INV_X1 U17 ( .A(S[0]), .ZN(n81) );
  NAND2_X1 U18 ( .A1(n87), .A2(n86), .ZN(Z[11]) );
  NAND2_X1 U19 ( .A1(n83), .A2(n82), .ZN(Z[0]) );
  AOI22_X1 U20 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n83) );
  AOI22_X1 U21 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n82) );
  NAND2_X1 U22 ( .A1(n135), .A2(n134), .ZN(Z[4]) );
  AOI22_X1 U23 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n135) );
  AOI22_X1 U24 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n134) );
  NAND2_X1 U25 ( .A1(n143), .A2(n142), .ZN(Z[8]) );
  AOI22_X1 U26 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n143) );
  AOI22_X1 U27 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n142) );
  NAND2_X1 U28 ( .A1(n89), .A2(n88), .ZN(Z[12]) );
  AOI22_X1 U29 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n89) );
  AOI22_X1 U30 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n88) );
  NAND2_X1 U31 ( .A1(n97), .A2(n96), .ZN(Z[16]) );
  AOI22_X1 U32 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n97) );
  AOI22_X1 U33 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n96) );
  NAND2_X1 U34 ( .A1(n137), .A2(n136), .ZN(Z[5]) );
  AOI22_X1 U35 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n137) );
  AOI22_X1 U36 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n136) );
  NAND2_X1 U37 ( .A1(n105), .A2(n104), .ZN(Z[1]) );
  AOI22_X1 U38 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n105) );
  AOI22_X1 U39 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n104) );
  NAND2_X1 U40 ( .A1(n91), .A2(n90), .ZN(Z[13]) );
  AOI22_X1 U41 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n91) );
  AOI22_X1 U42 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n90) );
  NAND2_X1 U43 ( .A1(n99), .A2(n98), .ZN(Z[17]) );
  AOI22_X1 U44 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n99) );
  AOI22_X1 U45 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n98) );
  NAND2_X1 U46 ( .A1(n117), .A2(n116), .ZN(Z[25]) );
  AOI22_X1 U47 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n117) );
  AOI22_X1 U48 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n116) );
  NAND2_X1 U49 ( .A1(n127), .A2(n126), .ZN(Z[2]) );
  AOI22_X1 U50 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n127) );
  AOI22_X1 U51 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n126) );
  NAND2_X1 U52 ( .A1(n139), .A2(n138), .ZN(Z[6]) );
  AOI22_X1 U53 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n139) );
  AOI22_X1 U54 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n138) );
  NAND2_X1 U55 ( .A1(n93), .A2(n92), .ZN(Z[14]) );
  AOI22_X1 U56 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n93) );
  AOI22_X1 U57 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n92) );
  NAND2_X1 U58 ( .A1(n101), .A2(n100), .ZN(Z[18]) );
  AOI22_X1 U59 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n101) );
  AOI22_X1 U60 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n100) );
  NAND2_X1 U61 ( .A1(n119), .A2(n118), .ZN(Z[26]) );
  AOI22_X1 U62 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n119) );
  AOI22_X1 U63 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n118) );
  NAND2_X1 U64 ( .A1(n111), .A2(n110), .ZN(Z[22]) );
  AOI22_X1 U65 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n111) );
  AOI22_X1 U66 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n110) );
  NAND2_X1 U67 ( .A1(n109), .A2(n108), .ZN(Z[21]) );
  AOI22_X1 U68 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n109) );
  AOI22_X1 U69 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n108) );
  NAND2_X1 U70 ( .A1(n129), .A2(n128), .ZN(Z[30]) );
  AOI22_X1 U71 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n129) );
  AOI22_X1 U72 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n128) );
  NAND2_X1 U73 ( .A1(n125), .A2(n124), .ZN(Z[29]) );
  AOI22_X1 U74 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n125) );
  AOI22_X1 U75 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n124) );
  NAND2_X1 U76 ( .A1(n123), .A2(n122), .ZN(Z[28]) );
  AOI22_X1 U77 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n123) );
  AOI22_X1 U78 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n122) );
  NAND2_X1 U79 ( .A1(n133), .A2(n132), .ZN(Z[3]) );
  AOI22_X1 U80 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n133) );
  AOI22_X1 U81 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n132) );
  NAND2_X1 U82 ( .A1(n141), .A2(n140), .ZN(Z[7]) );
  AOI22_X1 U83 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n141) );
  AOI22_X1 U84 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n140) );
  NAND2_X1 U85 ( .A1(n95), .A2(n94), .ZN(Z[15]) );
  AOI22_X1 U86 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n95) );
  AOI22_X1 U87 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n94) );
  NAND2_X1 U88 ( .A1(n103), .A2(n102), .ZN(Z[19]) );
  AOI22_X1 U89 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n103) );
  AOI22_X1 U90 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n102) );
  NAND2_X1 U91 ( .A1(n113), .A2(n112), .ZN(Z[23]) );
  AOI22_X1 U92 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n113) );
  AOI22_X1 U93 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n112) );
  NAND2_X1 U94 ( .A1(n121), .A2(n120), .ZN(Z[27]) );
  AOI22_X1 U95 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n121) );
  AOI22_X1 U96 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n120) );
  NAND2_X1 U97 ( .A1(n131), .A2(n130), .ZN(Z[31]) );
  AOI22_X1 U98 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n131) );
  AOI22_X1 U99 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n130) );
  NAND2_X1 U100 ( .A1(n115), .A2(n114), .ZN(Z[24]) );
  AOI22_X1 U101 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n115) );
  AOI22_X1 U102 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n114) );
  NAND2_X1 U103 ( .A1(n149), .A2(n148), .ZN(Z[9]) );
  AOI22_X1 U104 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n149) );
  AOI22_X1 U105 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n148) );
  NAND2_X1 U106 ( .A1(n85), .A2(n84), .ZN(Z[10]) );
  AOI22_X1 U107 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n85) );
  AOI22_X1 U108 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n84) );
  NAND2_X1 U109 ( .A1(n107), .A2(n106), .ZN(Z[20]) );
  AOI22_X1 U110 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n107) );
  AOI22_X1 U111 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n106) );
  AOI22_X1 U112 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n87) );
  AOI22_X1 U113 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n86) );
endmodule


module mux21_NBIT32_4 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100;

  BUF_X1 U1 ( .A(n68), .Z(n1) );
  BUF_X1 U2 ( .A(n68), .Z(n2) );
  BUF_X1 U3 ( .A(n68), .Z(n3) );
  INV_X1 U4 ( .A(n69), .ZN(Z[0]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n1), .B1(B[0]), .B2(S), .ZN(n69) );
  INV_X1 U6 ( .A(n81), .ZN(Z[20]) );
  AOI22_X1 U7 ( .A1(A[20]), .A2(n2), .B1(B[20]), .B2(S), .ZN(n81) );
  INV_X1 U8 ( .A(n85), .ZN(Z[24]) );
  AOI22_X1 U9 ( .A1(A[24]), .A2(n2), .B1(B[24]), .B2(S), .ZN(n85) );
  INV_X1 U10 ( .A(n97), .ZN(Z[6]) );
  AOI22_X1 U11 ( .A1(A[6]), .A2(n3), .B1(B[6]), .B2(S), .ZN(n97) );
  INV_X1 U12 ( .A(n70), .ZN(Z[10]) );
  AOI22_X1 U13 ( .A1(A[10]), .A2(n1), .B1(B[10]), .B2(S), .ZN(n70) );
  INV_X1 U14 ( .A(n73), .ZN(Z[13]) );
  AOI22_X1 U15 ( .A1(A[13]), .A2(n1), .B1(B[13]), .B2(S), .ZN(n73) );
  INV_X1 U16 ( .A(n77), .ZN(Z[17]) );
  AOI22_X1 U17 ( .A1(A[17]), .A2(n1), .B1(B[17]), .B2(S), .ZN(n77) );
  INV_X1 U18 ( .A(n89), .ZN(Z[28]) );
  AOI22_X1 U19 ( .A1(A[28]), .A2(n2), .B1(B[28]), .B2(S), .ZN(n89) );
  INV_X1 U20 ( .A(n93), .ZN(Z[31]) );
  AOI22_X1 U21 ( .A1(A[31]), .A2(n3), .B1(B[31]), .B2(S), .ZN(n93) );
  INV_X1 U22 ( .A(n94), .ZN(Z[3]) );
  AOI22_X1 U23 ( .A1(A[3]), .A2(n3), .B1(B[3]), .B2(S), .ZN(n94) );
  INV_X1 U24 ( .A(n98), .ZN(Z[7]) );
  AOI22_X1 U25 ( .A1(A[7]), .A2(n3), .B1(B[7]), .B2(S), .ZN(n98) );
  INV_X1 U26 ( .A(n74), .ZN(Z[14]) );
  AOI22_X1 U27 ( .A1(A[14]), .A2(n1), .B1(B[14]), .B2(S), .ZN(n74) );
  INV_X1 U28 ( .A(n78), .ZN(Z[18]) );
  AOI22_X1 U29 ( .A1(A[18]), .A2(n1), .B1(B[18]), .B2(S), .ZN(n78) );
  INV_X1 U30 ( .A(n82), .ZN(Z[21]) );
  AOI22_X1 U31 ( .A1(A[21]), .A2(n2), .B1(B[21]), .B2(S), .ZN(n82) );
  INV_X1 U32 ( .A(n86), .ZN(Z[25]) );
  AOI22_X1 U33 ( .A1(A[25]), .A2(n2), .B1(B[25]), .B2(S), .ZN(n86) );
  INV_X1 U34 ( .A(n90), .ZN(Z[29]) );
  AOI22_X1 U35 ( .A1(A[29]), .A2(n2), .B1(B[29]), .B2(S), .ZN(n90) );
  INV_X1 U36 ( .A(n71), .ZN(Z[11]) );
  AOI22_X1 U37 ( .A1(A[11]), .A2(n1), .B1(B[11]), .B2(S), .ZN(n71) );
  INV_X1 U38 ( .A(n91), .ZN(Z[2]) );
  AOI22_X1 U39 ( .A1(A[2]), .A2(n2), .B1(B[2]), .B2(S), .ZN(n91) );
  INV_X1 U40 ( .A(n95), .ZN(Z[4]) );
  AOI22_X1 U41 ( .A1(A[4]), .A2(n3), .B1(B[4]), .B2(S), .ZN(n95) );
  INV_X1 U42 ( .A(n99), .ZN(Z[8]) );
  AOI22_X1 U43 ( .A1(A[8]), .A2(n3), .B1(B[8]), .B2(S), .ZN(n99) );
  INV_X1 U44 ( .A(n75), .ZN(Z[15]) );
  AOI22_X1 U45 ( .A1(A[15]), .A2(n1), .B1(B[15]), .B2(S), .ZN(n75) );
  INV_X1 U46 ( .A(n79), .ZN(Z[19]) );
  AOI22_X1 U47 ( .A1(A[19]), .A2(n1), .B1(B[19]), .B2(S), .ZN(n79) );
  INV_X1 U48 ( .A(n83), .ZN(Z[22]) );
  AOI22_X1 U49 ( .A1(A[22]), .A2(n2), .B1(B[22]), .B2(S), .ZN(n83) );
  INV_X1 U50 ( .A(n87), .ZN(Z[26]) );
  AOI22_X1 U51 ( .A1(A[26]), .A2(n2), .B1(B[26]), .B2(S), .ZN(n87) );
  INV_X1 U52 ( .A(n80), .ZN(Z[1]) );
  AOI22_X1 U53 ( .A1(A[1]), .A2(n1), .B1(B[1]), .B2(S), .ZN(n80) );
  INV_X1 U54 ( .A(n96), .ZN(Z[5]) );
  AOI22_X1 U55 ( .A1(A[5]), .A2(n3), .B1(B[5]), .B2(S), .ZN(n96) );
  INV_X1 U56 ( .A(n72), .ZN(Z[12]) );
  AOI22_X1 U57 ( .A1(A[12]), .A2(n1), .B1(B[12]), .B2(S), .ZN(n72) );
  INV_X1 U58 ( .A(n76), .ZN(Z[16]) );
  AOI22_X1 U59 ( .A1(A[16]), .A2(n1), .B1(B[16]), .B2(S), .ZN(n76) );
  INV_X1 U60 ( .A(n84), .ZN(Z[23]) );
  AOI22_X1 U61 ( .A1(A[23]), .A2(n2), .B1(B[23]), .B2(S), .ZN(n84) );
  INV_X1 U62 ( .A(n88), .ZN(Z[27]) );
  AOI22_X1 U63 ( .A1(A[27]), .A2(n2), .B1(B[27]), .B2(S), .ZN(n88) );
  INV_X1 U64 ( .A(n92), .ZN(Z[30]) );
  AOI22_X1 U65 ( .A1(A[30]), .A2(n2), .B1(B[30]), .B2(S), .ZN(n92) );
  INV_X1 U66 ( .A(n100), .ZN(Z[9]) );
  AOI22_X1 U67 ( .A1(A[9]), .A2(n3), .B1(S), .B2(B[9]), .ZN(n100) );
  INV_X1 U68 ( .A(S), .ZN(n68) );
endmodule


module mux41_NBIT32_3 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149;

  BUF_X1 U1 ( .A(n145), .Z(n72) );
  BUF_X1 U2 ( .A(n147), .Z(n78) );
  BUF_X1 U3 ( .A(n145), .Z(n73) );
  BUF_X1 U4 ( .A(n147), .Z(n79) );
  BUF_X1 U5 ( .A(n144), .Z(n1) );
  BUF_X1 U6 ( .A(n146), .Z(n75) );
  BUF_X1 U7 ( .A(n144), .Z(n70) );
  BUF_X1 U8 ( .A(n146), .Z(n76) );
  BUF_X1 U9 ( .A(n145), .Z(n74) );
  BUF_X1 U10 ( .A(n147), .Z(n80) );
  BUF_X1 U11 ( .A(n144), .Z(n71) );
  BUF_X1 U12 ( .A(n146), .Z(n77) );
  NAND2_X1 U13 ( .A1(n83), .A2(n82), .ZN(Z[0]) );
  AOI22_X1 U14 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n82) );
  AOI22_X1 U15 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n83) );
  NAND2_X1 U16 ( .A1(n135), .A2(n134), .ZN(Z[4]) );
  AOI22_X1 U17 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n134) );
  AOI22_X1 U18 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n135) );
  NAND2_X1 U19 ( .A1(n143), .A2(n142), .ZN(Z[8]) );
  AOI22_X1 U20 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n142) );
  AOI22_X1 U21 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n143) );
  NAND2_X1 U22 ( .A1(n89), .A2(n88), .ZN(Z[12]) );
  AOI22_X1 U23 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n88) );
  AOI22_X1 U24 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n89) );
  NAND2_X1 U25 ( .A1(n97), .A2(n96), .ZN(Z[16]) );
  AOI22_X1 U26 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n96) );
  AOI22_X1 U27 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n97) );
  NAND2_X1 U28 ( .A1(n115), .A2(n114), .ZN(Z[24]) );
  AOI22_X1 U29 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n114) );
  AOI22_X1 U30 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n115) );
  NAND2_X1 U31 ( .A1(n137), .A2(n136), .ZN(Z[5]) );
  AOI22_X1 U32 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n136) );
  AOI22_X1 U33 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n137) );
  NAND2_X1 U34 ( .A1(n105), .A2(n104), .ZN(Z[1]) );
  AOI22_X1 U35 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n104) );
  AOI22_X1 U36 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n105) );
  NAND2_X1 U37 ( .A1(n149), .A2(n148), .ZN(Z[9]) );
  AOI22_X1 U38 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n148) );
  AOI22_X1 U39 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n149) );
  NAND2_X1 U40 ( .A1(n91), .A2(n90), .ZN(Z[13]) );
  AOI22_X1 U41 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n90) );
  AOI22_X1 U42 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n91) );
  NAND2_X1 U43 ( .A1(n99), .A2(n98), .ZN(Z[17]) );
  AOI22_X1 U44 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n98) );
  AOI22_X1 U45 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n99) );
  NAND2_X1 U46 ( .A1(n117), .A2(n116), .ZN(Z[25]) );
  AOI22_X1 U47 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n116) );
  AOI22_X1 U48 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n117) );
  NAND2_X1 U49 ( .A1(n127), .A2(n126), .ZN(Z[2]) );
  AOI22_X1 U50 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n126) );
  AOI22_X1 U51 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n127) );
  NAND2_X1 U52 ( .A1(n139), .A2(n138), .ZN(Z[6]) );
  AOI22_X1 U53 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n138) );
  AOI22_X1 U54 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n139) );
  NAND2_X1 U55 ( .A1(n85), .A2(n84), .ZN(Z[10]) );
  AOI22_X1 U56 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n84) );
  AOI22_X1 U57 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n85) );
  NAND2_X1 U58 ( .A1(n93), .A2(n92), .ZN(Z[14]) );
  AOI22_X1 U59 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n92) );
  AOI22_X1 U60 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n93) );
  NAND2_X1 U61 ( .A1(n101), .A2(n100), .ZN(Z[18]) );
  AOI22_X1 U62 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n100) );
  AOI22_X1 U63 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n101) );
  NAND2_X1 U64 ( .A1(n119), .A2(n118), .ZN(Z[26]) );
  AOI22_X1 U65 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n118) );
  AOI22_X1 U66 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n119) );
  NAND2_X1 U67 ( .A1(n111), .A2(n110), .ZN(Z[22]) );
  AOI22_X1 U68 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n110) );
  AOI22_X1 U69 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n111) );
  NAND2_X1 U70 ( .A1(n109), .A2(n108), .ZN(Z[21]) );
  AOI22_X1 U71 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n108) );
  AOI22_X1 U72 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n109) );
  NAND2_X1 U73 ( .A1(n107), .A2(n106), .ZN(Z[20]) );
  AOI22_X1 U74 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n106) );
  AOI22_X1 U75 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n107) );
  NAND2_X1 U76 ( .A1(n129), .A2(n128), .ZN(Z[30]) );
  AOI22_X1 U77 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n128) );
  AOI22_X1 U78 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n129) );
  NAND2_X1 U79 ( .A1(n125), .A2(n124), .ZN(Z[29]) );
  AOI22_X1 U80 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n124) );
  AOI22_X1 U81 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n125) );
  NAND2_X1 U82 ( .A1(n123), .A2(n122), .ZN(Z[28]) );
  AOI22_X1 U83 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n122) );
  AOI22_X1 U84 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n123) );
  NAND2_X1 U85 ( .A1(n133), .A2(n132), .ZN(Z[3]) );
  AOI22_X1 U86 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n132) );
  AOI22_X1 U87 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n133) );
  NAND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(Z[7]) );
  AOI22_X1 U89 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n140) );
  AOI22_X1 U90 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n141) );
  NAND2_X1 U91 ( .A1(n87), .A2(n86), .ZN(Z[11]) );
  AOI22_X1 U92 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n86) );
  AOI22_X1 U93 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n87) );
  NAND2_X1 U94 ( .A1(n95), .A2(n94), .ZN(Z[15]) );
  AOI22_X1 U95 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n94) );
  AOI22_X1 U96 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n95) );
  NAND2_X1 U97 ( .A1(n103), .A2(n102), .ZN(Z[19]) );
  AOI22_X1 U98 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n102) );
  AOI22_X1 U99 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n103) );
  NAND2_X1 U100 ( .A1(n113), .A2(n112), .ZN(Z[23]) );
  AOI22_X1 U101 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n112) );
  AOI22_X1 U102 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n113) );
  NAND2_X1 U103 ( .A1(n121), .A2(n120), .ZN(Z[27]) );
  AOI22_X1 U104 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n120) );
  AOI22_X1 U105 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n121) );
  NAND2_X1 U106 ( .A1(n131), .A2(n130), .ZN(Z[31]) );
  AOI22_X1 U107 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n130) );
  AOI22_X1 U108 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n131) );
  NOR2_X1 U109 ( .A1(n81), .A2(S[1]), .ZN(n145) );
  NOR2_X1 U110 ( .A1(S[0]), .A2(S[1]), .ZN(n144) );
  AND2_X1 U111 ( .A1(S[1]), .A2(S[0]), .ZN(n147) );
  AND2_X1 U112 ( .A1(S[1]), .A2(n81), .ZN(n146) );
  INV_X1 U113 ( .A(S[0]), .ZN(n81) );
endmodule


module comparator_NBIT32_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202;

  INV_X1 U1 ( .A(NE), .ZN(EQ) );
  INV_X1 U2 ( .A(n142), .ZN(n55) );
  INV_X1 U3 ( .A(n130), .ZN(n7) );
  INV_X1 U4 ( .A(n118), .ZN(n15) );
  INV_X1 U5 ( .A(n106), .ZN(n23) );
  INV_X1 U6 ( .A(n94), .ZN(n31) );
  INV_X1 U7 ( .A(n82), .ZN(n39) );
  INV_X1 U8 ( .A(n139), .ZN(n58) );
  INV_X1 U9 ( .A(n127), .ZN(n10) );
  INV_X1 U10 ( .A(n115), .ZN(n18) );
  INV_X1 U11 ( .A(n103), .ZN(n26) );
  INV_X1 U12 ( .A(n91), .ZN(n34) );
  INV_X1 U13 ( .A(n79), .ZN(n42) );
  INV_X1 U14 ( .A(GT), .ZN(LE) );
  INV_X1 U15 ( .A(n132), .ZN(n61) );
  INV_X1 U16 ( .A(n141), .ZN(n56) );
  INV_X1 U17 ( .A(n144), .ZN(n53) );
  INV_X1 U18 ( .A(n120), .ZN(n13) );
  INV_X1 U19 ( .A(n108), .ZN(n21) );
  INV_X1 U20 ( .A(n96), .ZN(n29) );
  INV_X1 U21 ( .A(n84), .ZN(n37) );
  INV_X1 U22 ( .A(n129), .ZN(n8) );
  INV_X1 U23 ( .A(n117), .ZN(n16) );
  INV_X1 U24 ( .A(n105), .ZN(n24) );
  INV_X1 U25 ( .A(n93), .ZN(n32) );
  INV_X1 U26 ( .A(n81), .ZN(n40) );
  INV_X1 U27 ( .A(n154), .ZN(n47) );
  INV_X1 U28 ( .A(n68), .ZN(n5) );
  INV_X1 U29 ( .A(A[30]), .ZN(n49) );
  INV_X1 U30 ( .A(n72), .ZN(n45) );
  INV_X1 U31 ( .A(n151), .ZN(n50) );
  INV_X1 U32 ( .A(B[30]), .ZN(n64) );
  INV_X1 U33 ( .A(n202), .ZN(n3) );
  INV_X1 U34 ( .A(B[1]), .ZN(n63) );
  INV_X1 U35 ( .A(A[0]), .ZN(n6) );
  INV_X1 U36 ( .A(A[3]), .ZN(n51) );
  INV_X1 U37 ( .A(A[5]), .ZN(n54) );
  INV_X1 U38 ( .A(A[7]), .ZN(n59) );
  INV_X1 U39 ( .A(A[9]), .ZN(n62) );
  INV_X1 U40 ( .A(A[11]), .ZN(n11) );
  INV_X1 U41 ( .A(A[13]), .ZN(n14) );
  INV_X1 U42 ( .A(A[15]), .ZN(n19) );
  INV_X1 U43 ( .A(B[31]), .ZN(n65) );
  INV_X1 U44 ( .A(A[17]), .ZN(n22) );
  INV_X1 U45 ( .A(A[19]), .ZN(n27) );
  INV_X1 U46 ( .A(A[21]), .ZN(n30) );
  INV_X1 U47 ( .A(A[23]), .ZN(n35) );
  INV_X1 U48 ( .A(A[25]), .ZN(n38) );
  INV_X1 U49 ( .A(A[27]), .ZN(n43) );
  INV_X1 U50 ( .A(A[29]), .ZN(n46) );
  INV_X1 U51 ( .A(A[4]), .ZN(n52) );
  INV_X1 U52 ( .A(A[8]), .ZN(n60) );
  INV_X1 U53 ( .A(A[12]), .ZN(n12) );
  INV_X1 U54 ( .A(A[2]), .ZN(n48) );
  INV_X1 U55 ( .A(A[6]), .ZN(n57) );
  INV_X1 U56 ( .A(A[10]), .ZN(n9) );
  INV_X1 U57 ( .A(A[14]), .ZN(n17) );
  INV_X1 U58 ( .A(A[16]), .ZN(n20) );
  INV_X1 U59 ( .A(A[20]), .ZN(n28) );
  INV_X1 U60 ( .A(A[24]), .ZN(n36) );
  INV_X1 U61 ( .A(A[28]), .ZN(n44) );
  INV_X1 U62 ( .A(A[18]), .ZN(n25) );
  INV_X1 U63 ( .A(A[22]), .ZN(n33) );
  INV_X1 U64 ( .A(A[26]), .ZN(n41) );
  INV_X1 U65 ( .A(GE), .ZN(LT) );
  NAND2_X1 U66 ( .A1(LE), .A2(GE), .ZN(NE) );
  AOI21_X1 U67 ( .B1(n66), .B2(n5), .A(n67), .ZN(GE) );
  AOI22_X1 U68 ( .A1(B[30]), .A2(n49), .B1(n69), .B2(n70), .ZN(n68) );
  AOI21_X1 U69 ( .B1(n71), .B2(n72), .A(n73), .ZN(n69) );
  AOI21_X1 U70 ( .B1(n74), .B2(n75), .A(n76), .ZN(n71) );
  AOI21_X1 U71 ( .B1(n77), .B2(n78), .A(n79), .ZN(n74) );
  AOI21_X1 U72 ( .B1(n80), .B2(n39), .A(n40), .ZN(n77) );
  AOI21_X1 U73 ( .B1(n83), .B2(n84), .A(n85), .ZN(n80) );
  AOI21_X1 U74 ( .B1(n86), .B2(n87), .A(n88), .ZN(n83) );
  AOI21_X1 U75 ( .B1(n89), .B2(n90), .A(n91), .ZN(n86) );
  AOI21_X1 U76 ( .B1(n92), .B2(n31), .A(n32), .ZN(n89) );
  AOI21_X1 U77 ( .B1(n95), .B2(n96), .A(n97), .ZN(n92) );
  AOI21_X1 U78 ( .B1(n98), .B2(n99), .A(n100), .ZN(n95) );
  AOI21_X1 U79 ( .B1(n101), .B2(n102), .A(n103), .ZN(n98) );
  AOI21_X1 U80 ( .B1(n104), .B2(n23), .A(n24), .ZN(n101) );
  AOI21_X1 U81 ( .B1(n107), .B2(n108), .A(n109), .ZN(n104) );
  AOI21_X1 U82 ( .B1(n110), .B2(n111), .A(n112), .ZN(n107) );
  AOI21_X1 U83 ( .B1(n113), .B2(n114), .A(n115), .ZN(n110) );
  AOI21_X1 U84 ( .B1(n116), .B2(n15), .A(n16), .ZN(n113) );
  AOI21_X1 U85 ( .B1(n119), .B2(n120), .A(n121), .ZN(n116) );
  AOI21_X1 U86 ( .B1(n122), .B2(n123), .A(n124), .ZN(n119) );
  AOI21_X1 U87 ( .B1(n125), .B2(n126), .A(n127), .ZN(n122) );
  AOI21_X1 U88 ( .B1(n128), .B2(n7), .A(n8), .ZN(n125) );
  AOI21_X1 U89 ( .B1(n131), .B2(n132), .A(n133), .ZN(n128) );
  AOI21_X1 U90 ( .B1(n134), .B2(n135), .A(n136), .ZN(n131) );
  AOI21_X1 U91 ( .B1(n137), .B2(n138), .A(n139), .ZN(n134) );
  AOI21_X1 U92 ( .B1(n140), .B2(n55), .A(n56), .ZN(n137) );
  AOI21_X1 U93 ( .B1(n143), .B2(n144), .A(n145), .ZN(n140) );
  AOI21_X1 U94 ( .B1(n146), .B2(n147), .A(n148), .ZN(n143) );
  AOI21_X1 U95 ( .B1(n149), .B2(n150), .A(n151), .ZN(n146) );
  AOI21_X1 U96 ( .B1(n152), .B2(n153), .A(n47), .ZN(n149) );
  AOI22_X1 U97 ( .A1(n155), .A2(n63), .B1(A[1]), .B2(n156), .ZN(n152) );
  OR2_X1 U98 ( .A1(n156), .A2(A[1]), .ZN(n155) );
  NAND2_X1 U99 ( .A1(B[0]), .A2(n6), .ZN(n156) );
  OAI21_X1 U100 ( .B1(n67), .B2(n157), .A(n66), .ZN(GT) );
  NAND2_X1 U101 ( .A1(A[31]), .A2(n65), .ZN(n66) );
  AOI22_X1 U102 ( .A1(A[30]), .A2(n64), .B1(n158), .B2(n70), .ZN(n157) );
  XOR2_X1 U103 ( .A(A[30]), .B(n64), .Z(n70) );
  AOI21_X1 U104 ( .B1(n159), .B2(n160), .A(n45), .ZN(n158) );
  NAND2_X1 U105 ( .A1(B[29]), .A2(n46), .ZN(n72) );
  OAI211_X1 U106 ( .C1(n161), .C2(n162), .A(n78), .B(n75), .ZN(n160) );
  NOR2_X1 U107 ( .A1(n163), .A2(n76), .ZN(n75) );
  AND2_X1 U108 ( .A1(B[28]), .A2(n44), .ZN(n76) );
  NAND2_X1 U109 ( .A1(B[27]), .A2(n43), .ZN(n78) );
  NAND2_X1 U110 ( .A1(n42), .A2(n164), .ZN(n162) );
  NOR2_X1 U111 ( .A1(n43), .A2(B[27]), .ZN(n79) );
  AOI211_X1 U112 ( .C1(n165), .C2(n166), .A(n82), .B(n37), .ZN(n161) );
  NAND2_X1 U113 ( .A1(B[25]), .A2(n38), .ZN(n84) );
  NAND2_X1 U114 ( .A1(n164), .A2(n81), .ZN(n82) );
  NAND2_X1 U115 ( .A1(B[26]), .A2(n41), .ZN(n81) );
  OR2_X1 U116 ( .A1(n41), .A2(B[26]), .ZN(n164) );
  OAI211_X1 U117 ( .C1(n167), .C2(n168), .A(n90), .B(n87), .ZN(n166) );
  NOR2_X1 U118 ( .A1(n169), .A2(n88), .ZN(n87) );
  AND2_X1 U119 ( .A1(B[24]), .A2(n36), .ZN(n88) );
  NAND2_X1 U120 ( .A1(B[23]), .A2(n35), .ZN(n90) );
  NAND2_X1 U121 ( .A1(n34), .A2(n170), .ZN(n168) );
  NOR2_X1 U122 ( .A1(n35), .A2(B[23]), .ZN(n91) );
  AOI211_X1 U123 ( .C1(n171), .C2(n172), .A(n94), .B(n29), .ZN(n167) );
  NAND2_X1 U124 ( .A1(B[21]), .A2(n30), .ZN(n96) );
  NAND2_X1 U125 ( .A1(n170), .A2(n93), .ZN(n94) );
  NAND2_X1 U126 ( .A1(B[22]), .A2(n33), .ZN(n93) );
  OR2_X1 U127 ( .A1(n33), .A2(B[22]), .ZN(n170) );
  OAI211_X1 U128 ( .C1(n173), .C2(n174), .A(n102), .B(n99), .ZN(n172) );
  NOR2_X1 U129 ( .A1(n175), .A2(n100), .ZN(n99) );
  AND2_X1 U130 ( .A1(B[20]), .A2(n28), .ZN(n100) );
  NAND2_X1 U131 ( .A1(B[19]), .A2(n27), .ZN(n102) );
  NAND2_X1 U132 ( .A1(n26), .A2(n176), .ZN(n174) );
  NOR2_X1 U133 ( .A1(n27), .A2(B[19]), .ZN(n103) );
  AOI211_X1 U134 ( .C1(n177), .C2(n178), .A(n106), .B(n21), .ZN(n173) );
  NAND2_X1 U135 ( .A1(B[17]), .A2(n22), .ZN(n108) );
  NAND2_X1 U136 ( .A1(n176), .A2(n105), .ZN(n106) );
  NAND2_X1 U137 ( .A1(B[18]), .A2(n25), .ZN(n105) );
  OR2_X1 U138 ( .A1(n25), .A2(B[18]), .ZN(n176) );
  OAI211_X1 U139 ( .C1(n179), .C2(n180), .A(n114), .B(n111), .ZN(n178) );
  NOR2_X1 U140 ( .A1(n181), .A2(n112), .ZN(n111) );
  AND2_X1 U141 ( .A1(B[16]), .A2(n20), .ZN(n112) );
  NAND2_X1 U142 ( .A1(B[15]), .A2(n19), .ZN(n114) );
  NAND2_X1 U143 ( .A1(n18), .A2(n182), .ZN(n180) );
  NOR2_X1 U144 ( .A1(n19), .A2(B[15]), .ZN(n115) );
  AOI211_X1 U145 ( .C1(n183), .C2(n184), .A(n118), .B(n13), .ZN(n179) );
  NAND2_X1 U146 ( .A1(B[13]), .A2(n14), .ZN(n120) );
  NAND2_X1 U147 ( .A1(n182), .A2(n117), .ZN(n118) );
  NAND2_X1 U148 ( .A1(B[14]), .A2(n17), .ZN(n117) );
  OR2_X1 U149 ( .A1(n17), .A2(B[14]), .ZN(n182) );
  OAI211_X1 U150 ( .C1(n185), .C2(n186), .A(n126), .B(n123), .ZN(n184) );
  NOR2_X1 U151 ( .A1(n187), .A2(n124), .ZN(n123) );
  AND2_X1 U152 ( .A1(B[12]), .A2(n12), .ZN(n124) );
  NAND2_X1 U153 ( .A1(B[11]), .A2(n11), .ZN(n126) );
  NAND2_X1 U154 ( .A1(n10), .A2(n188), .ZN(n186) );
  NOR2_X1 U155 ( .A1(n11), .A2(B[11]), .ZN(n127) );
  AOI211_X1 U156 ( .C1(n189), .C2(n190), .A(n130), .B(n61), .ZN(n185) );
  NAND2_X1 U157 ( .A1(B[9]), .A2(n62), .ZN(n132) );
  NAND2_X1 U158 ( .A1(n188), .A2(n129), .ZN(n130) );
  NAND2_X1 U159 ( .A1(B[10]), .A2(n9), .ZN(n129) );
  OR2_X1 U160 ( .A1(n9), .A2(B[10]), .ZN(n188) );
  OAI211_X1 U161 ( .C1(n191), .C2(n192), .A(n138), .B(n135), .ZN(n190) );
  NOR2_X1 U162 ( .A1(n193), .A2(n136), .ZN(n135) );
  AND2_X1 U163 ( .A1(B[8]), .A2(n60), .ZN(n136) );
  NAND2_X1 U164 ( .A1(B[7]), .A2(n59), .ZN(n138) );
  NAND2_X1 U165 ( .A1(n58), .A2(n194), .ZN(n192) );
  NOR2_X1 U166 ( .A1(n59), .A2(B[7]), .ZN(n139) );
  AOI211_X1 U167 ( .C1(n195), .C2(n196), .A(n142), .B(n53), .ZN(n191) );
  NAND2_X1 U168 ( .A1(B[5]), .A2(n54), .ZN(n144) );
  NAND2_X1 U169 ( .A1(n194), .A2(n141), .ZN(n142) );
  NAND2_X1 U170 ( .A1(B[6]), .A2(n57), .ZN(n141) );
  OR2_X1 U171 ( .A1(n57), .A2(B[6]), .ZN(n194) );
  NAND3_X1 U172 ( .A1(n197), .A2(n150), .A3(n147), .ZN(n196) );
  NOR2_X1 U173 ( .A1(n198), .A2(n148), .ZN(n147) );
  AND2_X1 U174 ( .A1(B[4]), .A2(n52), .ZN(n148) );
  NAND2_X1 U175 ( .A1(B[3]), .A2(n51), .ZN(n150) );
  NAND3_X1 U176 ( .A1(n50), .A2(n199), .A3(n200), .ZN(n197) );
  OAI211_X1 U177 ( .C1(A[1]), .C2(n201), .A(n3), .B(n153), .ZN(n200) );
  AND2_X1 U178 ( .A1(n199), .A2(n154), .ZN(n153) );
  NAND2_X1 U179 ( .A1(B[2]), .A2(n48), .ZN(n154) );
  AOI21_X1 U180 ( .B1(A[1]), .B2(n201), .A(n63), .ZN(n202) );
  NOR2_X1 U181 ( .A1(n6), .A2(B[0]), .ZN(n201) );
  OR2_X1 U182 ( .A1(n48), .A2(B[2]), .ZN(n199) );
  NOR2_X1 U183 ( .A1(n51), .A2(B[3]), .ZN(n151) );
  NOR2_X1 U184 ( .A1(n198), .A2(n145), .ZN(n195) );
  NOR2_X1 U185 ( .A1(n54), .A2(B[5]), .ZN(n145) );
  NOR2_X1 U186 ( .A1(n52), .A2(B[4]), .ZN(n198) );
  NOR2_X1 U187 ( .A1(n193), .A2(n133), .ZN(n189) );
  NOR2_X1 U188 ( .A1(n62), .A2(B[9]), .ZN(n133) );
  NOR2_X1 U189 ( .A1(n60), .A2(B[8]), .ZN(n193) );
  NOR2_X1 U190 ( .A1(n187), .A2(n121), .ZN(n183) );
  NOR2_X1 U191 ( .A1(n14), .A2(B[13]), .ZN(n121) );
  NOR2_X1 U192 ( .A1(n12), .A2(B[12]), .ZN(n187) );
  NOR2_X1 U193 ( .A1(n181), .A2(n109), .ZN(n177) );
  NOR2_X1 U194 ( .A1(n22), .A2(B[17]), .ZN(n109) );
  NOR2_X1 U195 ( .A1(n20), .A2(B[16]), .ZN(n181) );
  NOR2_X1 U196 ( .A1(n175), .A2(n97), .ZN(n171) );
  NOR2_X1 U197 ( .A1(n30), .A2(B[21]), .ZN(n97) );
  NOR2_X1 U198 ( .A1(n28), .A2(B[20]), .ZN(n175) );
  NOR2_X1 U199 ( .A1(n169), .A2(n85), .ZN(n165) );
  NOR2_X1 U200 ( .A1(n38), .A2(B[25]), .ZN(n85) );
  NOR2_X1 U201 ( .A1(n36), .A2(B[24]), .ZN(n169) );
  NOR2_X1 U202 ( .A1(n163), .A2(n73), .ZN(n159) );
  NOR2_X1 U203 ( .A1(n46), .A2(B[29]), .ZN(n73) );
  NOR2_X1 U204 ( .A1(n44), .A2(B[28]), .ZN(n163) );
  NOR2_X1 U205 ( .A1(n65), .A2(A[31]), .ZN(n67) );
endmodule


module comparator_NBIT32 ( A, B, .OPSel({\OPSel[2] , \OPSel[1] , \OPSel[0] }), 
        RES );
  input [31:0] A;
  input [31:0] B;
  output [31:0] RES;
  input \OPSel[2] , \OPSel[1] , \OPSel[0] ;
  wire   N26, N27, N28, N29, N30, N31, n15, n16, n17, n18, n19, n20, n2, n3,
         n4;
  wire   [2:0] OPSel;
  assign RES[1] = 1'b0;
  assign RES[2] = 1'b0;
  assign RES[3] = 1'b0;
  assign RES[4] = 1'b0;
  assign RES[5] = 1'b0;
  assign RES[6] = 1'b0;
  assign RES[7] = 1'b0;
  assign RES[8] = 1'b0;
  assign RES[9] = 1'b0;
  assign RES[10] = 1'b0;
  assign RES[11] = 1'b0;
  assign RES[12] = 1'b0;
  assign RES[13] = 1'b0;
  assign RES[14] = 1'b0;
  assign RES[15] = 1'b0;
  assign RES[16] = 1'b0;
  assign RES[17] = 1'b0;
  assign RES[18] = 1'b0;
  assign RES[19] = 1'b0;
  assign RES[20] = 1'b0;
  assign RES[21] = 1'b0;
  assign RES[22] = 1'b0;
  assign RES[23] = 1'b0;
  assign RES[24] = 1'b0;
  assign RES[25] = 1'b0;
  assign RES[26] = 1'b0;
  assign RES[27] = 1'b0;
  assign RES[28] = 1'b0;
  assign RES[29] = 1'b0;
  assign RES[30] = 1'b0;
  assign RES[31] = 1'b0;

  comparator_NBIT32_DW01_cmp6_0 r57 ( .A(A), .B(B), .TC(1'b0), .LT(N30), .GT(
        N28), .EQ(N26), .LE(N31), .GE(N29), .NE(N27) );
  INV_X1 U3 ( .A(n15), .ZN(RES[0]) );
  AOI21_X1 U4 ( .B1(n16), .B2(n4), .A(n17), .ZN(n15) );
  INV_X1 U5 ( .A(OPSel[0]), .ZN(n3) );
  OAI22_X1 U6 ( .A1(n19), .A2(n2), .B1(OPSel[1]), .B2(n20), .ZN(n16) );
  INV_X1 U7 ( .A(OPSel[1]), .ZN(n2) );
  AOI22_X1 U8 ( .A1(N28), .A2(n3), .B1(N29), .B2(OPSel[0]), .ZN(n19) );
  AOI22_X1 U9 ( .A1(N26), .A2(n3), .B1(N27), .B2(OPSel[0]), .ZN(n20) );
  NOR3_X1 U10 ( .A1(n4), .A2(OPSel[1]), .A3(n18), .ZN(n17) );
  AOI22_X1 U11 ( .A1(N30), .A2(n3), .B1(OPSel[0]), .B2(N31), .ZN(n18) );
  INV_X1 U12 ( .A(OPSel[2]), .ZN(n4) );
endmodule


module shifter_NBIT32 ( A, B, LOGIC_ARITH, LEFT_RIGHT, RES );
  input [31:0] A;
  input [31:0] B;
  output [31:0] RES;
  input LOGIC_ARITH, LEFT_RIGHT;
  wire   n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n266, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649;

  AOI21_X2 U264 ( .B1(A[31]), .B2(B[18]), .A(n483), .ZN(n282) );
  OAI21_X2 U267 ( .B1(n613), .B2(n629), .A(n486), .ZN(n285) );
  AOI21_X2 U269 ( .B1(A[31]), .B2(n39), .A(n487), .ZN(n288) );
  AOI221_X2 U388 ( .B1(n31), .B2(A[18]), .C1(n21), .C2(A[17]), .A(n568), .ZN(
        n196) );
  NOR2_X2 U428 ( .A1(n639), .A2(n39), .ZN(n165) );
  NOR2_X2 U461 ( .A1(n643), .A2(n39), .ZN(n199) );
  NAND3_X1 U637 ( .A1(n227), .A2(n647), .A3(n228), .ZN(n226) );
  NAND3_X1 U638 ( .A1(n227), .A2(n647), .A3(B[4]), .ZN(n428) );
  NAND3_X1 U639 ( .A1(n445), .A2(n199), .A3(LEFT_RIGHT), .ZN(n240) );
  NAND3_X1 U641 ( .A1(n489), .A2(n629), .A3(n579), .ZN(n255) );
  NAND3_X1 U642 ( .A1(n267), .A2(n199), .A3(n445), .ZN(n138) );
  NOR4_X1 U2 ( .A1(B[20]), .A2(B[21]), .A3(B[19]), .A4(n594), .ZN(n484) );
  NOR2_X2 U3 ( .A1(n640), .A2(B[3]), .ZN(n262) );
  NOR2_X2 U4 ( .A1(n490), .A2(B[11]), .ZN(n283) );
  NAND3_X1 U5 ( .A1(n445), .A2(n35), .A3(LEFT_RIGHT), .ZN(n269) );
  INV_X1 U6 ( .A(n167), .ZN(n636) );
  NOR2_X1 U7 ( .A1(n637), .A2(B[4]), .ZN(n167) );
  INV_X1 U8 ( .A(n169), .ZN(n645) );
  INV_X1 U9 ( .A(n165), .ZN(n638) );
  INV_X1 U10 ( .A(n199), .ZN(n642) );
  INV_X1 U11 ( .A(n32), .ZN(n28) );
  INV_X1 U12 ( .A(n32), .ZN(n26) );
  INV_X1 U13 ( .A(n32), .ZN(n27) );
  INV_X1 U14 ( .A(n22), .ZN(n14) );
  INV_X1 U15 ( .A(n22), .ZN(n15) );
  INV_X1 U16 ( .A(n21), .ZN(n16) );
  INV_X1 U17 ( .A(n505), .ZN(n644) );
  INV_X1 U18 ( .A(n31), .ZN(n29) );
  INV_X1 U19 ( .A(n493), .ZN(n641) );
  NOR2_X1 U20 ( .A1(n646), .A2(n39), .ZN(n169) );
  NAND2_X1 U21 ( .A1(n488), .A2(n454), .ZN(n161) );
  INV_X1 U22 ( .A(n42), .ZN(n39) );
  OAI222_X1 U23 ( .A1(n79), .A2(n645), .B1(n63), .B2(n636), .C1(n91), .C2(n638), .ZN(n371) );
  OAI222_X1 U24 ( .A1(n82), .A2(n645), .B1(n62), .B2(n636), .C1(n95), .C2(n638), .ZN(n360) );
  OAI222_X1 U25 ( .A1(n85), .A2(n645), .B1(n73), .B2(n636), .C1(n99), .C2(n638), .ZN(n349) );
  OAI222_X1 U26 ( .A1(n87), .A2(n645), .B1(n76), .B2(n636), .C1(n104), .C2(
        n638), .ZN(n338) );
  NOR2_X1 U27 ( .A1(n41), .A2(n643), .ZN(n493) );
  OAI22_X1 U28 ( .A1(n116), .A2(n643), .B1(n127), .B2(n639), .ZN(n383) );
  INV_X1 U29 ( .A(n454), .ZN(n637) );
  AOI21_X1 U30 ( .B1(n135), .B2(n2), .A(n519), .ZN(n286) );
  AOI21_X1 U31 ( .B1(n130), .B2(n3), .A(n519), .ZN(n312) );
  BUF_X1 U32 ( .A(n138), .Z(n34) );
  BUF_X1 U33 ( .A(n138), .Z(n33) );
  NOR2_X1 U34 ( .A1(n383), .A2(n359), .ZN(n197) );
  NOR2_X1 U35 ( .A1(n119), .A2(n359), .ZN(n181) );
  BUF_X1 U36 ( .A(n138), .Z(n35) );
  NAND2_X1 U37 ( .A1(n488), .A2(n5), .ZN(n505) );
  INV_X1 U38 ( .A(n182), .ZN(n119) );
  INV_X1 U39 ( .A(n238), .ZN(n107) );
  INV_X1 U40 ( .A(n214), .ZN(n56) );
  INV_X1 U41 ( .A(n202), .ZN(n50) );
  INV_X1 U42 ( .A(n188), .ZN(n48) );
  NOR2_X1 U43 ( .A1(n613), .A2(n148), .ZN(n150) );
  OAI21_X2 U44 ( .B1(n612), .B2(n633), .A(n481), .ZN(n279) );
  NOR2_X1 U45 ( .A1(n640), .A2(n647), .ZN(n454) );
  NAND2_X1 U46 ( .A1(n484), .A2(n631), .ZN(n281) );
  AOI222_X1 U47 ( .A1(n370), .A2(n262), .B1(n320), .B2(n260), .C1(n185), .C2(
        n3), .ZN(n238) );
  INV_X1 U48 ( .A(n356), .ZN(n643) );
  AOI222_X1 U49 ( .A1(n168), .A2(n262), .B1(n355), .B2(n260), .C1(n170), .C2(
        n3), .ZN(n471) );
  AOI222_X1 U50 ( .A1(n402), .A2(n262), .B1(n403), .B2(n260), .C1(n464), .C2(
        n2), .ZN(n461) );
  NAND2_X1 U51 ( .A1(n488), .A2(n262), .ZN(n157) );
  NAND2_X1 U52 ( .A1(n488), .A2(n260), .ZN(n158) );
  OAI222_X1 U53 ( .A1(n374), .A2(n639), .B1(n646), .B2(n375), .C1(n376), .C2(
        n643), .ZN(n172) );
  OAI222_X1 U54 ( .A1(n132), .A2(n639), .B1(n362), .B2(n646), .C1(n363), .C2(
        n643), .ZN(n139) );
  OAI222_X1 U55 ( .A1(n614), .A2(n639), .B1(n293), .B2(n646), .C1(n405), .C2(
        n643), .ZN(n348) );
  OAI222_X1 U56 ( .A1(n616), .A2(n639), .B1(n46), .B2(n646), .C1(n387), .C2(
        n643), .ZN(n337) );
  AOI221_X1 U57 ( .B1(n130), .B2(n262), .C1(n355), .C2(n2), .A(n359), .ZN(n159) );
  AOI221_X1 U58 ( .B1(n135), .B2(n262), .C1(n403), .C2(n3), .A(n359), .ZN(n347) );
  OAI221_X1 U59 ( .B1(n106), .B2(n639), .C1(n90), .C2(n643), .A(n607), .ZN(
        n480) );
  AOI22_X1 U60 ( .A1(n454), .A2(n320), .B1(n260), .B2(n370), .ZN(n607) );
  AOI222_X1 U61 ( .A1(n169), .A2(n185), .B1(n493), .B2(n320), .C1(n167), .C2(
        n370), .ZN(n550) );
  OAI222_X1 U62 ( .A1(n62), .A2(n645), .B1(n363), .B2(n636), .C1(n82), .C2(
        n638), .ZN(n418) );
  OAI222_X1 U63 ( .A1(n73), .A2(n645), .B1(n405), .B2(n636), .C1(n85), .C2(
        n638), .ZN(n404) );
  OAI222_X1 U64 ( .A1(n76), .A2(n645), .B1(n387), .B2(n636), .C1(n87), .C2(
        n638), .ZN(n386) );
  INV_X1 U65 ( .A(n260), .ZN(n646) );
  NOR2_X1 U66 ( .A1(n648), .A2(B[4]), .ZN(n488) );
  INV_X1 U67 ( .A(n262), .ZN(n639) );
  INV_X1 U68 ( .A(n332), .ZN(n628) );
  OAI222_X1 U69 ( .A1(n133), .A2(n14), .B1(n29), .B2(n615), .C1(n1), .C2(n103), 
        .ZN(n602) );
  OAI221_X1 U70 ( .B1(n363), .B2(n639), .C1(n62), .C2(n643), .A(n522), .ZN(
        n314) );
  AOI22_X1 U71 ( .A1(n454), .A2(n58), .B1(n260), .B2(n420), .ZN(n522) );
  OAI221_X1 U72 ( .B1(n405), .B2(n639), .C1(n73), .C2(n643), .A(n509), .ZN(
        n290) );
  AOI22_X1 U73 ( .A1(n454), .A2(n52), .B1(n260), .B2(n407), .ZN(n509) );
  OAI221_X1 U74 ( .B1(n387), .B2(n639), .C1(n76), .C2(n643), .A(n496), .ZN(
        n271) );
  AOI22_X1 U75 ( .A1(n454), .A2(n390), .B1(n260), .B2(n389), .ZN(n496) );
  OAI21_X1 U76 ( .B1(n613), .B2(n631), .A(n486), .ZN(n253) );
  NOR2_X1 U77 ( .A1(n613), .A2(n647), .ZN(n359) );
  NOR2_X1 U78 ( .A1(n613), .A2(n2), .ZN(n519) );
  AOI221_X1 U79 ( .B1(n219), .B2(n199), .C1(n223), .C2(n39), .A(n224), .ZN(
        n222) );
  OAI222_X1 U80 ( .A1(n638), .A2(n71), .B1(n636), .B2(n93), .C1(n645), .C2(n81), .ZN(n224) );
  AOI221_X1 U81 ( .B1(n207), .B2(n199), .C1(n211), .C2(n39), .A(n212), .ZN(
        n210) );
  OAI222_X1 U82 ( .A1(n638), .A2(n68), .B1(n636), .B2(n97), .C1(n645), .C2(n84), .ZN(n212) );
  AOI221_X1 U83 ( .B1(n193), .B2(n199), .C1(n115), .C2(n39), .A(n200), .ZN(
        n198) );
  OAI222_X1 U84 ( .A1(n638), .A2(n75), .B1(n636), .B2(n101), .C1(n645), .C2(
        n196), .ZN(n200) );
  OAI22_X1 U85 ( .A1(n8), .A2(n131), .B1(n1), .B2(n266), .ZN(n533) );
  OAI221_X1 U86 ( .B1(n618), .B2(n642), .C1(n238), .C2(n41), .A(n239), .ZN(
        n229) );
  AOI222_X1 U87 ( .A1(n165), .A2(n178), .B1(n167), .B2(n186), .C1(n169), .C2(
        n184), .ZN(n239) );
  OAI221_X1 U88 ( .B1(n65), .B2(n642), .C1(n182), .C2(n41), .A(n183), .ZN(n173) );
  AOI222_X1 U89 ( .A1(n165), .A2(n184), .B1(n167), .B2(n185), .C1(n169), .C2(
        n186), .ZN(n183) );
  OAI221_X1 U90 ( .B1(n71), .B2(n642), .C1(n163), .C2(n42), .A(n164), .ZN(n141) );
  AOI222_X1 U91 ( .A1(n165), .A2(n166), .B1(n167), .B2(n168), .C1(n169), .C2(
        n170), .ZN(n164) );
  OAI221_X1 U92 ( .B1(n68), .B2(n642), .C1(n344), .C2(n42), .A(n581), .ZN(n572) );
  AOI222_X1 U93 ( .A1(n165), .A2(n516), .B1(n167), .B2(n402), .C1(n169), .C2(
        n464), .ZN(n581) );
  OAI221_X1 U94 ( .B1(n93), .B2(n638), .C1(n81), .C2(n642), .A(n534), .ZN(n526) );
  AOI222_X1 U95 ( .A1(n169), .A2(n168), .B1(n493), .B2(n129), .C1(n167), .C2(
        n355), .ZN(n534) );
  OAI221_X1 U96 ( .B1(n97), .B2(n638), .C1(n84), .C2(n642), .A(n520), .ZN(n511) );
  AOI222_X1 U97 ( .A1(n169), .A2(n402), .B1(n493), .B2(n134), .C1(n167), .C2(
        n403), .ZN(n520) );
  OAI221_X1 U98 ( .B1(n101), .B2(n638), .C1(n196), .C2(n642), .A(n507), .ZN(
        n498) );
  AOI222_X1 U99 ( .A1(n169), .A2(n453), .B1(n493), .B2(n382), .C1(n167), .C2(
        n506), .ZN(n507) );
  NOR2_X1 U100 ( .A1(n613), .A2(n8), .ZN(n382) );
  OAI221_X1 U101 ( .B1(n127), .B2(n161), .C1(n116), .C2(n158), .A(n162), .ZN(
        n503) );
  OAI221_X1 U102 ( .B1(n237), .B2(n160), .C1(n90), .C2(n161), .A(n162), .ZN(
        n235) );
  OAI221_X1 U103 ( .B1(n110), .B2(n160), .C1(n93), .C2(n161), .A(n162), .ZN(
        n220) );
  OAI221_X1 U104 ( .B1(n113), .B2(n160), .C1(n97), .C2(n161), .A(n162), .ZN(
        n208) );
  OAI221_X1 U105 ( .B1(n197), .B2(n160), .C1(n101), .C2(n161), .A(n162), .ZN(
        n194) );
  OAI221_X1 U106 ( .B1(n181), .B2(n160), .C1(n106), .C2(n161), .A(n162), .ZN(
        n179) );
  OAI221_X1 U107 ( .B1(n159), .B2(n160), .C1(n109), .C2(n161), .A(n162), .ZN(
        n155) );
  OAI221_X1 U108 ( .B1(n347), .B2(n160), .C1(n112), .C2(n161), .A(n162), .ZN(
        n577) );
  OAI221_X1 U109 ( .B1(n336), .B2(n160), .C1(n116), .C2(n161), .A(n162), .ZN(
        n560) );
  OAI221_X1 U110 ( .B1(n323), .B2(n160), .C1(n118), .C2(n161), .A(n162), .ZN(
        n548) );
  INV_X1 U111 ( .A(n370), .ZN(n118) );
  OAI221_X1 U112 ( .B1(n312), .B2(n160), .C1(n121), .C2(n161), .A(n162), .ZN(
        n531) );
  INV_X1 U113 ( .A(n355), .ZN(n121) );
  OAI221_X1 U114 ( .B1(n286), .B2(n160), .C1(n124), .C2(n161), .A(n162), .ZN(
        n517) );
  INV_X1 U115 ( .A(n403), .ZN(n124) );
  AND2_X1 U116 ( .A1(n491), .A2(n633), .ZN(n276) );
  AOI22_X1 U117 ( .A1(n480), .A2(n39), .B1(n43), .B2(n64), .ZN(n587) );
  INV_X1 U118 ( .A(n601), .ZN(n64) );
  AOI221_X1 U119 ( .B1(n4), .B2(n602), .C1(n454), .C2(n184), .A(n603), .ZN(
        n601) );
  OAI22_X1 U120 ( .A1(n618), .A2(n639), .B1(n65), .B2(n646), .ZN(n603) );
  AOI22_X1 U121 ( .A1(n420), .A2(n2), .B1(n58), .B2(n262), .ZN(n214) );
  AOI22_X1 U122 ( .A1(n407), .A2(n5), .B1(n52), .B2(n262), .ZN(n202) );
  AOI22_X1 U123 ( .A1(n389), .A2(n3), .B1(n390), .B2(n262), .ZN(n188) );
  AOI22_X1 U124 ( .A1(n168), .A2(n3), .B1(n355), .B2(n262), .ZN(n413) );
  AOI22_X1 U125 ( .A1(n402), .A2(n5), .B1(n403), .B2(n262), .ZN(n396) );
  AOI22_X1 U126 ( .A1(n452), .A2(n4), .B1(n453), .B2(n262), .ZN(n449) );
  AOI22_X1 U127 ( .A1(n370), .A2(n4), .B1(n320), .B2(n262), .ZN(n182) );
  AOI22_X1 U128 ( .A1(n355), .A2(n2), .B1(n129), .B2(n262), .ZN(n163) );
  AOI22_X1 U129 ( .A1(n403), .A2(n4), .B1(n134), .B2(n262), .ZN(n344) );
  AOI21_X1 U130 ( .B1(n148), .B2(n232), .A(n150), .ZN(n231) );
  OAI21_X1 U131 ( .B1(n233), .B2(n152), .A(n153), .ZN(n232) );
  AOI211_X1 U132 ( .C1(n644), .C2(n234), .A(n235), .B(n236), .ZN(n233) );
  OAI22_X1 U133 ( .A1(n65), .A2(n157), .B1(n78), .B2(n158), .ZN(n236) );
  AOI21_X1 U134 ( .B1(n148), .B2(n217), .A(n150), .ZN(n216) );
  OAI21_X1 U135 ( .B1(n218), .B2(n152), .A(n153), .ZN(n217) );
  AOI211_X1 U136 ( .C1(n644), .C2(n219), .A(n220), .B(n221), .ZN(n218) );
  OAI22_X1 U137 ( .A1(n71), .A2(n157), .B1(n81), .B2(n158), .ZN(n221) );
  AOI21_X1 U138 ( .B1(n148), .B2(n205), .A(n150), .ZN(n204) );
  OAI21_X1 U139 ( .B1(n206), .B2(n152), .A(n153), .ZN(n205) );
  AOI211_X1 U140 ( .C1(n644), .C2(n207), .A(n208), .B(n209), .ZN(n206) );
  OAI22_X1 U141 ( .A1(n68), .A2(n157), .B1(n84), .B2(n158), .ZN(n209) );
  AOI21_X1 U142 ( .B1(n148), .B2(n191), .A(n150), .ZN(n190) );
  OAI21_X1 U143 ( .B1(n192), .B2(n152), .A(n153), .ZN(n191) );
  AOI211_X1 U144 ( .C1(n644), .C2(n193), .A(n194), .B(n195), .ZN(n192) );
  OAI22_X1 U145 ( .A1(n75), .A2(n157), .B1(n196), .B2(n158), .ZN(n195) );
  AOI21_X1 U146 ( .B1(n148), .B2(n176), .A(n150), .ZN(n175) );
  OAI21_X1 U147 ( .B1(n177), .B2(n152), .A(n153), .ZN(n176) );
  AOI211_X1 U148 ( .C1(n644), .C2(n178), .A(n179), .B(n180), .ZN(n177) );
  OAI22_X1 U149 ( .A1(n78), .A2(n157), .B1(n90), .B2(n158), .ZN(n180) );
  AOI21_X1 U150 ( .B1(n148), .B2(n149), .A(n150), .ZN(n145) );
  OAI21_X1 U151 ( .B1(n151), .B2(n152), .A(n153), .ZN(n149) );
  AOI211_X1 U152 ( .C1(n644), .C2(n154), .A(n155), .B(n156), .ZN(n151) );
  OAI22_X1 U153 ( .A1(n81), .A2(n157), .B1(n93), .B2(n158), .ZN(n156) );
  AOI21_X1 U154 ( .B1(n148), .B2(n575), .A(n150), .ZN(n574) );
  OAI21_X1 U155 ( .B1(n576), .B2(n152), .A(n153), .ZN(n575) );
  AOI211_X1 U156 ( .C1(n644), .C2(n305), .A(n577), .B(n578), .ZN(n576) );
  OAI22_X1 U157 ( .A1(n84), .A2(n157), .B1(n97), .B2(n158), .ZN(n578) );
  AOI21_X1 U158 ( .B1(n148), .B2(n558), .A(n150), .ZN(n557) );
  OAI21_X1 U159 ( .B1(n559), .B2(n152), .A(n153), .ZN(n558) );
  AOI211_X1 U160 ( .C1(n644), .C2(n261), .A(n560), .B(n561), .ZN(n559) );
  OAI22_X1 U161 ( .A1(n196), .A2(n157), .B1(n101), .B2(n158), .ZN(n561) );
  AOI21_X1 U162 ( .B1(n148), .B2(n546), .A(n150), .ZN(n545) );
  OAI21_X1 U163 ( .B1(n547), .B2(n152), .A(n153), .ZN(n546) );
  AOI211_X1 U164 ( .C1(n644), .C2(n184), .A(n548), .B(n549), .ZN(n547) );
  OAI22_X1 U165 ( .A1(n90), .A2(n157), .B1(n106), .B2(n158), .ZN(n549) );
  AOI21_X1 U166 ( .B1(n148), .B2(n529), .A(n150), .ZN(n528) );
  OAI21_X1 U167 ( .B1(n530), .B2(n152), .A(n153), .ZN(n529) );
  AOI211_X1 U168 ( .C1(n644), .C2(n166), .A(n531), .B(n532), .ZN(n530) );
  OAI22_X1 U169 ( .A1(n93), .A2(n157), .B1(n109), .B2(n158), .ZN(n532) );
  AOI21_X1 U170 ( .B1(n148), .B2(n514), .A(n150), .ZN(n513) );
  OAI21_X1 U171 ( .B1(n515), .B2(n152), .A(n153), .ZN(n514) );
  AOI211_X1 U172 ( .C1(n644), .C2(n516), .A(n517), .B(n518), .ZN(n515) );
  OAI22_X1 U173 ( .A1(n97), .A2(n157), .B1(n112), .B2(n158), .ZN(n518) );
  AOI21_X1 U174 ( .B1(n283), .B2(n415), .A(n285), .ZN(n414) );
  OAI21_X1 U175 ( .B1(n110), .B2(n287), .A(n288), .ZN(n415) );
  AOI21_X1 U176 ( .B1(n283), .B2(n398), .A(n285), .ZN(n397) );
  OAI21_X1 U177 ( .B1(n113), .B2(n287), .A(n288), .ZN(n398) );
  AOI21_X1 U178 ( .B1(n283), .B2(n385), .A(n285), .ZN(n384) );
  OAI21_X1 U179 ( .B1(n197), .B2(n287), .A(n288), .ZN(n385) );
  AOI21_X1 U180 ( .B1(n283), .B2(n369), .A(n285), .ZN(n368) );
  OAI21_X1 U181 ( .B1(n181), .B2(n287), .A(n288), .ZN(n369) );
  AOI21_X1 U182 ( .B1(n283), .B2(n335), .A(n285), .ZN(n334) );
  OAI21_X1 U183 ( .B1(n336), .B2(n287), .A(n288), .ZN(n335) );
  OAI211_X1 U184 ( .C1(n127), .C2(n646), .A(n401), .B(n449), .ZN(n257) );
  AOI21_X1 U185 ( .B1(n320), .B2(n4), .A(n519), .ZN(n323) );
  AOI21_X1 U186 ( .B1(n506), .B2(n5), .A(n519), .ZN(n336) );
  NAND2_X1 U187 ( .A1(n484), .A2(n633), .ZN(n249) );
  OAI21_X1 U188 ( .B1(n417), .B2(n637), .A(n471), .ZN(n440) );
  OAI21_X1 U189 ( .B1(n400), .B2(n637), .A(n461), .ZN(n302) );
  NOR2_X1 U190 ( .A1(n613), .A2(n484), .ZN(n483) );
  OAI21_X1 U191 ( .B1(n412), .B2(n637), .A(n471), .ZN(n434) );
  OAI21_X1 U192 ( .B1(n395), .B2(n637), .A(n461), .ZN(n297) );
  OAI21_X1 U193 ( .B1(n412), .B2(n646), .A(n413), .ZN(n223) );
  OAI21_X1 U194 ( .B1(n395), .B2(n646), .A(n396), .ZN(n211) );
  OAI21_X1 U195 ( .B1(n333), .B2(n647), .A(n449), .ZN(n246) );
  OAI21_X1 U196 ( .B1(n482), .B2(n281), .A(n282), .ZN(n479) );
  AOI21_X1 U197 ( .B1(n283), .B2(n485), .A(n285), .ZN(n482) );
  OAI21_X1 U198 ( .B1(n89), .B2(n287), .A(n288), .ZN(n485) );
  INV_X1 U199 ( .A(n480), .ZN(n89) );
  OAI21_X1 U200 ( .B1(n472), .B2(n281), .A(n282), .ZN(n470) );
  AOI21_X1 U201 ( .B1(n283), .B2(n473), .A(n285), .ZN(n472) );
  OAI21_X1 U202 ( .B1(n94), .B2(n287), .A(n288), .ZN(n473) );
  INV_X1 U203 ( .A(n440), .ZN(n94) );
  OAI21_X1 U204 ( .B1(n462), .B2(n281), .A(n282), .ZN(n460) );
  AOI21_X1 U205 ( .B1(n283), .B2(n463), .A(n285), .ZN(n462) );
  OAI21_X1 U206 ( .B1(n98), .B2(n287), .A(n288), .ZN(n463) );
  INV_X1 U207 ( .A(n302), .ZN(n98) );
  OAI21_X1 U208 ( .B1(n450), .B2(n281), .A(n282), .ZN(n448) );
  AOI21_X1 U209 ( .B1(n283), .B2(n451), .A(n285), .ZN(n450) );
  OAI21_X1 U210 ( .B1(n102), .B2(n287), .A(n288), .ZN(n451) );
  INV_X1 U211 ( .A(n257), .ZN(n102) );
  OAI21_X1 U212 ( .B1(n425), .B2(n281), .A(n282), .ZN(n424) );
  AOI21_X1 U213 ( .B1(n283), .B2(n426), .A(n285), .ZN(n425) );
  OAI21_X1 U214 ( .B1(n237), .B2(n287), .A(n288), .ZN(n426) );
  OAI21_X1 U215 ( .B1(n357), .B2(n281), .A(n282), .ZN(n354) );
  AOI21_X1 U216 ( .B1(n283), .B2(n358), .A(n285), .ZN(n357) );
  OAI21_X1 U217 ( .B1(n159), .B2(n287), .A(n288), .ZN(n358) );
  OAI21_X1 U218 ( .B1(n345), .B2(n281), .A(n282), .ZN(n343) );
  AOI21_X1 U219 ( .B1(n283), .B2(n346), .A(n285), .ZN(n345) );
  OAI21_X1 U220 ( .B1(n347), .B2(n287), .A(n288), .ZN(n346) );
  OAI21_X1 U221 ( .B1(n321), .B2(n281), .A(n282), .ZN(n319) );
  AOI21_X1 U222 ( .B1(n283), .B2(n322), .A(n285), .ZN(n321) );
  OAI21_X1 U223 ( .B1(n323), .B2(n287), .A(n288), .ZN(n322) );
  OAI21_X1 U224 ( .B1(n310), .B2(n281), .A(n282), .ZN(n309) );
  AOI21_X1 U225 ( .B1(n283), .B2(n311), .A(n285), .ZN(n310) );
  OAI21_X1 U226 ( .B1(n312), .B2(n287), .A(n288), .ZN(n311) );
  OAI21_X1 U227 ( .B1(n280), .B2(n281), .A(n282), .ZN(n277) );
  AOI21_X1 U228 ( .B1(n283), .B2(n284), .A(n285), .ZN(n280) );
  OAI21_X1 U229 ( .B1(n286), .B2(n287), .A(n288), .ZN(n284) );
  AOI22_X1 U230 ( .A1(n246), .A2(n39), .B1(n43), .B2(n247), .ZN(n245) );
  AOI22_X1 U231 ( .A1(n434), .A2(n39), .B1(n42), .B2(n435), .ZN(n433) );
  AOI22_X1 U232 ( .A1(n297), .A2(n39), .B1(n42), .B2(n298), .ZN(n296) );
  INV_X1 U233 ( .A(n452), .ZN(n101) );
  INV_X1 U234 ( .A(n464), .ZN(n97) );
  INV_X1 U235 ( .A(n170), .ZN(n93) );
  INV_X1 U236 ( .A(n186), .ZN(n90) );
  INV_X1 U237 ( .A(n516), .ZN(n84) );
  INV_X1 U238 ( .A(n166), .ZN(n81) );
  NOR2_X1 U239 ( .A1(n266), .A2(n8), .ZN(n580) );
  AOI21_X1 U240 ( .B1(n251), .B2(n438), .A(n253), .ZN(n437) );
  OAI21_X1 U241 ( .B1(n439), .B2(n255), .A(n256), .ZN(n438) );
  AOI22_X1 U242 ( .A1(n435), .A2(n40), .B1(B[4]), .B2(n440), .ZN(n439) );
  AOI21_X1 U243 ( .B1(n251), .B2(n300), .A(n253), .ZN(n299) );
  OAI21_X1 U244 ( .B1(n301), .B2(n255), .A(n256), .ZN(n300) );
  AOI22_X1 U245 ( .A1(n298), .A2(n40), .B1(B[4]), .B2(n302), .ZN(n301) );
  AOI21_X1 U246 ( .B1(n251), .B2(n252), .A(n253), .ZN(n248) );
  OAI21_X1 U247 ( .B1(n254), .B2(n255), .A(n256), .ZN(n252) );
  AOI22_X1 U248 ( .A1(n247), .A2(n40), .B1(B[4]), .B2(n257), .ZN(n254) );
  BUF_X1 U249 ( .A(n356), .Z(n2) );
  BUF_X1 U250 ( .A(n356), .Z(n3) );
  INV_X1 U251 ( .A(n293), .ZN(n52) );
  INV_X1 U252 ( .A(n184), .ZN(n78) );
  INV_X1 U253 ( .A(n506), .ZN(n127) );
  INV_X1 U254 ( .A(n185), .ZN(n106) );
  INV_X1 U255 ( .A(n412), .ZN(n129) );
  INV_X1 U256 ( .A(n395), .ZN(n134) );
  INV_X1 U257 ( .A(n390), .ZN(n46) );
  BUF_X1 U258 ( .A(n356), .Z(n4) );
  BUF_X1 U259 ( .A(n356), .Z(n5) );
  INV_X1 U260 ( .A(n453), .ZN(n116) );
  INV_X1 U261 ( .A(n154), .ZN(n71) );
  INV_X1 U262 ( .A(n305), .ZN(n68) );
  INV_X1 U263 ( .A(n178), .ZN(n65) );
  INV_X1 U265 ( .A(n168), .ZN(n109) );
  INV_X1 U266 ( .A(n402), .ZN(n112) );
  INV_X1 U268 ( .A(n261), .ZN(n75) );
  INV_X1 U270 ( .A(n419), .ZN(n82) );
  INV_X1 U271 ( .A(n406), .ZN(n85) );
  INV_X1 U272 ( .A(n388), .ZN(n87) );
  BUF_X1 U273 ( .A(n44), .Z(n42) );
  INV_X1 U274 ( .A(n362), .ZN(n58) );
  INV_X1 U275 ( .A(n474), .ZN(n62) );
  INV_X1 U276 ( .A(n465), .ZN(n73) );
  INV_X1 U277 ( .A(n455), .ZN(n76) );
  INV_X1 U278 ( .A(n267), .ZN(n8) );
  BUF_X1 U279 ( .A(n44), .Z(n43) );
  BUF_X1 U280 ( .A(n44), .Z(n40) );
  INV_X1 U281 ( .A(n417), .ZN(n130) );
  INV_X1 U282 ( .A(n400), .ZN(n135) );
  BUF_X1 U283 ( .A(n44), .Z(n41) );
  INV_X1 U284 ( .A(n373), .ZN(n79) );
  INV_X1 U285 ( .A(n420), .ZN(n132) );
  INV_X1 U286 ( .A(n407), .ZN(n614) );
  INV_X1 U287 ( .A(n389), .ZN(n616) );
  INV_X1 U288 ( .A(n429), .ZN(n63) );
  INV_X1 U289 ( .A(n372), .ZN(n91) );
  INV_X1 U290 ( .A(n361), .ZN(n95) );
  INV_X1 U291 ( .A(n350), .ZN(n99) );
  INV_X1 U292 ( .A(n339), .ZN(n104) );
  AND2_X1 U293 ( .A1(n238), .A2(n401), .ZN(n237) );
  INV_X1 U294 ( .A(n234), .ZN(n618) );
  INV_X1 U295 ( .A(n416), .ZN(n110) );
  OAI211_X1 U296 ( .C1(n417), .C2(n646), .A(n401), .B(n413), .ZN(n416) );
  INV_X1 U297 ( .A(n399), .ZN(n113) );
  OAI211_X1 U298 ( .C1(n400), .C2(n646), .A(n401), .B(n396), .ZN(n399) );
  INV_X1 U299 ( .A(n381), .ZN(n115) );
  AOI21_X1 U300 ( .B1(n260), .B2(n382), .A(n383), .ZN(n381) );
  OR4_X1 U301 ( .A1(B[21]), .A2(B[20]), .A3(B[19]), .A4(B[18]), .ZN(n598) );
  OAI22_X1 U302 ( .A1(n88), .A2(n1), .B1(n86), .B2(n8), .ZN(n568) );
  AOI222_X1 U303 ( .A1(n11), .A2(A[1]), .B1(A[0]), .B2(n18), .C1(n7), .C2(A[2]), .ZN(n293) );
  AOI221_X1 U304 ( .B1(n31), .B2(A[6]), .C1(n20), .C2(A[7]), .A(n525), .ZN(
        n363) );
  OAI22_X1 U305 ( .A1(n623), .A2(n1), .B1(n624), .B2(n8), .ZN(n525) );
  AOI221_X1 U306 ( .B1(n30), .B2(A[7]), .C1(n20), .C2(A[8]), .A(n570), .ZN(
        n405) );
  OAI22_X1 U307 ( .A1(n624), .A2(n1), .B1(n66), .B2(n8), .ZN(n570) );
  AOI221_X1 U308 ( .B1(n31), .B2(A[8]), .C1(n21), .C2(A[9]), .A(n552), .ZN(
        n387) );
  OAI22_X1 U309 ( .A1(n66), .A2(n1), .B1(n74), .B2(n8), .ZN(n552) );
  AOI221_X1 U310 ( .B1(n30), .B2(A[5]), .C1(n20), .C2(A[6]), .A(n541), .ZN(
        n376) );
  OAI22_X1 U311 ( .A1(n622), .A2(n1), .B1(n623), .B2(n8), .ZN(n541) );
  OAI221_X1 U312 ( .B1(n29), .B2(n613), .C1(n17), .C2(n266), .A(n609), .ZN(
        n320) );
  AOI22_X1 U313 ( .A1(A[29]), .A2(n10), .B1(A[28]), .B2(n267), .ZN(n609) );
  OAI221_X1 U314 ( .B1(n27), .B2(n128), .C1(n15), .C2(n126), .A(n535), .ZN(
        n355) );
  AOI22_X1 U315 ( .A1(A[26]), .A2(n11), .B1(A[25]), .B2(n6), .ZN(n535) );
  OAI221_X1 U316 ( .B1(n28), .B2(n131), .C1(n16), .C2(n128), .A(n585), .ZN(
        n403) );
  AOI22_X1 U317 ( .A1(A[27]), .A2(n9), .B1(A[26]), .B2(n267), .ZN(n585) );
  OR3_X1 U318 ( .A1(B[22]), .A2(B[24]), .A3(B[23]), .ZN(n594) );
  NAND3_X1 U319 ( .A1(n489), .A2(n629), .A3(n600), .ZN(n152) );
  NOR3_X1 U320 ( .A1(B[12]), .A2(B[14]), .A3(B[13]), .ZN(n600) );
  NAND3_X1 U321 ( .A1(n592), .A2(n632), .A3(n599), .ZN(n146) );
  INV_X1 U322 ( .A(B[22]), .ZN(n632) );
  NOR3_X1 U323 ( .A1(B[23]), .A2(B[25]), .A3(B[24]), .ZN(n599) );
  NAND2_X1 U324 ( .A1(A[31]), .A2(n648), .ZN(n162) );
  OAI221_X1 U325 ( .B1(n29), .B2(n86), .C1(n17), .C2(n83), .A(n606), .ZN(n184)
         );
  AOI22_X1 U326 ( .A1(A[13]), .A2(n10), .B1(A[12]), .B2(n267), .ZN(n606) );
  OAI221_X1 U327 ( .B1(n29), .B2(n126), .C1(n17), .C2(n123), .A(n608), .ZN(
        n370) );
  AOI22_X1 U328 ( .A1(A[25]), .A2(n10), .B1(A[24]), .B2(n267), .ZN(n608) );
  NAND2_X1 U329 ( .A1(n488), .A2(n489), .ZN(n287) );
  OAI221_X1 U330 ( .B1(n27), .B2(n117), .C1(n15), .C2(n114), .A(n536), .ZN(
        n168) );
  AOI22_X1 U331 ( .A1(A[22]), .A2(n9), .B1(A[21]), .B2(n7), .ZN(n536) );
  OAI221_X1 U332 ( .B1(n28), .B2(n120), .C1(n16), .C2(n117), .A(n583), .ZN(
        n402) );
  AOI22_X1 U333 ( .A1(A[23]), .A2(n9), .B1(A[22]), .B2(n267), .ZN(n583) );
  AOI221_X1 U334 ( .B1(A[1]), .B2(n32), .C1(A[2]), .C2(n18), .A(n540), .ZN(
        n374) );
  OAI22_X1 U335 ( .A1(n615), .A2(n1), .B1(n617), .B2(n8), .ZN(n540) );
  NAND2_X1 U336 ( .A1(A[31]), .A2(n152), .ZN(n153) );
  NAND2_X1 U337 ( .A1(A[31]), .A2(n146), .ZN(n147) );
  NOR2_X2 U338 ( .A1(n612), .A2(n591), .ZN(n144) );
  OAI221_X1 U339 ( .B1(n28), .B2(n266), .C1(n16), .C2(n131), .A(n564), .ZN(
        n506) );
  AOI22_X1 U340 ( .A1(A[28]), .A2(n9), .B1(A[27]), .B2(n7), .ZN(n564) );
  OAI221_X1 U341 ( .B1(n28), .B2(n123), .C1(n16), .C2(n120), .A(n565), .ZN(
        n453) );
  AOI22_X1 U342 ( .A1(A[24]), .A2(n9), .B1(A[23]), .B2(n7), .ZN(n565) );
  NOR2_X2 U343 ( .A1(n647), .A2(B[2]), .ZN(n260) );
  OAI221_X1 U344 ( .B1(n26), .B2(n114), .C1(n14), .C2(n111), .A(n611), .ZN(
        n185) );
  AOI22_X1 U345 ( .A1(A[21]), .A2(n11), .B1(A[20]), .B2(n6), .ZN(n611) );
  AOI222_X1 U346 ( .A1(n429), .A2(n5), .B1(n620), .B2(n262), .C1(n227), .C2(
        B[3]), .ZN(n327) );
  INV_X1 U347 ( .A(n376), .ZN(n620) );
  OAI221_X1 U348 ( .B1(n26), .B2(n77), .C1(n15), .C2(n74), .A(n444), .ZN(n154)
         );
  AOI22_X1 U349 ( .A1(A[10]), .A2(n11), .B1(A[9]), .B2(n6), .ZN(n444) );
  OAI221_X1 U350 ( .B1(n29), .B2(n80), .C1(n16), .C2(n77), .A(n586), .ZN(n305)
         );
  AOI22_X1 U351 ( .A1(A[11]), .A2(n10), .B1(A[10]), .B2(n267), .ZN(n586) );
  OAI221_X1 U352 ( .B1(n28), .B2(n83), .C1(n16), .C2(n80), .A(n567), .ZN(n261)
         );
  AOI22_X1 U353 ( .A1(A[12]), .A2(n9), .B1(A[11]), .B2(n7), .ZN(n567) );
  OAI221_X1 U354 ( .B1(n26), .B2(n623), .C1(n14), .C2(n622), .A(n443), .ZN(
        n219) );
  AOI22_X1 U355 ( .A1(A[6]), .A2(n11), .B1(A[5]), .B2(n7), .ZN(n443) );
  OAI221_X1 U356 ( .B1(n26), .B2(n624), .C1(n14), .C2(n623), .A(n306), .ZN(
        n207) );
  AOI22_X1 U357 ( .A1(A[7]), .A2(n11), .B1(A[6]), .B2(n6), .ZN(n306) );
  OAI221_X1 U358 ( .B1(n27), .B2(n66), .C1(n15), .C2(n624), .A(n265), .ZN(n193) );
  AOI22_X1 U359 ( .A1(A[8]), .A2(n10), .B1(A[7]), .B2(n6), .ZN(n265) );
  OAI221_X1 U360 ( .B1(n29), .B2(n100), .C1(n17), .C2(n96), .A(n610), .ZN(n186) );
  AOI22_X1 U361 ( .A1(A[17]), .A2(n10), .B1(A[16]), .B2(n267), .ZN(n610) );
  OAI221_X1 U362 ( .B1(n29), .B2(n74), .C1(n17), .C2(n66), .A(n604), .ZN(n178)
         );
  AOI22_X1 U363 ( .A1(A[9]), .A2(n10), .B1(A[8]), .B2(n267), .ZN(n604) );
  OAI221_X1 U364 ( .B1(n27), .B2(n88), .C1(n15), .C2(n86), .A(n537), .ZN(n166)
         );
  AOI22_X1 U365 ( .A1(A[14]), .A2(n11), .B1(A[13]), .B2(n7), .ZN(n537) );
  OAI221_X1 U366 ( .B1(n28), .B2(n92), .C1(n16), .C2(n88), .A(n584), .ZN(n516)
         );
  AOI22_X1 U367 ( .A1(A[15]), .A2(n9), .B1(A[14]), .B2(n7), .ZN(n584) );
  OAI221_X1 U368 ( .B1(n27), .B2(n80), .C1(n15), .C2(n83), .A(n494), .ZN(n373)
         );
  AOI22_X1 U369 ( .A1(A[15]), .A2(n9), .B1(A[16]), .B2(n6), .ZN(n494) );
  OAI221_X1 U370 ( .B1(n27), .B2(n133), .C1(n15), .C2(n615), .A(n523), .ZN(
        n420) );
  AOI22_X1 U371 ( .A1(A[4]), .A2(n10), .B1(A[5]), .B2(n7), .ZN(n523) );
  OAI221_X1 U372 ( .B1(n28), .B2(n615), .C1(n16), .C2(n617), .A(n571), .ZN(
        n407) );
  AOI22_X1 U373 ( .A1(A[5]), .A2(n9), .B1(A[6]), .B2(n7), .ZN(n571) );
  OAI221_X1 U374 ( .B1(n28), .B2(n617), .C1(n16), .C2(n619), .A(n554), .ZN(
        n389) );
  AOI22_X1 U375 ( .A1(A[6]), .A2(n9), .B1(A[7]), .B2(n7), .ZN(n554) );
  OAI221_X1 U376 ( .B1(n49), .B2(n29), .C1(n103), .C2(n14), .A(n553), .ZN(n390) );
  AOI22_X1 U377 ( .A1(A[2]), .A2(n9), .B1(A[3]), .B2(n7), .ZN(n553) );
  OAI221_X1 U378 ( .B1(n28), .B2(n624), .C1(n16), .C2(n66), .A(n542), .ZN(n429) );
  AOI22_X1 U379 ( .A1(A[11]), .A2(n9), .B1(A[12]), .B2(n7), .ZN(n542) );
  OAI221_X1 U380 ( .B1(n28), .B2(n111), .C1(n16), .C2(n108), .A(n566), .ZN(
        n452) );
  AOI22_X1 U381 ( .A1(A[20]), .A2(n9), .B1(A[19]), .B2(n7), .ZN(n566) );
  OAI221_X1 U382 ( .B1(n28), .B2(n105), .C1(n16), .C2(n100), .A(n538), .ZN(
        n170) );
  AOI22_X1 U383 ( .A1(A[18]), .A2(n9), .B1(A[17]), .B2(n7), .ZN(n538) );
  OAI221_X1 U384 ( .B1(n28), .B2(n108), .C1(n16), .C2(n105), .A(n582), .ZN(
        n464) );
  AOI22_X1 U385 ( .A1(A[19]), .A2(n10), .B1(A[18]), .B2(n7), .ZN(n582) );
  INV_X1 U386 ( .A(A[31]), .ZN(n613) );
  AOI22_X1 U387 ( .A1(n267), .A2(A[1]), .B1(n11), .B2(A[0]), .ZN(n362) );
  NAND2_X1 U389 ( .A1(B[4]), .A2(n579), .ZN(n160) );
  OAI222_X1 U390 ( .A1(n79), .A2(n636), .B1(n326), .B2(n642), .C1(n91), .C2(
        n645), .ZN(n325) );
  AOI222_X1 U391 ( .A1(A[27]), .A2(n10), .B1(A[25]), .B2(n30), .C1(A[26]), 
        .C2(n18), .ZN(n326) );
  AOI222_X1 U392 ( .A1(A[28]), .A2(n10), .B1(A[26]), .B2(n30), .C1(A[27]), 
        .C2(n19), .ZN(n316) );
  AOI222_X1 U393 ( .A1(A[29]), .A2(n11), .B1(A[27]), .B2(n32), .C1(A[28]), 
        .C2(n18), .ZN(n292) );
  AOI222_X1 U394 ( .A1(A[30]), .A2(n11), .B1(A[28]), .B2(n30), .C1(A[29]), 
        .C2(n22), .ZN(n273) );
  AOI21_X1 U395 ( .B1(A[31]), .B2(B[11]), .A(n487), .ZN(n256) );
  AOI21_X1 U396 ( .B1(A[31]), .B2(B[25]), .A(n483), .ZN(n250) );
  OAI222_X1 U397 ( .A1(n171), .A2(n36), .B1(n55), .B2(n626), .C1(n623), .C2(
        n33), .ZN(RES[8]) );
  INV_X1 U398 ( .A(n172), .ZN(n55) );
  AOI221_X1 U399 ( .B1(n140), .B2(n173), .C1(n142), .C2(n174), .A(n144), .ZN(
        n171) );
  OAI21_X1 U400 ( .B1(n175), .B2(n146), .A(n147), .ZN(n174) );
  OAI222_X1 U401 ( .A1(n187), .A2(n36), .B1(n188), .B2(n626), .C1(n622), .C2(
        n33), .ZN(RES[7]) );
  AOI221_X1 U402 ( .B1(n140), .B2(n61), .C1(n142), .C2(n189), .A(n144), .ZN(
        n187) );
  INV_X1 U403 ( .A(n198), .ZN(n61) );
  OAI21_X1 U404 ( .B1(n190), .B2(n146), .A(n147), .ZN(n189) );
  OAI222_X1 U405 ( .A1(n136), .A2(n36), .B1(n59), .B2(n626), .C1(n624), .C2(
        n33), .ZN(RES[9]) );
  INV_X1 U406 ( .A(n139), .ZN(n59) );
  AOI221_X1 U407 ( .B1(n140), .B2(n141), .C1(n142), .C2(n143), .A(n144), .ZN(
        n136) );
  OAI21_X1 U408 ( .B1(n145), .B2(n146), .A(n147), .ZN(n143) );
  OAI222_X1 U409 ( .A1(n539), .A2(n36), .B1(n327), .B2(n626), .C1(n77), .C2(
        n35), .ZN(RES[12]) );
  AOI221_X1 U410 ( .B1(n140), .B2(n543), .C1(n142), .C2(n544), .A(n144), .ZN(
        n539) );
  OAI21_X1 U411 ( .B1(n545), .B2(n146), .A(n147), .ZN(n544) );
  OAI221_X1 U412 ( .B1(n90), .B2(n638), .C1(n78), .C2(n642), .A(n550), .ZN(
        n543) );
  OAI222_X1 U413 ( .A1(n521), .A2(n36), .B1(n57), .B2(n626), .C1(n80), .C2(n35), .ZN(RES[13]) );
  INV_X1 U414 ( .A(n314), .ZN(n57) );
  AOI221_X1 U415 ( .B1(n140), .B2(n526), .C1(n142), .C2(n527), .A(n144), .ZN(
        n521) );
  OAI21_X1 U416 ( .B1(n528), .B2(n146), .A(n147), .ZN(n527) );
  OAI222_X1 U417 ( .A1(n508), .A2(n36), .B1(n51), .B2(n626), .C1(n83), .C2(n35), .ZN(RES[14]) );
  INV_X1 U418 ( .A(n290), .ZN(n51) );
  AOI221_X1 U419 ( .B1(n140), .B2(n511), .C1(n142), .C2(n512), .A(n144), .ZN(
        n508) );
  OAI21_X1 U420 ( .B1(n513), .B2(n146), .A(n147), .ZN(n512) );
  OAI222_X1 U421 ( .A1(n551), .A2(n36), .B1(n45), .B2(n626), .C1(n74), .C2(n35), .ZN(RES[11]) );
  INV_X1 U422 ( .A(n337), .ZN(n45) );
  AOI221_X1 U423 ( .B1(n140), .B2(n555), .C1(n142), .C2(n556), .A(n144), .ZN(
        n551) );
  OAI21_X1 U424 ( .B1(n557), .B2(n146), .A(n147), .ZN(n556) );
  OAI222_X1 U425 ( .A1(n495), .A2(n36), .B1(n47), .B2(n626), .C1(n86), .C2(n35), .ZN(RES[15]) );
  INV_X1 U426 ( .A(n271), .ZN(n47) );
  AOI221_X1 U427 ( .B1(n140), .B2(n498), .C1(n142), .C2(n499), .A(n144), .ZN(
        n495) );
  OAI21_X1 U429 ( .B1(n500), .B2(n146), .A(n147), .ZN(n499) );
  OAI222_X1 U430 ( .A1(n569), .A2(n36), .B1(n53), .B2(n626), .C1(n66), .C2(n35), .ZN(RES[10]) );
  INV_X1 U431 ( .A(n348), .ZN(n53) );
  AOI221_X1 U432 ( .B1(n140), .B2(n572), .C1(n142), .C2(n573), .A(n144), .ZN(
        n569) );
  OAI21_X1 U433 ( .B1(n574), .B2(n146), .A(n147), .ZN(n573) );
  OAI222_X1 U434 ( .A1(n201), .A2(n36), .B1(n202), .B2(n626), .C1(n621), .C2(
        n33), .ZN(RES[6]) );
  AOI221_X1 U435 ( .B1(n140), .B2(n67), .C1(n142), .C2(n203), .A(n144), .ZN(
        n201) );
  INV_X1 U436 ( .A(n210), .ZN(n67) );
  OAI21_X1 U437 ( .B1(n204), .B2(n146), .A(n147), .ZN(n203) );
  OAI222_X1 U438 ( .A1(n213), .A2(n36), .B1(n214), .B2(n626), .C1(n619), .C2(
        n33), .ZN(RES[5]) );
  AOI221_X1 U439 ( .B1(n140), .B2(n70), .C1(n142), .C2(n215), .A(n144), .ZN(
        n213) );
  INV_X1 U440 ( .A(n222), .ZN(n70) );
  OAI21_X1 U441 ( .B1(n216), .B2(n146), .A(n147), .ZN(n215) );
  OAI221_X1 U442 ( .B1(n27), .B2(n83), .C1(n15), .C2(n86), .A(n476), .ZN(n419)
         );
  AOI22_X1 U443 ( .A1(A[16]), .A2(n11), .B1(A[17]), .B2(n6), .ZN(n476) );
  OAI221_X1 U444 ( .B1(n27), .B2(n86), .C1(n15), .C2(n88), .A(n467), .ZN(n406)
         );
  AOI22_X1 U445 ( .A1(A[17]), .A2(n9), .B1(A[18]), .B2(n7), .ZN(n467) );
  OAI221_X1 U446 ( .B1(n27), .B2(n88), .C1(n15), .C2(n92), .A(n457), .ZN(n388)
         );
  AOI22_X1 U447 ( .A1(A[18]), .A2(n10), .B1(A[19]), .B2(n6), .ZN(n457) );
  OAI221_X1 U448 ( .B1(n26), .B2(n92), .C1(n14), .C2(n96), .A(n430), .ZN(n372)
         );
  AOI22_X1 U449 ( .A1(A[19]), .A2(n11), .B1(A[20]), .B2(n6), .ZN(n430) );
  OAI221_X1 U450 ( .B1(n29), .B2(n622), .C1(n17), .C2(n621), .A(n605), .ZN(
        n234) );
  AOI22_X1 U451 ( .A1(A[5]), .A2(n10), .B1(A[4]), .B2(n267), .ZN(n605) );
  OAI221_X1 U452 ( .B1(n258), .B2(n643), .C1(n196), .C2(n637), .A(n259), .ZN(
        n247) );
  AOI22_X1 U453 ( .A1(n260), .A2(n261), .B1(n262), .B2(n193), .ZN(n259) );
  AOI222_X1 U454 ( .A1(A[4]), .A2(n11), .B1(A[6]), .B2(n31), .C1(A[5]), .C2(
        n19), .ZN(n258) );
  OAI221_X1 U455 ( .B1(n303), .B2(n643), .C1(n84), .C2(n637), .A(n304), .ZN(
        n298) );
  AOI22_X1 U456 ( .A1(n260), .A2(n305), .B1(n262), .B2(n207), .ZN(n304) );
  AOI222_X1 U457 ( .A1(A[3]), .A2(n10), .B1(A[5]), .B2(n32), .C1(A[4]), .C2(
        n19), .ZN(n303) );
  OAI221_X1 U458 ( .B1(n441), .B2(n643), .C1(n81), .C2(n637), .A(n442), .ZN(
        n435) );
  AOI22_X1 U459 ( .A1(n260), .A2(n154), .B1(n262), .B2(n219), .ZN(n442) );
  AOI222_X1 U460 ( .A1(A[2]), .A2(n10), .B1(A[4]), .B2(n30), .C1(A[3]), .C2(
        n20), .ZN(n441) );
  INV_X1 U462 ( .A(n228), .ZN(n626) );
  OAI221_X1 U463 ( .B1(n27), .B2(n66), .C1(n15), .C2(n74), .A(n524), .ZN(n474)
         );
  AOI22_X1 U464 ( .A1(A[12]), .A2(n11), .B1(A[13]), .B2(n7), .ZN(n524) );
  OAI221_X1 U465 ( .B1(n27), .B2(n74), .C1(n15), .C2(n77), .A(n510), .ZN(n465)
         );
  AOI22_X1 U466 ( .A1(A[13]), .A2(n9), .B1(A[14]), .B2(n6), .ZN(n510) );
  OAI221_X1 U467 ( .B1(n27), .B2(n77), .C1(n15), .C2(n80), .A(n497), .ZN(n455)
         );
  AOI22_X1 U468 ( .A1(A[14]), .A2(n10), .B1(A[15]), .B2(n7), .ZN(n497) );
  OAI221_X1 U469 ( .B1(n26), .B2(n96), .C1(n14), .C2(n100), .A(n421), .ZN(n361) );
  AOI22_X1 U470 ( .A1(A[20]), .A2(n11), .B1(A[21]), .B2(n6), .ZN(n421) );
  OAI221_X1 U471 ( .B1(n26), .B2(n100), .C1(n14), .C2(n105), .A(n408), .ZN(
        n350) );
  AOI22_X1 U472 ( .A1(A[21]), .A2(n11), .B1(A[22]), .B2(n6), .ZN(n408) );
  OAI221_X1 U473 ( .B1(n26), .B2(n105), .C1(n14), .C2(n108), .A(n391), .ZN(
        n339) );
  AOI22_X1 U474 ( .A1(A[22]), .A2(n9), .B1(A[23]), .B2(n6), .ZN(n391) );
  OAI221_X1 U475 ( .B1(n26), .B2(n108), .C1(n14), .C2(n111), .A(n377), .ZN(
        n324) );
  AOI22_X1 U476 ( .A1(A[23]), .A2(n9), .B1(A[24]), .B2(n6), .ZN(n377) );
  OAI221_X1 U477 ( .B1(n26), .B2(n111), .C1(n14), .C2(n114), .A(n364), .ZN(
        n313) );
  AOI22_X1 U478 ( .A1(A[24]), .A2(n10), .B1(A[25]), .B2(n6), .ZN(n364) );
  OAI221_X1 U479 ( .B1(n26), .B2(n114), .C1(n14), .C2(n117), .A(n351), .ZN(
        n289) );
  AOI22_X1 U480 ( .A1(A[25]), .A2(n11), .B1(A[26]), .B2(n6), .ZN(n351) );
  OAI221_X1 U481 ( .B1(n26), .B2(n117), .C1(n14), .C2(n120), .A(n340), .ZN(
        n270) );
  AOI22_X1 U482 ( .A1(A[26]), .A2(n10), .B1(A[27]), .B2(n6), .ZN(n340) );
  AOI22_X1 U483 ( .A1(n640), .A2(n506), .B1(B[2]), .B2(n382), .ZN(n333) );
  AOI21_X1 U484 ( .B1(n22), .B2(A[31]), .A(n533), .ZN(n412) );
  AOI21_X1 U485 ( .B1(n11), .B2(A[31]), .A(n580), .ZN(n395) );
  AOI21_X1 U486 ( .B1(B[1]), .B2(A[31]), .A(n533), .ZN(n417) );
  AOI21_X1 U487 ( .B1(n8), .B2(A[31]), .A(n580), .ZN(n400) );
  NOR2_X1 U488 ( .A1(n490), .A2(B[18]), .ZN(n251) );
  OAI22_X1 U489 ( .A1(B[2]), .A2(n374), .B1(n640), .B2(n375), .ZN(n227) );
  OAI221_X1 U490 ( .B1(n196), .B2(n638), .C1(n75), .C2(n642), .A(n562), .ZN(
        n555) );
  AOI221_X1 U491 ( .B1(n169), .B2(n452), .C1(n167), .C2(n453), .A(n563), .ZN(
        n562) );
  NOR3_X1 U492 ( .A1(n41), .A2(B[3]), .A3(n333), .ZN(n563) );
  NOR2_X1 U493 ( .A1(B[0]), .A2(B[1]), .ZN(n267) );
  AOI21_X1 U494 ( .B1(n634), .B2(n590), .A(n144), .ZN(n481) );
  INV_X1 U495 ( .A(n592), .ZN(n634) );
  NAND2_X1 U496 ( .A1(A[31]), .A2(n490), .ZN(n486) );
  OAI221_X1 U497 ( .B1(n225), .B2(n36), .C1(n617), .C2(n33), .A(n226), .ZN(
        RES[4]) );
  AOI221_X1 U498 ( .B1(n140), .B2(n229), .C1(n142), .C2(n230), .A(n144), .ZN(
        n225) );
  OAI21_X1 U499 ( .B1(n231), .B2(n146), .A(n147), .ZN(n230) );
  NAND2_X1 U500 ( .A1(n454), .A2(A[31]), .ZN(n401) );
  NOR2_X1 U501 ( .A1(B[2]), .A2(B[3]), .ZN(n356) );
  AOI21_X1 U502 ( .B1(n148), .B2(n501), .A(n150), .ZN(n500) );
  OAI21_X1 U503 ( .B1(n502), .B2(n152), .A(n153), .ZN(n501) );
  AOI211_X1 U504 ( .C1(B[4]), .C2(A[31]), .A(n503), .B(n504), .ZN(n502) );
  OAI22_X1 U505 ( .A1(n196), .A2(n505), .B1(n101), .B2(n157), .ZN(n504) );
  INV_X1 U506 ( .A(A[10]), .ZN(n66) );
  OAI21_X1 U507 ( .B1(n489), .B2(n613), .A(n162), .ZN(n487) );
  NOR3_X1 U508 ( .A1(n332), .A2(B[3]), .A3(n333), .ZN(n331) );
  INV_X1 U509 ( .A(B[3]), .ZN(n647) );
  INV_X1 U510 ( .A(A[11]), .ZN(n74) );
  INV_X1 U511 ( .A(A[15]), .ZN(n86) );
  INV_X1 U512 ( .A(A[9]), .ZN(n624) );
  INV_X1 U513 ( .A(A[16]), .ZN(n88) );
  BUF_X1 U514 ( .A(n137), .Z(n36) );
  BUF_X1 U515 ( .A(n137), .Z(n37) );
  NAND2_X1 U516 ( .A1(A[0]), .A2(n6), .ZN(n375) );
  INV_X1 U517 ( .A(A[23]), .ZN(n114) );
  INV_X1 U518 ( .A(A[19]), .ZN(n100) );
  INV_X1 U519 ( .A(A[24]), .ZN(n117) );
  INV_X1 U520 ( .A(A[20]), .ZN(n105) );
  INV_X1 U521 ( .A(A[21]), .ZN(n108) );
  INV_X1 U522 ( .A(A[22]), .ZN(n111) );
  INV_X1 U523 ( .A(A[8]), .ZN(n623) );
  INV_X1 U524 ( .A(A[12]), .ZN(n77) );
  INV_X1 U525 ( .A(A[13]), .ZN(n80) );
  INV_X1 U526 ( .A(A[14]), .ZN(n83) );
  INV_X1 U527 ( .A(A[30]), .ZN(n266) );
  INV_X1 U528 ( .A(A[3]), .ZN(n615) );
  OR4_X1 U529 ( .A1(B[13]), .A2(B[14]), .A3(B[12]), .A4(n596), .ZN(n490) );
  OR3_X1 U530 ( .A1(B[15]), .A2(B[17]), .A3(B[16]), .ZN(n596) );
  INV_X1 U531 ( .A(B[2]), .ZN(n640) );
  INV_X1 U532 ( .A(A[17]), .ZN(n92) );
  INV_X1 U533 ( .A(A[7]), .ZN(n622) );
  INV_X1 U534 ( .A(A[18]), .ZN(n96) );
  INV_X1 U535 ( .A(A[25]), .ZN(n120) );
  AND3_X1 U536 ( .A1(n579), .A2(n591), .A3(n597), .ZN(n445) );
  NOR3_X1 U537 ( .A1(n152), .A2(n146), .A3(n630), .ZN(n597) );
  INV_X1 U538 ( .A(n148), .ZN(n630) );
  INV_X1 U539 ( .A(A[4]), .ZN(n617) );
  INV_X1 U540 ( .A(n590), .ZN(n612) );
  INV_X1 U541 ( .A(A[27]), .ZN(n126) );
  INV_X1 U542 ( .A(A[26]), .ZN(n123) );
  INV_X1 U543 ( .A(A[6]), .ZN(n621) );
  INV_X1 U544 ( .A(A[5]), .ZN(n619) );
  INV_X1 U545 ( .A(A[28]), .ZN(n128) );
  INV_X1 U546 ( .A(A[29]), .ZN(n131) );
  INV_X1 U547 ( .A(B[25]), .ZN(n633) );
  INV_X1 U548 ( .A(A[2]), .ZN(n133) );
  AND2_X1 U549 ( .A1(n140), .A2(n199), .ZN(n278) );
  INV_X1 U550 ( .A(A[1]), .ZN(n103) );
  INV_X1 U551 ( .A(n579), .ZN(n648) );
  INV_X1 U552 ( .A(A[0]), .ZN(n49) );
  OR2_X1 U553 ( .A1(n625), .A2(B[1]), .ZN(n1) );
  NAND2_X1 U554 ( .A1(n140), .A2(n40), .ZN(n332) );
  INV_X1 U555 ( .A(n436), .ZN(n627) );
  NAND2_X1 U556 ( .A1(B[1]), .A2(B[0]), .ZN(n263) );
  NAND2_X1 U557 ( .A1(B[1]), .A2(n625), .ZN(n264) );
  INV_X1 U558 ( .A(B[11]), .ZN(n629) );
  INV_X1 U559 ( .A(B[18]), .ZN(n631) );
  AND2_X1 U560 ( .A1(n142), .A2(n592), .ZN(n491) );
  BUF_X1 U561 ( .A(n137), .Z(n38) );
  INV_X1 U562 ( .A(B[0]), .ZN(n625) );
  INV_X1 U563 ( .A(B[4]), .ZN(n44) );
  NOR2_X2 U564 ( .A1(n635), .A2(LOGIC_ARITH), .ZN(n142) );
  INV_X1 U565 ( .A(n591), .ZN(n635) );
  NOR3_X1 U566 ( .A1(B[9]), .A2(B[8]), .A3(B[10]), .ZN(n489) );
  NOR3_X1 U567 ( .A1(B[7]), .A2(B[6]), .A3(B[5]), .ZN(n579) );
  NOR3_X1 U568 ( .A1(B[28]), .A2(B[27]), .A3(B[26]), .ZN(n592) );
  OAI222_X1 U569 ( .A1(n468), .A2(n269), .B1(n469), .B2(n37), .C1(n92), .C2(
        n34), .ZN(RES[17]) );
  AOI221_X1 U570 ( .B1(n165), .B2(n474), .C1(n199), .C2(n419), .A(n475), .ZN(
        n468) );
  AOI221_X1 U571 ( .B1(n276), .B2(n470), .C1(n628), .C2(n434), .A(n279), .ZN(
        n469) );
  OAI222_X1 U572 ( .A1(n132), .A2(n636), .B1(n362), .B2(n641), .C1(n363), .C2(
        n645), .ZN(n475) );
  OAI222_X1 U573 ( .A1(n458), .A2(n269), .B1(n459), .B2(n38), .C1(n96), .C2(
        n34), .ZN(RES[18]) );
  AOI221_X1 U574 ( .B1(n165), .B2(n465), .C1(n199), .C2(n406), .A(n466), .ZN(
        n458) );
  AOI221_X1 U575 ( .B1(n276), .B2(n460), .C1(n628), .C2(n297), .A(n279), .ZN(
        n459) );
  OAI222_X1 U576 ( .A1(n614), .A2(n636), .B1(n293), .B2(n641), .C1(n405), .C2(
        n645), .ZN(n466) );
  OAI222_X1 U577 ( .A1(n446), .A2(n269), .B1(n447), .B2(n37), .C1(n100), .C2(
        n34), .ZN(RES[19]) );
  AOI221_X1 U578 ( .B1(n165), .B2(n455), .C1(n199), .C2(n388), .A(n456), .ZN(
        n446) );
  AOI221_X1 U579 ( .B1(n276), .B2(n448), .C1(n628), .C2(n246), .A(n279), .ZN(
        n447) );
  OAI222_X1 U580 ( .A1(n616), .A2(n636), .B1(n46), .B2(n641), .C1(n387), .C2(
        n645), .ZN(n456) );
  OAI222_X1 U581 ( .A1(n422), .A2(n269), .B1(n423), .B2(n37), .C1(n105), .C2(
        n34), .ZN(RES[20]) );
  AOI221_X1 U582 ( .B1(n165), .B2(n373), .C1(n199), .C2(n372), .A(n427), .ZN(
        n422) );
  AOI221_X1 U583 ( .B1(n276), .B2(n424), .C1(n628), .C2(n107), .A(n279), .ZN(
        n423) );
  OAI221_X1 U584 ( .B1(n376), .B2(n636), .C1(n63), .C2(n645), .A(n428), .ZN(
        n427) );
  OAI222_X1 U585 ( .A1(n409), .A2(n269), .B1(n410), .B2(n37), .C1(n108), .C2(
        n34), .ZN(RES[21]) );
  AOI221_X1 U586 ( .B1(n276), .B2(n411), .C1(n628), .C2(n223), .A(n279), .ZN(
        n410) );
  AOI221_X1 U587 ( .B1(n199), .B2(n361), .C1(B[4]), .C2(n56), .A(n418), .ZN(
        n409) );
  OAI21_X1 U588 ( .B1(n414), .B2(n281), .A(n282), .ZN(n411) );
  OAI222_X1 U589 ( .A1(n392), .A2(n269), .B1(n393), .B2(n37), .C1(n111), .C2(
        n34), .ZN(RES[22]) );
  AOI221_X1 U590 ( .B1(n276), .B2(n394), .C1(n628), .C2(n211), .A(n279), .ZN(
        n393) );
  AOI221_X1 U591 ( .B1(n199), .B2(n350), .C1(B[4]), .C2(n50), .A(n404), .ZN(
        n392) );
  OAI21_X1 U592 ( .B1(n397), .B2(n281), .A(n282), .ZN(n394) );
  OAI222_X1 U593 ( .A1(n378), .A2(n269), .B1(n379), .B2(n37), .C1(n114), .C2(
        n34), .ZN(RES[23]) );
  AOI221_X1 U594 ( .B1(n276), .B2(n380), .C1(n628), .C2(n115), .A(n279), .ZN(
        n379) );
  AOI221_X1 U595 ( .B1(n199), .B2(n339), .C1(B[4]), .C2(n48), .A(n386), .ZN(
        n378) );
  OAI21_X1 U596 ( .B1(n384), .B2(n281), .A(n282), .ZN(n380) );
  OAI222_X1 U597 ( .A1(n365), .A2(n269), .B1(n366), .B2(n37), .C1(n117), .C2(
        n34), .ZN(RES[24]) );
  AOI221_X1 U598 ( .B1(n276), .B2(n367), .C1(n628), .C2(n119), .A(n279), .ZN(
        n366) );
  AOI221_X1 U599 ( .B1(n199), .B2(n324), .C1(n39), .C2(n172), .A(n371), .ZN(
        n365) );
  OAI21_X1 U600 ( .B1(n368), .B2(n281), .A(n282), .ZN(n367) );
  OAI222_X1 U601 ( .A1(n352), .A2(n269), .B1(n353), .B2(n37), .C1(n120), .C2(
        n34), .ZN(RES[25]) );
  AOI221_X1 U602 ( .B1(n276), .B2(n354), .C1(n628), .C2(n122), .A(n279), .ZN(
        n353) );
  AOI221_X1 U603 ( .B1(n199), .B2(n313), .C1(n39), .C2(n139), .A(n360), .ZN(
        n352) );
  INV_X1 U604 ( .A(n163), .ZN(n122) );
  OAI222_X1 U605 ( .A1(n477), .A2(n269), .B1(n478), .B2(n38), .C1(n88), .C2(
        n35), .ZN(RES[16]) );
  AOI221_X1 U606 ( .B1(n165), .B2(n429), .C1(n199), .C2(n373), .A(n492), .ZN(
        n477) );
  AOI221_X1 U607 ( .B1(n276), .B2(n479), .C1(n628), .C2(n480), .A(n279), .ZN(
        n478) );
  OAI222_X1 U608 ( .A1(n374), .A2(n636), .B1(n375), .B2(n641), .C1(n376), .C2(
        n645), .ZN(n492) );
  OAI222_X1 U609 ( .A1(n341), .A2(n269), .B1(n342), .B2(n37), .C1(n123), .C2(
        n34), .ZN(RES[26]) );
  AOI221_X1 U610 ( .B1(n276), .B2(n343), .C1(n628), .C2(n125), .A(n279), .ZN(
        n342) );
  AOI221_X1 U611 ( .B1(n199), .B2(n289), .C1(n39), .C2(n348), .A(n349), .ZN(
        n341) );
  INV_X1 U612 ( .A(n344), .ZN(n125) );
  OAI222_X1 U613 ( .A1(n328), .A2(n269), .B1(n329), .B2(n37), .C1(n126), .C2(
        n34), .ZN(RES[27]) );
  AOI211_X1 U614 ( .C1(n276), .C2(n330), .A(n279), .B(n331), .ZN(n329) );
  AOI221_X1 U615 ( .B1(n199), .B2(n270), .C1(n39), .C2(n337), .A(n338), .ZN(
        n328) );
  OAI21_X1 U616 ( .B1(n334), .B2(n281), .A(n282), .ZN(n330) );
  OAI222_X1 U617 ( .A1(n317), .A2(n269), .B1(n318), .B2(n37), .C1(n128), .C2(
        n34), .ZN(RES[28]) );
  AOI221_X1 U618 ( .B1(n165), .B2(n324), .C1(n39), .C2(n54), .A(n325), .ZN(
        n317) );
  AOI221_X1 U619 ( .B1(n276), .B2(n319), .C1(n278), .C2(n320), .A(n279), .ZN(
        n318) );
  INV_X1 U620 ( .A(n327), .ZN(n54) );
  OAI222_X1 U621 ( .A1(n307), .A2(n269), .B1(n308), .B2(n37), .C1(n131), .C2(
        n33), .ZN(RES[29]) );
  AOI221_X1 U622 ( .B1(n165), .B2(n313), .C1(n39), .C2(n314), .A(n315), .ZN(
        n307) );
  AOI221_X1 U623 ( .B1(n276), .B2(n309), .C1(n278), .C2(n129), .A(n279), .ZN(
        n308) );
  OAI222_X1 U624 ( .A1(n82), .A2(n636), .B1(n316), .B2(n642), .C1(n95), .C2(
        n645), .ZN(n315) );
  OAI222_X1 U625 ( .A1(n274), .A2(n269), .B1(n275), .B2(n38), .C1(n266), .C2(
        n33), .ZN(RES[30]) );
  AOI221_X1 U626 ( .B1(n165), .B2(n289), .C1(n39), .C2(n290), .A(n291), .ZN(
        n274) );
  AOI221_X1 U627 ( .B1(n276), .B2(n277), .C1(n278), .C2(n134), .A(n279), .ZN(
        n275) );
  OAI222_X1 U628 ( .A1(n85), .A2(n636), .B1(n292), .B2(n642), .C1(n99), .C2(
        n645), .ZN(n291) );
  OAI221_X1 U629 ( .B1(n293), .B2(n240), .C1(n133), .C2(n33), .A(n294), .ZN(
        RES[2]) );
  AOI221_X1 U630 ( .B1(n242), .B2(n295), .C1(n627), .C2(n69), .A(n244), .ZN(
        n294) );
  INV_X1 U631 ( .A(n296), .ZN(n69) );
  OAI21_X1 U632 ( .B1(n299), .B2(n249), .A(n250), .ZN(n295) );
  OAI221_X1 U633 ( .B1(n362), .B2(n240), .C1(n103), .C2(n33), .A(n431), .ZN(
        RES[1]) );
  AOI221_X1 U634 ( .B1(n242), .B2(n432), .C1(n627), .C2(n72), .A(n244), .ZN(
        n431) );
  INV_X1 U635 ( .A(n433), .ZN(n72) );
  OAI21_X1 U636 ( .B1(n437), .B2(n249), .A(n250), .ZN(n432) );
  OAI221_X1 U640 ( .B1(n46), .B2(n240), .C1(n615), .C2(n33), .A(n241), .ZN(
        RES[3]) );
  AOI221_X1 U643 ( .B1(n242), .B2(n243), .C1(n627), .C2(n60), .A(n244), .ZN(
        n241) );
  INV_X1 U644 ( .A(n245), .ZN(n60) );
  OAI21_X1 U645 ( .B1(n248), .B2(n249), .A(n250), .ZN(n243) );
  NOR2_X1 U646 ( .A1(B[29]), .A2(B[30]), .ZN(n591) );
  AND2_X1 U647 ( .A1(LOGIC_ARITH), .A2(n445), .ZN(n140) );
  NOR2_X1 U648 ( .A1(n613), .A2(LOGIC_ARITH), .ZN(n590) );
  OAI221_X1 U649 ( .B1(n587), .B2(n436), .C1(n49), .C2(n33), .A(n588), .ZN(
        RES[0]) );
  NOR2_X1 U650 ( .A1(n269), .A2(n39), .ZN(n228) );
  AOI21_X1 U651 ( .B1(n242), .B2(n589), .A(n244), .ZN(n588) );
  OAI21_X1 U652 ( .B1(n593), .B2(n249), .A(n250), .ZN(n589) );
  AOI21_X1 U653 ( .B1(n251), .B2(n595), .A(n253), .ZN(n593) );
  OAI21_X1 U654 ( .B1(n587), .B2(n255), .A(n256), .ZN(n595) );
  AND2_X1 U655 ( .A1(n491), .A2(n649), .ZN(n242) );
  NAND2_X1 U656 ( .A1(n35), .A2(n649), .ZN(n137) );
  NAND2_X1 U657 ( .A1(n140), .A2(n649), .ZN(n436) );
  NOR2_X1 U658 ( .A1(n481), .A2(LEFT_RIGHT), .ZN(n244) );
  INV_X1 U659 ( .A(LEFT_RIGHT), .ZN(n649) );
  OAI222_X1 U660 ( .A1(n268), .A2(n269), .B1(LEFT_RIGHT), .B2(n612), .C1(n613), 
        .C2(n34), .ZN(RES[31]) );
  AOI221_X1 U661 ( .B1(n165), .B2(n270), .C1(n39), .C2(n271), .A(n272), .ZN(
        n268) );
  OAI222_X1 U662 ( .A1(n87), .A2(n636), .B1(n273), .B2(n642), .C1(n104), .C2(
        n645), .ZN(n272) );
  NOR4_X4 U663 ( .A1(B[16]), .A2(B[17]), .A3(B[15]), .A4(n598), .ZN(n148) );
  INV_X1 U664 ( .A(n8), .ZN(n6) );
  INV_X1 U665 ( .A(n8), .ZN(n7) );
  INV_X1 U666 ( .A(n1), .ZN(n9) );
  INV_X1 U667 ( .A(n1), .ZN(n10) );
  INV_X1 U668 ( .A(n1), .ZN(n11) );
  CLKBUF_X1 U669 ( .A(n264), .Z(n12) );
  CLKBUF_X1 U670 ( .A(n264), .Z(n13) );
  INV_X1 U671 ( .A(n19), .ZN(n17) );
  INV_X1 U672 ( .A(n12), .ZN(n18) );
  INV_X1 U673 ( .A(n12), .ZN(n19) );
  INV_X1 U674 ( .A(n264), .ZN(n20) );
  INV_X1 U675 ( .A(n13), .ZN(n21) );
  INV_X1 U676 ( .A(n13), .ZN(n22) );
  CLKBUF_X1 U677 ( .A(n263), .Z(n23) );
  CLKBUF_X1 U678 ( .A(n263), .Z(n24) );
  CLKBUF_X1 U679 ( .A(n263), .Z(n25) );
  INV_X1 U680 ( .A(n23), .ZN(n30) );
  INV_X1 U681 ( .A(n24), .ZN(n31) );
  INV_X1 U682 ( .A(n25), .ZN(n32) );
endmodule


module PG_net_0 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_30 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_29 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_28 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_27 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_26 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_25 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_24 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_23 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_22 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_21 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_20 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_19 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_18 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_17 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_16 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_15 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_14 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_13 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_12 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_11 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_10 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_9 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_8 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_7 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_6 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_5 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_4 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_3 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_2 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_1 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module Gblock_0 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n2) );
endmodule


module Gblock_8 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_7 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_6 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_5 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_4 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_3 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_2 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_1 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module PGblock_0 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n2) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_26 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_25 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_24 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_23 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_22 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_21 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_20 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_19 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_18 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_17 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_16 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_15 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_14 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_13 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_12 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_11 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_10 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_9 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_8 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_7 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_6 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_5 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_4 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_3 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_2 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_1 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module carry_generator_NBIT32_NBIT_PER_BLOCK4 ( A, B, Cin, Co );
  input [32:1] A;
  input [32:1] B;
  output [7:0] Co;
  input Cin;
  wire   \G[16][16] , \G[16][15] , \G[16][13] , \G[16][9] , \G[15][15] ,
         \G[14][14] , \G[14][13] , \G[13][13] , \G[12][12] , \G[12][11] ,
         \G[12][9] , \G[11][11] , \G[10][10] , \G[10][9] , \G[9][9] ,
         \G[8][8] , \G[8][7] , \G[8][5] , \G[7][7] , \G[6][6] , \G[6][5] ,
         \G[5][5] , \G[4][4] , \G[4][3] , \G[3][3] , \G[2][2] , \G[2][1] ,
         \G[1][1] , \P[16][16] , \P[16][15] , \P[16][13] , \P[16][9] ,
         \P[15][15] , \P[14][14] , \P[14][13] , \P[13][13] , \P[12][12] ,
         \P[12][11] , \P[12][9] , \P[11][11] , \P[10][10] , \P[10][9] ,
         \P[9][9] , \P[8][8] , \P[8][7] , \P[8][5] , \P[7][7] , \P[6][6] ,
         \P[6][5] , \P[5][5] , \P[4][4] , \P[4][3] , \P[3][3] , \P[2][2] ,
         \G[32][32] , \G[32][31] , \G[32][29] , \G[32][25] , \G[32][17] ,
         \G[31][31] , \G[30][30] , \G[30][29] , \G[29][29] , \G[28][28] ,
         \G[28][27] , \G[28][25] , \G[28][17] , \G[27][27] , \G[26][26] ,
         \G[26][25] , \G[25][25] , \G[24][24] , \G[24][23] , \G[24][21] ,
         \G[24][17] , \G[23][23] , \G[22][22] , \G[22][21] , \G[21][21] ,
         \G[20][20] , \G[20][19] , \G[20][17] , \G[19][19] , \G[18][18] ,
         \G[18][17] , \G[17][17] , \P[32][32] , \P[32][31] , \P[32][29] ,
         \P[32][25] , \P[32][17] , \P[31][31] , \P[30][30] , \P[30][29] ,
         \P[29][29] , \P[28][28] , \P[28][27] , \P[28][25] , \P[28][17] ,
         \P[27][27] , \P[26][26] , \P[26][25] , \P[25][25] , \P[24][24] ,
         \P[24][23] , \P[24][21] , \P[24][17] , \P[23][23] , \P[22][22] ,
         \P[22][21] , \P[21][21] , \P[20][20] , \P[20][19] , \P[20][17] ,
         \P[19][19] , \P[18][18] , \P[18][17] , \P[17][17] , n3, n1, n2;

  PG_net_0 PGnetblock_2 ( .a(A[2]), .b(B[2]), .p(\P[2][2] ), .g(\G[2][2] ) );
  PG_net_30 PGnetblock_3 ( .a(A[3]), .b(B[3]), .p(\P[3][3] ), .g(\G[3][3] ) );
  PG_net_29 PGnetblock_4 ( .a(A[4]), .b(B[4]), .p(\P[4][4] ), .g(\G[4][4] ) );
  PG_net_28 PGnetblock_5 ( .a(A[5]), .b(B[5]), .p(\P[5][5] ), .g(\G[5][5] ) );
  PG_net_27 PGnetblock_6 ( .a(A[6]), .b(B[6]), .p(\P[6][6] ), .g(\G[6][6] ) );
  PG_net_26 PGnetblock_7 ( .a(A[7]), .b(B[7]), .p(\P[7][7] ), .g(\G[7][7] ) );
  PG_net_25 PGnetblock_8 ( .a(A[8]), .b(B[8]), .p(\P[8][8] ), .g(\G[8][8] ) );
  PG_net_24 PGnetblock_9 ( .a(A[9]), .b(B[9]), .p(\P[9][9] ), .g(\G[9][9] ) );
  PG_net_23 PGnetblock_10 ( .a(A[10]), .b(B[10]), .p(\P[10][10] ), .g(
        \G[10][10] ) );
  PG_net_22 PGnetblock_11 ( .a(A[11]), .b(B[11]), .p(\P[11][11] ), .g(
        \G[11][11] ) );
  PG_net_21 PGnetblock_12 ( .a(A[12]), .b(B[12]), .p(\P[12][12] ), .g(
        \G[12][12] ) );
  PG_net_20 PGnetblock_13 ( .a(A[13]), .b(B[13]), .p(\P[13][13] ), .g(
        \G[13][13] ) );
  PG_net_19 PGnetblock_14 ( .a(A[14]), .b(B[14]), .p(\P[14][14] ), .g(
        \G[14][14] ) );
  PG_net_18 PGnetblock_15 ( .a(A[15]), .b(B[15]), .p(\P[15][15] ), .g(
        \G[15][15] ) );
  PG_net_17 PGnetblock_16 ( .a(A[16]), .b(B[16]), .p(\P[16][16] ), .g(
        \G[16][16] ) );
  PG_net_16 PGnetblock_17 ( .a(A[17]), .b(B[17]), .p(\P[17][17] ), .g(
        \G[17][17] ) );
  PG_net_15 PGnetblock_18 ( .a(A[18]), .b(B[18]), .p(\P[18][18] ), .g(
        \G[18][18] ) );
  PG_net_14 PGnetblock_19 ( .a(A[19]), .b(B[19]), .p(\P[19][19] ), .g(
        \G[19][19] ) );
  PG_net_13 PGnetblock_20 ( .a(A[20]), .b(B[20]), .p(\P[20][20] ), .g(
        \G[20][20] ) );
  PG_net_12 PGnetblock_21 ( .a(A[21]), .b(B[21]), .p(\P[21][21] ), .g(
        \G[21][21] ) );
  PG_net_11 PGnetblock_22 ( .a(A[22]), .b(B[22]), .p(\P[22][22] ), .g(
        \G[22][22] ) );
  PG_net_10 PGnetblock_23 ( .a(A[23]), .b(B[23]), .p(\P[23][23] ), .g(
        \G[23][23] ) );
  PG_net_9 PGnetblock_24 ( .a(A[24]), .b(B[24]), .p(\P[24][24] ), .g(
        \G[24][24] ) );
  PG_net_8 PGnetblock_25 ( .a(A[25]), .b(B[25]), .p(\P[25][25] ), .g(
        \G[25][25] ) );
  PG_net_7 PGnetblock_26 ( .a(A[26]), .b(B[26]), .p(\P[26][26] ), .g(
        \G[26][26] ) );
  PG_net_6 PGnetblock_27 ( .a(A[27]), .b(B[27]), .p(\P[27][27] ), .g(
        \G[27][27] ) );
  PG_net_5 PGnetblock_28 ( .a(A[28]), .b(B[28]), .p(\P[28][28] ), .g(
        \G[28][28] ) );
  PG_net_4 PGnetblock_29 ( .a(A[29]), .b(B[29]), .p(\P[29][29] ), .g(
        \G[29][29] ) );
  PG_net_3 PGnetblock_30 ( .a(A[30]), .b(B[30]), .p(\P[30][30] ), .g(
        \G[30][30] ) );
  PG_net_2 PGnetblock_31 ( .a(A[31]), .b(B[31]), .p(\P[31][31] ), .g(
        \G[31][31] ) );
  PG_net_1 PGnetblock_32 ( .a(A[32]), .b(B[32]), .p(\P[32][32] ), .g(
        \G[32][32] ) );
  Gblock_0 GB_low_1_2 ( .Pik(\P[2][2] ), .Gik(\G[2][2] ), .Gk_1j(\G[1][1] ), 
        .Gij(\G[2][1] ) );
  Gblock_8 GB_low_2_4 ( .Pik(\P[4][3] ), .Gik(\G[4][3] ), .Gk_1j(\G[2][1] ), 
        .Gij(Co[0]) );
  Gblock_7 GB_low_3_8 ( .Pik(\P[8][5] ), .Gik(\G[8][5] ), .Gk_1j(Co[0]), .Gij(
        Co[1]) );
  Gblock_6 GB_high_4_16_0 ( .Pik(\P[16][9] ), .Gik(\G[16][9] ), .Gk_1j(Co[1]), 
        .Gij(Co[3]) );
  Gblock_5 GB_high_4_16_1 ( .Pik(\P[12][9] ), .Gik(\G[12][9] ), .Gk_1j(Co[1]), 
        .Gij(Co[2]) );
  Gblock_4 GB_high_5_32_0 ( .Pik(\P[32][17] ), .Gik(\G[32][17] ), .Gk_1j(Co[3]), .Gij(Co[7]) );
  Gblock_3 GB_high_5_32_1 ( .Pik(\P[28][17] ), .Gik(\G[28][17] ), .Gk_1j(Co[3]), .Gij(Co[6]) );
  Gblock_2 GB_high_5_32_2 ( .Pik(\P[24][17] ), .Gik(\G[24][17] ), .Gk_1j(Co[3]), .Gij(Co[5]) );
  Gblock_1 GB_high_5_32_3 ( .Pik(\P[20][17] ), .Gik(\G[20][17] ), .Gk_1j(Co[3]), .Gij(Co[4]) );
  PGblock_0 PGB_low_1_4 ( .Pik(\P[4][4] ), .Gik(\G[4][4] ), .Pk_1j(\P[3][3] ), 
        .Gk_1j(\G[3][3] ), .Pij(\P[4][3] ), .Gij(\G[4][3] ) );
  PGblock_26 PGB_low_1_6 ( .Pik(\P[6][6] ), .Gik(\G[6][6] ), .Pk_1j(\P[5][5] ), 
        .Gk_1j(\G[5][5] ), .Pij(\P[6][5] ), .Gij(\G[6][5] ) );
  PGblock_25 PGB_low_1_8 ( .Pik(\P[8][8] ), .Gik(\G[8][8] ), .Pk_1j(\P[7][7] ), 
        .Gk_1j(\G[7][7] ), .Pij(\P[8][7] ), .Gij(\G[8][7] ) );
  PGblock_24 PGB_low_1_10 ( .Pik(\P[10][10] ), .Gik(\G[10][10] ), .Pk_1j(
        \P[9][9] ), .Gk_1j(\G[9][9] ), .Pij(\P[10][9] ), .Gij(\G[10][9] ) );
  PGblock_23 PGB_low_1_12 ( .Pik(\P[12][12] ), .Gik(\G[12][12] ), .Pk_1j(
        \P[11][11] ), .Gk_1j(\G[11][11] ), .Pij(\P[12][11] ), .Gij(\G[12][11] ) );
  PGblock_22 PGB_low_1_14 ( .Pik(\P[14][14] ), .Gik(\G[14][14] ), .Pk_1j(
        \P[13][13] ), .Gk_1j(\G[13][13] ), .Pij(\P[14][13] ), .Gij(\G[14][13] ) );
  PGblock_21 PGB_low_1_16 ( .Pik(\P[16][16] ), .Gik(\G[16][16] ), .Pk_1j(
        \P[15][15] ), .Gk_1j(\G[15][15] ), .Pij(\P[16][15] ), .Gij(\G[16][15] ) );
  PGblock_20 PGB_low_1_18 ( .Pik(\P[18][18] ), .Gik(\G[18][18] ), .Pk_1j(
        \P[17][17] ), .Gk_1j(\G[17][17] ), .Pij(\P[18][17] ), .Gij(\G[18][17] ) );
  PGblock_19 PGB_low_1_20 ( .Pik(\P[20][20] ), .Gik(\G[20][20] ), .Pk_1j(
        \P[19][19] ), .Gk_1j(\G[19][19] ), .Pij(\P[20][19] ), .Gij(\G[20][19] ) );
  PGblock_18 PGB_low_1_22 ( .Pik(\P[22][22] ), .Gik(\G[22][22] ), .Pk_1j(
        \P[21][21] ), .Gk_1j(\G[21][21] ), .Pij(\P[22][21] ), .Gij(\G[22][21] ) );
  PGblock_17 PGB_low_1_24 ( .Pik(\P[24][24] ), .Gik(\G[24][24] ), .Pk_1j(
        \P[23][23] ), .Gk_1j(\G[23][23] ), .Pij(\P[24][23] ), .Gij(\G[24][23] ) );
  PGblock_16 PGB_low_1_26 ( .Pik(\P[26][26] ), .Gik(\G[26][26] ), .Pk_1j(
        \P[25][25] ), .Gk_1j(\G[25][25] ), .Pij(\P[26][25] ), .Gij(\G[26][25] ) );
  PGblock_15 PGB_low_1_28 ( .Pik(\P[28][28] ), .Gik(\G[28][28] ), .Pk_1j(
        \P[27][27] ), .Gk_1j(\G[27][27] ), .Pij(\P[28][27] ), .Gij(\G[28][27] ) );
  PGblock_14 PGB_low_1_30 ( .Pik(\P[30][30] ), .Gik(\G[30][30] ), .Pk_1j(
        \P[29][29] ), .Gk_1j(\G[29][29] ), .Pij(\P[30][29] ), .Gij(\G[30][29] ) );
  PGblock_13 PGB_low_1_32 ( .Pik(\P[32][32] ), .Gik(\G[32][32] ), .Pk_1j(
        \P[31][31] ), .Gk_1j(\G[31][31] ), .Pij(\P[32][31] ), .Gij(\G[32][31] ) );
  PGblock_12 PGB_low_2_8 ( .Pik(\P[8][7] ), .Gik(\G[8][7] ), .Pk_1j(\P[6][5] ), 
        .Gk_1j(\G[6][5] ), .Pij(\P[8][5] ), .Gij(\G[8][5] ) );
  PGblock_11 PGB_low_2_12 ( .Pik(\P[12][11] ), .Gik(\G[12][11] ), .Pk_1j(
        \P[10][9] ), .Gk_1j(\G[10][9] ), .Pij(\P[12][9] ), .Gij(\G[12][9] ) );
  PGblock_10 PGB_low_2_16 ( .Pik(\P[16][15] ), .Gik(\G[16][15] ), .Pk_1j(
        \P[14][13] ), .Gk_1j(\G[14][13] ), .Pij(\P[16][13] ), .Gij(\G[16][13] ) );
  PGblock_9 PGB_low_2_20 ( .Pik(\P[20][19] ), .Gik(\G[20][19] ), .Pk_1j(
        \P[18][17] ), .Gk_1j(\G[18][17] ), .Pij(\P[20][17] ), .Gij(\G[20][17] ) );
  PGblock_8 PGB_low_2_24 ( .Pik(\P[24][23] ), .Gik(\G[24][23] ), .Pk_1j(
        \P[22][21] ), .Gk_1j(\G[22][21] ), .Pij(\P[24][21] ), .Gij(\G[24][21] ) );
  PGblock_7 PGB_low_2_28 ( .Pik(\P[28][27] ), .Gik(\G[28][27] ), .Pk_1j(
        \P[26][25] ), .Gk_1j(\G[26][25] ), .Pij(\P[28][25] ), .Gij(\G[28][25] ) );
  PGblock_6 PGB_low_2_32 ( .Pik(\P[32][31] ), .Gik(\G[32][31] ), .Pk_1j(
        \P[30][29] ), .Gk_1j(\G[30][29] ), .Pij(\P[32][29] ), .Gij(\G[32][29] ) );
  PGblock_5 PGB_low_3_16 ( .Pik(\P[16][13] ), .Gik(\G[16][13] ), .Pk_1j(
        \P[12][9] ), .Gk_1j(\G[12][9] ), .Pij(\P[16][9] ), .Gij(\G[16][9] ) );
  PGblock_4 PGB_low_3_24 ( .Pik(\P[24][21] ), .Gik(\G[24][21] ), .Pk_1j(
        \P[20][17] ), .Gk_1j(\G[20][17] ), .Pij(\P[24][17] ), .Gij(\G[24][17] ) );
  PGblock_3 PGB_low_3_32 ( .Pik(\P[32][29] ), .Gik(\G[32][29] ), .Pk_1j(
        \P[28][25] ), .Gk_1j(\G[28][25] ), .Pij(\P[32][25] ), .Gij(\G[32][25] ) );
  PGblock_2 PGB_high_4_32_0 ( .Pik(\P[32][25] ), .Gik(\G[32][25] ), .Pk_1j(
        \P[24][17] ), .Gk_1j(\G[24][17] ), .Pij(\P[32][17] ), .Gij(\G[32][17] ) );
  PGblock_1 PGB_high_4_32_1 ( .Pik(\P[28][25] ), .Gik(\G[28][25] ), .Pk_1j(
        \P[24][17] ), .Gk_1j(\G[24][17] ), .Pij(\P[28][17] ), .Gij(\G[28][17] ) );
  INV_X1 U1 ( .A(A[1]), .ZN(n1) );
  OAI21_X1 U2 ( .B1(n1), .B2(n2), .A(n3), .ZN(\G[1][1] ) );
  INV_X1 U3 ( .A(B[1]), .ZN(n2) );
  OAI21_X1 U4 ( .B1(A[1]), .B2(B[1]), .A(Cin), .ZN(n3) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_0 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n6, n7, n8, n9, n5;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_0 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_15 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n6), .ZN(S[3]) );
  AOI22_X1 U5 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n6) );
  INV_X1 U6 ( .A(n8), .ZN(S[1]) );
  AOI22_X1 U7 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n8) );
  INV_X1 U8 ( .A(n7), .ZN(S[2]) );
  AOI22_X1 U9 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n7) );
  INV_X1 U10 ( .A(n9), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n9) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_7 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_14 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_13 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U9 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_6 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_12 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_11 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U9 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_5 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_10 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_9 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U9 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_4 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_8 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_7 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U9 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_3 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_6 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_5 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U9 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_2 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_4 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_3 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U9 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_1 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_2 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_1 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U5 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U6 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U7 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U8 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U9 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_select_basic_N4_0 CSBI_1 ( .A(A[3:0]), .B(B[3:0]), .C_i(Ci[0]), .S(
        S[3:0]) );
  carry_select_basic_N4_7 CSBI_2 ( .A(A[7:4]), .B(B[7:4]), .C_i(Ci[1]), .S(
        S[7:4]) );
  carry_select_basic_N4_6 CSBI_3 ( .A(A[11:8]), .B(B[11:8]), .C_i(Ci[2]), .S(
        S[11:8]) );
  carry_select_basic_N4_5 CSBI_4 ( .A(A[15:12]), .B(B[15:12]), .C_i(Ci[3]), 
        .S(S[15:12]) );
  carry_select_basic_N4_4 CSBI_5 ( .A(A[19:16]), .B(B[19:16]), .C_i(Ci[4]), 
        .S(S[19:16]) );
  carry_select_basic_N4_3 CSBI_6 ( .A(A[23:20]), .B(B[23:20]), .C_i(Ci[5]), 
        .S(S[23:20]) );
  carry_select_basic_N4_2 CSBI_7 ( .A(A[27:24]), .B(B[27:24]), .C_i(Ci[6]), 
        .S(S[27:24]) );
  carry_select_basic_N4_1 CSBI_8 ( .A(A[31:28]), .B(B[31:28]), .C_i(Ci[7]), 
        .S(S[31:28]) );
endmodule


module P4Adder_NBIT32 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;

  wire   [7:1] Csum;

  carry_generator_NBIT32_NBIT_PER_BLOCK4 Carrygen0 ( .A(A), .B(B), .Cin(Cin), 
        .Co({Cout, Csum}) );
  SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 Sumgen0 ( .A(A), .B(B), .Ci({Csum, 
        Cin}), .S(S) );
endmodule


module booth_encoder_numBit16 ( B, SEL_out );
  input [15:0] B;
  output [23:0] SEL_out;
  wire   \B[15] , \B[14] , \B[13] , SEL_out_19, SEL_out_18, SEL_out_16,
         SEL_out_15, SEL_out_13, SEL_out_12, SEL_out_10, SEL_out_9, SEL_out_7,
         SEL_out_6, SEL_out_4, SEL_out_3, SEL_out_1;
  assign SEL_out[0] = 1'b0;
  assign SEL_out[23] = \B[15] ;
  assign \B[15]  = B[15];
  assign SEL_out[22] = \B[14] ;
  assign \B[14]  = B[14];
  assign SEL_out[20] = \B[13] ;
  assign SEL_out[21] = \B[13] ;
  assign \B[13]  = B[13];
  assign SEL_out[19] = SEL_out_19;
  assign SEL_out_19 = B[12];
  assign SEL_out[17] = SEL_out_18;
  assign SEL_out[18] = SEL_out_18;
  assign SEL_out_18 = B[11];
  assign SEL_out[16] = SEL_out_16;
  assign SEL_out_16 = B[10];
  assign SEL_out[14] = SEL_out_15;
  assign SEL_out[15] = SEL_out_15;
  assign SEL_out_15 = B[9];
  assign SEL_out[13] = SEL_out_13;
  assign SEL_out_13 = B[8];
  assign SEL_out[11] = SEL_out_12;
  assign SEL_out[12] = SEL_out_12;
  assign SEL_out_12 = B[7];
  assign SEL_out[10] = SEL_out_10;
  assign SEL_out_10 = B[6];
  assign SEL_out[8] = SEL_out_9;
  assign SEL_out[9] = SEL_out_9;
  assign SEL_out_9 = B[5];
  assign SEL_out[7] = SEL_out_7;
  assign SEL_out_7 = B[4];
  assign SEL_out[5] = SEL_out_6;
  assign SEL_out[6] = SEL_out_6;
  assign SEL_out_6 = B[3];
  assign SEL_out[4] = SEL_out_4;
  assign SEL_out_4 = B[2];
  assign SEL_out[2] = SEL_out_3;
  assign SEL_out[3] = SEL_out_3;
  assign SEL_out_3 = B[1];
  assign SEL_out[1] = SEL_out_1;
  assign SEL_out_1 = B[0];

endmodule


module mux5to1_numBit32_0 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  OAI33_X1 U109 ( .A1(n91), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n90), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n8) );
  BUF_X1 U2 ( .A(n10), .Z(n4) );
  BUF_X1 U3 ( .A(n10), .Z(n77) );
  BUF_X1 U4 ( .A(n10), .Z(n78) );
  INV_X1 U5 ( .A(SEL_in[1]), .ZN(n90) );
  AOI222_X1 U6 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n68) );
  AOI222_X1 U7 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n66) );
  AOI222_X1 U8 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n64) );
  AOI222_X1 U9 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n62) );
  AOI222_X1 U10 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n60) );
  AOI222_X1 U11 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n58) );
  AOI222_X1 U12 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n56) );
  AOI222_X1 U13 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n54) );
  AOI222_X1 U14 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), 
        .C2(n79), .ZN(n52) );
  AOI222_X1 U15 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), 
        .C2(n79), .ZN(n50) );
  AOI222_X1 U16 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), 
        .C2(n80), .ZN(n48) );
  AOI222_X1 U17 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), 
        .C2(n80), .ZN(n46) );
  AOI222_X1 U18 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n44) );
  AOI222_X1 U19 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n42) );
  AOI222_X1 U20 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n22) );
  AOI222_X1 U21 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n20) );
  AOI222_X1 U22 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n18) );
  AOI222_X1 U23 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), 
        .C2(n81), .ZN(n16) );
  AOI222_X1 U24 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), 
        .C2(n81), .ZN(n14) );
  AOI222_X1 U25 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), 
        .C2(n81), .ZN(n12) );
  AOI222_X1 U26 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n70) );
  AOI222_X1 U27 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n40) );
  AOI222_X1 U28 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n38) );
  AOI222_X1 U29 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n36) );
  AOI222_X1 U30 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n34) );
  AOI222_X1 U31 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n32) );
  AOI222_X1 U32 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n30) );
  AOI222_X1 U33 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n28) );
  AOI222_X1 U34 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n26) );
  AOI222_X1 U35 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n24) );
  BUF_X1 U36 ( .A(n9), .Z(n79) );
  BUF_X1 U37 ( .A(n9), .Z(n80) );
  BUF_X1 U38 ( .A(n7), .Z(n85) );
  BUF_X1 U39 ( .A(n7), .Z(n86) );
  BUF_X1 U40 ( .A(n89), .Z(n1) );
  BUF_X1 U41 ( .A(n89), .Z(n2) );
  NOR2_X1 U42 ( .A1(n88), .A2(n75), .ZN(n10) );
  INV_X1 U43 ( .A(n74), .ZN(n88) );
  BUF_X1 U44 ( .A(n89), .Z(n3) );
  BUF_X1 U45 ( .A(n9), .Z(n81) );
  BUF_X1 U46 ( .A(n7), .Z(n87) );
  NOR4_X1 U47 ( .A1(n76), .A2(n85), .A3(n79), .A4(n82), .ZN(n74) );
  NOR3_X1 U48 ( .A1(n90), .A2(SEL_in[2]), .A3(n91), .ZN(n7) );
  BUF_X1 U49 ( .A(n8), .Z(n82) );
  BUF_X1 U50 ( .A(n8), .Z(n83) );
  BUF_X1 U51 ( .A(n8), .Z(n84) );
  NOR2_X1 U52 ( .A1(n90), .A2(n91), .ZN(n75) );
  AND3_X1 U53 ( .A1(n91), .A2(n90), .A3(SEL_in[2]), .ZN(n9) );
  NAND2_X1 U54 ( .A1(n65), .A2(n66), .ZN(Z[3]) );
  INV_X1 U55 ( .A(n73), .ZN(n89) );
  AOI21_X1 U56 ( .B1(n74), .B2(n75), .A(n76), .ZN(n73) );
  AOI22_X1 U57 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n69) );
  AOI22_X1 U58 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n67) );
  AOI22_X1 U59 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n65) );
  AOI22_X1 U60 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n63) );
  AOI22_X1 U61 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n61) );
  AOI22_X1 U62 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n59) );
  AOI22_X1 U63 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n57) );
  AOI22_X1 U64 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n55) );
  AOI22_X1 U65 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n53) );
  AOI22_X1 U66 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n51) );
  AOI22_X1 U67 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n49) );
  AOI22_X1 U68 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n47) );
  AOI22_X1 U69 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n45) );
  AOI22_X1 U70 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n43) );
  NOR3_X1 U71 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n76) );
  AOI222_X1 U72 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n72) );
  AOI22_X1 U73 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n41) );
  AOI22_X1 U74 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n23) );
  AOI22_X1 U75 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n21) );
  AOI22_X1 U76 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n19) );
  AOI22_X1 U77 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n17) );
  AOI22_X1 U78 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n15) );
  AOI22_X1 U79 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n13) );
  AOI22_X1 U80 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n11) );
  AOI22_X1 U81 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n71) );
  AOI22_X1 U82 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n33) );
  AOI22_X1 U83 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n31) );
  AOI22_X1 U84 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n29) );
  AOI22_X1 U85 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n27) );
  AOI22_X1 U86 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n25) );
  NAND2_X1 U87 ( .A1(n63), .A2(n64), .ZN(Z[4]) );
  NAND2_X1 U88 ( .A1(n61), .A2(n62), .ZN(Z[5]) );
  NAND2_X1 U89 ( .A1(n59), .A2(n60), .ZN(Z[6]) );
  NAND2_X1 U90 ( .A1(n57), .A2(n58), .ZN(Z[7]) );
  NAND2_X1 U91 ( .A1(n55), .A2(n56), .ZN(Z[8]) );
  NAND2_X1 U92 ( .A1(n53), .A2(n54), .ZN(Z[9]) );
  NAND2_X1 U93 ( .A1(n51), .A2(n52), .ZN(Z[10]) );
  NAND2_X1 U94 ( .A1(n49), .A2(n50), .ZN(Z[11]) );
  NAND2_X1 U95 ( .A1(n47), .A2(n48), .ZN(Z[12]) );
  NAND2_X1 U96 ( .A1(n45), .A2(n46), .ZN(Z[13]) );
  NAND2_X1 U97 ( .A1(n43), .A2(n44), .ZN(Z[14]) );
  NAND2_X1 U98 ( .A1(n41), .A2(n42), .ZN(Z[15]) );
  NAND2_X1 U99 ( .A1(n39), .A2(n40), .ZN(Z[16]) );
  AOI22_X1 U100 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n39) );
  NAND2_X1 U101 ( .A1(n37), .A2(n38), .ZN(Z[17]) );
  AOI22_X1 U102 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n37) );
  NAND2_X1 U103 ( .A1(n35), .A2(n36), .ZN(Z[18]) );
  AOI22_X1 U104 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n35) );
  NAND2_X1 U105 ( .A1(n33), .A2(n34), .ZN(Z[19]) );
  NAND2_X1 U106 ( .A1(n31), .A2(n32), .ZN(Z[20]) );
  NAND2_X1 U107 ( .A1(n29), .A2(n30), .ZN(Z[21]) );
  NAND2_X1 U108 ( .A1(n27), .A2(n28), .ZN(Z[22]) );
  NAND2_X1 U110 ( .A1(n25), .A2(n26), .ZN(Z[23]) );
  NAND2_X1 U111 ( .A1(n23), .A2(n24), .ZN(Z[24]) );
  NAND2_X1 U112 ( .A1(n21), .A2(n22), .ZN(Z[25]) );
  NAND2_X1 U113 ( .A1(n19), .A2(n20), .ZN(Z[26]) );
  NAND2_X1 U114 ( .A1(n17), .A2(n18), .ZN(Z[27]) );
  NAND2_X1 U115 ( .A1(n15), .A2(n16), .ZN(Z[28]) );
  NAND2_X1 U116 ( .A1(n13), .A2(n14), .ZN(Z[29]) );
  NAND2_X1 U117 ( .A1(n11), .A2(n12), .ZN(Z[30]) );
  NAND2_X1 U118 ( .A1(n67), .A2(n68), .ZN(Z[2]) );
  NAND2_X1 U119 ( .A1(n71), .A2(n72), .ZN(Z[0]) );
  NAND2_X1 U120 ( .A1(n69), .A2(n70), .ZN(Z[1]) );
  NAND2_X1 U121 ( .A1(n5), .A2(n6), .ZN(Z[31]) );
  AOI22_X1 U122 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n5) );
  AOI222_X1 U123 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), .C2(n81), .ZN(n6) );
  INV_X1 U124 ( .A(SEL_in[0]), .ZN(n91) );
endmodule


module mux5to1_numBit32_7 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  OAI33_X1 U109 ( .A1(n90), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n91), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n160) );
  BUF_X1 U2 ( .A(n158), .Z(n4) );
  BUF_X1 U3 ( .A(n158), .Z(n77) );
  BUF_X1 U4 ( .A(n158), .Z(n78) );
  AOI222_X1 U5 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n146) );
  AOI222_X1 U6 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n148) );
  AOI222_X1 U7 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n150) );
  AOI222_X1 U8 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), 
        .C2(n81), .ZN(n152) );
  AOI222_X1 U9 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), 
        .C2(n81), .ZN(n154) );
  AOI222_X1 U10 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), 
        .C2(n81), .ZN(n156) );
  AOI222_X1 U11 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n132) );
  AOI222_X1 U12 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n134) );
  AOI222_X1 U13 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n136) );
  AOI222_X1 U14 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n138) );
  AOI222_X1 U15 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n140) );
  AOI222_X1 U16 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n142) );
  AOI222_X1 U17 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n144) );
  BUF_X1 U18 ( .A(n89), .Z(n1) );
  BUF_X1 U19 ( .A(n89), .Z(n2) );
  NOR2_X1 U20 ( .A1(n88), .A2(n93), .ZN(n158) );
  INV_X1 U21 ( .A(n94), .ZN(n88) );
  BUF_X1 U22 ( .A(n89), .Z(n3) );
  NOR4_X1 U23 ( .A1(n92), .A2(n85), .A3(n79), .A4(n82), .ZN(n94) );
  BUF_X1 U24 ( .A(n160), .Z(n82) );
  BUF_X1 U25 ( .A(n160), .Z(n83) );
  BUF_X1 U26 ( .A(n159), .Z(n79) );
  BUF_X1 U27 ( .A(n159), .Z(n80) );
  BUF_X1 U28 ( .A(n161), .Z(n85) );
  BUF_X1 U29 ( .A(n161), .Z(n86) );
  BUF_X1 U30 ( .A(n160), .Z(n84) );
  NOR2_X1 U31 ( .A1(n91), .A2(n90), .ZN(n93) );
  BUF_X1 U32 ( .A(n159), .Z(n81) );
  BUF_X1 U33 ( .A(n161), .Z(n87) );
  INV_X1 U34 ( .A(n95), .ZN(n89) );
  AOI21_X1 U35 ( .B1(n94), .B2(n93), .A(n92), .ZN(n95) );
  AOI222_X1 U36 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n104) );
  AOI222_X1 U37 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n106) );
  AOI222_X1 U38 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n108) );
  AOI222_X1 U39 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n110) );
  AOI222_X1 U40 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n112) );
  AOI222_X1 U41 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n114) );
  AOI222_X1 U42 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), 
        .C2(n79), .ZN(n116) );
  AOI222_X1 U43 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), 
        .C2(n79), .ZN(n118) );
  AOI222_X1 U44 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), 
        .C2(n80), .ZN(n120) );
  AOI222_X1 U45 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), 
        .C2(n80), .ZN(n122) );
  AOI222_X1 U46 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n124) );
  AOI222_X1 U47 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n126) );
  AOI222_X1 U48 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n128) );
  AOI222_X1 U49 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n130) );
  NOR3_X1 U50 ( .A1(n91), .A2(SEL_in[2]), .A3(n90), .ZN(n161) );
  NOR3_X1 U51 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n92) );
  INV_X1 U52 ( .A(SEL_in[0]), .ZN(n90) );
  AND3_X1 U53 ( .A1(n90), .A2(n91), .A3(SEL_in[2]), .ZN(n159) );
  INV_X1 U54 ( .A(SEL_in[1]), .ZN(n91) );
  NAND2_X1 U55 ( .A1(n103), .A2(n102), .ZN(Z[3]) );
  AOI222_X1 U56 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n102) );
  AOI22_X1 U57 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n103) );
  AOI22_X1 U58 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n129) );
  AOI222_X1 U59 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n100) );
  AOI22_X1 U60 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n131) );
  AOI22_X1 U61 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n133) );
  NAND2_X1 U62 ( .A1(n105), .A2(n104), .ZN(Z[4]) );
  AOI22_X1 U63 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n105) );
  NAND2_X1 U64 ( .A1(n107), .A2(n106), .ZN(Z[5]) );
  AOI22_X1 U65 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n107) );
  NAND2_X1 U66 ( .A1(n109), .A2(n108), .ZN(Z[6]) );
  AOI22_X1 U67 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n109) );
  NAND2_X1 U68 ( .A1(n111), .A2(n110), .ZN(Z[7]) );
  AOI22_X1 U69 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n111) );
  NAND2_X1 U70 ( .A1(n113), .A2(n112), .ZN(Z[8]) );
  AOI22_X1 U71 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n113) );
  NAND2_X1 U72 ( .A1(n115), .A2(n114), .ZN(Z[9]) );
  AOI22_X1 U73 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n115) );
  NAND2_X1 U74 ( .A1(n117), .A2(n116), .ZN(Z[10]) );
  AOI22_X1 U75 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n117) );
  NAND2_X1 U76 ( .A1(n119), .A2(n118), .ZN(Z[11]) );
  AOI22_X1 U77 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n119) );
  NAND2_X1 U78 ( .A1(n121), .A2(n120), .ZN(Z[12]) );
  AOI22_X1 U79 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n121) );
  NAND2_X1 U80 ( .A1(n123), .A2(n122), .ZN(Z[13]) );
  AOI22_X1 U81 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n123) );
  NAND2_X1 U82 ( .A1(n125), .A2(n124), .ZN(Z[14]) );
  AOI22_X1 U83 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n125) );
  NAND2_X1 U84 ( .A1(n127), .A2(n126), .ZN(Z[15]) );
  AOI22_X1 U85 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n127) );
  NAND2_X1 U86 ( .A1(n129), .A2(n128), .ZN(Z[16]) );
  NAND2_X1 U87 ( .A1(n131), .A2(n130), .ZN(Z[17]) );
  NAND2_X1 U88 ( .A1(n133), .A2(n132), .ZN(Z[18]) );
  NAND2_X1 U89 ( .A1(n135), .A2(n134), .ZN(Z[19]) );
  AOI22_X1 U90 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n135) );
  NAND2_X1 U91 ( .A1(n137), .A2(n136), .ZN(Z[20]) );
  AOI22_X1 U92 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n137) );
  NAND2_X1 U93 ( .A1(n139), .A2(n138), .ZN(Z[21]) );
  AOI22_X1 U94 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n139) );
  NAND2_X1 U95 ( .A1(n141), .A2(n140), .ZN(Z[22]) );
  AOI22_X1 U96 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n141) );
  NAND2_X1 U97 ( .A1(n143), .A2(n142), .ZN(Z[23]) );
  AOI22_X1 U98 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n143) );
  NAND2_X1 U99 ( .A1(n145), .A2(n144), .ZN(Z[24]) );
  AOI22_X1 U100 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n145) );
  NAND2_X1 U101 ( .A1(n147), .A2(n146), .ZN(Z[25]) );
  AOI22_X1 U102 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n147) );
  NAND2_X1 U103 ( .A1(n149), .A2(n148), .ZN(Z[26]) );
  AOI22_X1 U104 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n149) );
  NAND2_X1 U105 ( .A1(n151), .A2(n150), .ZN(Z[27]) );
  AOI22_X1 U106 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n151) );
  NAND2_X1 U107 ( .A1(n153), .A2(n152), .ZN(Z[28]) );
  AOI22_X1 U108 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n153) );
  NAND2_X1 U110 ( .A1(n155), .A2(n154), .ZN(Z[29]) );
  AOI22_X1 U111 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n155) );
  NAND2_X1 U112 ( .A1(n157), .A2(n156), .ZN(Z[30]) );
  AOI22_X1 U113 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n157) );
  NAND2_X1 U114 ( .A1(n101), .A2(n100), .ZN(Z[2]) );
  AOI22_X1 U115 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n101) );
  NAND2_X1 U116 ( .A1(n97), .A2(n96), .ZN(Z[0]) );
  AOI22_X1 U117 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n97) );
  NAND2_X1 U118 ( .A1(n99), .A2(n98), .ZN(Z[1]) );
  AOI22_X1 U119 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n99) );
  NAND2_X1 U120 ( .A1(n163), .A2(n162), .ZN(Z[31]) );
  AOI22_X1 U121 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n163) );
  AOI222_X1 U122 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), .C2(n81), .ZN(n162) );
  AOI222_X1 U123 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n96) );
  AOI222_X1 U124 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n98) );
endmodule


module mux5to1_numBit32_6 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  OAI33_X1 U109 ( .A1(n90), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n91), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n160) );
  BUF_X1 U2 ( .A(n158), .Z(n4) );
  BUF_X1 U3 ( .A(n158), .Z(n77) );
  BUF_X1 U4 ( .A(n158), .Z(n78) );
  AOI222_X1 U5 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), 
        .C2(n81), .ZN(n162) );
  BUF_X1 U6 ( .A(n89), .Z(n1) );
  BUF_X1 U7 ( .A(n89), .Z(n2) );
  NOR2_X1 U8 ( .A1(n88), .A2(n93), .ZN(n158) );
  INV_X1 U9 ( .A(n94), .ZN(n88) );
  BUF_X1 U10 ( .A(n89), .Z(n3) );
  NOR4_X1 U11 ( .A1(n92), .A2(n85), .A3(n79), .A4(n82), .ZN(n94) );
  BUF_X1 U12 ( .A(n160), .Z(n82) );
  BUF_X1 U13 ( .A(n160), .Z(n83) );
  BUF_X1 U14 ( .A(n159), .Z(n79) );
  BUF_X1 U15 ( .A(n159), .Z(n80) );
  BUF_X1 U16 ( .A(n161), .Z(n85) );
  BUF_X1 U17 ( .A(n161), .Z(n86) );
  BUF_X1 U18 ( .A(n160), .Z(n84) );
  NOR2_X1 U19 ( .A1(n91), .A2(n90), .ZN(n93) );
  BUF_X1 U20 ( .A(n159), .Z(n81) );
  BUF_X1 U21 ( .A(n161), .Z(n87) );
  INV_X1 U22 ( .A(n95), .ZN(n89) );
  AOI21_X1 U23 ( .B1(n94), .B2(n93), .A(n92), .ZN(n95) );
  NOR3_X1 U24 ( .A1(n91), .A2(SEL_in[2]), .A3(n90), .ZN(n161) );
  NOR3_X1 U25 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n92) );
  INV_X1 U26 ( .A(SEL_in[0]), .ZN(n90) );
  AND3_X1 U27 ( .A1(n90), .A2(n91), .A3(SEL_in[2]), .ZN(n159) );
  INV_X1 U28 ( .A(SEL_in[1]), .ZN(n91) );
  NAND2_X1 U29 ( .A1(n107), .A2(n106), .ZN(Z[5]) );
  AOI222_X1 U30 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n106) );
  AOI22_X1 U31 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n107) );
  NAND2_X1 U32 ( .A1(n109), .A2(n108), .ZN(Z[6]) );
  AOI22_X1 U33 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n109) );
  AOI222_X1 U34 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n108) );
  NAND2_X1 U35 ( .A1(n111), .A2(n110), .ZN(Z[7]) );
  AOI22_X1 U36 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n111) );
  AOI222_X1 U37 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n110) );
  NAND2_X1 U38 ( .A1(n113), .A2(n112), .ZN(Z[8]) );
  AOI22_X1 U39 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n113) );
  AOI222_X1 U40 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n112) );
  NAND2_X1 U41 ( .A1(n115), .A2(n114), .ZN(Z[9]) );
  AOI22_X1 U42 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n115) );
  AOI222_X1 U43 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n114) );
  NAND2_X1 U44 ( .A1(n117), .A2(n116), .ZN(Z[10]) );
  AOI22_X1 U45 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n117) );
  AOI222_X1 U46 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), 
        .C2(n79), .ZN(n116) );
  NAND2_X1 U47 ( .A1(n119), .A2(n118), .ZN(Z[11]) );
  AOI22_X1 U48 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n119) );
  AOI222_X1 U49 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), 
        .C2(n79), .ZN(n118) );
  NAND2_X1 U50 ( .A1(n121), .A2(n120), .ZN(Z[12]) );
  AOI22_X1 U51 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n121) );
  AOI222_X1 U52 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), 
        .C2(n80), .ZN(n120) );
  NAND2_X1 U53 ( .A1(n123), .A2(n122), .ZN(Z[13]) );
  AOI22_X1 U54 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n123) );
  AOI222_X1 U55 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), 
        .C2(n80), .ZN(n122) );
  NAND2_X1 U56 ( .A1(n125), .A2(n124), .ZN(Z[14]) );
  AOI22_X1 U57 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n125) );
  AOI222_X1 U58 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n124) );
  NAND2_X1 U59 ( .A1(n127), .A2(n126), .ZN(Z[15]) );
  AOI22_X1 U60 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n127) );
  AOI222_X1 U61 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n126) );
  NAND2_X1 U62 ( .A1(n129), .A2(n128), .ZN(Z[16]) );
  AOI22_X1 U63 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n129) );
  AOI222_X1 U64 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n128) );
  NAND2_X1 U65 ( .A1(n131), .A2(n130), .ZN(Z[17]) );
  AOI22_X1 U66 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n131) );
  AOI222_X1 U67 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n130) );
  NAND2_X1 U68 ( .A1(n133), .A2(n132), .ZN(Z[18]) );
  AOI22_X1 U69 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n133) );
  AOI222_X1 U70 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n132) );
  NAND2_X1 U71 ( .A1(n135), .A2(n134), .ZN(Z[19]) );
  AOI22_X1 U72 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n135) );
  AOI222_X1 U73 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n134) );
  NAND2_X1 U74 ( .A1(n137), .A2(n136), .ZN(Z[20]) );
  AOI22_X1 U75 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n137) );
  AOI222_X1 U76 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n136) );
  NAND2_X1 U77 ( .A1(n139), .A2(n138), .ZN(Z[21]) );
  AOI22_X1 U78 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n139) );
  AOI222_X1 U79 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n138) );
  NAND2_X1 U80 ( .A1(n141), .A2(n140), .ZN(Z[22]) );
  AOI22_X1 U81 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n141) );
  AOI222_X1 U82 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n140) );
  NAND2_X1 U83 ( .A1(n143), .A2(n142), .ZN(Z[23]) );
  AOI22_X1 U84 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n143) );
  AOI222_X1 U85 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n142) );
  NAND2_X1 U86 ( .A1(n145), .A2(n144), .ZN(Z[24]) );
  AOI22_X1 U87 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n145) );
  AOI222_X1 U88 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n144) );
  NAND2_X1 U89 ( .A1(n147), .A2(n146), .ZN(Z[25]) );
  AOI22_X1 U90 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n147) );
  AOI222_X1 U91 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n146) );
  NAND2_X1 U92 ( .A1(n149), .A2(n148), .ZN(Z[26]) );
  AOI22_X1 U93 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n149) );
  AOI222_X1 U94 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n148) );
  NAND2_X1 U95 ( .A1(n151), .A2(n150), .ZN(Z[27]) );
  AOI22_X1 U96 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n151) );
  AOI222_X1 U97 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n150) );
  NAND2_X1 U98 ( .A1(n153), .A2(n152), .ZN(Z[28]) );
  AOI22_X1 U99 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n153) );
  AOI222_X1 U100 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), .C2(n81), .ZN(n152) );
  NAND2_X1 U101 ( .A1(n155), .A2(n154), .ZN(Z[29]) );
  AOI22_X1 U102 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n155) );
  AOI222_X1 U103 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), .C2(n81), .ZN(n154) );
  NAND2_X1 U104 ( .A1(n157), .A2(n156), .ZN(Z[30]) );
  AOI22_X1 U105 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n157) );
  AOI222_X1 U106 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), .C2(n81), .ZN(n156) );
  NAND2_X1 U107 ( .A1(n105), .A2(n104), .ZN(Z[4]) );
  AOI22_X1 U108 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n105) );
  AOI222_X1 U110 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n104) );
  NAND2_X1 U111 ( .A1(n97), .A2(n96), .ZN(Z[0]) );
  AOI22_X1 U112 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n97) );
  AOI222_X1 U113 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n96) );
  NAND2_X1 U114 ( .A1(n99), .A2(n98), .ZN(Z[1]) );
  AOI22_X1 U115 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n99) );
  AOI222_X1 U116 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n98) );
  NAND2_X1 U117 ( .A1(n101), .A2(n100), .ZN(Z[2]) );
  AOI22_X1 U118 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n101) );
  AOI222_X1 U119 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n100) );
  NAND2_X1 U120 ( .A1(n103), .A2(n102), .ZN(Z[3]) );
  AOI22_X1 U121 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n103) );
  AOI222_X1 U122 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n102) );
  NAND2_X1 U123 ( .A1(n163), .A2(n162), .ZN(Z[31]) );
  AOI22_X1 U124 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n163) );
endmodule


module mux5to1_numBit32_5 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  OAI33_X1 U109 ( .A1(n90), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n91), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n160) );
  BUF_X1 U2 ( .A(n158), .Z(n4) );
  BUF_X1 U3 ( .A(n158), .Z(n77) );
  BUF_X1 U4 ( .A(n158), .Z(n78) );
  BUF_X1 U5 ( .A(n89), .Z(n1) );
  BUF_X1 U6 ( .A(n89), .Z(n2) );
  NOR2_X1 U7 ( .A1(n88), .A2(n93), .ZN(n158) );
  INV_X1 U8 ( .A(n94), .ZN(n88) );
  BUF_X1 U9 ( .A(n89), .Z(n3) );
  NOR4_X1 U10 ( .A1(n92), .A2(n85), .A3(n79), .A4(n82), .ZN(n94) );
  BUF_X1 U11 ( .A(n160), .Z(n82) );
  BUF_X1 U12 ( .A(n160), .Z(n83) );
  BUF_X1 U13 ( .A(n159), .Z(n79) );
  BUF_X1 U14 ( .A(n159), .Z(n80) );
  BUF_X1 U15 ( .A(n161), .Z(n85) );
  BUF_X1 U16 ( .A(n161), .Z(n86) );
  BUF_X1 U17 ( .A(n160), .Z(n84) );
  NOR2_X1 U18 ( .A1(n91), .A2(n90), .ZN(n93) );
  BUF_X1 U19 ( .A(n159), .Z(n81) );
  BUF_X1 U20 ( .A(n161), .Z(n87) );
  INV_X1 U21 ( .A(n95), .ZN(n89) );
  AOI21_X1 U22 ( .B1(n94), .B2(n93), .A(n92), .ZN(n95) );
  NOR3_X1 U23 ( .A1(n91), .A2(SEL_in[2]), .A3(n90), .ZN(n161) );
  NOR3_X1 U24 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n92) );
  INV_X1 U25 ( .A(SEL_in[0]), .ZN(n90) );
  AND3_X1 U26 ( .A1(n90), .A2(n91), .A3(SEL_in[2]), .ZN(n159) );
  INV_X1 U27 ( .A(SEL_in[1]), .ZN(n91) );
  NAND2_X1 U28 ( .A1(n111), .A2(n110), .ZN(Z[7]) );
  AOI222_X1 U29 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n110) );
  AOI22_X1 U30 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n111) );
  NAND2_X1 U31 ( .A1(n113), .A2(n112), .ZN(Z[8]) );
  AOI22_X1 U32 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n113) );
  AOI222_X1 U33 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n112) );
  NAND2_X1 U34 ( .A1(n115), .A2(n114), .ZN(Z[9]) );
  AOI22_X1 U35 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n115) );
  AOI222_X1 U36 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n114) );
  NAND2_X1 U37 ( .A1(n117), .A2(n116), .ZN(Z[10]) );
  AOI22_X1 U38 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n117) );
  AOI222_X1 U39 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), 
        .C2(n79), .ZN(n116) );
  NAND2_X1 U40 ( .A1(n119), .A2(n118), .ZN(Z[11]) );
  AOI22_X1 U41 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n119) );
  AOI222_X1 U42 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), 
        .C2(n79), .ZN(n118) );
  NAND2_X1 U43 ( .A1(n121), .A2(n120), .ZN(Z[12]) );
  AOI22_X1 U44 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n121) );
  AOI222_X1 U45 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), 
        .C2(n80), .ZN(n120) );
  NAND2_X1 U46 ( .A1(n123), .A2(n122), .ZN(Z[13]) );
  AOI22_X1 U47 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n123) );
  AOI222_X1 U48 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), 
        .C2(n80), .ZN(n122) );
  NAND2_X1 U49 ( .A1(n125), .A2(n124), .ZN(Z[14]) );
  AOI22_X1 U50 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n125) );
  AOI222_X1 U51 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n124) );
  NAND2_X1 U52 ( .A1(n127), .A2(n126), .ZN(Z[15]) );
  AOI22_X1 U53 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n127) );
  AOI222_X1 U54 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n126) );
  NAND2_X1 U55 ( .A1(n129), .A2(n128), .ZN(Z[16]) );
  AOI22_X1 U56 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n129) );
  AOI222_X1 U57 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n128) );
  NAND2_X1 U58 ( .A1(n131), .A2(n130), .ZN(Z[17]) );
  AOI22_X1 U59 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n131) );
  AOI222_X1 U60 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n130) );
  NAND2_X1 U61 ( .A1(n133), .A2(n132), .ZN(Z[18]) );
  AOI22_X1 U62 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n133) );
  AOI222_X1 U63 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n132) );
  NAND2_X1 U64 ( .A1(n135), .A2(n134), .ZN(Z[19]) );
  AOI22_X1 U65 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n135) );
  AOI222_X1 U66 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n134) );
  NAND2_X1 U67 ( .A1(n137), .A2(n136), .ZN(Z[20]) );
  AOI22_X1 U68 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n137) );
  AOI222_X1 U69 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n136) );
  NAND2_X1 U70 ( .A1(n139), .A2(n138), .ZN(Z[21]) );
  AOI22_X1 U71 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n139) );
  AOI222_X1 U72 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n138) );
  NAND2_X1 U73 ( .A1(n141), .A2(n140), .ZN(Z[22]) );
  AOI22_X1 U74 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n141) );
  AOI222_X1 U75 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n140) );
  NAND2_X1 U76 ( .A1(n143), .A2(n142), .ZN(Z[23]) );
  AOI22_X1 U77 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n143) );
  AOI222_X1 U78 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n142) );
  NAND2_X1 U79 ( .A1(n145), .A2(n144), .ZN(Z[24]) );
  AOI22_X1 U80 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n145) );
  AOI222_X1 U81 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n144) );
  NAND2_X1 U82 ( .A1(n147), .A2(n146), .ZN(Z[25]) );
  AOI22_X1 U83 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n147) );
  AOI222_X1 U84 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n146) );
  NAND2_X1 U85 ( .A1(n149), .A2(n148), .ZN(Z[26]) );
  AOI22_X1 U86 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n149) );
  AOI222_X1 U87 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n148) );
  NAND2_X1 U88 ( .A1(n151), .A2(n150), .ZN(Z[27]) );
  AOI22_X1 U89 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n151) );
  AOI222_X1 U90 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n150) );
  NAND2_X1 U91 ( .A1(n153), .A2(n152), .ZN(Z[28]) );
  AOI22_X1 U92 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n153) );
  AOI222_X1 U93 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), 
        .C2(n81), .ZN(n152) );
  NAND2_X1 U94 ( .A1(n155), .A2(n154), .ZN(Z[29]) );
  AOI22_X1 U95 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n155) );
  AOI222_X1 U96 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), 
        .C2(n81), .ZN(n154) );
  NAND2_X1 U97 ( .A1(n157), .A2(n156), .ZN(Z[30]) );
  AOI22_X1 U98 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n157) );
  AOI222_X1 U99 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), 
        .C2(n81), .ZN(n156) );
  NAND2_X1 U100 ( .A1(n109), .A2(n108), .ZN(Z[6]) );
  AOI22_X1 U101 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n109) );
  AOI222_X1 U102 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n108) );
  NAND2_X1 U103 ( .A1(n97), .A2(n96), .ZN(Z[0]) );
  AOI22_X1 U104 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n97) );
  AOI222_X1 U105 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n96) );
  NAND2_X1 U106 ( .A1(n99), .A2(n98), .ZN(Z[1]) );
  AOI22_X1 U107 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n99) );
  AOI222_X1 U108 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n98) );
  NAND2_X1 U110 ( .A1(n101), .A2(n100), .ZN(Z[2]) );
  AOI22_X1 U111 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n101) );
  AOI222_X1 U112 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n100) );
  NAND2_X1 U113 ( .A1(n103), .A2(n102), .ZN(Z[3]) );
  AOI22_X1 U114 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n103) );
  AOI222_X1 U115 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n102) );
  NAND2_X1 U116 ( .A1(n105), .A2(n104), .ZN(Z[4]) );
  AOI22_X1 U117 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n105) );
  AOI222_X1 U118 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n104) );
  NAND2_X1 U119 ( .A1(n107), .A2(n106), .ZN(Z[5]) );
  AOI22_X1 U120 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n107) );
  AOI222_X1 U121 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n106) );
  NAND2_X1 U122 ( .A1(n163), .A2(n162), .ZN(Z[31]) );
  AOI22_X1 U123 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n163) );
  AOI222_X1 U124 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), .C2(n81), .ZN(n162) );
endmodule


module mux5to1_numBit32_4 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  OAI33_X1 U109 ( .A1(n90), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n91), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n160) );
  BUF_X1 U2 ( .A(n158), .Z(n4) );
  BUF_X1 U3 ( .A(n158), .Z(n77) );
  BUF_X1 U4 ( .A(n158), .Z(n78) );
  AOI222_X1 U5 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), 
        .C2(n81), .ZN(n162) );
  BUF_X1 U6 ( .A(n89), .Z(n1) );
  BUF_X1 U7 ( .A(n89), .Z(n2) );
  NOR2_X1 U8 ( .A1(n88), .A2(n93), .ZN(n158) );
  INV_X1 U9 ( .A(n94), .ZN(n88) );
  BUF_X1 U10 ( .A(n89), .Z(n3) );
  NOR4_X1 U11 ( .A1(n92), .A2(n85), .A3(n79), .A4(n82), .ZN(n94) );
  BUF_X1 U12 ( .A(n160), .Z(n82) );
  BUF_X1 U13 ( .A(n160), .Z(n83) );
  BUF_X1 U14 ( .A(n159), .Z(n79) );
  BUF_X1 U15 ( .A(n159), .Z(n80) );
  BUF_X1 U16 ( .A(n161), .Z(n85) );
  BUF_X1 U17 ( .A(n161), .Z(n86) );
  BUF_X1 U18 ( .A(n160), .Z(n84) );
  NOR2_X1 U19 ( .A1(n91), .A2(n90), .ZN(n93) );
  BUF_X1 U20 ( .A(n159), .Z(n81) );
  BUF_X1 U21 ( .A(n161), .Z(n87) );
  INV_X1 U22 ( .A(n95), .ZN(n89) );
  AOI21_X1 U23 ( .B1(n94), .B2(n93), .A(n92), .ZN(n95) );
  NOR3_X1 U24 ( .A1(n91), .A2(SEL_in[2]), .A3(n90), .ZN(n161) );
  NOR3_X1 U25 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n92) );
  INV_X1 U26 ( .A(SEL_in[0]), .ZN(n90) );
  AND3_X1 U27 ( .A1(n90), .A2(n91), .A3(SEL_in[2]), .ZN(n159) );
  INV_X1 U28 ( .A(SEL_in[1]), .ZN(n91) );
  NAND2_X1 U29 ( .A1(n115), .A2(n114), .ZN(Z[9]) );
  AOI222_X1 U30 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n114) );
  AOI22_X1 U31 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n115) );
  NAND2_X1 U32 ( .A1(n117), .A2(n116), .ZN(Z[10]) );
  AOI22_X1 U33 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n117) );
  AOI222_X1 U34 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), 
        .C2(n79), .ZN(n116) );
  NAND2_X1 U35 ( .A1(n119), .A2(n118), .ZN(Z[11]) );
  AOI22_X1 U36 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n119) );
  AOI222_X1 U37 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), 
        .C2(n79), .ZN(n118) );
  NAND2_X1 U38 ( .A1(n121), .A2(n120), .ZN(Z[12]) );
  AOI22_X1 U39 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n121) );
  AOI222_X1 U40 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), 
        .C2(n80), .ZN(n120) );
  NAND2_X1 U41 ( .A1(n123), .A2(n122), .ZN(Z[13]) );
  AOI22_X1 U42 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n123) );
  AOI222_X1 U43 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), 
        .C2(n80), .ZN(n122) );
  NAND2_X1 U44 ( .A1(n125), .A2(n124), .ZN(Z[14]) );
  AOI22_X1 U45 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n125) );
  AOI222_X1 U46 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n124) );
  NAND2_X1 U47 ( .A1(n127), .A2(n126), .ZN(Z[15]) );
  AOI22_X1 U48 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n127) );
  AOI222_X1 U49 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n126) );
  NAND2_X1 U50 ( .A1(n129), .A2(n128), .ZN(Z[16]) );
  AOI22_X1 U51 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n129) );
  AOI222_X1 U52 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n128) );
  NAND2_X1 U53 ( .A1(n131), .A2(n130), .ZN(Z[17]) );
  AOI22_X1 U54 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n131) );
  AOI222_X1 U55 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n130) );
  NAND2_X1 U56 ( .A1(n133), .A2(n132), .ZN(Z[18]) );
  AOI22_X1 U57 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n133) );
  AOI222_X1 U58 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n132) );
  NAND2_X1 U59 ( .A1(n135), .A2(n134), .ZN(Z[19]) );
  AOI22_X1 U60 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n135) );
  AOI222_X1 U61 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n134) );
  NAND2_X1 U62 ( .A1(n137), .A2(n136), .ZN(Z[20]) );
  AOI22_X1 U63 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n137) );
  AOI222_X1 U64 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n136) );
  NAND2_X1 U65 ( .A1(n139), .A2(n138), .ZN(Z[21]) );
  AOI22_X1 U66 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n139) );
  AOI222_X1 U67 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n138) );
  NAND2_X1 U68 ( .A1(n141), .A2(n140), .ZN(Z[22]) );
  AOI22_X1 U69 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n141) );
  AOI222_X1 U70 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n140) );
  NAND2_X1 U71 ( .A1(n143), .A2(n142), .ZN(Z[23]) );
  AOI22_X1 U72 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n143) );
  AOI222_X1 U73 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n142) );
  NAND2_X1 U74 ( .A1(n145), .A2(n144), .ZN(Z[24]) );
  AOI22_X1 U75 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n145) );
  AOI222_X1 U76 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n144) );
  NAND2_X1 U77 ( .A1(n147), .A2(n146), .ZN(Z[25]) );
  AOI22_X1 U78 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n147) );
  AOI222_X1 U79 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n146) );
  NAND2_X1 U80 ( .A1(n149), .A2(n148), .ZN(Z[26]) );
  AOI22_X1 U81 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n149) );
  AOI222_X1 U82 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n148) );
  NAND2_X1 U83 ( .A1(n151), .A2(n150), .ZN(Z[27]) );
  AOI22_X1 U84 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n151) );
  AOI222_X1 U85 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n150) );
  NAND2_X1 U86 ( .A1(n153), .A2(n152), .ZN(Z[28]) );
  AOI22_X1 U87 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n153) );
  AOI222_X1 U88 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), 
        .C2(n81), .ZN(n152) );
  NAND2_X1 U89 ( .A1(n155), .A2(n154), .ZN(Z[29]) );
  AOI22_X1 U90 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n155) );
  AOI222_X1 U91 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), 
        .C2(n81), .ZN(n154) );
  NAND2_X1 U92 ( .A1(n157), .A2(n156), .ZN(Z[30]) );
  AOI22_X1 U93 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n157) );
  AOI222_X1 U94 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), 
        .C2(n81), .ZN(n156) );
  NAND2_X1 U95 ( .A1(n113), .A2(n112), .ZN(Z[8]) );
  AOI22_X1 U96 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n113) );
  AOI222_X1 U97 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n112) );
  NAND2_X1 U98 ( .A1(n97), .A2(n96), .ZN(Z[0]) );
  AOI22_X1 U99 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n97) );
  AOI222_X1 U100 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n96) );
  NAND2_X1 U101 ( .A1(n99), .A2(n98), .ZN(Z[1]) );
  AOI22_X1 U102 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n99) );
  AOI222_X1 U103 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n98) );
  NAND2_X1 U104 ( .A1(n101), .A2(n100), .ZN(Z[2]) );
  AOI22_X1 U105 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n101) );
  AOI222_X1 U106 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n100) );
  NAND2_X1 U107 ( .A1(n103), .A2(n102), .ZN(Z[3]) );
  AOI22_X1 U108 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n103) );
  AOI222_X1 U110 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n102) );
  NAND2_X1 U111 ( .A1(n105), .A2(n104), .ZN(Z[4]) );
  AOI22_X1 U112 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n105) );
  AOI222_X1 U113 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n104) );
  NAND2_X1 U114 ( .A1(n107), .A2(n106), .ZN(Z[5]) );
  AOI22_X1 U115 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n107) );
  AOI222_X1 U116 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n106) );
  NAND2_X1 U117 ( .A1(n109), .A2(n108), .ZN(Z[6]) );
  AOI22_X1 U118 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n109) );
  AOI222_X1 U119 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n108) );
  NAND2_X1 U120 ( .A1(n111), .A2(n110), .ZN(Z[7]) );
  AOI22_X1 U121 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n111) );
  AOI222_X1 U122 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n110) );
  NAND2_X1 U123 ( .A1(n163), .A2(n162), .ZN(Z[31]) );
  AOI22_X1 U124 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n163) );
endmodule


module mux5to1_numBit32_3 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  OAI33_X1 U109 ( .A1(n91), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n90), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n160) );
  BUF_X1 U2 ( .A(n158), .Z(n4) );
  BUF_X1 U3 ( .A(n158), .Z(n77) );
  BUF_X1 U4 ( .A(n158), .Z(n78) );
  BUF_X1 U5 ( .A(n89), .Z(n1) );
  BUF_X1 U6 ( .A(n89), .Z(n2) );
  NOR2_X1 U7 ( .A1(n88), .A2(n93), .ZN(n158) );
  INV_X1 U8 ( .A(n94), .ZN(n88) );
  BUF_X1 U9 ( .A(n89), .Z(n3) );
  NOR4_X1 U10 ( .A1(n92), .A2(n85), .A3(n79), .A4(n82), .ZN(n94) );
  BUF_X1 U11 ( .A(n160), .Z(n82) );
  BUF_X1 U12 ( .A(n160), .Z(n83) );
  BUF_X1 U13 ( .A(n159), .Z(n79) );
  BUF_X1 U14 ( .A(n159), .Z(n80) );
  BUF_X1 U15 ( .A(n161), .Z(n85) );
  BUF_X1 U16 ( .A(n161), .Z(n86) );
  BUF_X1 U17 ( .A(n160), .Z(n84) );
  NOR2_X1 U18 ( .A1(n90), .A2(n91), .ZN(n93) );
  BUF_X1 U19 ( .A(n159), .Z(n81) );
  BUF_X1 U20 ( .A(n161), .Z(n87) );
  INV_X1 U21 ( .A(n95), .ZN(n89) );
  AOI21_X1 U22 ( .B1(n94), .B2(n93), .A(n92), .ZN(n95) );
  NOR3_X1 U23 ( .A1(n90), .A2(SEL_in[2]), .A3(n91), .ZN(n161) );
  NOR3_X1 U24 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n92) );
  INV_X1 U25 ( .A(SEL_in[0]), .ZN(n91) );
  AND3_X1 U26 ( .A1(n91), .A2(n90), .A3(SEL_in[2]), .ZN(n159) );
  INV_X1 U27 ( .A(SEL_in[1]), .ZN(n90) );
  NAND2_X1 U28 ( .A1(n119), .A2(n118), .ZN(Z[11]) );
  AOI222_X1 U29 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), 
        .C2(n79), .ZN(n118) );
  AOI22_X1 U30 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n119) );
  NAND2_X1 U31 ( .A1(n121), .A2(n120), .ZN(Z[12]) );
  AOI22_X1 U32 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n121) );
  AOI222_X1 U33 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), 
        .C2(n80), .ZN(n120) );
  NAND2_X1 U34 ( .A1(n123), .A2(n122), .ZN(Z[13]) );
  AOI22_X1 U35 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n123) );
  AOI222_X1 U36 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), 
        .C2(n80), .ZN(n122) );
  NAND2_X1 U37 ( .A1(n125), .A2(n124), .ZN(Z[14]) );
  AOI22_X1 U38 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n125) );
  AOI222_X1 U39 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n124) );
  NAND2_X1 U40 ( .A1(n127), .A2(n126), .ZN(Z[15]) );
  AOI22_X1 U41 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n127) );
  AOI222_X1 U42 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n126) );
  NAND2_X1 U43 ( .A1(n129), .A2(n128), .ZN(Z[16]) );
  AOI22_X1 U44 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n129) );
  AOI222_X1 U45 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n128) );
  NAND2_X1 U46 ( .A1(n131), .A2(n130), .ZN(Z[17]) );
  AOI22_X1 U47 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n131) );
  AOI222_X1 U48 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n130) );
  NAND2_X1 U49 ( .A1(n133), .A2(n132), .ZN(Z[18]) );
  AOI22_X1 U50 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n133) );
  AOI222_X1 U51 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n132) );
  NAND2_X1 U52 ( .A1(n135), .A2(n134), .ZN(Z[19]) );
  AOI22_X1 U53 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n135) );
  AOI222_X1 U54 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n134) );
  NAND2_X1 U55 ( .A1(n137), .A2(n136), .ZN(Z[20]) );
  AOI22_X1 U56 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n137) );
  AOI222_X1 U57 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n136) );
  NAND2_X1 U58 ( .A1(n139), .A2(n138), .ZN(Z[21]) );
  AOI22_X1 U59 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n139) );
  AOI222_X1 U60 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n138) );
  NAND2_X1 U61 ( .A1(n141), .A2(n140), .ZN(Z[22]) );
  AOI22_X1 U62 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n141) );
  AOI222_X1 U63 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n140) );
  NAND2_X1 U64 ( .A1(n143), .A2(n142), .ZN(Z[23]) );
  AOI22_X1 U65 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n143) );
  AOI222_X1 U66 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n142) );
  NAND2_X1 U67 ( .A1(n145), .A2(n144), .ZN(Z[24]) );
  AOI22_X1 U68 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n145) );
  AOI222_X1 U69 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n144) );
  NAND2_X1 U70 ( .A1(n147), .A2(n146), .ZN(Z[25]) );
  AOI22_X1 U71 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n147) );
  AOI222_X1 U72 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n146) );
  NAND2_X1 U73 ( .A1(n149), .A2(n148), .ZN(Z[26]) );
  AOI22_X1 U74 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n149) );
  AOI222_X1 U75 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n148) );
  NAND2_X1 U76 ( .A1(n151), .A2(n150), .ZN(Z[27]) );
  AOI22_X1 U77 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n151) );
  AOI222_X1 U78 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n150) );
  NAND2_X1 U79 ( .A1(n153), .A2(n152), .ZN(Z[28]) );
  AOI22_X1 U80 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n153) );
  AOI222_X1 U81 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), 
        .C2(n81), .ZN(n152) );
  NAND2_X1 U82 ( .A1(n155), .A2(n154), .ZN(Z[29]) );
  AOI22_X1 U83 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n155) );
  AOI222_X1 U84 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), 
        .C2(n81), .ZN(n154) );
  NAND2_X1 U85 ( .A1(n157), .A2(n156), .ZN(Z[30]) );
  AOI22_X1 U86 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n157) );
  AOI222_X1 U87 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), 
        .C2(n81), .ZN(n156) );
  NAND2_X1 U88 ( .A1(n117), .A2(n116), .ZN(Z[10]) );
  AOI22_X1 U89 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n117) );
  AOI222_X1 U90 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), 
        .C2(n79), .ZN(n116) );
  NAND2_X1 U91 ( .A1(n97), .A2(n96), .ZN(Z[0]) );
  AOI22_X1 U92 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n97) );
  AOI222_X1 U93 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n96) );
  NAND2_X1 U94 ( .A1(n99), .A2(n98), .ZN(Z[1]) );
  AOI22_X1 U95 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n99) );
  AOI222_X1 U96 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n98) );
  NAND2_X1 U97 ( .A1(n101), .A2(n100), .ZN(Z[2]) );
  AOI22_X1 U98 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n101) );
  AOI222_X1 U99 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n100) );
  NAND2_X1 U100 ( .A1(n103), .A2(n102), .ZN(Z[3]) );
  AOI22_X1 U101 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n103) );
  AOI222_X1 U102 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n102) );
  NAND2_X1 U103 ( .A1(n105), .A2(n104), .ZN(Z[4]) );
  AOI22_X1 U104 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n105) );
  AOI222_X1 U105 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n104) );
  NAND2_X1 U106 ( .A1(n107), .A2(n106), .ZN(Z[5]) );
  AOI22_X1 U107 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n107) );
  AOI222_X1 U108 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n106) );
  NAND2_X1 U110 ( .A1(n109), .A2(n108), .ZN(Z[6]) );
  AOI22_X1 U111 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n109) );
  AOI222_X1 U112 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n108) );
  NAND2_X1 U113 ( .A1(n111), .A2(n110), .ZN(Z[7]) );
  AOI22_X1 U114 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n111) );
  AOI222_X1 U115 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n110) );
  NAND2_X1 U116 ( .A1(n113), .A2(n112), .ZN(Z[8]) );
  AOI22_X1 U117 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n113) );
  AOI222_X1 U118 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n112) );
  NAND2_X1 U119 ( .A1(n115), .A2(n114), .ZN(Z[9]) );
  AOI22_X1 U120 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n115) );
  AOI222_X1 U121 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n114) );
  NAND2_X1 U122 ( .A1(n163), .A2(n162), .ZN(Z[31]) );
  AOI22_X1 U123 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n163) );
  AOI222_X1 U124 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), .C2(n81), .ZN(n162) );
endmodule


module mux5to1_numBit32_2 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  OAI33_X1 U109 ( .A1(n90), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n91), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n160) );
  BUF_X1 U2 ( .A(n158), .Z(n4) );
  BUF_X1 U3 ( .A(n158), .Z(n77) );
  BUF_X1 U4 ( .A(n158), .Z(n78) );
  AOI222_X1 U5 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), 
        .C2(n81), .ZN(n162) );
  BUF_X1 U6 ( .A(n89), .Z(n1) );
  BUF_X1 U7 ( .A(n89), .Z(n2) );
  NOR2_X1 U8 ( .A1(n88), .A2(n93), .ZN(n158) );
  INV_X1 U9 ( .A(n94), .ZN(n88) );
  BUF_X1 U10 ( .A(n89), .Z(n3) );
  NOR4_X1 U11 ( .A1(n92), .A2(n85), .A3(n79), .A4(n82), .ZN(n94) );
  BUF_X1 U12 ( .A(n160), .Z(n82) );
  BUF_X1 U13 ( .A(n160), .Z(n83) );
  BUF_X1 U14 ( .A(n159), .Z(n79) );
  BUF_X1 U15 ( .A(n159), .Z(n80) );
  BUF_X1 U16 ( .A(n161), .Z(n85) );
  BUF_X1 U17 ( .A(n161), .Z(n86) );
  BUF_X1 U18 ( .A(n160), .Z(n84) );
  NOR2_X1 U19 ( .A1(n91), .A2(n90), .ZN(n93) );
  BUF_X1 U20 ( .A(n159), .Z(n81) );
  BUF_X1 U21 ( .A(n161), .Z(n87) );
  INV_X1 U22 ( .A(n95), .ZN(n89) );
  AOI21_X1 U23 ( .B1(n94), .B2(n93), .A(n92), .ZN(n95) );
  NOR3_X1 U24 ( .A1(n91), .A2(SEL_in[2]), .A3(n90), .ZN(n161) );
  NOR3_X1 U25 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n92) );
  INV_X1 U26 ( .A(SEL_in[0]), .ZN(n90) );
  AND3_X1 U27 ( .A1(n90), .A2(n91), .A3(SEL_in[2]), .ZN(n159) );
  INV_X1 U28 ( .A(SEL_in[1]), .ZN(n91) );
  NAND2_X1 U29 ( .A1(n123), .A2(n122), .ZN(Z[13]) );
  AOI222_X1 U30 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), 
        .C2(n80), .ZN(n122) );
  AOI22_X1 U31 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n123) );
  NAND2_X1 U32 ( .A1(n125), .A2(n124), .ZN(Z[14]) );
  AOI22_X1 U33 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n125) );
  AOI222_X1 U34 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n124) );
  NAND2_X1 U35 ( .A1(n127), .A2(n126), .ZN(Z[15]) );
  AOI22_X1 U36 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n127) );
  AOI222_X1 U37 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n126) );
  NAND2_X1 U38 ( .A1(n129), .A2(n128), .ZN(Z[16]) );
  AOI22_X1 U39 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n129) );
  AOI222_X1 U40 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n128) );
  NAND2_X1 U41 ( .A1(n131), .A2(n130), .ZN(Z[17]) );
  AOI22_X1 U42 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n131) );
  AOI222_X1 U43 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n130) );
  NAND2_X1 U44 ( .A1(n133), .A2(n132), .ZN(Z[18]) );
  AOI22_X1 U45 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n133) );
  AOI222_X1 U46 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n132) );
  NAND2_X1 U47 ( .A1(n135), .A2(n134), .ZN(Z[19]) );
  AOI22_X1 U48 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n135) );
  AOI222_X1 U49 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n134) );
  NAND2_X1 U50 ( .A1(n137), .A2(n136), .ZN(Z[20]) );
  AOI22_X1 U51 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n137) );
  AOI222_X1 U52 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n136) );
  NAND2_X1 U53 ( .A1(n139), .A2(n138), .ZN(Z[21]) );
  AOI22_X1 U54 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n139) );
  AOI222_X1 U55 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n138) );
  NAND2_X1 U56 ( .A1(n141), .A2(n140), .ZN(Z[22]) );
  AOI22_X1 U57 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n141) );
  AOI222_X1 U58 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n140) );
  NAND2_X1 U59 ( .A1(n143), .A2(n142), .ZN(Z[23]) );
  AOI22_X1 U60 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n143) );
  AOI222_X1 U61 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n142) );
  NAND2_X1 U62 ( .A1(n145), .A2(n144), .ZN(Z[24]) );
  AOI22_X1 U63 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n145) );
  AOI222_X1 U64 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n144) );
  NAND2_X1 U65 ( .A1(n147), .A2(n146), .ZN(Z[25]) );
  AOI22_X1 U66 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n147) );
  AOI222_X1 U67 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n146) );
  NAND2_X1 U68 ( .A1(n149), .A2(n148), .ZN(Z[26]) );
  AOI22_X1 U69 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n149) );
  AOI222_X1 U70 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n148) );
  NAND2_X1 U71 ( .A1(n151), .A2(n150), .ZN(Z[27]) );
  AOI22_X1 U72 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n151) );
  AOI222_X1 U73 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n150) );
  NAND2_X1 U74 ( .A1(n153), .A2(n152), .ZN(Z[28]) );
  AOI22_X1 U75 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n153) );
  AOI222_X1 U76 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), 
        .C2(n81), .ZN(n152) );
  NAND2_X1 U77 ( .A1(n155), .A2(n154), .ZN(Z[29]) );
  AOI22_X1 U78 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n155) );
  AOI222_X1 U79 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), 
        .C2(n81), .ZN(n154) );
  NAND2_X1 U80 ( .A1(n157), .A2(n156), .ZN(Z[30]) );
  AOI22_X1 U81 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n157) );
  AOI222_X1 U82 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), 
        .C2(n81), .ZN(n156) );
  NAND2_X1 U83 ( .A1(n121), .A2(n120), .ZN(Z[12]) );
  AOI22_X1 U84 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n121) );
  AOI222_X1 U85 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), 
        .C2(n80), .ZN(n120) );
  NAND2_X1 U86 ( .A1(n97), .A2(n96), .ZN(Z[0]) );
  AOI22_X1 U87 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n97) );
  AOI222_X1 U88 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n96) );
  NAND2_X1 U89 ( .A1(n99), .A2(n98), .ZN(Z[1]) );
  AOI22_X1 U90 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n99) );
  AOI222_X1 U91 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n98) );
  NAND2_X1 U92 ( .A1(n101), .A2(n100), .ZN(Z[2]) );
  AOI22_X1 U93 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n101) );
  AOI222_X1 U94 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n100) );
  NAND2_X1 U95 ( .A1(n103), .A2(n102), .ZN(Z[3]) );
  AOI22_X1 U96 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n103) );
  AOI222_X1 U97 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n102) );
  NAND2_X1 U98 ( .A1(n105), .A2(n104), .ZN(Z[4]) );
  AOI22_X1 U99 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n105) );
  AOI222_X1 U100 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n104) );
  NAND2_X1 U101 ( .A1(n107), .A2(n106), .ZN(Z[5]) );
  AOI22_X1 U102 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n107) );
  AOI222_X1 U103 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n106) );
  NAND2_X1 U104 ( .A1(n109), .A2(n108), .ZN(Z[6]) );
  AOI22_X1 U105 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n109) );
  AOI222_X1 U106 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n108) );
  NAND2_X1 U107 ( .A1(n111), .A2(n110), .ZN(Z[7]) );
  AOI22_X1 U108 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n111) );
  AOI222_X1 U110 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n110) );
  NAND2_X1 U111 ( .A1(n113), .A2(n112), .ZN(Z[8]) );
  AOI22_X1 U112 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n113) );
  AOI222_X1 U113 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n112) );
  NAND2_X1 U114 ( .A1(n115), .A2(n114), .ZN(Z[9]) );
  AOI22_X1 U115 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n115) );
  AOI222_X1 U116 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n114) );
  NAND2_X1 U117 ( .A1(n117), .A2(n116), .ZN(Z[10]) );
  AOI22_X1 U118 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n117) );
  AOI222_X1 U119 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), .C2(n79), .ZN(n116) );
  NAND2_X1 U120 ( .A1(n119), .A2(n118), .ZN(Z[11]) );
  AOI22_X1 U121 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n119) );
  AOI222_X1 U122 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), .C2(n79), .ZN(n118) );
  NAND2_X1 U123 ( .A1(n163), .A2(n162), .ZN(Z[31]) );
  AOI22_X1 U124 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n163) );
endmodule


module mux5to1_numBit32_1 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  OAI33_X1 U109 ( .A1(n90), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n91), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n160) );
  BUF_X1 U2 ( .A(n158), .Z(n4) );
  BUF_X1 U3 ( .A(n158), .Z(n77) );
  BUF_X1 U4 ( .A(n158), .Z(n78) );
  BUF_X1 U5 ( .A(n89), .Z(n1) );
  BUF_X1 U6 ( .A(n89), .Z(n2) );
  NOR2_X1 U7 ( .A1(n88), .A2(n93), .ZN(n158) );
  INV_X1 U8 ( .A(n94), .ZN(n88) );
  BUF_X1 U9 ( .A(n89), .Z(n3) );
  NOR4_X1 U10 ( .A1(n92), .A2(n85), .A3(n79), .A4(n82), .ZN(n94) );
  BUF_X1 U11 ( .A(n160), .Z(n82) );
  BUF_X1 U12 ( .A(n160), .Z(n83) );
  BUF_X1 U13 ( .A(n159), .Z(n79) );
  BUF_X1 U14 ( .A(n159), .Z(n80) );
  BUF_X1 U15 ( .A(n161), .Z(n85) );
  BUF_X1 U16 ( .A(n161), .Z(n86) );
  BUF_X1 U17 ( .A(n160), .Z(n84) );
  NOR2_X1 U18 ( .A1(n91), .A2(n90), .ZN(n93) );
  BUF_X1 U19 ( .A(n159), .Z(n81) );
  BUF_X1 U20 ( .A(n161), .Z(n87) );
  INV_X1 U21 ( .A(n95), .ZN(n89) );
  AOI21_X1 U22 ( .B1(n94), .B2(n93), .A(n92), .ZN(n95) );
  NOR3_X1 U23 ( .A1(n91), .A2(SEL_in[2]), .A3(n90), .ZN(n161) );
  NOR3_X1 U24 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n92) );
  INV_X1 U25 ( .A(SEL_in[0]), .ZN(n90) );
  AND3_X1 U26 ( .A1(n90), .A2(n91), .A3(SEL_in[2]), .ZN(n159) );
  INV_X1 U27 ( .A(SEL_in[1]), .ZN(n91) );
  NAND2_X1 U28 ( .A1(n127), .A2(n126), .ZN(Z[15]) );
  AOI222_X1 U29 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n126) );
  AOI22_X1 U30 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n127) );
  NAND2_X1 U31 ( .A1(n129), .A2(n128), .ZN(Z[16]) );
  AOI22_X1 U32 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n129) );
  AOI222_X1 U33 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n128) );
  NAND2_X1 U34 ( .A1(n131), .A2(n130), .ZN(Z[17]) );
  AOI22_X1 U35 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n131) );
  AOI222_X1 U36 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n130) );
  NAND2_X1 U37 ( .A1(n133), .A2(n132), .ZN(Z[18]) );
  AOI22_X1 U38 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n133) );
  AOI222_X1 U39 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n132) );
  NAND2_X1 U40 ( .A1(n135), .A2(n134), .ZN(Z[19]) );
  AOI22_X1 U41 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n135) );
  AOI222_X1 U42 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n134) );
  NAND2_X1 U43 ( .A1(n137), .A2(n136), .ZN(Z[20]) );
  AOI22_X1 U44 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n137) );
  AOI222_X1 U45 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n136) );
  NAND2_X1 U46 ( .A1(n139), .A2(n138), .ZN(Z[21]) );
  AOI22_X1 U47 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n139) );
  AOI222_X1 U48 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n138) );
  NAND2_X1 U49 ( .A1(n141), .A2(n140), .ZN(Z[22]) );
  AOI22_X1 U50 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n141) );
  AOI222_X1 U51 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n140) );
  NAND2_X1 U52 ( .A1(n143), .A2(n142), .ZN(Z[23]) );
  AOI22_X1 U53 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n143) );
  AOI222_X1 U54 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n142) );
  NAND2_X1 U55 ( .A1(n145), .A2(n144), .ZN(Z[24]) );
  AOI22_X1 U56 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n145) );
  AOI222_X1 U57 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n144) );
  NAND2_X1 U58 ( .A1(n147), .A2(n146), .ZN(Z[25]) );
  AOI22_X1 U59 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n147) );
  AOI222_X1 U60 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n146) );
  NAND2_X1 U61 ( .A1(n149), .A2(n148), .ZN(Z[26]) );
  AOI22_X1 U62 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n149) );
  AOI222_X1 U63 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n148) );
  NAND2_X1 U64 ( .A1(n151), .A2(n150), .ZN(Z[27]) );
  AOI22_X1 U65 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n151) );
  AOI222_X1 U66 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n150) );
  NAND2_X1 U67 ( .A1(n153), .A2(n152), .ZN(Z[28]) );
  AOI22_X1 U68 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n153) );
  AOI222_X1 U69 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), 
        .C2(n81), .ZN(n152) );
  NAND2_X1 U70 ( .A1(n155), .A2(n154), .ZN(Z[29]) );
  AOI22_X1 U71 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n155) );
  AOI222_X1 U72 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), 
        .C2(n81), .ZN(n154) );
  NAND2_X1 U73 ( .A1(n157), .A2(n156), .ZN(Z[30]) );
  AOI22_X1 U74 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n157) );
  AOI222_X1 U75 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), 
        .C2(n81), .ZN(n156) );
  NAND2_X1 U76 ( .A1(n125), .A2(n124), .ZN(Z[14]) );
  AOI22_X1 U77 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n125) );
  AOI222_X1 U78 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n124) );
  NAND2_X1 U79 ( .A1(n97), .A2(n96), .ZN(Z[0]) );
  AOI22_X1 U80 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n97) );
  AOI222_X1 U81 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n96) );
  NAND2_X1 U82 ( .A1(n99), .A2(n98), .ZN(Z[1]) );
  AOI22_X1 U83 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n99) );
  AOI222_X1 U84 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n98) );
  NAND2_X1 U85 ( .A1(n101), .A2(n100), .ZN(Z[2]) );
  AOI22_X1 U86 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n101) );
  AOI222_X1 U87 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n100) );
  NAND2_X1 U88 ( .A1(n103), .A2(n102), .ZN(Z[3]) );
  AOI22_X1 U89 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n103) );
  AOI222_X1 U90 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n102) );
  NAND2_X1 U91 ( .A1(n105), .A2(n104), .ZN(Z[4]) );
  AOI22_X1 U92 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n105) );
  AOI222_X1 U93 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n104) );
  NAND2_X1 U94 ( .A1(n107), .A2(n106), .ZN(Z[5]) );
  AOI22_X1 U95 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n107) );
  AOI222_X1 U96 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n106) );
  NAND2_X1 U97 ( .A1(n109), .A2(n108), .ZN(Z[6]) );
  AOI22_X1 U98 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n109) );
  AOI222_X1 U99 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n108) );
  NAND2_X1 U100 ( .A1(n111), .A2(n110), .ZN(Z[7]) );
  AOI22_X1 U101 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n111) );
  AOI222_X1 U102 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n110) );
  NAND2_X1 U103 ( .A1(n113), .A2(n112), .ZN(Z[8]) );
  AOI22_X1 U104 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n113) );
  AOI222_X1 U105 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n112) );
  NAND2_X1 U106 ( .A1(n115), .A2(n114), .ZN(Z[9]) );
  AOI22_X1 U107 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n115) );
  AOI222_X1 U108 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n114) );
  NAND2_X1 U110 ( .A1(n117), .A2(n116), .ZN(Z[10]) );
  AOI22_X1 U111 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n117) );
  AOI222_X1 U112 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), .C2(n79), .ZN(n116) );
  NAND2_X1 U113 ( .A1(n119), .A2(n118), .ZN(Z[11]) );
  AOI22_X1 U114 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n119) );
  AOI222_X1 U115 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), .C2(n79), .ZN(n118) );
  NAND2_X1 U116 ( .A1(n121), .A2(n120), .ZN(Z[12]) );
  AOI22_X1 U117 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n121) );
  AOI222_X1 U118 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), .C2(n80), .ZN(n120) );
  NAND2_X1 U119 ( .A1(n123), .A2(n122), .ZN(Z[13]) );
  AOI22_X1 U120 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n123) );
  AOI222_X1 U121 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), .C2(n80), .ZN(n122) );
  NAND2_X1 U122 ( .A1(n163), .A2(n162), .ZN(Z[31]) );
  AOI22_X1 U123 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n163) );
  AOI222_X1 U124 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), .C2(n81), .ZN(n162) );
endmodule


module rca_bhv_numBit32_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;

  wire   [32:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module rca_bhv_numBit32_0 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;


  rca_bhv_numBit32_0_DW01_add_0 add_1_root_add_35_2 ( .A({A[31], A}), .B({
        B[31], B}), .CI(Ci), .SUM({Co, S}) );
endmodule


module rca_bhv_numBit32_6_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;

  wire   [32:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module rca_bhv_numBit32_6 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;


  rca_bhv_numBit32_6_DW01_add_0 add_1_root_add_35_2 ( .A({A[31], A}), .B({
        B[31], B}), .CI(Ci), .SUM({Co, S}) );
endmodule


module rca_bhv_numBit32_5_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;

  wire   [32:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module rca_bhv_numBit32_5 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;


  rca_bhv_numBit32_5_DW01_add_0 add_1_root_add_35_2 ( .A({A[31], A}), .B({
        B[31], B}), .CI(Ci), .SUM({Co, S}) );
endmodule


module rca_bhv_numBit32_4_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;

  wire   [32:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module rca_bhv_numBit32_4 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;


  rca_bhv_numBit32_4_DW01_add_0 add_1_root_add_35_2 ( .A({A[31], A}), .B({
        B[31], B}), .CI(Ci), .SUM({Co, S}) );
endmodule


module rca_bhv_numBit32_3_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;

  wire   [32:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module rca_bhv_numBit32_3 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;


  rca_bhv_numBit32_3_DW01_add_0 add_1_root_add_35_2 ( .A({A[31], A}), .B({
        B[31], B}), .CI(Ci), .SUM({Co, S}) );
endmodule


module rca_bhv_numBit32_2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;

  wire   [32:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module rca_bhv_numBit32_2 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;


  rca_bhv_numBit32_2_DW01_add_0 add_1_root_add_35_2 ( .A({A[31], A}), .B({
        B[31], B}), .CI(Ci), .SUM({Co, S}) );
endmodule


module rca_bhv_numBit32_1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;

  wire   [32:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module rca_bhv_numBit32_1 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;


  rca_bhv_numBit32_1_DW01_add_0 add_1_root_add_35_2 ( .A({A[31], A}), .B({
        B[31], B}), .CI(Ci), .SUM({Co, S}) );
endmodule


module BOOTHMUL_numBit16 ( A, B, P );
  input [15:0] A;
  input [15:0] B;
  output [31:0] P;
  wire   \sum_op[7][31] , \sum_op[7][30] , \sum_op[7][29] , \sum_op[7][28] ,
         \sum_op[7][27] , \sum_op[7][26] , \sum_op[7][25] , \sum_op[7][24] ,
         \sum_op[7][23] , \sum_op[7][22] , \sum_op[7][21] , \sum_op[7][20] ,
         \sum_op[7][19] , \sum_op[7][18] , \sum_op[7][17] , \sum_op[7][16] ,
         \sum_op[7][15] , \sum_op[7][14] , \sum_op[7][13] , \sum_op[7][12] ,
         \sum_op[7][11] , \sum_op[7][10] , \sum_op[7][9] , \sum_op[7][8] ,
         \sum_op[7][7] , \sum_op[7][6] , \sum_op[7][5] , \sum_op[7][4] ,
         \sum_op[7][3] , \sum_op[7][2] , \sum_op[7][1] , \sum_op[7][0] ,
         \sum_op[6][31] , \sum_op[6][30] , \sum_op[6][29] , \sum_op[6][28] ,
         \sum_op[6][27] , \sum_op[6][26] , \sum_op[6][25] , \sum_op[6][24] ,
         \sum_op[6][23] , \sum_op[6][22] , \sum_op[6][21] , \sum_op[6][20] ,
         \sum_op[6][19] , \sum_op[6][18] , \sum_op[6][17] , \sum_op[6][16] ,
         \sum_op[6][15] , \sum_op[6][14] , \sum_op[6][13] , \sum_op[6][12] ,
         \sum_op[6][11] , \sum_op[6][10] , \sum_op[6][9] , \sum_op[6][8] ,
         \sum_op[6][7] , \sum_op[6][6] , \sum_op[6][5] , \sum_op[6][4] ,
         \sum_op[6][3] , \sum_op[6][2] , \sum_op[6][1] , \sum_op[6][0] ,
         \sum_op[5][31] , \sum_op[5][30] , \sum_op[5][29] , \sum_op[5][28] ,
         \sum_op[5][27] , \sum_op[5][26] , \sum_op[5][25] , \sum_op[5][24] ,
         \sum_op[5][23] , \sum_op[5][22] , \sum_op[5][21] , \sum_op[5][20] ,
         \sum_op[5][19] , \sum_op[5][18] , \sum_op[5][17] , \sum_op[5][16] ,
         \sum_op[5][15] , \sum_op[5][14] , \sum_op[5][13] , \sum_op[5][12] ,
         \sum_op[5][11] , \sum_op[5][10] , \sum_op[5][9] , \sum_op[5][8] ,
         \sum_op[5][7] , \sum_op[5][6] , \sum_op[5][5] , \sum_op[5][4] ,
         \sum_op[5][3] , \sum_op[5][2] , \sum_op[5][1] , \sum_op[5][0] ,
         \sum_op[4][31] , \sum_op[4][30] , \sum_op[4][29] , \sum_op[4][28] ,
         \sum_op[4][27] , \sum_op[4][26] , \sum_op[4][25] , \sum_op[4][24] ,
         \sum_op[4][23] , \sum_op[4][22] , \sum_op[4][21] , \sum_op[4][20] ,
         \sum_op[4][19] , \sum_op[4][18] , \sum_op[4][17] , \sum_op[4][16] ,
         \sum_op[4][15] , \sum_op[4][14] , \sum_op[4][13] , \sum_op[4][12] ,
         \sum_op[4][11] , \sum_op[4][10] , \sum_op[4][9] , \sum_op[4][8] ,
         \sum_op[4][7] , \sum_op[4][6] , \sum_op[4][5] , \sum_op[4][4] ,
         \sum_op[4][3] , \sum_op[4][2] , \sum_op[4][1] , \sum_op[4][0] ,
         \sum_op[3][31] , \sum_op[3][30] , \sum_op[3][29] , \sum_op[3][28] ,
         \sum_op[3][27] , \sum_op[3][26] , \sum_op[3][25] , \sum_op[3][24] ,
         \sum_op[3][23] , \sum_op[3][22] , \sum_op[3][21] , \sum_op[3][20] ,
         \sum_op[3][19] , \sum_op[3][18] , \sum_op[3][17] , \sum_op[3][16] ,
         \sum_op[3][15] , \sum_op[3][14] , \sum_op[3][13] , \sum_op[3][12] ,
         \sum_op[3][11] , \sum_op[3][10] , \sum_op[3][9] , \sum_op[3][8] ,
         \sum_op[3][7] , \sum_op[3][6] , \sum_op[3][5] , \sum_op[3][4] ,
         \sum_op[3][3] , \sum_op[3][2] , \sum_op[3][1] , \sum_op[3][0] ,
         \sum_op[2][31] , \sum_op[2][30] , \sum_op[2][29] , \sum_op[2][28] ,
         \sum_op[2][27] , \sum_op[2][26] , \sum_op[2][25] , \sum_op[2][24] ,
         \sum_op[2][23] , \sum_op[2][22] , \sum_op[2][21] , \sum_op[2][20] ,
         \sum_op[2][19] , \sum_op[2][18] , \sum_op[2][17] , \sum_op[2][16] ,
         \sum_op[2][15] , \sum_op[2][14] , \sum_op[2][13] , \sum_op[2][12] ,
         \sum_op[2][11] , \sum_op[2][10] , \sum_op[2][9] , \sum_op[2][8] ,
         \sum_op[2][7] , \sum_op[2][6] , \sum_op[2][5] , \sum_op[2][4] ,
         \sum_op[2][3] , \sum_op[2][2] , \sum_op[2][1] , \sum_op[2][0] ,
         \sum_op[1][31] , \sum_op[1][30] , \sum_op[1][29] , \sum_op[1][28] ,
         \sum_op[1][27] , \sum_op[1][26] , \sum_op[1][25] , \sum_op[1][24] ,
         \sum_op[1][23] , \sum_op[1][22] , \sum_op[1][21] , \sum_op[1][20] ,
         \sum_op[1][19] , \sum_op[1][18] , \sum_op[1][17] , \sum_op[1][16] ,
         \sum_op[1][15] , \sum_op[1][14] , \sum_op[1][13] , \sum_op[1][12] ,
         \sum_op[1][11] , \sum_op[1][10] , \sum_op[1][9] , \sum_op[1][8] ,
         \sum_op[1][7] , \sum_op[1][6] , \sum_op[1][5] , \sum_op[1][4] ,
         \sum_op[1][3] , \sum_op[1][2] , \sum_op[1][1] , \sum_op[1][0] ,
         \sum_op[0][31] , \sum_op[0][30] , \sum_op[0][29] , \sum_op[0][28] ,
         \sum_op[0][27] , \sum_op[0][26] , \sum_op[0][25] , \sum_op[0][24] ,
         \sum_op[0][23] , \sum_op[0][22] , \sum_op[0][21] , \sum_op[0][20] ,
         \sum_op[0][19] , \sum_op[0][18] , \sum_op[0][17] , \sum_op[0][16] ,
         \sum_op[0][15] , \sum_op[0][14] , \sum_op[0][13] , \sum_op[0][12] ,
         \sum_op[0][11] , \sum_op[0][10] , \sum_op[0][9] , \sum_op[0][8] ,
         \sum_op[0][7] , \sum_op[0][6] , \sum_op[0][5] , \sum_op[0][4] ,
         \sum_op[0][3] , \sum_op[0][2] , \sum_op[0][1] , \sum_op[0][0] ,
         \rca_out[5][31] , \rca_out[5][30] , \rca_out[5][29] ,
         \rca_out[5][28] , \rca_out[5][27] , \rca_out[5][26] ,
         \rca_out[5][25] , \rca_out[5][24] , \rca_out[5][23] ,
         \rca_out[5][22] , \rca_out[5][21] , \rca_out[5][20] ,
         \rca_out[5][19] , \rca_out[5][18] , \rca_out[5][17] ,
         \rca_out[5][16] , \rca_out[5][15] , \rca_out[5][14] ,
         \rca_out[5][13] , \rca_out[5][12] , \rca_out[5][11] ,
         \rca_out[5][10] , \rca_out[5][9] , \rca_out[5][8] , \rca_out[5][7] ,
         \rca_out[5][6] , \rca_out[5][5] , \rca_out[5][4] , \rca_out[5][3] ,
         \rca_out[5][2] , \rca_out[5][1] , \rca_out[5][0] , \rca_out[4][31] ,
         \rca_out[4][30] , \rca_out[4][29] , \rca_out[4][28] ,
         \rca_out[4][27] , \rca_out[4][26] , \rca_out[4][25] ,
         \rca_out[4][24] , \rca_out[4][23] , \rca_out[4][22] ,
         \rca_out[4][21] , \rca_out[4][20] , \rca_out[4][19] ,
         \rca_out[4][18] , \rca_out[4][17] , \rca_out[4][16] ,
         \rca_out[4][15] , \rca_out[4][14] , \rca_out[4][13] ,
         \rca_out[4][12] , \rca_out[4][11] , \rca_out[4][10] , \rca_out[4][9] ,
         \rca_out[4][8] , \rca_out[4][7] , \rca_out[4][6] , \rca_out[4][5] ,
         \rca_out[4][4] , \rca_out[4][3] , \rca_out[4][2] , \rca_out[4][1] ,
         \rca_out[4][0] , \rca_out[3][31] , \rca_out[3][30] , \rca_out[3][29] ,
         \rca_out[3][28] , \rca_out[3][27] , \rca_out[3][26] ,
         \rca_out[3][25] , \rca_out[3][24] , \rca_out[3][23] ,
         \rca_out[3][22] , \rca_out[3][21] , \rca_out[3][20] ,
         \rca_out[3][19] , \rca_out[3][18] , \rca_out[3][17] ,
         \rca_out[3][16] , \rca_out[3][15] , \rca_out[3][14] ,
         \rca_out[3][13] , \rca_out[3][12] , \rca_out[3][11] ,
         \rca_out[3][10] , \rca_out[3][9] , \rca_out[3][8] , \rca_out[3][7] ,
         \rca_out[3][6] , \rca_out[3][5] , \rca_out[3][4] , \rca_out[3][3] ,
         \rca_out[3][2] , \rca_out[3][1] , \rca_out[3][0] , \rca_out[2][31] ,
         \rca_out[2][30] , \rca_out[2][29] , \rca_out[2][28] ,
         \rca_out[2][27] , \rca_out[2][26] , \rca_out[2][25] ,
         \rca_out[2][24] , \rca_out[2][23] , \rca_out[2][22] ,
         \rca_out[2][21] , \rca_out[2][20] , \rca_out[2][19] ,
         \rca_out[2][18] , \rca_out[2][17] , \rca_out[2][16] ,
         \rca_out[2][15] , \rca_out[2][14] , \rca_out[2][13] ,
         \rca_out[2][12] , \rca_out[2][11] , \rca_out[2][10] , \rca_out[2][9] ,
         \rca_out[2][8] , \rca_out[2][7] , \rca_out[2][6] , \rca_out[2][5] ,
         \rca_out[2][4] , \rca_out[2][3] , \rca_out[2][2] , \rca_out[2][1] ,
         \rca_out[2][0] , \rca_out[1][31] , \rca_out[1][30] , \rca_out[1][29] ,
         \rca_out[1][28] , \rca_out[1][27] , \rca_out[1][26] ,
         \rca_out[1][25] , \rca_out[1][24] , \rca_out[1][23] ,
         \rca_out[1][22] , \rca_out[1][21] , \rca_out[1][20] ,
         \rca_out[1][19] , \rca_out[1][18] , \rca_out[1][17] ,
         \rca_out[1][16] , \rca_out[1][15] , \rca_out[1][14] ,
         \rca_out[1][13] , \rca_out[1][12] , \rca_out[1][11] ,
         \rca_out[1][10] , \rca_out[1][9] , \rca_out[1][8] , \rca_out[1][7] ,
         \rca_out[1][6] , \rca_out[1][5] , \rca_out[1][4] , \rca_out[1][3] ,
         \rca_out[1][2] , \rca_out[1][1] , \rca_out[1][0] , \rca_out[0][31] ,
         \rca_out[0][30] , \rca_out[0][29] , \rca_out[0][28] ,
         \rca_out[0][27] , \rca_out[0][26] , \rca_out[0][25] ,
         \rca_out[0][24] , \rca_out[0][23] , \rca_out[0][22] ,
         \rca_out[0][21] , \rca_out[0][20] , \rca_out[0][19] ,
         \rca_out[0][18] , \rca_out[0][17] , \rca_out[0][16] ,
         \rca_out[0][15] , \rca_out[0][14] , \rca_out[0][13] ,
         \rca_out[0][12] , \rca_out[0][11] , \rca_out[0][10] , \rca_out[0][9] ,
         \rca_out[0][8] , \rca_out[0][7] , \rca_out[0][6] , \rca_out[0][5] ,
         \rca_out[0][4] , \rca_out[0][3] , \rca_out[0][2] , \rca_out[0][1] ,
         \rca_out[0][0] , \add_65/carry[2] , \add_65/carry[3] ,
         \add_65/carry[4] , \add_65/carry[5] , \add_65/carry[6] ,
         \add_65/carry[7] , \add_65/carry[8] , \add_65/carry[9] ,
         \add_65/carry[10] , \add_65/carry[11] , \add_65/carry[12] ,
         \add_65/carry[13] , \add_65/carry[14] , \add_65/carry[15] ,
         \add_65/A[0] , \add_65/A[1] , \add_65/A[2] , \add_65/A[3] ,
         \add_65/A[4] , \add_65/A[5] , \add_65/A[6] , \add_65/A[7] ,
         \add_65/A[8] , \add_65/A[9] , \add_65/A[10] , \add_65/A[11] ,
         \add_65/A[12] , \add_65/A[13] , \add_65/A[14] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54;
  wire   [23:0] encoder_out;
  wire   [31:0] A_minus;
  wire   SYNOPSYS_UNCONNECTED__0;

  booth_encoder_numBit16 encode ( .B(B), .SEL_out({encoder_out[23:1], 
        SYNOPSYS_UNCONNECTED__0}) );
  mux5to1_numBit32_0 mux0_0 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({n48, n48, n49, n48, n48, n49, n48, n49, n48, n48, n48, 
        n49, n48, n49, n48, n49, n48, A[14:0]}), .IN3({n35, n31, n31, n36, n31, 
        n35, n31, n36, n31, n36, n32, n35, n32, n35, n33, n34, A_minus[15], n2, 
        n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, 
        A_minus[0]}), .IN4({n42, n42, n42, n42, n42, n42, n42, n42, n42, n42, 
        n42, n43, n43, n43, n43, n43, A[14:0], 1'b0}), .IN5({n41, n41, n41, 
        n41, n41, n41, n40, n40, n39, n40, n38, n39, n38, n38, n39, 
        A_minus[15], n2, n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, 
        n26, n28, A_minus[0], 1'b0}), .SEL_in({encoder_out[2:1], 1'b0}), .Z({
        \sum_op[0][31] , \sum_op[0][30] , \sum_op[0][29] , \sum_op[0][28] , 
        \sum_op[0][27] , \sum_op[0][26] , \sum_op[0][25] , \sum_op[0][24] , 
        \sum_op[0][23] , \sum_op[0][22] , \sum_op[0][21] , \sum_op[0][20] , 
        \sum_op[0][19] , \sum_op[0][18] , \sum_op[0][17] , \sum_op[0][16] , 
        \sum_op[0][15] , \sum_op[0][14] , \sum_op[0][13] , \sum_op[0][12] , 
        \sum_op[0][11] , \sum_op[0][10] , \sum_op[0][9] , \sum_op[0][8] , 
        \sum_op[0][7] , \sum_op[0][6] , \sum_op[0][5] , \sum_op[0][4] , 
        \sum_op[0][3] , \sum_op[0][2] , \sum_op[0][1] , \sum_op[0][0] }) );
  mux5to1_numBit32_7 mux_i_1 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({n52, n51, n51, n51, n51, n51, n50, n50, n50, n50, n50, 
        n49, n49, n49, n49, A[14:0], 1'b0, 1'b0}), .IN3({n31, n36, n31, n35, 
        n31, n35, n32, n36, n32, n35, n33, n34, n33, n34, A_minus[15], n2, n4, 
        n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, A_minus[0], 
        1'b0, 1'b0}), .IN4({n47, n47, n47, n47, n46, n47, n47, n47, n46, n46, 
        n46, n46, n46, n42, A[14:0], 1'b0, 1'b0, 1'b0}), .IN5({n41, n41, n40, 
        n40, n40, n40, n40, n41, n37, n39, n37, n39, n37, A_minus[15], n2, n4, 
        n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, A_minus[0], 
        1'b0, 1'b0, 1'b0}), .SEL_in(encoder_out[5:3]), .Z({\sum_op[1][31] , 
        \sum_op[1][30] , \sum_op[1][29] , \sum_op[1][28] , \sum_op[1][27] , 
        \sum_op[1][26] , \sum_op[1][25] , \sum_op[1][24] , \sum_op[1][23] , 
        \sum_op[1][22] , \sum_op[1][21] , \sum_op[1][20] , \sum_op[1][19] , 
        \sum_op[1][18] , \sum_op[1][17] , \sum_op[1][16] , \sum_op[1][15] , 
        \sum_op[1][14] , \sum_op[1][13] , \sum_op[1][12] , \sum_op[1][11] , 
        \sum_op[1][10] , \sum_op[1][9] , \sum_op[1][8] , \sum_op[1][7] , 
        \sum_op[1][6] , \sum_op[1][5] , \sum_op[1][4] , \sum_op[1][3] , 
        \sum_op[1][2] , \sum_op[1][1] , \sum_op[1][0] }) );
  mux5to1_numBit32_6 mux_i_2 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({A[15], A[15], A[15], A[15], A[15], A[15], n48, A[15], 
        A[15], n53, n53, n53, n53, A[14:0], 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({
        n31, n36, n31, n36, n32, n36, n32, n36, n33, n34, n33, n34, 
        A_minus[15], n2, n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, 
        n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({n46, n46, n46, 
        n46, n46, n47, n46, n47, n45, n47, n47, n47, A[14:0], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN5({n41, n41, n40, n40, n39, n39, n38, n38, n37, n37, 
        n38, A_minus[15], n2, n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, 
        n24, n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL_in(
        encoder_out[8:6]), .Z({\sum_op[2][31] , \sum_op[2][30] , 
        \sum_op[2][29] , \sum_op[2][28] , \sum_op[2][27] , \sum_op[2][26] , 
        \sum_op[2][25] , \sum_op[2][24] , \sum_op[2][23] , \sum_op[2][22] , 
        \sum_op[2][21] , \sum_op[2][20] , \sum_op[2][19] , \sum_op[2][18] , 
        \sum_op[2][17] , \sum_op[2][16] , \sum_op[2][15] , \sum_op[2][14] , 
        \sum_op[2][13] , \sum_op[2][12] , \sum_op[2][11] , \sum_op[2][10] , 
        \sum_op[2][9] , \sum_op[2][8] , \sum_op[2][7] , \sum_op[2][6] , 
        \sum_op[2][5] , \sum_op[2][4] , \sum_op[2][3] , \sum_op[2][2] , 
        \sum_op[2][1] , \sum_op[2][0] }) );
  mux5to1_numBit32_5 mux_i_3 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({n52, n52, n50, n53, n53, n53, n53, n53, n53, n53, n53, 
        A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({n31, n35, n32, 
        n35, n32, n36, n33, n34, n33, n34, A_minus[15], n2, n4, n6, n8, n10, 
        n12, n14, n16, n18, n20, n22, n24, n26, n28, A_minus[0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .IN4({n45, n45, n45, n45, n45, n45, n45, n45, 
        n45, n45, A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5({
        n40, n40, n39, n39, n37, n38, n38, n37, n38, A_minus[15], n2, n4, n6, 
        n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, A_minus[0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL_in(encoder_out[11:9]), .Z({
        \sum_op[3][31] , \sum_op[3][30] , \sum_op[3][29] , \sum_op[3][28] , 
        \sum_op[3][27] , \sum_op[3][26] , \sum_op[3][25] , \sum_op[3][24] , 
        \sum_op[3][23] , \sum_op[3][22] , \sum_op[3][21] , \sum_op[3][20] , 
        \sum_op[3][19] , \sum_op[3][18] , \sum_op[3][17] , \sum_op[3][16] , 
        \sum_op[3][15] , \sum_op[3][14] , \sum_op[3][13] , \sum_op[3][12] , 
        \sum_op[3][11] , \sum_op[3][10] , \sum_op[3][9] , \sum_op[3][8] , 
        \sum_op[3][7] , \sum_op[3][6] , \sum_op[3][5] , \sum_op[3][4] , 
        \sum_op[3][3] , \sum_op[3][2] , \sum_op[3][1] , \sum_op[3][0] }) );
  mux5to1_numBit32_4 mux_i_4 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({n52, n52, n52, n52, n52, n52, n52, n52, n52, A[14:0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({n31, n36, n32, 
        n36, n33, n34, n33, n34, A_minus[15], n2, n4, n6, n8, n10, n12, n14, 
        n16, n18, n20, n22, n24, n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .IN4({n44, n44, n44, n44, n44, n44, n44, n44, 
        A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5(
        {n39, n39, n38, n41, n37, n38, n39, A_minus[15], n2, n4, n6, n8, n10, 
        n12, n14, n16, n18, n20, n22, n24, n26, n28, A_minus[0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL_in(encoder_out[14:12]), .Z({\sum_op[4][31] , \sum_op[4][30] , \sum_op[4][29] , \sum_op[4][28] , 
        \sum_op[4][27] , \sum_op[4][26] , \sum_op[4][25] , \sum_op[4][24] , 
        \sum_op[4][23] , \sum_op[4][22] , \sum_op[4][21] , \sum_op[4][20] , 
        \sum_op[4][19] , \sum_op[4][18] , \sum_op[4][17] , \sum_op[4][16] , 
        \sum_op[4][15] , \sum_op[4][14] , \sum_op[4][13] , \sum_op[4][12] , 
        \sum_op[4][11] , \sum_op[4][10] , \sum_op[4][9] , \sum_op[4][8] , 
        \sum_op[4][7] , \sum_op[4][6] , \sum_op[4][5] , \sum_op[4][4] , 
        \sum_op[4][3] , \sum_op[4][2] , \sum_op[4][1] , \sum_op[4][0] }) );
  mux5to1_numBit32_3 mux_i_5 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({n51, n51, n51, n51, n51, n51, n51, A[14:0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({n32, n35, n32, 
        n35, n33, n34, A_minus[15], n2, n4, n6, n8, n10, n12, n14, n16, n18, 
        n20, n22, n24, n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({n43, n43, n44, n44, n44, n44, 
        A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN5({n40, n39, n37, n38, n37, A_minus[15], n2, n4, n6, n8, 
        n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, A_minus[0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL_in(
        encoder_out[17:15]), .Z({\sum_op[5][31] , \sum_op[5][30] , 
        \sum_op[5][29] , \sum_op[5][28] , \sum_op[5][27] , \sum_op[5][26] , 
        \sum_op[5][25] , \sum_op[5][24] , \sum_op[5][23] , \sum_op[5][22] , 
        \sum_op[5][21] , \sum_op[5][20] , \sum_op[5][19] , \sum_op[5][18] , 
        \sum_op[5][17] , \sum_op[5][16] , \sum_op[5][15] , \sum_op[5][14] , 
        \sum_op[5][13] , \sum_op[5][12] , \sum_op[5][11] , \sum_op[5][10] , 
        \sum_op[5][9] , \sum_op[5][8] , \sum_op[5][7] , \sum_op[5][6] , 
        \sum_op[5][5] , \sum_op[5][4] , \sum_op[5][3] , \sum_op[5][2] , 
        \sum_op[5][1] , \sum_op[5][0] }) );
  mux5to1_numBit32_2 mux_i_6 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({n50, n50, n50, n50, n50, A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({n32, n35, n33, 
        n34, A_minus[15], n2, n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, 
        n24, n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({n43, n43, n43, n43, A[14:0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN5({n37, n38, n37, A_minus[15], n2, n4, n6, n8, n10, n12, 
        n14, n16, n18, n20, n22, n24, n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL_in(
        encoder_out[20:18]), .Z({\sum_op[6][31] , \sum_op[6][30] , 
        \sum_op[6][29] , \sum_op[6][28] , \sum_op[6][27] , \sum_op[6][26] , 
        \sum_op[6][25] , \sum_op[6][24] , \sum_op[6][23] , \sum_op[6][22] , 
        \sum_op[6][21] , \sum_op[6][20] , \sum_op[6][19] , \sum_op[6][18] , 
        \sum_op[6][17] , \sum_op[6][16] , \sum_op[6][15] , \sum_op[6][14] , 
        \sum_op[6][13] , \sum_op[6][12] , \sum_op[6][11] , \sum_op[6][10] , 
        \sum_op[6][9] , \sum_op[6][8] , \sum_op[6][7] , \sum_op[6][6] , 
        \sum_op[6][5] , \sum_op[6][4] , \sum_op[6][3] , \sum_op[6][2] , 
        \sum_op[6][1] , \sum_op[6][0] }) );
  mux5to1_numBit32_1 mux_i_7 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({n49, n49, n50, A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({n33, n34, 
        A_minus[15], n2, n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, 
        n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({n43, n45, A[14:0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN5({n37, A_minus[15], n2, n4, n6, n8, n10, n12, n14, 
        n16, n18, n20, n22, n24, n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL_in(encoder_out[23:21]), .Z({\sum_op[7][31] , \sum_op[7][30] , 
        \sum_op[7][29] , \sum_op[7][28] , \sum_op[7][27] , \sum_op[7][26] , 
        \sum_op[7][25] , \sum_op[7][24] , \sum_op[7][23] , \sum_op[7][22] , 
        \sum_op[7][21] , \sum_op[7][20] , \sum_op[7][19] , \sum_op[7][18] , 
        \sum_op[7][17] , \sum_op[7][16] , \sum_op[7][15] , \sum_op[7][14] , 
        \sum_op[7][13] , \sum_op[7][12] , \sum_op[7][11] , \sum_op[7][10] , 
        \sum_op[7][9] , \sum_op[7][8] , \sum_op[7][7] , \sum_op[7][6] , 
        \sum_op[7][5] , \sum_op[7][4] , \sum_op[7][3] , \sum_op[7][2] , 
        \sum_op[7][1] , \sum_op[7][0] }) );
  rca_bhv_numBit32_0 rca0_0 ( .A({\sum_op[0][31] , \sum_op[0][30] , 
        \sum_op[0][29] , \sum_op[0][28] , \sum_op[0][27] , \sum_op[0][26] , 
        \sum_op[0][25] , \sum_op[0][24] , \sum_op[0][23] , \sum_op[0][22] , 
        \sum_op[0][21] , \sum_op[0][20] , \sum_op[0][19] , \sum_op[0][18] , 
        \sum_op[0][17] , \sum_op[0][16] , \sum_op[0][15] , \sum_op[0][14] , 
        \sum_op[0][13] , \sum_op[0][12] , \sum_op[0][11] , \sum_op[0][10] , 
        \sum_op[0][9] , \sum_op[0][8] , \sum_op[0][7] , \sum_op[0][6] , 
        \sum_op[0][5] , \sum_op[0][4] , \sum_op[0][3] , \sum_op[0][2] , 
        \sum_op[0][1] , \sum_op[0][0] }), .B({\sum_op[1][31] , \sum_op[1][30] , 
        \sum_op[1][29] , \sum_op[1][28] , \sum_op[1][27] , \sum_op[1][26] , 
        \sum_op[1][25] , \sum_op[1][24] , \sum_op[1][23] , \sum_op[1][22] , 
        \sum_op[1][21] , \sum_op[1][20] , \sum_op[1][19] , \sum_op[1][18] , 
        \sum_op[1][17] , \sum_op[1][16] , \sum_op[1][15] , \sum_op[1][14] , 
        \sum_op[1][13] , \sum_op[1][12] , \sum_op[1][11] , \sum_op[1][10] , 
        \sum_op[1][9] , \sum_op[1][8] , \sum_op[1][7] , \sum_op[1][6] , 
        \sum_op[1][5] , \sum_op[1][4] , \sum_op[1][3] , \sum_op[1][2] , 
        \sum_op[1][1] , \sum_op[1][0] }), .Ci(1'b0), .S({\rca_out[0][31] , 
        \rca_out[0][30] , \rca_out[0][29] , \rca_out[0][28] , \rca_out[0][27] , 
        \rca_out[0][26] , \rca_out[0][25] , \rca_out[0][24] , \rca_out[0][23] , 
        \rca_out[0][22] , \rca_out[0][21] , \rca_out[0][20] , \rca_out[0][19] , 
        \rca_out[0][18] , \rca_out[0][17] , \rca_out[0][16] , \rca_out[0][15] , 
        \rca_out[0][14] , \rca_out[0][13] , \rca_out[0][12] , \rca_out[0][11] , 
        \rca_out[0][10] , \rca_out[0][9] , \rca_out[0][8] , \rca_out[0][7] , 
        \rca_out[0][6] , \rca_out[0][5] , \rca_out[0][4] , \rca_out[0][3] , 
        \rca_out[0][2] , \rca_out[0][1] , \rca_out[0][0] }) );
  rca_bhv_numBit32_6 rca_i_1 ( .A({\rca_out[0][31] , \rca_out[0][30] , 
        \rca_out[0][29] , \rca_out[0][28] , \rca_out[0][27] , \rca_out[0][26] , 
        \rca_out[0][25] , \rca_out[0][24] , \rca_out[0][23] , \rca_out[0][22] , 
        \rca_out[0][21] , \rca_out[0][20] , \rca_out[0][19] , \rca_out[0][18] , 
        \rca_out[0][17] , \rca_out[0][16] , \rca_out[0][15] , \rca_out[0][14] , 
        \rca_out[0][13] , \rca_out[0][12] , \rca_out[0][11] , \rca_out[0][10] , 
        \rca_out[0][9] , \rca_out[0][8] , \rca_out[0][7] , \rca_out[0][6] , 
        \rca_out[0][5] , \rca_out[0][4] , \rca_out[0][3] , \rca_out[0][2] , 
        \rca_out[0][1] , \rca_out[0][0] }), .B({\sum_op[2][31] , 
        \sum_op[2][30] , \sum_op[2][29] , \sum_op[2][28] , \sum_op[2][27] , 
        \sum_op[2][26] , \sum_op[2][25] , \sum_op[2][24] , \sum_op[2][23] , 
        \sum_op[2][22] , \sum_op[2][21] , \sum_op[2][20] , \sum_op[2][19] , 
        \sum_op[2][18] , \sum_op[2][17] , \sum_op[2][16] , \sum_op[2][15] , 
        \sum_op[2][14] , \sum_op[2][13] , \sum_op[2][12] , \sum_op[2][11] , 
        \sum_op[2][10] , \sum_op[2][9] , \sum_op[2][8] , \sum_op[2][7] , 
        \sum_op[2][6] , \sum_op[2][5] , \sum_op[2][4] , \sum_op[2][3] , 
        \sum_op[2][2] , \sum_op[2][1] , \sum_op[2][0] }), .Ci(1'b0), .S({
        \rca_out[1][31] , \rca_out[1][30] , \rca_out[1][29] , \rca_out[1][28] , 
        \rca_out[1][27] , \rca_out[1][26] , \rca_out[1][25] , \rca_out[1][24] , 
        \rca_out[1][23] , \rca_out[1][22] , \rca_out[1][21] , \rca_out[1][20] , 
        \rca_out[1][19] , \rca_out[1][18] , \rca_out[1][17] , \rca_out[1][16] , 
        \rca_out[1][15] , \rca_out[1][14] , \rca_out[1][13] , \rca_out[1][12] , 
        \rca_out[1][11] , \rca_out[1][10] , \rca_out[1][9] , \rca_out[1][8] , 
        \rca_out[1][7] , \rca_out[1][6] , \rca_out[1][5] , \rca_out[1][4] , 
        \rca_out[1][3] , \rca_out[1][2] , \rca_out[1][1] , \rca_out[1][0] })
         );
  rca_bhv_numBit32_5 rca_i_2 ( .A({\rca_out[1][31] , \rca_out[1][30] , 
        \rca_out[1][29] , \rca_out[1][28] , \rca_out[1][27] , \rca_out[1][26] , 
        \rca_out[1][25] , \rca_out[1][24] , \rca_out[1][23] , \rca_out[1][22] , 
        \rca_out[1][21] , \rca_out[1][20] , \rca_out[1][19] , \rca_out[1][18] , 
        \rca_out[1][17] , \rca_out[1][16] , \rca_out[1][15] , \rca_out[1][14] , 
        \rca_out[1][13] , \rca_out[1][12] , \rca_out[1][11] , \rca_out[1][10] , 
        \rca_out[1][9] , \rca_out[1][8] , \rca_out[1][7] , \rca_out[1][6] , 
        \rca_out[1][5] , \rca_out[1][4] , \rca_out[1][3] , \rca_out[1][2] , 
        \rca_out[1][1] , \rca_out[1][0] }), .B({\sum_op[3][31] , 
        \sum_op[3][30] , \sum_op[3][29] , \sum_op[3][28] , \sum_op[3][27] , 
        \sum_op[3][26] , \sum_op[3][25] , \sum_op[3][24] , \sum_op[3][23] , 
        \sum_op[3][22] , \sum_op[3][21] , \sum_op[3][20] , \sum_op[3][19] , 
        \sum_op[3][18] , \sum_op[3][17] , \sum_op[3][16] , \sum_op[3][15] , 
        \sum_op[3][14] , \sum_op[3][13] , \sum_op[3][12] , \sum_op[3][11] , 
        \sum_op[3][10] , \sum_op[3][9] , \sum_op[3][8] , \sum_op[3][7] , 
        \sum_op[3][6] , \sum_op[3][5] , \sum_op[3][4] , \sum_op[3][3] , 
        \sum_op[3][2] , \sum_op[3][1] , \sum_op[3][0] }), .Ci(1'b0), .S({
        \rca_out[2][31] , \rca_out[2][30] , \rca_out[2][29] , \rca_out[2][28] , 
        \rca_out[2][27] , \rca_out[2][26] , \rca_out[2][25] , \rca_out[2][24] , 
        \rca_out[2][23] , \rca_out[2][22] , \rca_out[2][21] , \rca_out[2][20] , 
        \rca_out[2][19] , \rca_out[2][18] , \rca_out[2][17] , \rca_out[2][16] , 
        \rca_out[2][15] , \rca_out[2][14] , \rca_out[2][13] , \rca_out[2][12] , 
        \rca_out[2][11] , \rca_out[2][10] , \rca_out[2][9] , \rca_out[2][8] , 
        \rca_out[2][7] , \rca_out[2][6] , \rca_out[2][5] , \rca_out[2][4] , 
        \rca_out[2][3] , \rca_out[2][2] , \rca_out[2][1] , \rca_out[2][0] })
         );
  rca_bhv_numBit32_4 rca_i_3 ( .A({\rca_out[2][31] , \rca_out[2][30] , 
        \rca_out[2][29] , \rca_out[2][28] , \rca_out[2][27] , \rca_out[2][26] , 
        \rca_out[2][25] , \rca_out[2][24] , \rca_out[2][23] , \rca_out[2][22] , 
        \rca_out[2][21] , \rca_out[2][20] , \rca_out[2][19] , \rca_out[2][18] , 
        \rca_out[2][17] , \rca_out[2][16] , \rca_out[2][15] , \rca_out[2][14] , 
        \rca_out[2][13] , \rca_out[2][12] , \rca_out[2][11] , \rca_out[2][10] , 
        \rca_out[2][9] , \rca_out[2][8] , \rca_out[2][7] , \rca_out[2][6] , 
        \rca_out[2][5] , \rca_out[2][4] , \rca_out[2][3] , \rca_out[2][2] , 
        \rca_out[2][1] , \rca_out[2][0] }), .B({\sum_op[4][31] , 
        \sum_op[4][30] , \sum_op[4][29] , \sum_op[4][28] , \sum_op[4][27] , 
        \sum_op[4][26] , \sum_op[4][25] , \sum_op[4][24] , \sum_op[4][23] , 
        \sum_op[4][22] , \sum_op[4][21] , \sum_op[4][20] , \sum_op[4][19] , 
        \sum_op[4][18] , \sum_op[4][17] , \sum_op[4][16] , \sum_op[4][15] , 
        \sum_op[4][14] , \sum_op[4][13] , \sum_op[4][12] , \sum_op[4][11] , 
        \sum_op[4][10] , \sum_op[4][9] , \sum_op[4][8] , \sum_op[4][7] , 
        \sum_op[4][6] , \sum_op[4][5] , \sum_op[4][4] , \sum_op[4][3] , 
        \sum_op[4][2] , \sum_op[4][1] , \sum_op[4][0] }), .Ci(1'b0), .S({
        \rca_out[3][31] , \rca_out[3][30] , \rca_out[3][29] , \rca_out[3][28] , 
        \rca_out[3][27] , \rca_out[3][26] , \rca_out[3][25] , \rca_out[3][24] , 
        \rca_out[3][23] , \rca_out[3][22] , \rca_out[3][21] , \rca_out[3][20] , 
        \rca_out[3][19] , \rca_out[3][18] , \rca_out[3][17] , \rca_out[3][16] , 
        \rca_out[3][15] , \rca_out[3][14] , \rca_out[3][13] , \rca_out[3][12] , 
        \rca_out[3][11] , \rca_out[3][10] , \rca_out[3][9] , \rca_out[3][8] , 
        \rca_out[3][7] , \rca_out[3][6] , \rca_out[3][5] , \rca_out[3][4] , 
        \rca_out[3][3] , \rca_out[3][2] , \rca_out[3][1] , \rca_out[3][0] })
         );
  rca_bhv_numBit32_3 rca_i_4 ( .A({\rca_out[3][31] , \rca_out[3][30] , 
        \rca_out[3][29] , \rca_out[3][28] , \rca_out[3][27] , \rca_out[3][26] , 
        \rca_out[3][25] , \rca_out[3][24] , \rca_out[3][23] , \rca_out[3][22] , 
        \rca_out[3][21] , \rca_out[3][20] , \rca_out[3][19] , \rca_out[3][18] , 
        \rca_out[3][17] , \rca_out[3][16] , \rca_out[3][15] , \rca_out[3][14] , 
        \rca_out[3][13] , \rca_out[3][12] , \rca_out[3][11] , \rca_out[3][10] , 
        \rca_out[3][9] , \rca_out[3][8] , \rca_out[3][7] , \rca_out[3][6] , 
        \rca_out[3][5] , \rca_out[3][4] , \rca_out[3][3] , \rca_out[3][2] , 
        \rca_out[3][1] , \rca_out[3][0] }), .B({\sum_op[5][31] , 
        \sum_op[5][30] , \sum_op[5][29] , \sum_op[5][28] , \sum_op[5][27] , 
        \sum_op[5][26] , \sum_op[5][25] , \sum_op[5][24] , \sum_op[5][23] , 
        \sum_op[5][22] , \sum_op[5][21] , \sum_op[5][20] , \sum_op[5][19] , 
        \sum_op[5][18] , \sum_op[5][17] , \sum_op[5][16] , \sum_op[5][15] , 
        \sum_op[5][14] , \sum_op[5][13] , \sum_op[5][12] , \sum_op[5][11] , 
        \sum_op[5][10] , \sum_op[5][9] , \sum_op[5][8] , \sum_op[5][7] , 
        \sum_op[5][6] , \sum_op[5][5] , \sum_op[5][4] , \sum_op[5][3] , 
        \sum_op[5][2] , \sum_op[5][1] , \sum_op[5][0] }), .Ci(1'b0), .S({
        \rca_out[4][31] , \rca_out[4][30] , \rca_out[4][29] , \rca_out[4][28] , 
        \rca_out[4][27] , \rca_out[4][26] , \rca_out[4][25] , \rca_out[4][24] , 
        \rca_out[4][23] , \rca_out[4][22] , \rca_out[4][21] , \rca_out[4][20] , 
        \rca_out[4][19] , \rca_out[4][18] , \rca_out[4][17] , \rca_out[4][16] , 
        \rca_out[4][15] , \rca_out[4][14] , \rca_out[4][13] , \rca_out[4][12] , 
        \rca_out[4][11] , \rca_out[4][10] , \rca_out[4][9] , \rca_out[4][8] , 
        \rca_out[4][7] , \rca_out[4][6] , \rca_out[4][5] , \rca_out[4][4] , 
        \rca_out[4][3] , \rca_out[4][2] , \rca_out[4][1] , \rca_out[4][0] })
         );
  rca_bhv_numBit32_2 rca_i_5 ( .A({\rca_out[4][31] , \rca_out[4][30] , 
        \rca_out[4][29] , \rca_out[4][28] , \rca_out[4][27] , \rca_out[4][26] , 
        \rca_out[4][25] , \rca_out[4][24] , \rca_out[4][23] , \rca_out[4][22] , 
        \rca_out[4][21] , \rca_out[4][20] , \rca_out[4][19] , \rca_out[4][18] , 
        \rca_out[4][17] , \rca_out[4][16] , \rca_out[4][15] , \rca_out[4][14] , 
        \rca_out[4][13] , \rca_out[4][12] , \rca_out[4][11] , \rca_out[4][10] , 
        \rca_out[4][9] , \rca_out[4][8] , \rca_out[4][7] , \rca_out[4][6] , 
        \rca_out[4][5] , \rca_out[4][4] , \rca_out[4][3] , \rca_out[4][2] , 
        \rca_out[4][1] , \rca_out[4][0] }), .B({\sum_op[6][31] , 
        \sum_op[6][30] , \sum_op[6][29] , \sum_op[6][28] , \sum_op[6][27] , 
        \sum_op[6][26] , \sum_op[6][25] , \sum_op[6][24] , \sum_op[6][23] , 
        \sum_op[6][22] , \sum_op[6][21] , \sum_op[6][20] , \sum_op[6][19] , 
        \sum_op[6][18] , \sum_op[6][17] , \sum_op[6][16] , \sum_op[6][15] , 
        \sum_op[6][14] , \sum_op[6][13] , \sum_op[6][12] , \sum_op[6][11] , 
        \sum_op[6][10] , \sum_op[6][9] , \sum_op[6][8] , \sum_op[6][7] , 
        \sum_op[6][6] , \sum_op[6][5] , \sum_op[6][4] , \sum_op[6][3] , 
        \sum_op[6][2] , \sum_op[6][1] , \sum_op[6][0] }), .Ci(1'b0), .S({
        \rca_out[5][31] , \rca_out[5][30] , \rca_out[5][29] , \rca_out[5][28] , 
        \rca_out[5][27] , \rca_out[5][26] , \rca_out[5][25] , \rca_out[5][24] , 
        \rca_out[5][23] , \rca_out[5][22] , \rca_out[5][21] , \rca_out[5][20] , 
        \rca_out[5][19] , \rca_out[5][18] , \rca_out[5][17] , \rca_out[5][16] , 
        \rca_out[5][15] , \rca_out[5][14] , \rca_out[5][13] , \rca_out[5][12] , 
        \rca_out[5][11] , \rca_out[5][10] , \rca_out[5][9] , \rca_out[5][8] , 
        \rca_out[5][7] , \rca_out[5][6] , \rca_out[5][5] , \rca_out[5][4] , 
        \rca_out[5][3] , \rca_out[5][2] , \rca_out[5][1] , \rca_out[5][0] })
         );
  rca_bhv_numBit32_1 rca_i_6 ( .A({\rca_out[5][31] , \rca_out[5][30] , 
        \rca_out[5][29] , \rca_out[5][28] , \rca_out[5][27] , \rca_out[5][26] , 
        \rca_out[5][25] , \rca_out[5][24] , \rca_out[5][23] , \rca_out[5][22] , 
        \rca_out[5][21] , \rca_out[5][20] , \rca_out[5][19] , \rca_out[5][18] , 
        \rca_out[5][17] , \rca_out[5][16] , \rca_out[5][15] , \rca_out[5][14] , 
        \rca_out[5][13] , \rca_out[5][12] , \rca_out[5][11] , \rca_out[5][10] , 
        \rca_out[5][9] , \rca_out[5][8] , \rca_out[5][7] , \rca_out[5][6] , 
        \rca_out[5][5] , \rca_out[5][4] , \rca_out[5][3] , \rca_out[5][2] , 
        \rca_out[5][1] , \rca_out[5][0] }), .B({\sum_op[7][31] , 
        \sum_op[7][30] , \sum_op[7][29] , \sum_op[7][28] , \sum_op[7][27] , 
        \sum_op[7][26] , \sum_op[7][25] , \sum_op[7][24] , \sum_op[7][23] , 
        \sum_op[7][22] , \sum_op[7][21] , \sum_op[7][20] , \sum_op[7][19] , 
        \sum_op[7][18] , \sum_op[7][17] , \sum_op[7][16] , \sum_op[7][15] , 
        \sum_op[7][14] , \sum_op[7][13] , \sum_op[7][12] , \sum_op[7][11] , 
        \sum_op[7][10] , \sum_op[7][9] , \sum_op[7][8] , \sum_op[7][7] , 
        \sum_op[7][6] , \sum_op[7][5] , \sum_op[7][4] , \sum_op[7][3] , 
        \sum_op[7][2] , \sum_op[7][1] , \sum_op[7][0] }), .Ci(1'b0), .S(P) );
  HA_X1 \add_65/U1_1_1  ( .A(\add_65/A[1] ), .B(\add_65/A[0] ), .CO(
        \add_65/carry[2] ), .S(A_minus[1]) );
  HA_X1 \add_65/U1_1_2  ( .A(\add_65/A[2] ), .B(\add_65/carry[2] ), .CO(
        \add_65/carry[3] ), .S(A_minus[2]) );
  HA_X1 \add_65/U1_1_3  ( .A(\add_65/A[3] ), .B(\add_65/carry[3] ), .CO(
        \add_65/carry[4] ), .S(A_minus[3]) );
  HA_X1 \add_65/U1_1_4  ( .A(\add_65/A[4] ), .B(\add_65/carry[4] ), .CO(
        \add_65/carry[5] ), .S(A_minus[4]) );
  HA_X1 \add_65/U1_1_5  ( .A(\add_65/A[5] ), .B(\add_65/carry[5] ), .CO(
        \add_65/carry[6] ), .S(A_minus[5]) );
  HA_X1 \add_65/U1_1_6  ( .A(\add_65/A[6] ), .B(\add_65/carry[6] ), .CO(
        \add_65/carry[7] ), .S(A_minus[6]) );
  HA_X1 \add_65/U1_1_7  ( .A(\add_65/A[7] ), .B(\add_65/carry[7] ), .CO(
        \add_65/carry[8] ), .S(A_minus[7]) );
  HA_X1 \add_65/U1_1_8  ( .A(\add_65/A[8] ), .B(\add_65/carry[8] ), .CO(
        \add_65/carry[9] ), .S(A_minus[8]) );
  HA_X1 \add_65/U1_1_9  ( .A(\add_65/A[9] ), .B(\add_65/carry[9] ), .CO(
        \add_65/carry[10] ), .S(A_minus[9]) );
  HA_X1 \add_65/U1_1_10  ( .A(\add_65/A[10] ), .B(\add_65/carry[10] ), .CO(
        \add_65/carry[11] ), .S(A_minus[10]) );
  HA_X1 \add_65/U1_1_11  ( .A(\add_65/A[11] ), .B(\add_65/carry[11] ), .CO(
        \add_65/carry[12] ), .S(A_minus[11]) );
  HA_X1 \add_65/U1_1_12  ( .A(\add_65/A[12] ), .B(\add_65/carry[12] ), .CO(
        \add_65/carry[13] ), .S(A_minus[12]) );
  HA_X1 \add_65/U1_1_13  ( .A(\add_65/A[13] ), .B(\add_65/carry[13] ), .CO(
        \add_65/carry[14] ), .S(A_minus[13]) );
  HA_X1 \add_65/U1_1_14  ( .A(\add_65/A[14] ), .B(\add_65/carry[14] ), .CO(
        \add_65/carry[15] ), .S(A_minus[14]) );
  INV_X1 U3 ( .A(A_minus[14]), .ZN(n1) );
  INV_X1 U4 ( .A(n1), .ZN(n2) );
  INV_X1 U5 ( .A(A_minus[13]), .ZN(n3) );
  INV_X1 U6 ( .A(n3), .ZN(n4) );
  INV_X1 U7 ( .A(A_minus[12]), .ZN(n5) );
  INV_X1 U8 ( .A(n5), .ZN(n6) );
  INV_X1 U9 ( .A(A_minus[11]), .ZN(n7) );
  INV_X1 U10 ( .A(n7), .ZN(n8) );
  INV_X1 U11 ( .A(A_minus[10]), .ZN(n9) );
  INV_X1 U12 ( .A(n9), .ZN(n10) );
  INV_X1 U13 ( .A(A_minus[9]), .ZN(n11) );
  INV_X1 U14 ( .A(n11), .ZN(n12) );
  INV_X1 U15 ( .A(A_minus[8]), .ZN(n13) );
  INV_X1 U16 ( .A(n13), .ZN(n14) );
  INV_X1 U17 ( .A(A_minus[7]), .ZN(n15) );
  INV_X1 U18 ( .A(n15), .ZN(n16) );
  INV_X1 U19 ( .A(A_minus[6]), .ZN(n17) );
  INV_X1 U20 ( .A(n17), .ZN(n18) );
  INV_X1 U21 ( .A(A_minus[5]), .ZN(n19) );
  INV_X1 U22 ( .A(n19), .ZN(n20) );
  INV_X1 U23 ( .A(A_minus[4]), .ZN(n21) );
  INV_X1 U24 ( .A(n21), .ZN(n22) );
  INV_X1 U25 ( .A(A_minus[3]), .ZN(n23) );
  INV_X1 U26 ( .A(n23), .ZN(n24) );
  INV_X1 U27 ( .A(A_minus[2]), .ZN(n25) );
  INV_X1 U28 ( .A(n25), .ZN(n26) );
  INV_X1 U29 ( .A(A_minus[1]), .ZN(n27) );
  INV_X1 U30 ( .A(n27), .ZN(n28) );
  BUF_X1 U31 ( .A(n30), .Z(n40) );
  BUF_X1 U32 ( .A(n30), .Z(n39) );
  BUF_X1 U33 ( .A(n30), .Z(n37) );
  BUF_X1 U34 ( .A(n30), .Z(n38) );
  BUF_X1 U35 ( .A(n29), .Z(n36) );
  BUF_X1 U36 ( .A(n29), .Z(n31) );
  BUF_X1 U37 ( .A(n29), .Z(n33) );
  BUF_X1 U38 ( .A(n29), .Z(n35) );
  BUF_X1 U39 ( .A(n29), .Z(n32) );
  BUF_X1 U40 ( .A(n29), .Z(n34) );
  BUF_X1 U41 ( .A(n30), .Z(n41) );
  BUF_X1 U42 ( .A(A_minus[31]), .Z(n29) );
  BUF_X1 U43 ( .A(A_minus[31]), .Z(n30) );
  INV_X1 U44 ( .A(n54), .ZN(n42) );
  INV_X1 U45 ( .A(n54), .ZN(n43) );
  INV_X1 U46 ( .A(n54), .ZN(n47) );
  INV_X1 U47 ( .A(n54), .ZN(n46) );
  INV_X1 U48 ( .A(n54), .ZN(n44) );
  INV_X1 U49 ( .A(n54), .ZN(n45) );
  INV_X1 U50 ( .A(n54), .ZN(n48) );
  INV_X1 U51 ( .A(n54), .ZN(n53) );
  INV_X1 U52 ( .A(n54), .ZN(n52) );
  INV_X1 U53 ( .A(n54), .ZN(n51) );
  INV_X1 U54 ( .A(n54), .ZN(n50) );
  INV_X1 U55 ( .A(n54), .ZN(n49) );
  INV_X1 U56 ( .A(\add_65/A[0] ), .ZN(A_minus[0]) );
  INV_X1 U57 ( .A(A[0]), .ZN(\add_65/A[0] ) );
  INV_X1 U58 ( .A(A[14]), .ZN(\add_65/A[14] ) );
  INV_X1 U59 ( .A(A[1]), .ZN(\add_65/A[1] ) );
  INV_X1 U60 ( .A(A[2]), .ZN(\add_65/A[2] ) );
  INV_X1 U61 ( .A(A[3]), .ZN(\add_65/A[3] ) );
  INV_X1 U62 ( .A(A[4]), .ZN(\add_65/A[4] ) );
  INV_X1 U63 ( .A(A[5]), .ZN(\add_65/A[5] ) );
  INV_X1 U64 ( .A(A[6]), .ZN(\add_65/A[6] ) );
  INV_X1 U65 ( .A(A[7]), .ZN(\add_65/A[7] ) );
  INV_X1 U66 ( .A(A[8]), .ZN(\add_65/A[8] ) );
  INV_X1 U67 ( .A(A[9]), .ZN(\add_65/A[9] ) );
  INV_X1 U68 ( .A(A[10]), .ZN(\add_65/A[10] ) );
  INV_X1 U69 ( .A(A[11]), .ZN(\add_65/A[11] ) );
  INV_X1 U70 ( .A(A[12]), .ZN(\add_65/A[12] ) );
  INV_X1 U71 ( .A(A[13]), .ZN(\add_65/A[13] ) );
  XOR2_X2 U72 ( .A(\add_65/carry[15] ), .B(n54), .Z(A_minus[15]) );
  INV_X1 U73 ( .A(A[15]), .ZN(n54) );
  NOR2_X1 U74 ( .A1(\add_65/carry[15] ), .A2(A[15]), .ZN(A_minus[31]) );
endmodule


module mux41_NBIT32_1 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149;

  BUF_X1 U1 ( .A(n145), .Z(n72) );
  BUF_X1 U2 ( .A(n145), .Z(n73) );
  BUF_X1 U3 ( .A(n146), .Z(n75) );
  BUF_X1 U4 ( .A(n146), .Z(n76) );
  BUF_X1 U5 ( .A(n145), .Z(n74) );
  BUF_X1 U6 ( .A(n146), .Z(n77) );
  NOR2_X1 U7 ( .A1(n81), .A2(S[1]), .ZN(n145) );
  BUF_X1 U8 ( .A(n147), .Z(n78) );
  BUF_X1 U9 ( .A(n147), .Z(n79) );
  BUF_X1 U10 ( .A(n144), .Z(n1) );
  BUF_X1 U11 ( .A(n144), .Z(n70) );
  BUF_X1 U12 ( .A(n147), .Z(n80) );
  BUF_X1 U13 ( .A(n144), .Z(n71) );
  AND2_X1 U14 ( .A1(S[1]), .A2(n81), .ZN(n146) );
  NOR2_X1 U15 ( .A1(S[0]), .A2(S[1]), .ZN(n144) );
  AOI22_X1 U16 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n82) );
  AOI22_X1 U17 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n137) );
  AOI22_X1 U18 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n139) );
  AOI22_X1 U19 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n141) );
  AOI22_X1 U20 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n149) );
  AOI22_X1 U21 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n131) );
  AOI22_X1 U22 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n85) );
  AOI22_X1 U23 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n87) );
  AOI22_X1 U24 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n91) );
  AOI22_X1 U25 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n93) );
  AOI22_X1 U26 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n95) );
  AOI22_X1 U27 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n99) );
  AOI22_X1 U28 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n101) );
  AOI22_X1 U29 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n103) );
  AOI22_X1 U30 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n109) );
  AOI22_X1 U31 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n111) );
  AOI22_X1 U32 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n113) );
  AOI22_X1 U33 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n117) );
  AOI22_X1 U34 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n119) );
  AOI22_X1 U35 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n121) );
  AOI22_X1 U36 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n125) );
  AOI22_X1 U37 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n129) );
  AND2_X1 U38 ( .A1(S[1]), .A2(S[0]), .ZN(n147) );
  INV_X1 U39 ( .A(S[0]), .ZN(n81) );
  AOI22_X1 U40 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n133) );
  AOI22_X1 U41 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n135) );
  AOI22_X1 U42 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n143) );
  AOI22_X1 U43 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n105) );
  AOI22_X1 U44 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n127) );
  AOI22_X1 U45 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n89) );
  AOI22_X1 U46 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n97) );
  AOI22_X1 U47 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n107) );
  AOI22_X1 U48 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n115) );
  AOI22_X1 U49 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n123) );
  NAND2_X1 U50 ( .A1(n131), .A2(n130), .ZN(Z[31]) );
  NAND2_X1 U51 ( .A1(n83), .A2(n82), .ZN(Z[0]) );
  AOI22_X1 U52 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n83) );
  AOI22_X1 U53 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n130) );
  NAND2_X1 U54 ( .A1(n133), .A2(n132), .ZN(Z[3]) );
  AOI22_X1 U55 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n132) );
  NAND2_X1 U56 ( .A1(n135), .A2(n134), .ZN(Z[4]) );
  AOI22_X1 U57 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n134) );
  NAND2_X1 U58 ( .A1(n137), .A2(n136), .ZN(Z[5]) );
  AOI22_X1 U59 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n136) );
  NAND2_X1 U60 ( .A1(n139), .A2(n138), .ZN(Z[6]) );
  AOI22_X1 U61 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n138) );
  NAND2_X1 U62 ( .A1(n141), .A2(n140), .ZN(Z[7]) );
  AOI22_X1 U63 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n140) );
  NAND2_X1 U64 ( .A1(n143), .A2(n142), .ZN(Z[8]) );
  AOI22_X1 U65 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n142) );
  NAND2_X1 U66 ( .A1(n149), .A2(n148), .ZN(Z[9]) );
  AOI22_X1 U67 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n148) );
  NAND2_X1 U68 ( .A1(n95), .A2(n94), .ZN(Z[15]) );
  AOI22_X1 U69 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n94) );
  NAND2_X1 U70 ( .A1(n97), .A2(n96), .ZN(Z[16]) );
  AOI22_X1 U71 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n96) );
  NAND2_X1 U72 ( .A1(n99), .A2(n98), .ZN(Z[17]) );
  AOI22_X1 U73 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n98) );
  NAND2_X1 U74 ( .A1(n101), .A2(n100), .ZN(Z[18]) );
  AOI22_X1 U75 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n100) );
  NAND2_X1 U76 ( .A1(n103), .A2(n102), .ZN(Z[19]) );
  AOI22_X1 U77 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n102) );
  NAND2_X1 U78 ( .A1(n107), .A2(n106), .ZN(Z[20]) );
  AOI22_X1 U79 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n106) );
  NAND2_X1 U80 ( .A1(n109), .A2(n108), .ZN(Z[21]) );
  AOI22_X1 U81 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n108) );
  NAND2_X1 U82 ( .A1(n111), .A2(n110), .ZN(Z[22]) );
  AOI22_X1 U83 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n110) );
  NAND2_X1 U84 ( .A1(n113), .A2(n112), .ZN(Z[23]) );
  AOI22_X1 U85 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n112) );
  NAND2_X1 U86 ( .A1(n115), .A2(n114), .ZN(Z[24]) );
  AOI22_X1 U87 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n114) );
  NAND2_X1 U88 ( .A1(n117), .A2(n116), .ZN(Z[25]) );
  AOI22_X1 U89 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n116) );
  NAND2_X1 U90 ( .A1(n119), .A2(n118), .ZN(Z[26]) );
  AOI22_X1 U91 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n118) );
  NAND2_X1 U92 ( .A1(n121), .A2(n120), .ZN(Z[27]) );
  AOI22_X1 U93 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n120) );
  NAND2_X1 U94 ( .A1(n123), .A2(n122), .ZN(Z[28]) );
  AOI22_X1 U95 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n122) );
  NAND2_X1 U96 ( .A1(n125), .A2(n124), .ZN(Z[29]) );
  AOI22_X1 U97 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n124) );
  NAND2_X1 U98 ( .A1(n129), .A2(n128), .ZN(Z[30]) );
  AOI22_X1 U99 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n128) );
  NAND2_X1 U100 ( .A1(n93), .A2(n92), .ZN(Z[14]) );
  AOI22_X1 U101 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n92) );
  NAND2_X1 U102 ( .A1(n105), .A2(n104), .ZN(Z[1]) );
  AOI22_X1 U103 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n104) );
  NAND2_X1 U104 ( .A1(n127), .A2(n126), .ZN(Z[2]) );
  AOI22_X1 U105 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n126) );
  NAND2_X1 U106 ( .A1(n85), .A2(n84), .ZN(Z[10]) );
  AOI22_X1 U107 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n84) );
  NAND2_X1 U108 ( .A1(n87), .A2(n86), .ZN(Z[11]) );
  AOI22_X1 U109 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n86) );
  NAND2_X1 U110 ( .A1(n89), .A2(n88), .ZN(Z[12]) );
  AOI22_X1 U111 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n88) );
  NAND2_X1 U112 ( .A1(n91), .A2(n90), .ZN(Z[13]) );
  AOI22_X1 U113 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n90) );
endmodule


module mux21_NBIT32_2 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n11) );
  BUF_X1 U6 ( .A(n2), .Z(n9) );
  BUF_X1 U7 ( .A(n1), .Z(n8) );
  BUF_X1 U8 ( .A(n2), .Z(n10) );
  BUF_X1 U9 ( .A(n1), .Z(n7) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  INV_X1 U12 ( .A(n103), .ZN(Z[31]) );
  AOI22_X1 U13 ( .A1(A[31]), .A2(n4), .B1(B[31]), .B2(n7), .ZN(n103) );
  BUF_X1 U14 ( .A(S), .Z(n3) );
  BUF_X1 U15 ( .A(S), .Z(n2) );
  BUF_X1 U16 ( .A(S), .Z(n1) );
  INV_X1 U17 ( .A(n79), .ZN(Z[0]) );
  AOI22_X1 U18 ( .A1(A[0]), .A2(n4), .B1(B[0]), .B2(n13), .ZN(n79) );
  INV_X1 U19 ( .A(n104), .ZN(Z[3]) );
  AOI22_X1 U20 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n7), .ZN(n104) );
  INV_X1 U21 ( .A(n105), .ZN(Z[4]) );
  AOI22_X1 U22 ( .A1(A[4]), .A2(n4), .B1(B[4]), .B2(n7), .ZN(n105) );
  INV_X1 U23 ( .A(n106), .ZN(Z[5]) );
  AOI22_X1 U24 ( .A1(A[5]), .A2(n5), .B1(B[5]), .B2(n6), .ZN(n106) );
  INV_X1 U25 ( .A(n107), .ZN(Z[6]) );
  AOI22_X1 U26 ( .A1(A[6]), .A2(n4), .B1(B[6]), .B2(n6), .ZN(n107) );
  INV_X1 U27 ( .A(n108), .ZN(Z[7]) );
  AOI22_X1 U28 ( .A1(A[7]), .A2(n5), .B1(B[7]), .B2(n6), .ZN(n108) );
  INV_X1 U29 ( .A(n109), .ZN(Z[8]) );
  AOI22_X1 U30 ( .A1(A[8]), .A2(n4), .B1(B[8]), .B2(n6), .ZN(n109) );
  INV_X1 U31 ( .A(n110), .ZN(Z[9]) );
  AOI22_X1 U32 ( .A1(A[9]), .A2(n5), .B1(n13), .B2(B[9]), .ZN(n110) );
  INV_X1 U33 ( .A(n85), .ZN(Z[15]) );
  AOI22_X1 U34 ( .A1(A[15]), .A2(n4), .B1(B[15]), .B2(n12), .ZN(n85) );
  INV_X1 U35 ( .A(n86), .ZN(Z[16]) );
  AOI22_X1 U36 ( .A1(A[16]), .A2(n4), .B1(B[16]), .B2(n11), .ZN(n86) );
  INV_X1 U37 ( .A(n87), .ZN(Z[17]) );
  AOI22_X1 U38 ( .A1(A[17]), .A2(n4), .B1(B[17]), .B2(n11), .ZN(n87) );
  INV_X1 U39 ( .A(n88), .ZN(Z[18]) );
  AOI22_X1 U40 ( .A1(A[18]), .A2(n4), .B1(B[18]), .B2(n11), .ZN(n88) );
  INV_X1 U41 ( .A(n89), .ZN(Z[19]) );
  AOI22_X1 U42 ( .A1(A[19]), .A2(n4), .B1(B[19]), .B2(n11), .ZN(n89) );
  INV_X1 U43 ( .A(n91), .ZN(Z[20]) );
  AOI22_X1 U44 ( .A1(A[20]), .A2(n5), .B1(B[20]), .B2(n10), .ZN(n91) );
  INV_X1 U45 ( .A(n92), .ZN(Z[21]) );
  AOI22_X1 U46 ( .A1(A[21]), .A2(n5), .B1(B[21]), .B2(n10), .ZN(n92) );
  INV_X1 U47 ( .A(n93), .ZN(Z[22]) );
  AOI22_X1 U48 ( .A1(A[22]), .A2(n5), .B1(B[22]), .B2(n9), .ZN(n93) );
  INV_X1 U49 ( .A(n94), .ZN(Z[23]) );
  AOI22_X1 U50 ( .A1(A[23]), .A2(n5), .B1(B[23]), .B2(n9), .ZN(n94) );
  INV_X1 U51 ( .A(n95), .ZN(Z[24]) );
  AOI22_X1 U52 ( .A1(A[24]), .A2(n5), .B1(B[24]), .B2(n9), .ZN(n95) );
  INV_X1 U53 ( .A(n96), .ZN(Z[25]) );
  AOI22_X1 U54 ( .A1(A[25]), .A2(n5), .B1(B[25]), .B2(n9), .ZN(n96) );
  INV_X1 U55 ( .A(n97), .ZN(Z[26]) );
  AOI22_X1 U56 ( .A1(A[26]), .A2(n5), .B1(B[26]), .B2(n8), .ZN(n97) );
  INV_X1 U57 ( .A(n98), .ZN(Z[27]) );
  AOI22_X1 U58 ( .A1(A[27]), .A2(n5), .B1(B[27]), .B2(n8), .ZN(n98) );
  INV_X1 U59 ( .A(n99), .ZN(Z[28]) );
  AOI22_X1 U60 ( .A1(A[28]), .A2(n5), .B1(B[28]), .B2(n8), .ZN(n99) );
  INV_X1 U61 ( .A(n100), .ZN(Z[29]) );
  AOI22_X1 U62 ( .A1(A[29]), .A2(n5), .B1(B[29]), .B2(n8), .ZN(n100) );
  INV_X1 U63 ( .A(n102), .ZN(Z[30]) );
  AOI22_X1 U64 ( .A1(A[30]), .A2(n5), .B1(B[30]), .B2(n10), .ZN(n102) );
  INV_X1 U65 ( .A(n84), .ZN(Z[14]) );
  AOI22_X1 U66 ( .A1(A[14]), .A2(n4), .B1(B[14]), .B2(n12), .ZN(n84) );
  INV_X1 U67 ( .A(n90), .ZN(Z[1]) );
  AOI22_X1 U68 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(n10), .ZN(n90) );
  INV_X1 U69 ( .A(n101), .ZN(Z[2]) );
  AOI22_X1 U70 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n7), .ZN(n101) );
  INV_X1 U71 ( .A(n80), .ZN(Z[10]) );
  AOI22_X1 U72 ( .A1(A[10]), .A2(n4), .B1(B[10]), .B2(n13), .ZN(n80) );
  INV_X1 U73 ( .A(n81), .ZN(Z[11]) );
  AOI22_X1 U74 ( .A1(A[11]), .A2(n4), .B1(B[11]), .B2(n13), .ZN(n81) );
  INV_X1 U75 ( .A(n82), .ZN(Z[12]) );
  AOI22_X1 U76 ( .A1(A[12]), .A2(n4), .B1(B[12]), .B2(n12), .ZN(n82) );
  INV_X1 U77 ( .A(n83), .ZN(Z[13]) );
  AOI22_X1 U78 ( .A1(A[13]), .A2(n4), .B1(B[13]), .B2(n12), .ZN(n83) );
endmodule


module mux21_NBIT32_1 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n11) );
  BUF_X1 U6 ( .A(n2), .Z(n9) );
  BUF_X1 U7 ( .A(n1), .Z(n8) );
  BUF_X1 U8 ( .A(n2), .Z(n10) );
  BUF_X1 U9 ( .A(n1), .Z(n7) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(S), .Z(n3) );
  BUF_X1 U13 ( .A(S), .Z(n2) );
  BUF_X1 U14 ( .A(S), .Z(n1) );
  INV_X1 U15 ( .A(n79), .ZN(Z[0]) );
  AOI22_X1 U16 ( .A1(A[0]), .A2(n4), .B1(B[0]), .B2(n13), .ZN(n79) );
  INV_X1 U17 ( .A(n90), .ZN(Z[1]) );
  AOI22_X1 U18 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(n10), .ZN(n90) );
  INV_X1 U19 ( .A(n101), .ZN(Z[2]) );
  AOI22_X1 U20 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n7), .ZN(n101) );
  INV_X1 U21 ( .A(n104), .ZN(Z[3]) );
  AOI22_X1 U22 ( .A1(A[3]), .A2(n4), .B1(B[3]), .B2(n7), .ZN(n104) );
  INV_X1 U23 ( .A(n105), .ZN(Z[4]) );
  AOI22_X1 U24 ( .A1(A[4]), .A2(n5), .B1(B[4]), .B2(n7), .ZN(n105) );
  INV_X1 U25 ( .A(n106), .ZN(Z[5]) );
  AOI22_X1 U26 ( .A1(A[5]), .A2(n4), .B1(B[5]), .B2(n6), .ZN(n106) );
  INV_X1 U27 ( .A(n107), .ZN(Z[6]) );
  AOI22_X1 U28 ( .A1(A[6]), .A2(n5), .B1(B[6]), .B2(n6), .ZN(n107) );
  INV_X1 U29 ( .A(n108), .ZN(Z[7]) );
  AOI22_X1 U30 ( .A1(A[7]), .A2(n4), .B1(B[7]), .B2(n6), .ZN(n108) );
  INV_X1 U31 ( .A(n109), .ZN(Z[8]) );
  AOI22_X1 U32 ( .A1(A[8]), .A2(n5), .B1(B[8]), .B2(n6), .ZN(n109) );
  INV_X1 U33 ( .A(n110), .ZN(Z[9]) );
  AOI22_X1 U34 ( .A1(A[9]), .A2(n4), .B1(n13), .B2(B[9]), .ZN(n110) );
  INV_X1 U35 ( .A(n80), .ZN(Z[10]) );
  AOI22_X1 U36 ( .A1(A[10]), .A2(n4), .B1(B[10]), .B2(n13), .ZN(n80) );
  INV_X1 U37 ( .A(n81), .ZN(Z[11]) );
  AOI22_X1 U38 ( .A1(A[11]), .A2(n4), .B1(B[11]), .B2(n13), .ZN(n81) );
  INV_X1 U39 ( .A(n82), .ZN(Z[12]) );
  AOI22_X1 U40 ( .A1(A[12]), .A2(n4), .B1(B[12]), .B2(n12), .ZN(n82) );
  INV_X1 U41 ( .A(n83), .ZN(Z[13]) );
  AOI22_X1 U42 ( .A1(A[13]), .A2(n4), .B1(B[13]), .B2(n12), .ZN(n83) );
  INV_X1 U43 ( .A(n84), .ZN(Z[14]) );
  AOI22_X1 U44 ( .A1(A[14]), .A2(n4), .B1(B[14]), .B2(n12), .ZN(n84) );
  INV_X1 U45 ( .A(n85), .ZN(Z[15]) );
  AOI22_X1 U46 ( .A1(A[15]), .A2(n4), .B1(B[15]), .B2(n12), .ZN(n85) );
  INV_X1 U47 ( .A(n86), .ZN(Z[16]) );
  AOI22_X1 U48 ( .A1(A[16]), .A2(n4), .B1(B[16]), .B2(n11), .ZN(n86) );
  INV_X1 U49 ( .A(n87), .ZN(Z[17]) );
  AOI22_X1 U50 ( .A1(A[17]), .A2(n4), .B1(B[17]), .B2(n11), .ZN(n87) );
  INV_X1 U51 ( .A(n88), .ZN(Z[18]) );
  AOI22_X1 U52 ( .A1(A[18]), .A2(n4), .B1(B[18]), .B2(n11), .ZN(n88) );
  INV_X1 U53 ( .A(n89), .ZN(Z[19]) );
  AOI22_X1 U54 ( .A1(A[19]), .A2(n4), .B1(B[19]), .B2(n11), .ZN(n89) );
  INV_X1 U55 ( .A(n91), .ZN(Z[20]) );
  AOI22_X1 U56 ( .A1(A[20]), .A2(n5), .B1(B[20]), .B2(n10), .ZN(n91) );
  INV_X1 U57 ( .A(n92), .ZN(Z[21]) );
  AOI22_X1 U58 ( .A1(A[21]), .A2(n5), .B1(B[21]), .B2(n10), .ZN(n92) );
  INV_X1 U59 ( .A(n93), .ZN(Z[22]) );
  AOI22_X1 U60 ( .A1(A[22]), .A2(n5), .B1(B[22]), .B2(n9), .ZN(n93) );
  INV_X1 U61 ( .A(n94), .ZN(Z[23]) );
  AOI22_X1 U62 ( .A1(A[23]), .A2(n5), .B1(B[23]), .B2(n9), .ZN(n94) );
  INV_X1 U63 ( .A(n95), .ZN(Z[24]) );
  AOI22_X1 U64 ( .A1(A[24]), .A2(n5), .B1(B[24]), .B2(n9), .ZN(n95) );
  INV_X1 U65 ( .A(n96), .ZN(Z[25]) );
  AOI22_X1 U66 ( .A1(A[25]), .A2(n5), .B1(B[25]), .B2(n9), .ZN(n96) );
  INV_X1 U67 ( .A(n97), .ZN(Z[26]) );
  AOI22_X1 U68 ( .A1(A[26]), .A2(n5), .B1(B[26]), .B2(n8), .ZN(n97) );
  INV_X1 U69 ( .A(n98), .ZN(Z[27]) );
  AOI22_X1 U70 ( .A1(A[27]), .A2(n5), .B1(B[27]), .B2(n8), .ZN(n98) );
  INV_X1 U71 ( .A(n99), .ZN(Z[28]) );
  AOI22_X1 U72 ( .A1(A[28]), .A2(n5), .B1(B[28]), .B2(n8), .ZN(n99) );
  INV_X1 U73 ( .A(n100), .ZN(Z[29]) );
  AOI22_X1 U74 ( .A1(A[29]), .A2(n5), .B1(B[29]), .B2(n8), .ZN(n100) );
  INV_X1 U75 ( .A(n102), .ZN(Z[30]) );
  AOI22_X1 U76 ( .A1(A[30]), .A2(n5), .B1(B[30]), .B2(n10), .ZN(n102) );
  INV_X1 U77 ( .A(n103), .ZN(Z[31]) );
  AOI22_X1 U78 ( .A1(A[31]), .A2(n5), .B1(B[31]), .B2(n7), .ZN(n103) );
endmodule


module ALU_NBIT32 ( OP1, OP2, .ALU_OPC({\ALU_OPC[4] , \ALU_OPC[3] , 
        \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), ALU_RES );
  input [31:0] OP1;
  input [31:0] OP2;
  output [31:0] ALU_RES;
  input \ALU_OPC[4] , \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] ;
  wire   select_zero_sig, LOGIC_ARITH, LEFT_RIGHT, ADD_SUB, n78, n79, n80, n81,
         n82, n83, n84, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n85,
         n86, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212;
  wire   [4:0] ALU_OPC;
  wire   [1:0] select_type_sig;
  wire   [31:0] A_CMP;
  wire   [31:0] B_CMP;
  wire   [31:0] A_SHF;
  wire   [31:0] B_SHF;
  wire   [31:0] A_ADD;
  wire   [31:0] B_ADD;
  wire   [15:0] A_MUL;
  wire   [15:0] B_MUL;
  wire   [2:0] OPSel;
  wire   [31:0] LOGIC_RES;
  wire   [31:0] COMP_RES;
  wire   [31:0] SHIFT_RES;
  wire   [31:0] ADD_SUB_RES;
  wire   [31:0] MUL_RES;
  wire   [31:0] sig_intraMux;
  wire   [31:0] sig_ALU_RES;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  OAI22_X2 U227 ( .A1(n195), .A2(n39), .B1(n45), .B2(n72), .ZN(A_SHF[31]) );
  NOR2_X2 U257 ( .A1(n86), .A2(n30), .ZN(A_MUL[9]) );
  NOR2_X2 U258 ( .A1(n85), .A2(n30), .ZN(A_MUL[8]) );
  NOR2_X2 U259 ( .A1(n77), .A2(n30), .ZN(A_MUL[7]) );
  NOR2_X2 U260 ( .A1(n76), .A2(n30), .ZN(A_MUL[6]) );
  NOR2_X2 U261 ( .A1(n75), .A2(n29), .ZN(A_MUL[5]) );
  NOR2_X2 U262 ( .A1(n74), .A2(n29), .ZN(A_MUL[4]) );
  NOR2_X2 U263 ( .A1(n73), .A2(n29), .ZN(A_MUL[3]) );
  NOR2_X2 U264 ( .A1(n70), .A2(n29), .ZN(A_MUL[2]) );
  NOR2_X2 U265 ( .A1(n59), .A2(n29), .ZN(A_MUL[1]) );
  NOR2_X2 U267 ( .A1(n53), .A2(n29), .ZN(A_MUL[14]) );
  NOR2_X2 U268 ( .A1(n52), .A2(n29), .ZN(A_MUL[13]) );
  NOR2_X2 U269 ( .A1(n51), .A2(n29), .ZN(A_MUL[12]) );
  NOR2_X2 U270 ( .A1(n50), .A2(n29), .ZN(A_MUL[11]) );
  NOR2_X2 U271 ( .A1(n49), .A2(n29), .ZN(A_MUL[10]) );
  NOR2_X2 U272 ( .A1(n48), .A2(n29), .ZN(A_MUL[0]) );
  NAND3_X1 U427 ( .A1(n212), .A2(n211), .A3(n80), .ZN(n79) );
  NAND3_X1 U428 ( .A1(n47), .A2(n41), .A3(n38), .ZN(select_type_sig[1]) );
  NAND3_X1 U429 ( .A1(n84), .A2(n7), .A3(n38), .ZN(select_type_sig[0]) );
  NAND3_X1 U430 ( .A1(ALU_OPC[3]), .A2(n212), .A3(n156), .ZN(n84) );
  NAND3_X1 U431 ( .A1(ALU_OPC[0]), .A2(ALU_OPC[3]), .A3(n156), .ZN(n158) );
  NAND3_X1 U432 ( .A1(ALU_OPC[4]), .A2(ALU_OPC[1]), .A3(n162), .ZN(n82) );
  NAND3_X1 U434 ( .A1(n211), .A2(n209), .A3(ALU_OPC[4]), .ZN(n164) );
  NAND3_X1 U436 ( .A1(n209), .A2(n204), .A3(n211), .ZN(n170) );
  comparator_NBIT32 Comp ( .A(A_CMP), .B(B_CMP), .OPSel({n206, OPSel[1:0]}), 
        .RES({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, COMP_RES[0]}) );
  shifter_NBIT32 Shift ( .A(A_SHF), .B(B_SHF), .LOGIC_ARITH(LOGIC_ARITH), 
        .LEFT_RIGHT(LEFT_RIGHT), .RES(SHIFT_RES) );
  P4Adder_NBIT32 Add_Sub_unit ( .A(A_ADD), .B(B_ADD), .Cin(ADD_SUB), .S(
        ADD_SUB_RES) );
  BOOTHMUL_numBit16 Booth_mul ( .A(A_MUL), .B(B_MUL), .P(MUL_RES) );
  mux41_NBIT32_1 Res_mux ( .A(ADD_SUB_RES), .B(LOGIC_RES), .C(SHIFT_RES), .D({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, COMP_RES[0]}), .S(
        select_type_sig), .Z(sig_intraMux) );
  mux21_NBIT32_2 Mul_mux ( .A(sig_intraMux), .B(MUL_RES), .S(n1), .Z(
        sig_ALU_RES) );
  mux21_NBIT32_1 Zeros_mux ( .A(sig_ALU_RES), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .S(select_zero_sig), .Z(ALU_RES) );
  OAI22_X1 U3 ( .A1(n198), .A2(n39), .B1(n44), .B2(n75), .ZN(A_SHF[5]) );
  OAI22_X1 U4 ( .A1(n199), .A2(n39), .B1(n44), .B2(n76), .ZN(A_SHF[6]) );
  OAI22_X1 U5 ( .A1(n189), .A2(n40), .B1(n45), .B2(n66), .ZN(A_SHF[26]) );
  OAI22_X1 U6 ( .A1(n190), .A2(n40), .B1(n45), .B2(n67), .ZN(A_SHF[27]) );
  AND3_X1 U7 ( .A1(ALU_OPC[0]), .A2(ALU_OPC[2]), .A3(n163), .ZN(n1) );
  OR2_X1 U8 ( .A1(n211), .A2(n205), .ZN(n2) );
  OR2_X1 U9 ( .A1(n170), .A2(ALU_OPC[0]), .ZN(n3) );
  INV_X1 U10 ( .A(n4), .ZN(ADD_SUB) );
  NOR2_X1 U11 ( .A1(n210), .A2(n3), .ZN(n5) );
  NOR2_X1 U12 ( .A1(n212), .A2(n2), .ZN(n6) );
  NOR2_X1 U13 ( .A1(n5), .A2(n6), .ZN(n4) );
  BUF_X1 U14 ( .A(n168), .Z(n17) );
  BUF_X1 U15 ( .A(n168), .Z(n18) );
  BUF_X1 U16 ( .A(n168), .Z(n19) );
  OAI22_X1 U17 ( .A1(n179), .A2(n41), .B1(n46), .B2(n56), .ZN(A_SHF[17]) );
  OAI22_X1 U18 ( .A1(n200), .A2(n39), .B1(n44), .B2(n77), .ZN(A_SHF[7]) );
  OAI22_X1 U19 ( .A1(n180), .A2(n41), .B1(n46), .B2(n57), .ZN(A_SHF[18]) );
  OAI22_X1 U20 ( .A1(n188), .A2(n40), .B1(n45), .B2(n65), .ZN(A_SHF[25]) );
  OAI22_X1 U21 ( .A1(n191), .A2(n40), .B1(n45), .B2(n68), .ZN(A_SHF[28]) );
  OAI22_X1 U22 ( .A1(n197), .A2(n40), .B1(n45), .B2(n74), .ZN(A_SHF[4]) );
  NOR2_X1 U23 ( .A1(n42), .A2(n196), .ZN(B_SHF[3]) );
  OAI22_X1 U24 ( .A1(n201), .A2(n39), .B1(n44), .B2(n85), .ZN(A_SHF[8]) );
  OAI22_X1 U25 ( .A1(n193), .A2(n39), .B1(n45), .B2(n70), .ZN(A_SHF[2]) );
  OAI22_X1 U26 ( .A1(n186), .A2(n40), .B1(n45), .B2(n63), .ZN(A_SHF[23]) );
  OAI22_X1 U27 ( .A1(n187), .A2(n40), .B1(n45), .B2(n64), .ZN(A_SHF[24]) );
  OAI22_X1 U28 ( .A1(n181), .A2(n40), .B1(n46), .B2(n58), .ZN(A_SHF[19]) );
  OAI22_X1 U29 ( .A1(n183), .A2(n40), .B1(n46), .B2(n60), .ZN(A_SHF[20]) );
  OAI22_X1 U30 ( .A1(n184), .A2(n40), .B1(n46), .B2(n61), .ZN(A_SHF[21]) );
  OAI22_X1 U31 ( .A1(n185), .A2(n40), .B1(n46), .B2(n62), .ZN(A_SHF[22]) );
  OAI22_X1 U32 ( .A1(n174), .A2(n41), .B1(n47), .B2(n51), .ZN(A_SHF[12]) );
  OAI22_X1 U33 ( .A1(n175), .A2(n41), .B1(n46), .B2(n52), .ZN(A_SHF[13]) );
  OAI22_X1 U34 ( .A1(n176), .A2(n41), .B1(n46), .B2(n53), .ZN(A_SHF[14]) );
  NOR2_X1 U35 ( .A1(n196), .A2(n30), .ZN(B_MUL[3]) );
  NOR2_X1 U36 ( .A1(n198), .A2(n30), .ZN(B_MUL[5]) );
  NOR2_X1 U37 ( .A1(n200), .A2(n30), .ZN(B_MUL[7]) );
  NOR2_X1 U38 ( .A1(n202), .A2(n30), .ZN(B_MUL[9]) );
  NOR2_X1 U39 ( .A1(n182), .A2(n30), .ZN(B_MUL[1]) );
  NOR2_X1 U40 ( .A1(n173), .A2(n30), .ZN(B_MUL[11]) );
  NOR2_X1 U41 ( .A1(n175), .A2(n30), .ZN(B_MUL[13]) );
  NOR2_X1 U42 ( .A1(n42), .A2(n202), .ZN(B_SHF[9]) );
  NOR2_X1 U43 ( .A1(n42), .A2(n201), .ZN(B_SHF[8]) );
  NOR2_X1 U44 ( .A1(n44), .A2(n172), .ZN(B_SHF[10]) );
  OAI22_X1 U45 ( .A1(n182), .A2(n40), .B1(n46), .B2(n59), .ZN(A_SHF[1]) );
  NOR2_X1 U46 ( .A1(n42), .A2(n193), .ZN(B_SHF[2]) );
  OAI22_X1 U47 ( .A1(n202), .A2(n39), .B1(n44), .B2(n86), .ZN(A_SHF[9]) );
  OAI22_X1 U48 ( .A1(n171), .A2(n39), .B1(n46), .B2(n48), .ZN(A_SHF[0]) );
  NOR2_X1 U49 ( .A1(n42), .A2(n200), .ZN(B_SHF[7]) );
  NOR2_X1 U50 ( .A1(n42), .A2(n199), .ZN(B_SHF[6]) );
  NOR2_X1 U51 ( .A1(n42), .A2(n198), .ZN(B_SHF[5]) );
  OAI22_X1 U52 ( .A1(n173), .A2(n41), .B1(n47), .B2(n50), .ZN(A_SHF[11]) );
  OAI22_X1 U53 ( .A1(n177), .A2(n41), .B1(n46), .B2(n54), .ZN(A_SHF[15]) );
  OAI22_X1 U54 ( .A1(n192), .A2(n39), .B1(n45), .B2(n69), .ZN(A_SHF[29]) );
  OAI22_X1 U55 ( .A1(n178), .A2(n41), .B1(n46), .B2(n55), .ZN(A_SHF[16]) );
  OAI22_X1 U56 ( .A1(n196), .A2(n39), .B1(n45), .B2(n73), .ZN(A_SHF[3]) );
  NOR2_X1 U57 ( .A1(n17), .A2(n48), .ZN(A_ADD[0]) );
  NOR2_X1 U58 ( .A1(n19), .A2(n74), .ZN(A_ADD[4]) );
  NOR2_X1 U59 ( .A1(n19), .A2(n85), .ZN(A_ADD[8]) );
  NOR2_X1 U60 ( .A1(n19), .A2(n75), .ZN(A_ADD[5]) );
  NOR2_X1 U61 ( .A1(n19), .A2(n86), .ZN(A_ADD[9]) );
  NOR2_X1 U62 ( .A1(n19), .A2(n76), .ZN(A_ADD[6]) );
  NOR2_X1 U63 ( .A1(n19), .A2(n73), .ZN(A_ADD[3]) );
  NOR2_X1 U64 ( .A1(n19), .A2(n77), .ZN(A_ADD[7]) );
  NOR2_X1 U65 ( .A1(n19), .A2(n72), .ZN(A_ADD[31]) );
  NOR2_X1 U66 ( .A1(n17), .A2(n51), .ZN(A_ADD[12]) );
  NOR2_X1 U67 ( .A1(n17), .A2(n55), .ZN(A_ADD[16]) );
  NOR2_X1 U68 ( .A1(n18), .A2(n64), .ZN(A_ADD[24]) );
  NOR2_X1 U69 ( .A1(n17), .A2(n59), .ZN(A_ADD[1]) );
  NOR2_X1 U70 ( .A1(n17), .A2(n52), .ZN(A_ADD[13]) );
  NOR2_X1 U71 ( .A1(n17), .A2(n56), .ZN(A_ADD[17]) );
  NOR2_X1 U72 ( .A1(n18), .A2(n65), .ZN(A_ADD[25]) );
  NOR2_X1 U73 ( .A1(n18), .A2(n70), .ZN(A_ADD[2]) );
  NOR2_X1 U74 ( .A1(n17), .A2(n49), .ZN(A_ADD[10]) );
  NOR2_X1 U75 ( .A1(n17), .A2(n53), .ZN(A_ADD[14]) );
  NOR2_X1 U76 ( .A1(n17), .A2(n57), .ZN(A_ADD[18]) );
  NOR2_X1 U77 ( .A1(n18), .A2(n66), .ZN(A_ADD[26]) );
  NOR2_X1 U78 ( .A1(n18), .A2(n62), .ZN(A_ADD[22]) );
  NOR2_X1 U79 ( .A1(n18), .A2(n61), .ZN(A_ADD[21]) );
  NOR2_X1 U80 ( .A1(n18), .A2(n60), .ZN(A_ADD[20]) );
  NOR2_X1 U81 ( .A1(n18), .A2(n71), .ZN(A_ADD[30]) );
  NOR2_X1 U82 ( .A1(n18), .A2(n69), .ZN(A_ADD[29]) );
  NOR2_X1 U83 ( .A1(n18), .A2(n68), .ZN(A_ADD[28]) );
  NOR2_X1 U84 ( .A1(n17), .A2(n50), .ZN(A_ADD[11]) );
  NOR2_X1 U85 ( .A1(n17), .A2(n54), .ZN(A_ADD[15]) );
  NOR2_X1 U86 ( .A1(n17), .A2(n58), .ZN(A_ADD[19]) );
  NOR2_X1 U87 ( .A1(n18), .A2(n63), .ZN(A_ADD[23]) );
  NOR2_X1 U88 ( .A1(n18), .A2(n67), .ZN(A_ADD[27]) );
  NOR2_X1 U89 ( .A1(n43), .A2(n182), .ZN(B_SHF[1]) );
  NOR2_X1 U90 ( .A1(n42), .A2(n191), .ZN(B_SHF[28]) );
  NOR2_X1 U91 ( .A1(n42), .A2(n190), .ZN(B_SHF[27]) );
  NOR2_X1 U92 ( .A1(n43), .A2(n189), .ZN(B_SHF[26]) );
  OAI22_X1 U93 ( .A1(n172), .A2(n41), .B1(n47), .B2(n49), .ZN(A_SHF[10]) );
  NOR2_X1 U94 ( .A1(n44), .A2(n173), .ZN(B_SHF[11]) );
  NOR2_X1 U95 ( .A1(n177), .A2(n30), .ZN(B_MUL[15]) );
  OAI22_X1 U96 ( .A1(n194), .A2(n39), .B1(n45), .B2(n71), .ZN(A_SHF[30]) );
  NOR2_X1 U97 ( .A1(n43), .A2(n180), .ZN(B_SHF[18]) );
  NOR2_X1 U98 ( .A1(n42), .A2(n192), .ZN(B_SHF[29]) );
  NOR2_X1 U99 ( .A1(n42), .A2(n194), .ZN(B_SHF[30]) );
  BUF_X1 U100 ( .A(n208), .Z(n11) );
  BUF_X1 U101 ( .A(n208), .Z(n12) );
  BUF_X1 U102 ( .A(n208), .Z(n13) );
  BUF_X1 U103 ( .A(n208), .Z(n15) );
  BUF_X1 U104 ( .A(n208), .Z(n14) );
  NOR2_X1 U105 ( .A1(n43), .A2(n188), .ZN(B_SHF[25]) );
  NOR2_X1 U106 ( .A1(n44), .A2(n171), .ZN(B_SHF[0]) );
  NOR2_X1 U107 ( .A1(n43), .A2(n178), .ZN(B_SHF[16]) );
  NOR2_X1 U108 ( .A1(n43), .A2(n179), .ZN(B_SHF[17]) );
  NOR2_X1 U109 ( .A1(n44), .A2(n177), .ZN(B_SHF[15]) );
  NOR2_X1 U110 ( .A1(n54), .A2(n29), .ZN(A_MUL[15]) );
  NOR2_X1 U111 ( .A1(n193), .A2(n30), .ZN(B_MUL[2]) );
  NOR2_X1 U112 ( .A1(n197), .A2(n29), .ZN(B_MUL[4]) );
  NOR2_X1 U113 ( .A1(n199), .A2(n30), .ZN(B_MUL[6]) );
  NOR2_X1 U114 ( .A1(n201), .A2(n29), .ZN(B_MUL[8]) );
  NOR2_X1 U115 ( .A1(n171), .A2(n30), .ZN(B_MUL[0]) );
  NOR2_X1 U116 ( .A1(n172), .A2(n30), .ZN(B_MUL[10]) );
  NOR2_X1 U117 ( .A1(n174), .A2(n30), .ZN(B_MUL[12]) );
  NOR2_X1 U118 ( .A1(n176), .A2(n30), .ZN(B_MUL[14]) );
  BUF_X1 U119 ( .A(n4), .Z(n9) );
  BUF_X1 U120 ( .A(n4), .Z(n8) );
  OAI21_X1 U121 ( .B1(n47), .B2(n197), .A(n41), .ZN(B_SHF[4]) );
  BUF_X1 U122 ( .A(n4), .Z(n10) );
  NOR2_X1 U123 ( .A1(n43), .A2(n187), .ZN(B_SHF[24]) );
  NOR2_X1 U124 ( .A1(n43), .A2(n186), .ZN(B_SHF[23]) );
  NOR2_X1 U125 ( .A1(n43), .A2(n185), .ZN(B_SHF[22]) );
  NOR2_X1 U126 ( .A1(n34), .A2(n71), .ZN(A_CMP[30]) );
  OAI22_X1 U127 ( .A1(n99), .A2(n198), .B1(n100), .B2(n75), .ZN(LOGIC_RES[5])
         );
  OAI22_X1 U128 ( .A1(n97), .A2(n199), .B1(n98), .B2(n76), .ZN(LOGIC_RES[6])
         );
  OAI22_X1 U129 ( .A1(n95), .A2(n200), .B1(n96), .B2(n77), .ZN(LOGIC_RES[7])
         );
  OAI22_X1 U130 ( .A1(n90), .A2(n202), .B1(n91), .B2(n86), .ZN(LOGIC_RES[9])
         );
  OAI22_X1 U131 ( .A1(n105), .A2(n195), .B1(n106), .B2(n72), .ZN(LOGIC_RES[31]) );
  NOR2_X1 U132 ( .A1(n33), .A2(n59), .ZN(A_CMP[1]) );
  OAI22_X1 U133 ( .A1(n151), .A2(n172), .B1(n152), .B2(n49), .ZN(LOGIC_RES[10]) );
  OAI22_X1 U134 ( .A1(n149), .A2(n173), .B1(n150), .B2(n50), .ZN(LOGIC_RES[11]) );
  OAI22_X1 U135 ( .A1(n145), .A2(n175), .B1(n146), .B2(n52), .ZN(LOGIC_RES[13]) );
  OAI22_X1 U136 ( .A1(n143), .A2(n176), .B1(n144), .B2(n53), .ZN(LOGIC_RES[14]) );
  OAI22_X1 U137 ( .A1(n141), .A2(n177), .B1(n142), .B2(n54), .ZN(LOGIC_RES[15]) );
  OAI22_X1 U138 ( .A1(n137), .A2(n179), .B1(n138), .B2(n56), .ZN(LOGIC_RES[17]) );
  OAI22_X1 U139 ( .A1(n135), .A2(n180), .B1(n136), .B2(n57), .ZN(LOGIC_RES[18]) );
  OAI22_X1 U140 ( .A1(n133), .A2(n181), .B1(n134), .B2(n58), .ZN(LOGIC_RES[19]) );
  OAI22_X1 U141 ( .A1(n127), .A2(n184), .B1(n128), .B2(n61), .ZN(LOGIC_RES[21]) );
  OAI22_X1 U142 ( .A1(n125), .A2(n185), .B1(n126), .B2(n62), .ZN(LOGIC_RES[22]) );
  OAI22_X1 U143 ( .A1(n123), .A2(n186), .B1(n124), .B2(n63), .ZN(LOGIC_RES[23]) );
  OAI22_X1 U144 ( .A1(n119), .A2(n188), .B1(n120), .B2(n65), .ZN(LOGIC_RES[25]) );
  OAI22_X1 U145 ( .A1(n117), .A2(n189), .B1(n118), .B2(n66), .ZN(LOGIC_RES[26]) );
  OAI22_X1 U146 ( .A1(n115), .A2(n190), .B1(n116), .B2(n67), .ZN(LOGIC_RES[27]) );
  OAI22_X1 U147 ( .A1(n111), .A2(n192), .B1(n112), .B2(n69), .ZN(LOGIC_RES[29]) );
  OAI22_X1 U148 ( .A1(n107), .A2(n194), .B1(n108), .B2(n71), .ZN(LOGIC_RES[30]) );
  NOR2_X1 U149 ( .A1(n43), .A2(n181), .ZN(B_SHF[19]) );
  NOR2_X1 U150 ( .A1(n43), .A2(n184), .ZN(B_SHF[21]) );
  NOR2_X1 U151 ( .A1(n44), .A2(n175), .ZN(B_SHF[13]) );
  NOR2_X1 U152 ( .A1(n43), .A2(n183), .ZN(B_SHF[20]) );
  NOR2_X1 U153 ( .A1(n44), .A2(n176), .ZN(B_SHF[14]) );
  NOR2_X1 U154 ( .A1(n44), .A2(n174), .ZN(B_SHF[12]) );
  NOR2_X1 U155 ( .A1(n38), .A2(n200), .ZN(B_CMP[7]) );
  NOR2_X1 U156 ( .A1(n38), .A2(n202), .ZN(B_CMP[9]) );
  AOI21_X1 U157 ( .B1(n13), .B2(n198), .A(n25), .ZN(n100) );
  AOI21_X1 U158 ( .B1(n13), .B2(n199), .A(n25), .ZN(n98) );
  AOI21_X1 U159 ( .B1(n13), .B2(n201), .A(n25), .ZN(n94) );
  AOI21_X1 U160 ( .B1(n15), .B2(n182), .A(n27), .ZN(n132) );
  AOI21_X1 U161 ( .B1(n14), .B2(n193), .A(n26), .ZN(n110) );
  AOI21_X1 U162 ( .B1(n14), .B2(n196), .A(n26), .ZN(n104) );
  AOI21_X1 U163 ( .B1(n14), .B2(n197), .A(n26), .ZN(n102) );
  AOI21_X1 U164 ( .B1(n14), .B2(n200), .A(n26), .ZN(n96) );
  AOI21_X1 U165 ( .B1(n14), .B2(n202), .A(n26), .ZN(n91) );
  AOI21_X1 U166 ( .B1(n15), .B2(n176), .A(n27), .ZN(n144) );
  AOI21_X1 U167 ( .B1(n15), .B2(n177), .A(n27), .ZN(n142) );
  AOI21_X1 U168 ( .B1(n15), .B2(n178), .A(n27), .ZN(n140) );
  AOI21_X1 U169 ( .B1(n15), .B2(n179), .A(n27), .ZN(n138) );
  AOI21_X1 U170 ( .B1(n15), .B2(n180), .A(n27), .ZN(n136) );
  AOI21_X1 U171 ( .B1(n15), .B2(n181), .A(n27), .ZN(n134) );
  AOI21_X1 U172 ( .B1(n15), .B2(n183), .A(n27), .ZN(n130) );
  AOI21_X1 U173 ( .B1(n15), .B2(n184), .A(n27), .ZN(n128) );
  AOI21_X1 U174 ( .B1(n15), .B2(n185), .A(n27), .ZN(n126) );
  AOI21_X1 U175 ( .B1(n15), .B2(n186), .A(n27), .ZN(n124) );
  AOI21_X1 U176 ( .B1(n15), .B2(n187), .A(n26), .ZN(n122) );
  AOI21_X1 U177 ( .B1(n14), .B2(n188), .A(n26), .ZN(n120) );
  AOI21_X1 U178 ( .B1(n14), .B2(n189), .A(n26), .ZN(n118) );
  AOI21_X1 U179 ( .B1(n14), .B2(n190), .A(n26), .ZN(n116) );
  AOI21_X1 U180 ( .B1(n14), .B2(n191), .A(n26), .ZN(n114) );
  AOI21_X1 U181 ( .B1(n14), .B2(n192), .A(n26), .ZN(n112) );
  AOI21_X1 U182 ( .B1(n14), .B2(n194), .A(n26), .ZN(n108) );
  AOI21_X1 U183 ( .B1(n14), .B2(n195), .A(n26), .ZN(n106) );
  AOI21_X1 U184 ( .B1(n16), .B2(n172), .A(n28), .ZN(n152) );
  AOI21_X1 U185 ( .B1(n16), .B2(n173), .A(n28), .ZN(n150) );
  AOI21_X1 U186 ( .B1(n16), .B2(n174), .A(n27), .ZN(n148) );
  AOI21_X1 U187 ( .B1(n16), .B2(n175), .A(n27), .ZN(n146) );
  NOR2_X1 U188 ( .A1(n38), .A2(n201), .ZN(B_CMP[8]) );
  NOR2_X1 U189 ( .A1(n38), .A2(n199), .ZN(B_CMP[6]) );
  NOR2_X1 U190 ( .A1(n37), .A2(n194), .ZN(B_CMP[30]) );
  NOR2_X1 U191 ( .A1(n35), .A2(n171), .ZN(B_CMP[0]) );
  NOR2_X1 U192 ( .A1(n37), .A2(n196), .ZN(B_CMP[3]) );
  NOR2_X1 U193 ( .A1(n37), .A2(n198), .ZN(B_CMP[5]) );
  NOR2_X1 U194 ( .A1(n35), .A2(n173), .ZN(B_CMP[11]) );
  NOR2_X1 U195 ( .A1(n36), .A2(n175), .ZN(B_CMP[13]) );
  NOR2_X1 U196 ( .A1(n36), .A2(n177), .ZN(B_CMP[15]) );
  NOR2_X1 U197 ( .A1(n36), .A2(n179), .ZN(B_CMP[17]) );
  NOR2_X1 U198 ( .A1(n36), .A2(n181), .ZN(B_CMP[19]) );
  NOR2_X1 U199 ( .A1(n36), .A2(n184), .ZN(B_CMP[21]) );
  NOR2_X1 U200 ( .A1(n36), .A2(n186), .ZN(B_CMP[23]) );
  NOR2_X1 U201 ( .A1(n37), .A2(n188), .ZN(B_CMP[25]) );
  NOR2_X1 U202 ( .A1(n37), .A2(n190), .ZN(B_CMP[27]) );
  NOR2_X1 U203 ( .A1(n37), .A2(n192), .ZN(B_CMP[29]) );
  NOR2_X1 U204 ( .A1(n35), .A2(n72), .ZN(A_CMP[31]) );
  NOR2_X1 U205 ( .A1(n37), .A2(n197), .ZN(B_CMP[4]) );
  NOR2_X1 U206 ( .A1(n35), .A2(n174), .ZN(B_CMP[12]) );
  NOR2_X1 U207 ( .A1(n36), .A2(n178), .ZN(B_CMP[16]) );
  NOR2_X1 U208 ( .A1(n36), .A2(n183), .ZN(B_CMP[20]) );
  NOR2_X1 U209 ( .A1(n37), .A2(n187), .ZN(B_CMP[24]) );
  NOR2_X1 U210 ( .A1(n37), .A2(n191), .ZN(B_CMP[28]) );
  NOR2_X1 U211 ( .A1(n37), .A2(n193), .ZN(B_CMP[2]) );
  NOR2_X1 U212 ( .A1(n35), .A2(n172), .ZN(B_CMP[10]) );
  NOR2_X1 U213 ( .A1(n36), .A2(n176), .ZN(B_CMP[14]) );
  NOR2_X1 U214 ( .A1(n36), .A2(n180), .ZN(B_CMP[18]) );
  NOR2_X1 U215 ( .A1(n36), .A2(n185), .ZN(B_CMP[22]) );
  NOR2_X1 U216 ( .A1(n37), .A2(n189), .ZN(B_CMP[26]) );
  AND2_X1 U217 ( .A1(n22), .A2(n10), .ZN(n168) );
  NOR2_X1 U218 ( .A1(n42), .A2(n195), .ZN(B_SHF[31]) );
  NOR2_X1 U219 ( .A1(n36), .A2(n182), .ZN(B_CMP[1]) );
  NOR2_X1 U220 ( .A1(n33), .A2(n48), .ZN(A_CMP[0]) );
  NOR2_X1 U221 ( .A1(n35), .A2(n73), .ZN(A_CMP[3]) );
  NOR2_X1 U222 ( .A1(n35), .A2(n75), .ZN(A_CMP[5]) );
  NOR2_X1 U223 ( .A1(n35), .A2(n77), .ZN(A_CMP[7]) );
  NOR2_X1 U224 ( .A1(n35), .A2(n86), .ZN(A_CMP[9]) );
  NOR2_X1 U225 ( .A1(n33), .A2(n50), .ZN(A_CMP[11]) );
  NOR2_X1 U226 ( .A1(n33), .A2(n52), .ZN(A_CMP[13]) );
  NOR2_X1 U228 ( .A1(n33), .A2(n54), .ZN(A_CMP[15]) );
  NOR2_X1 U229 ( .A1(n37), .A2(n195), .ZN(B_CMP[31]) );
  NOR2_X1 U230 ( .A1(n33), .A2(n56), .ZN(A_CMP[17]) );
  NOR2_X1 U231 ( .A1(n33), .A2(n58), .ZN(A_CMP[19]) );
  NOR2_X1 U232 ( .A1(n34), .A2(n61), .ZN(A_CMP[21]) );
  NOR2_X1 U233 ( .A1(n34), .A2(n63), .ZN(A_CMP[23]) );
  NOR2_X1 U234 ( .A1(n34), .A2(n65), .ZN(A_CMP[25]) );
  NOR2_X1 U235 ( .A1(n34), .A2(n67), .ZN(A_CMP[27]) );
  NOR2_X1 U236 ( .A1(n34), .A2(n69), .ZN(A_CMP[29]) );
  NOR2_X1 U237 ( .A1(n35), .A2(n74), .ZN(A_CMP[4]) );
  NOR2_X1 U238 ( .A1(n35), .A2(n85), .ZN(A_CMP[8]) );
  NOR2_X1 U239 ( .A1(n33), .A2(n51), .ZN(A_CMP[12]) );
  NOR2_X1 U240 ( .A1(n34), .A2(n70), .ZN(A_CMP[2]) );
  NOR2_X1 U241 ( .A1(n35), .A2(n76), .ZN(A_CMP[6]) );
  NOR2_X1 U242 ( .A1(n33), .A2(n49), .ZN(A_CMP[10]) );
  NOR2_X1 U243 ( .A1(n33), .A2(n53), .ZN(A_CMP[14]) );
  NOR2_X1 U244 ( .A1(n33), .A2(n55), .ZN(A_CMP[16]) );
  NOR2_X1 U245 ( .A1(n34), .A2(n60), .ZN(A_CMP[20]) );
  NOR2_X1 U246 ( .A1(n34), .A2(n64), .ZN(A_CMP[24]) );
  NOR2_X1 U247 ( .A1(n34), .A2(n68), .ZN(A_CMP[28]) );
  NOR2_X1 U248 ( .A1(n33), .A2(n57), .ZN(A_CMP[18]) );
  NOR2_X1 U249 ( .A1(n34), .A2(n62), .ZN(A_CMP[22]) );
  NOR2_X1 U250 ( .A1(n34), .A2(n66), .ZN(A_CMP[26]) );
  OAI22_X1 U251 ( .A1(OP2[0]), .A2(n10), .B1(n171), .B2(n22), .ZN(B_ADD[0]) );
  OAI22_X1 U252 ( .A1(OP2[4]), .A2(n8), .B1(n197), .B2(n20), .ZN(B_ADD[4]) );
  OAI22_X1 U253 ( .A1(OP2[8]), .A2(n8), .B1(n201), .B2(n20), .ZN(B_ADD[8]) );
  OAI22_X1 U254 ( .A1(OP2[12]), .A2(n10), .B1(n174), .B2(n22), .ZN(B_ADD[12])
         );
  OAI22_X1 U255 ( .A1(OP2[16]), .A2(n10), .B1(n178), .B2(n22), .ZN(B_ADD[16])
         );
  OAI22_X1 U256 ( .A1(OP2[24]), .A2(n9), .B1(n187), .B2(n21), .ZN(B_ADD[24])
         );
  OAI22_X1 U266 ( .A1(OP2[5]), .A2(n8), .B1(n198), .B2(n20), .ZN(B_ADD[5]) );
  OAI22_X1 U273 ( .A1(OP2[1]), .A2(n9), .B1(n182), .B2(n21), .ZN(B_ADD[1]) );
  OAI22_X1 U274 ( .A1(OP2[9]), .A2(n8), .B1(n202), .B2(n20), .ZN(B_ADD[9]) );
  OAI22_X1 U275 ( .A1(OP2[13]), .A2(n10), .B1(n175), .B2(n22), .ZN(B_ADD[13])
         );
  OAI22_X1 U276 ( .A1(OP2[17]), .A2(n9), .B1(n179), .B2(n21), .ZN(B_ADD[17])
         );
  OAI22_X1 U277 ( .A1(OP2[25]), .A2(n9), .B1(n188), .B2(n21), .ZN(B_ADD[25])
         );
  OAI22_X1 U278 ( .A1(OP2[2]), .A2(n8), .B1(n193), .B2(n20), .ZN(B_ADD[2]) );
  OAI22_X1 U279 ( .A1(OP2[6]), .A2(n8), .B1(n199), .B2(n20), .ZN(B_ADD[6]) );
  OAI22_X1 U280 ( .A1(OP2[10]), .A2(n10), .B1(n172), .B2(n22), .ZN(B_ADD[10])
         );
  OAI22_X1 U281 ( .A1(OP2[14]), .A2(n10), .B1(n176), .B2(n22), .ZN(B_ADD[14])
         );
  OAI22_X1 U282 ( .A1(OP2[18]), .A2(n9), .B1(n180), .B2(n21), .ZN(B_ADD[18])
         );
  OAI22_X1 U283 ( .A1(OP2[26]), .A2(n9), .B1(n189), .B2(n21), .ZN(B_ADD[26])
         );
  OAI22_X1 U284 ( .A1(OP2[22]), .A2(n9), .B1(n185), .B2(n21), .ZN(B_ADD[22])
         );
  OAI22_X1 U285 ( .A1(OP2[21]), .A2(n9), .B1(n184), .B2(n21), .ZN(B_ADD[21])
         );
  OAI22_X1 U286 ( .A1(OP2[20]), .A2(n9), .B1(n183), .B2(n21), .ZN(B_ADD[20])
         );
  OAI22_X1 U287 ( .A1(OP2[30]), .A2(n8), .B1(n194), .B2(n20), .ZN(B_ADD[30])
         );
  OAI22_X1 U288 ( .A1(OP2[29]), .A2(n8), .B1(n192), .B2(n20), .ZN(B_ADD[29])
         );
  OAI22_X1 U289 ( .A1(OP2[28]), .A2(n8), .B1(n191), .B2(n20), .ZN(B_ADD[28])
         );
  OAI22_X1 U290 ( .A1(OP2[3]), .A2(n8), .B1(n196), .B2(n20), .ZN(B_ADD[3]) );
  OAI22_X1 U291 ( .A1(OP2[7]), .A2(n8), .B1(n200), .B2(n20), .ZN(B_ADD[7]) );
  OAI22_X1 U292 ( .A1(OP2[11]), .A2(n10), .B1(n173), .B2(n22), .ZN(B_ADD[11])
         );
  OAI22_X1 U293 ( .A1(OP2[15]), .A2(n10), .B1(n177), .B2(n22), .ZN(B_ADD[15])
         );
  OAI22_X1 U294 ( .A1(OP2[19]), .A2(n9), .B1(n181), .B2(n21), .ZN(B_ADD[19])
         );
  OAI22_X1 U295 ( .A1(OP2[23]), .A2(n9), .B1(n186), .B2(n21), .ZN(B_ADD[23])
         );
  OAI22_X1 U296 ( .A1(OP2[27]), .A2(n9), .B1(n190), .B2(n21), .ZN(B_ADD[27])
         );
  OAI22_X1 U297 ( .A1(OP2[31]), .A2(n8), .B1(n195), .B2(n20), .ZN(B_ADD[31])
         );
  INV_X1 U298 ( .A(n1), .ZN(n30) );
  INV_X1 U299 ( .A(n1), .ZN(n29) );
  INV_X1 U300 ( .A(n7), .ZN(n31) );
  INV_X1 U301 ( .A(n7), .ZN(n32) );
  AOI221_X1 U302 ( .B1(OP1[10]), .B2(n31), .C1(n11), .C2(n49), .A(n23), .ZN(
        n151) );
  AOI221_X1 U303 ( .B1(OP1[11]), .B2(n32), .C1(n11), .C2(n50), .A(n23), .ZN(
        n149) );
  AOI221_X1 U304 ( .B1(OP1[12]), .B2(n31), .C1(n11), .C2(n51), .A(n23), .ZN(
        n147) );
  AOI221_X1 U305 ( .B1(OP1[13]), .B2(n32), .C1(n11), .C2(n52), .A(n23), .ZN(
        n145) );
  AOI221_X1 U306 ( .B1(OP1[14]), .B2(n31), .C1(n11), .C2(n53), .A(n23), .ZN(
        n143) );
  AOI221_X1 U307 ( .B1(OP1[15]), .B2(n32), .C1(n11), .C2(n54), .A(n23), .ZN(
        n141) );
  AOI221_X1 U308 ( .B1(OP1[16]), .B2(n31), .C1(n11), .C2(n55), .A(n23), .ZN(
        n139) );
  AOI221_X1 U309 ( .B1(OP1[1]), .B2(n32), .C1(n12), .C2(n59), .A(n24), .ZN(
        n131) );
  AOI221_X1 U310 ( .B1(OP1[2]), .B2(n31), .C1(n13), .C2(n70), .A(n25), .ZN(
        n109) );
  AOI221_X1 U311 ( .B1(OP1[3]), .B2(n31), .C1(n12), .C2(n73), .A(n24), .ZN(
        n103) );
  AOI221_X1 U312 ( .B1(OP1[4]), .B2(n31), .C1(n12), .C2(n74), .A(n24), .ZN(
        n101) );
  AOI221_X1 U313 ( .B1(OP1[5]), .B2(n31), .C1(n12), .C2(n75), .A(n24), .ZN(n99) );
  AOI221_X1 U314 ( .B1(OP1[6]), .B2(n31), .C1(n11), .C2(n76), .A(n23), .ZN(n97) );
  AOI221_X1 U315 ( .B1(OP1[7]), .B2(n31), .C1(n11), .C2(n77), .A(n23), .ZN(n95) );
  AOI221_X1 U316 ( .B1(OP1[8]), .B2(n31), .C1(n11), .C2(n85), .A(n23), .ZN(n93) );
  AOI221_X1 U317 ( .B1(OP1[17]), .B2(n32), .C1(n12), .C2(n56), .A(n24), .ZN(
        n137) );
  AOI221_X1 U318 ( .B1(OP1[18]), .B2(n32), .C1(n12), .C2(n57), .A(n24), .ZN(
        n135) );
  AOI221_X1 U319 ( .B1(OP1[19]), .B2(n32), .C1(n12), .C2(n58), .A(n24), .ZN(
        n133) );
  AOI221_X1 U320 ( .B1(OP1[20]), .B2(n32), .C1(n12), .C2(n60), .A(n24), .ZN(
        n129) );
  AOI221_X1 U321 ( .B1(OP1[21]), .B2(n32), .C1(n12), .C2(n61), .A(n24), .ZN(
        n127) );
  AOI221_X1 U322 ( .B1(OP1[22]), .B2(n32), .C1(n12), .C2(n62), .A(n24), .ZN(
        n125) );
  AOI221_X1 U323 ( .B1(OP1[23]), .B2(n32), .C1(n12), .C2(n63), .A(n24), .ZN(
        n123) );
  AOI221_X1 U324 ( .B1(OP1[24]), .B2(n32), .C1(n13), .C2(n64), .A(n25), .ZN(
        n121) );
  AOI221_X1 U325 ( .B1(OP1[25]), .B2(n32), .C1(n13), .C2(n65), .A(n25), .ZN(
        n119) );
  AOI221_X1 U326 ( .B1(OP1[26]), .B2(n32), .C1(n12), .C2(n66), .A(n24), .ZN(
        n117) );
  AOI221_X1 U327 ( .B1(OP1[27]), .B2(n32), .C1(n13), .C2(n67), .A(n25), .ZN(
        n115) );
  AOI221_X1 U328 ( .B1(OP1[28]), .B2(n31), .C1(n13), .C2(n68), .A(n25), .ZN(
        n113) );
  AOI221_X1 U329 ( .B1(OP1[29]), .B2(n31), .C1(n13), .C2(n69), .A(n25), .ZN(
        n111) );
  AOI221_X1 U330 ( .B1(OP1[30]), .B2(n31), .C1(n13), .C2(n71), .A(n25), .ZN(
        n107) );
  AOI221_X1 U331 ( .B1(OP1[31]), .B2(n31), .C1(n13), .C2(n72), .A(n25), .ZN(
        n105) );
  AOI221_X1 U332 ( .B1(n31), .B2(OP1[9]), .C1(n11), .C2(n86), .A(n23), .ZN(n90) );
  BUF_X1 U333 ( .A(n81), .Z(n43) );
  BUF_X1 U334 ( .A(n81), .Z(n44) );
  BUF_X1 U335 ( .A(n81), .Z(n45) );
  BUF_X1 U336 ( .A(n81), .Z(n46) );
  INV_X1 U337 ( .A(OP2[0]), .ZN(n171) );
  INV_X1 U338 ( .A(OP2[1]), .ZN(n182) );
  INV_X1 U339 ( .A(OP2[2]), .ZN(n193) );
  INV_X1 U340 ( .A(OP2[3]), .ZN(n196) );
  INV_X1 U341 ( .A(OP2[5]), .ZN(n198) );
  INV_X1 U342 ( .A(OP2[6]), .ZN(n199) );
  INV_X1 U343 ( .A(OP2[7]), .ZN(n200) );
  INV_X1 U344 ( .A(OP2[8]), .ZN(n201) );
  INV_X1 U345 ( .A(OP2[9]), .ZN(n202) );
  INV_X1 U346 ( .A(OP2[10]), .ZN(n172) );
  INV_X1 U347 ( .A(OP2[11]), .ZN(n173) );
  INV_X1 U348 ( .A(OP2[12]), .ZN(n174) );
  INV_X1 U349 ( .A(OP2[13]), .ZN(n175) );
  INV_X1 U350 ( .A(OP2[14]), .ZN(n176) );
  INV_X1 U351 ( .A(OP2[15]), .ZN(n177) );
  INV_X1 U352 ( .A(OP2[4]), .ZN(n197) );
  BUF_X1 U353 ( .A(n92), .Z(n23) );
  BUF_X1 U354 ( .A(n92), .Z(n24) );
  OAI22_X1 U355 ( .A1(n153), .A2(n171), .B1(n154), .B2(n48), .ZN(LOGIC_RES[0])
         );
  AOI21_X1 U356 ( .B1(n13), .B2(n171), .A(n25), .ZN(n154) );
  AOI221_X1 U357 ( .B1(OP1[0]), .B2(n32), .C1(n11), .C2(n48), .A(n23), .ZN(
        n153) );
  BUF_X1 U358 ( .A(n92), .Z(n27) );
  BUF_X1 U359 ( .A(n92), .Z(n26) );
  BUF_X1 U360 ( .A(n82), .Z(n39) );
  BUF_X1 U361 ( .A(n82), .Z(n40) );
  BUF_X1 U362 ( .A(n92), .Z(n25) );
  BUF_X1 U363 ( .A(n159), .Z(n21) );
  BUF_X1 U364 ( .A(n159), .Z(n20) );
  BUF_X1 U365 ( .A(n83), .Z(n37) );
  BUF_X1 U366 ( .A(n83), .Z(n35) );
  BUF_X1 U367 ( .A(n83), .Z(n33) );
  BUF_X1 U368 ( .A(n83), .Z(n36) );
  BUF_X1 U369 ( .A(n83), .Z(n34) );
  BUF_X1 U370 ( .A(n81), .Z(n42) );
  INV_X1 U371 ( .A(OP1[0]), .ZN(n48) );
  INV_X1 U372 ( .A(OP1[1]), .ZN(n59) );
  INV_X1 U373 ( .A(OP1[2]), .ZN(n70) );
  INV_X1 U374 ( .A(OP1[3]), .ZN(n73) );
  INV_X1 U375 ( .A(OP1[4]), .ZN(n74) );
  INV_X1 U376 ( .A(OP1[5]), .ZN(n75) );
  INV_X1 U377 ( .A(OP1[6]), .ZN(n76) );
  INV_X1 U378 ( .A(OP1[7]), .ZN(n77) );
  INV_X1 U379 ( .A(OP1[8]), .ZN(n85) );
  INV_X1 U380 ( .A(OP1[9]), .ZN(n86) );
  INV_X1 U381 ( .A(OP1[10]), .ZN(n49) );
  INV_X1 U382 ( .A(OP1[11]), .ZN(n50) );
  INV_X1 U383 ( .A(OP1[12]), .ZN(n51) );
  INV_X1 U384 ( .A(OP1[13]), .ZN(n52) );
  INV_X1 U385 ( .A(OP1[14]), .ZN(n53) );
  INV_X1 U386 ( .A(OP1[15]), .ZN(n54) );
  BUF_X1 U387 ( .A(n159), .Z(n22) );
  INV_X1 U388 ( .A(OP2[16]), .ZN(n178) );
  INV_X1 U389 ( .A(OP2[17]), .ZN(n179) );
  INV_X1 U390 ( .A(OP2[18]), .ZN(n180) );
  INV_X1 U391 ( .A(OP2[19]), .ZN(n181) );
  INV_X1 U392 ( .A(OP2[20]), .ZN(n183) );
  INV_X1 U393 ( .A(OP2[21]), .ZN(n184) );
  INV_X1 U394 ( .A(OP2[22]), .ZN(n185) );
  INV_X1 U395 ( .A(OP2[23]), .ZN(n186) );
  INV_X1 U396 ( .A(OP2[24]), .ZN(n187) );
  INV_X1 U397 ( .A(OP2[25]), .ZN(n188) );
  INV_X1 U398 ( .A(OP2[26]), .ZN(n189) );
  INV_X1 U399 ( .A(OP2[27]), .ZN(n190) );
  INV_X1 U400 ( .A(OP2[28]), .ZN(n191) );
  INV_X1 U401 ( .A(OP2[29]), .ZN(n192) );
  INV_X1 U402 ( .A(OP2[30]), .ZN(n194) );
  INV_X1 U403 ( .A(OP2[31]), .ZN(n195) );
  BUF_X1 U404 ( .A(n82), .Z(n41) );
  NAND2_X1 U405 ( .A1(n88), .A2(n89), .ZN(OPSel[0]) );
  OAI22_X1 U406 ( .A1(n103), .A2(n196), .B1(n104), .B2(n73), .ZN(LOGIC_RES[3])
         );
  OAI22_X1 U407 ( .A1(n101), .A2(n197), .B1(n102), .B2(n74), .ZN(LOGIC_RES[4])
         );
  OAI22_X1 U408 ( .A1(n93), .A2(n201), .B1(n94), .B2(n85), .ZN(LOGIC_RES[8])
         );
  OAI22_X1 U409 ( .A1(n131), .A2(n182), .B1(n132), .B2(n59), .ZN(LOGIC_RES[1])
         );
  OAI22_X1 U410 ( .A1(n109), .A2(n193), .B1(n110), .B2(n70), .ZN(LOGIC_RES[2])
         );
  OAI22_X1 U411 ( .A1(n147), .A2(n174), .B1(n148), .B2(n51), .ZN(LOGIC_RES[12]) );
  OAI22_X1 U412 ( .A1(n139), .A2(n178), .B1(n140), .B2(n55), .ZN(LOGIC_RES[16]) );
  OAI22_X1 U413 ( .A1(n129), .A2(n183), .B1(n130), .B2(n60), .ZN(LOGIC_RES[20]) );
  OAI22_X1 U414 ( .A1(n121), .A2(n187), .B1(n122), .B2(n64), .ZN(LOGIC_RES[24]) );
  OAI22_X1 U415 ( .A1(n113), .A2(n191), .B1(n114), .B2(n68), .ZN(LOGIC_RES[28]) );
  INV_X1 U416 ( .A(OP1[16]), .ZN(n55) );
  INV_X1 U417 ( .A(OP1[17]), .ZN(n56) );
  INV_X1 U418 ( .A(OP1[18]), .ZN(n57) );
  INV_X1 U419 ( .A(OP1[19]), .ZN(n58) );
  INV_X1 U420 ( .A(OP1[20]), .ZN(n60) );
  INV_X1 U421 ( .A(OP1[21]), .ZN(n61) );
  INV_X1 U422 ( .A(OP1[22]), .ZN(n62) );
  INV_X1 U423 ( .A(OP1[23]), .ZN(n63) );
  INV_X1 U424 ( .A(OP1[24]), .ZN(n64) );
  INV_X1 U425 ( .A(OP1[25]), .ZN(n65) );
  INV_X1 U426 ( .A(OP1[26]), .ZN(n66) );
  INV_X1 U433 ( .A(OP1[27]), .ZN(n67) );
  INV_X1 U435 ( .A(OP1[28]), .ZN(n68) );
  INV_X1 U437 ( .A(OP1[29]), .ZN(n69) );
  INV_X1 U438 ( .A(OP1[30]), .ZN(n71) );
  INV_X1 U439 ( .A(OP1[31]), .ZN(n72) );
  NAND2_X1 U440 ( .A1(n157), .A2(n207), .ZN(LOGIC_ARITH) );
  INV_X1 U441 ( .A(LEFT_RIGHT), .ZN(n207) );
  INV_X1 U442 ( .A(n84), .ZN(n208) );
  INV_X1 U443 ( .A(n87), .ZN(n206) );
  INV_X1 U444 ( .A(n80), .ZN(n205) );
  NOR3_X1 U445 ( .A1(n212), .A2(ALU_OPC[3]), .A3(n210), .ZN(n162) );
  NOR3_X1 U446 ( .A1(ALU_OPC[3]), .A2(ALU_OPC[4]), .A3(ALU_OPC[2]), .ZN(n80)
         );
  NAND4_X1 U447 ( .A1(ALU_OPC[4]), .A2(ALU_OPC[1]), .A3(n212), .A4(n209), .ZN(
        n88) );
  NAND4_X1 U448 ( .A1(ALU_OPC[1]), .A2(ALU_OPC[3]), .A3(ALU_OPC[2]), .A4(n204), 
        .ZN(n89) );
  INV_X1 U449 ( .A(ALU_OPC[1]), .ZN(n211) );
  NAND2_X1 U450 ( .A1(n158), .A2(n39), .ZN(LEFT_RIGHT) );
  NOR3_X1 U451 ( .A1(ALU_OPC[1]), .A2(ALU_OPC[4]), .A3(ALU_OPC[2]), .ZN(n156)
         );
  NAND4_X1 U452 ( .A1(ALU_OPC[1]), .A2(ALU_OPC[3]), .A3(n161), .A4(n212), .ZN(
        n157) );
  NOR2_X1 U453 ( .A1(ALU_OPC[4]), .A2(ALU_OPC[2]), .ZN(n161) );
  INV_X1 U454 ( .A(ALU_OPC[2]), .ZN(n210) );
  INV_X1 U455 ( .A(ALU_OPC[3]), .ZN(n209) );
  OAI211_X1 U456 ( .C1(n166), .C2(n167), .A(n209), .B(ALU_OPC[4]), .ZN(n87) );
  NOR2_X1 U457 ( .A1(ALU_OPC[2]), .A2(n211), .ZN(n167) );
  NOR3_X1 U458 ( .A1(n210), .A2(ALU_OPC[1]), .A3(ALU_OPC[0]), .ZN(n166) );
  AND3_X1 U459 ( .A1(ALU_OPC[1]), .A2(ALU_OPC[0]), .A3(n155), .ZN(n92) );
  NOR3_X1 U460 ( .A1(n210), .A2(ALU_OPC[4]), .A3(ALU_OPC[3]), .ZN(n155) );
  INV_X1 U461 ( .A(ALU_OPC[4]), .ZN(n204) );
  INV_X1 U462 ( .A(ALU_OPC[0]), .ZN(n212) );
  OAI21_X1 U463 ( .B1(n78), .B2(n209), .A(n79), .ZN(select_zero_sig) );
  AOI21_X1 U464 ( .B1(ALU_OPC[2]), .B2(n211), .A(ALU_OPC[4]), .ZN(n78) );
  NAND2_X1 U465 ( .A1(n165), .A2(n89), .ZN(OPSel[1]) );
  NAND4_X1 U466 ( .A1(ALU_OPC[4]), .A2(n211), .A3(n210), .A4(n209), .ZN(n165)
         );
  NAND2_X1 U467 ( .A1(n80), .A2(n169), .ZN(n159) );
  XNOR2_X1 U468 ( .A(n211), .B(ALU_OPC[0]), .ZN(n169) );
  AND4_X1 U469 ( .A1(n164), .A2(n88), .A3(n87), .A4(n203), .ZN(n83) );
  INV_X1 U470 ( .A(OPSel[1]), .ZN(n203) );
  OR4_X1 U471 ( .A1(n211), .A2(n210), .A3(ALU_OPC[3]), .A4(ALU_OPC[4]), .ZN(n7) );
  AND2_X1 U472 ( .A1(n160), .A2(n157), .ZN(n81) );
  NAND4_X1 U473 ( .A1(ALU_OPC[0]), .A2(ALU_OPC[3]), .A3(n210), .A4(n204), .ZN(
        n160) );
  NOR3_X1 U474 ( .A1(ALU_OPC[1]), .A2(ALU_OPC[4]), .A3(ALU_OPC[3]), .ZN(n163)
         );
  CLKBUF_X1 U475 ( .A(n208), .Z(n16) );
  CLKBUF_X1 U476 ( .A(n92), .Z(n28) );
  CLKBUF_X1 U477 ( .A(n83), .Z(n38) );
  CLKBUF_X1 U478 ( .A(n81), .Z(n47) );
endmodule


module regn_N32_5 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
endmodule


module regn_N32_4 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
endmodule


module regn_N5_2 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 \DOUT_reg[4]  ( .D(n16), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n21)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n17), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n22)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n18), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n23)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n19), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n24)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n20), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n25)
         );
  OAI21_X1 U2 ( .B1(n25), .B2(EN), .A(n30), .ZN(n20) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n30) );
  OAI21_X1 U4 ( .B1(n24), .B2(EN), .A(n29), .ZN(n19) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n29) );
  OAI21_X1 U6 ( .B1(n22), .B2(EN), .A(n27), .ZN(n17) );
  NAND2_X1 U7 ( .A1(DIN[3]), .A2(EN), .ZN(n27) );
  OAI21_X1 U8 ( .B1(n23), .B2(EN), .A(n28), .ZN(n18) );
  NAND2_X1 U9 ( .A1(DIN[2]), .A2(EN), .ZN(n28) );
  OAI21_X1 U10 ( .B1(n21), .B2(EN), .A(n26), .ZN(n16) );
  NAND2_X1 U11 ( .A1(DIN[4]), .A2(EN), .ZN(n26) );
endmodule


module regn_N32_3 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
endmodule


module regn_N32_2 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
endmodule


module Execute_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \B[0] , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57;
  assign SUM[1] = B[1];
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR2_X1 U1 ( .A(B[31]), .B(n57), .ZN(SUM[31]) );
  NAND2_X1 U2 ( .A1(B[30]), .A2(n56), .ZN(n57) );
  INV_X1 U3 ( .A(B[2]), .ZN(SUM[2]) );
  XOR2_X1 U4 ( .A(B[3]), .B(B[2]), .Z(SUM[3]) );
  XOR2_X1 U5 ( .A(B[4]), .B(n30), .Z(SUM[4]) );
  XOR2_X1 U6 ( .A(B[5]), .B(n31), .Z(SUM[5]) );
  XOR2_X1 U7 ( .A(B[6]), .B(n32), .Z(SUM[6]) );
  XOR2_X1 U8 ( .A(B[7]), .B(n33), .Z(SUM[7]) );
  XOR2_X1 U9 ( .A(B[8]), .B(n34), .Z(SUM[8]) );
  XOR2_X1 U10 ( .A(B[9]), .B(n35), .Z(SUM[9]) );
  XOR2_X1 U11 ( .A(B[10]), .B(n36), .Z(SUM[10]) );
  XOR2_X1 U12 ( .A(B[11]), .B(n37), .Z(SUM[11]) );
  XOR2_X1 U13 ( .A(B[12]), .B(n38), .Z(SUM[12]) );
  XOR2_X1 U14 ( .A(B[13]), .B(n39), .Z(SUM[13]) );
  XOR2_X1 U15 ( .A(B[14]), .B(n40), .Z(SUM[14]) );
  XOR2_X1 U16 ( .A(B[15]), .B(n41), .Z(SUM[15]) );
  XOR2_X1 U17 ( .A(B[16]), .B(n42), .Z(SUM[16]) );
  XOR2_X1 U18 ( .A(B[17]), .B(n43), .Z(SUM[17]) );
  XOR2_X1 U19 ( .A(B[18]), .B(n44), .Z(SUM[18]) );
  XOR2_X1 U20 ( .A(B[19]), .B(n45), .Z(SUM[19]) );
  XOR2_X1 U21 ( .A(B[20]), .B(n46), .Z(SUM[20]) );
  XOR2_X1 U22 ( .A(B[21]), .B(n47), .Z(SUM[21]) );
  XOR2_X1 U23 ( .A(B[22]), .B(n48), .Z(SUM[22]) );
  XOR2_X1 U24 ( .A(B[23]), .B(n49), .Z(SUM[23]) );
  XOR2_X1 U25 ( .A(B[24]), .B(n50), .Z(SUM[24]) );
  XOR2_X1 U26 ( .A(B[25]), .B(n51), .Z(SUM[25]) );
  XOR2_X1 U27 ( .A(B[26]), .B(n52), .Z(SUM[26]) );
  XOR2_X1 U28 ( .A(B[27]), .B(n53), .Z(SUM[27]) );
  XOR2_X1 U29 ( .A(B[28]), .B(n54), .Z(SUM[28]) );
  XOR2_X1 U30 ( .A(B[29]), .B(n55), .Z(SUM[29]) );
  XOR2_X1 U31 ( .A(B[30]), .B(n56), .Z(SUM[30]) );
  AND2_X1 U32 ( .A1(B[3]), .A2(B[2]), .ZN(n30) );
  AND2_X1 U33 ( .A1(B[4]), .A2(n30), .ZN(n31) );
  AND2_X1 U34 ( .A1(B[5]), .A2(n31), .ZN(n32) );
  AND2_X1 U35 ( .A1(B[6]), .A2(n32), .ZN(n33) );
  AND2_X1 U36 ( .A1(B[7]), .A2(n33), .ZN(n34) );
  AND2_X1 U37 ( .A1(B[8]), .A2(n34), .ZN(n35) );
  AND2_X1 U38 ( .A1(B[9]), .A2(n35), .ZN(n36) );
  AND2_X1 U39 ( .A1(B[10]), .A2(n36), .ZN(n37) );
  AND2_X1 U40 ( .A1(B[11]), .A2(n37), .ZN(n38) );
  AND2_X1 U41 ( .A1(B[12]), .A2(n38), .ZN(n39) );
  AND2_X1 U42 ( .A1(B[13]), .A2(n39), .ZN(n40) );
  AND2_X1 U43 ( .A1(B[14]), .A2(n40), .ZN(n41) );
  AND2_X1 U44 ( .A1(B[15]), .A2(n41), .ZN(n42) );
  AND2_X1 U45 ( .A1(B[16]), .A2(n42), .ZN(n43) );
  AND2_X1 U46 ( .A1(B[17]), .A2(n43), .ZN(n44) );
  AND2_X1 U47 ( .A1(B[18]), .A2(n44), .ZN(n45) );
  AND2_X1 U48 ( .A1(B[19]), .A2(n45), .ZN(n46) );
  AND2_X1 U49 ( .A1(B[20]), .A2(n46), .ZN(n47) );
  AND2_X1 U50 ( .A1(B[21]), .A2(n47), .ZN(n48) );
  AND2_X1 U51 ( .A1(B[22]), .A2(n48), .ZN(n49) );
  AND2_X1 U52 ( .A1(B[23]), .A2(n49), .ZN(n50) );
  AND2_X1 U53 ( .A1(B[24]), .A2(n50), .ZN(n51) );
  AND2_X1 U54 ( .A1(B[25]), .A2(n51), .ZN(n52) );
  AND2_X1 U55 ( .A1(B[26]), .A2(n52), .ZN(n53) );
  AND2_X1 U56 ( .A1(B[27]), .A2(n53), .ZN(n54) );
  AND2_X1 U57 ( .A1(B[28]), .A2(n54), .ZN(n55) );
  AND2_X1 U58 ( .A1(B[29]), .A2(n55), .ZN(n56) );
endmodule


module Execute_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module Execute ( CLK, RST, MUX_A_SEL, MUX_B_SEL, .ALU_OPC({\ALU_OPC[4] , 
        \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), 
        ALU_OUTREG_EN, JUMP_TYPE, PC_IN, A_IN, B_IN, IMM_IN, ADD_WR_IN, 
        ADD_RS1_IN, ADD_RS2_IN, ADD_WR_MEM, ADD_WR_WB, RF_WE_MEM, RF_WE_WB, 
        OP_MEM, OP_WB, PC_SEL, ZERO_FLAG, NPC_ABS, NPC_REL, ALU_RES, B_OUT, 
        ADD_WR_OUT );
  input [1:0] MUX_B_SEL;
  input [1:0] JUMP_TYPE;
  input [31:0] PC_IN;
  input [31:0] A_IN;
  input [31:0] B_IN;
  input [31:0] IMM_IN;
  input [4:0] ADD_WR_IN;
  input [4:0] ADD_RS1_IN;
  input [4:0] ADD_RS2_IN;
  input [4:0] ADD_WR_MEM;
  input [4:0] ADD_WR_WB;
  input [31:0] OP_MEM;
  input [31:0] OP_WB;
  output [1:0] PC_SEL;
  output [31:0] NPC_ABS;
  output [31:0] NPC_REL;
  output [31:0] ALU_RES;
  output [31:0] B_OUT;
  output [4:0] ADD_WR_OUT;
  input CLK, RST, MUX_A_SEL, \ALU_OPC[4] , \ALU_OPC[3] , \ALU_OPC[2] ,
         \ALU_OPC[1] , \ALU_OPC[0] , ALU_OUTREG_EN, RF_WE_MEM, RF_WE_WB;
  output ZERO_FLAG;
  wire   sig_RST, sig_ZERO_FLAG, N9, N8, N7, N6, N5, N4, N31, N30, N3, N29,
         N28, N27, N26, N25, N24, N23, N22, N21, N20, N2, N19, N18, N17, N16,
         N15, N14, N13, N12, N11, N10, N1, N0, n1;
  wire   [4:0] ALU_OPC;
  wire   [31:0] sig_NPC_ABS;
  wire   [31:0] sig_NPC_REL;
  wire   [1:0] sig_PC_SEL;
  wire   [1:0] FWDA;
  wire   [1:0] FWDB;
  wire   [31:0] OP2_FW;
  wire   [31:0] sig_OP1;
  wire   [31:0] sig_OP2;
  wire   [31:0] sig_ALU_RES;

  Branch_Cond_Unit_NBIT32 Branch_Cond ( .RST(sig_RST), .A(sig_NPC_ABS), 
        .ALU_OPC({\ALU_OPC[4] , \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , 
        \ALU_OPC[0] }), .JUMP_TYPE(JUMP_TYPE), .PC_SEL(sig_PC_SEL), .ZERO(
        sig_ZERO_FLAG) );
  ff_1 ff0 ( .D(sig_ZERO_FLAG), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(ZERO_FLAG)
         );
  regn_N2 reg0 ( .DIN(sig_PC_SEL), .CLK(CLK), .EN(1'b1), .RST(RST), .DOUT(
        PC_SEL) );
  FWD_Unit FWD ( .RST(sig_RST), .ADD_RS1(ADD_RS1_IN), .ADD_RS2(ADD_RS2_IN), 
        .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_WB(ADD_WR_WB), .RF_WE_MEM(RF_WE_MEM), 
        .RF_WE_WB(RF_WE_WB), .FWDA(FWDA), .FWDB(FWDB) );
  mux41_NBIT32_0 FW1 ( .A(A_IN), .B(OP_WB), .C(OP_MEM), .D(A_IN), .S(FWDA), 
        .Z(sig_NPC_ABS) );
  mux41_NBIT32_4 FW2 ( .A(B_IN), .B(OP_WB), .C(OP_MEM), .D(B_IN), .S(FWDB), 
        .Z(OP2_FW) );
  mux21_NBIT32_4 muxA ( .A(sig_NPC_ABS), .B(PC_IN), .S(MUX_A_SEL), .Z(sig_OP1)
         );
  mux41_NBIT32_3 muxB ( .A(OP2_FW), .B(IMM_IN), .C({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(MUX_B_SEL), .Z(sig_OP2) );
  ALU_NBIT32 alu0 ( .OP1(sig_OP1), .OP2(sig_OP2), .ALU_OPC({\ALU_OPC[4] , 
        \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), .ALU_RES(
        sig_ALU_RES) );
  regn_N32_5 alureg ( .DIN(sig_ALU_RES), .CLK(CLK), .EN(ALU_OUTREG_EN), .RST(
        RST), .DOUT(ALU_RES) );
  regn_N32_4 B_reg ( .DIN(OP2_FW), .CLK(CLK), .EN(ALU_OUTREG_EN), .RST(RST), 
        .DOUT(B_OUT) );
  regn_N5_2 ADD_WR_reg ( .DIN(ADD_WR_IN), .CLK(CLK), .EN(1'b1), .RST(RST), 
        .DOUT(ADD_WR_OUT) );
  regn_N32_3 NPC_ABS_reg ( .DIN(sig_NPC_ABS), .CLK(CLK), .EN(ALU_OUTREG_EN), 
        .RST(RST), .DOUT(NPC_ABS) );
  regn_N32_2 NPC_REL_reg ( .DIN(sig_NPC_REL), .CLK(CLK), .EN(ALU_OUTREG_EN), 
        .RST(RST), .DOUT(NPC_REL) );
  Execute_DW01_add_1 add_1_root_add_0_root_add_122_2 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .B(IMM_IN), .CI(1'b0), .SUM({N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0})
         );
  Execute_DW01_add_0 add_0_root_add_0_root_add_122_2 ( .A(PC_IN), .B({N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}), 
        .CI(1'b0), .SUM(sig_NPC_REL) );
  NOR2_X1 U3 ( .A1(ZERO_FLAG), .A2(n1), .ZN(sig_RST) );
  INV_X1 U4 ( .A(RST), .ZN(n1) );
endmodule


module ff_0 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n2, n3;

  DFFR_X1 Q_reg ( .D(n3), .CK(CLK), .RN(RST), .Q(Q), .QN(n2) );
  OAI21_X1 U2 ( .B1(n2), .B2(EN), .A(n1), .ZN(n3) );
  NAND2_X1 U3 ( .A1(EN), .A2(D), .ZN(n1) );
endmodule


module regn_N5_1 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 \DOUT_reg[4]  ( .D(n16), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n21)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n17), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n22)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n18), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n23)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n19), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n24)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n20), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n25)
         );
  OAI21_X1 U2 ( .B1(n25), .B2(EN), .A(n30), .ZN(n20) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n30) );
  OAI21_X1 U4 ( .B1(n24), .B2(EN), .A(n29), .ZN(n19) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n29) );
  OAI21_X1 U6 ( .B1(n23), .B2(EN), .A(n28), .ZN(n18) );
  NAND2_X1 U7 ( .A1(DIN[2]), .A2(EN), .ZN(n28) );
  OAI21_X1 U8 ( .B1(n22), .B2(EN), .A(n27), .ZN(n17) );
  NAND2_X1 U9 ( .A1(DIN[3]), .A2(EN), .ZN(n27) );
  OAI21_X1 U10 ( .B1(n21), .B2(EN), .A(n26), .ZN(n16) );
  NAND2_X1 U11 ( .A1(DIN[4]), .A2(EN), .ZN(n26) );
endmodule


module regn_N32_1 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  OAI21_X1 U2 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U4 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U6 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U7 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U8 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U9 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U10 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U11 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U12 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U13 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U14 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U15 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U16 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U17 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U18 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U19 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U20 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U21 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U22 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U23 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U24 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U25 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U26 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U27 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U28 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U29 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U30 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U31 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U32 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U33 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U34 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U35 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U36 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U37 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U38 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U39 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U40 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U41 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U42 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U43 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U44 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U45 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U46 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U47 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U48 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U49 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U50 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U51 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U52 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U53 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U54 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U55 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U56 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U57 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U58 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U59 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U60 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U61 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U62 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U63 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U64 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U65 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
  BUF_X1 U66 ( .A(RST), .Z(n97) );
  BUF_X1 U67 ( .A(RST), .Z(n98) );
  BUF_X1 U68 ( .A(RST), .Z(n99) );
endmodule


module mux41_NBIT32_2 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n20, n21, n22, n23, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94;

  BUF_X1 U1 ( .A(n1), .Z(n20) );
  BUF_X1 U2 ( .A(n1), .Z(n9) );
  BUF_X1 U3 ( .A(n3), .Z(n22) );
  BUF_X1 U4 ( .A(n2), .Z(n6) );
  BUF_X1 U5 ( .A(n3), .Z(n21) );
  BUF_X1 U6 ( .A(n2), .Z(n5) );
  AND2_X1 U7 ( .A1(n23), .A2(n26), .ZN(n1) );
  BUF_X1 U8 ( .A(n4), .Z(n8) );
  BUF_X1 U9 ( .A(n4), .Z(n7) );
  NAND2_X1 U10 ( .A1(n80), .A2(n79), .ZN(Z[0]) );
  AOI22_X1 U11 ( .A1(D[0]), .A2(n7), .B1(C[0]), .B2(n5), .ZN(n79) );
  AOI22_X1 U12 ( .A1(B[0]), .A2(n21), .B1(A[0]), .B2(n9), .ZN(n80) );
  NAND2_X1 U13 ( .A1(n94), .A2(n93), .ZN(Z[7]) );
  AOI22_X1 U14 ( .A1(D[7]), .A2(n7), .B1(C[7]), .B2(n5), .ZN(n93) );
  AOI22_X1 U15 ( .A1(B[7]), .A2(n21), .B1(A[7]), .B2(n9), .ZN(n94) );
  AND2_X1 U16 ( .A1(S[1]), .A2(n26), .ZN(n2) );
  AND2_X1 U17 ( .A1(S[0]), .A2(n23), .ZN(n3) );
  NAND2_X1 U18 ( .A1(n82), .A2(n81), .ZN(Z[1]) );
  AOI22_X1 U19 ( .A1(D[1]), .A2(n7), .B1(C[1]), .B2(n5), .ZN(n81) );
  AOI22_X1 U20 ( .A1(B[1]), .A2(n21), .B1(A[1]), .B2(n9), .ZN(n82) );
  NAND2_X1 U21 ( .A1(n84), .A2(n83), .ZN(Z[2]) );
  AOI22_X1 U22 ( .A1(D[2]), .A2(n7), .B1(C[2]), .B2(n5), .ZN(n83) );
  AOI22_X1 U23 ( .A1(B[2]), .A2(n21), .B1(A[2]), .B2(n9), .ZN(n84) );
  NAND2_X1 U24 ( .A1(n86), .A2(n85), .ZN(Z[3]) );
  AOI22_X1 U25 ( .A1(D[3]), .A2(n7), .B1(C[3]), .B2(n5), .ZN(n85) );
  AOI22_X1 U26 ( .A1(B[3]), .A2(n21), .B1(A[3]), .B2(n9), .ZN(n86) );
  NAND2_X1 U27 ( .A1(n92), .A2(n91), .ZN(Z[6]) );
  AOI22_X1 U28 ( .A1(D[6]), .A2(n7), .B1(C[6]), .B2(n5), .ZN(n91) );
  AOI22_X1 U29 ( .A1(B[6]), .A2(n21), .B1(A[6]), .B2(n9), .ZN(n92) );
  NAND2_X1 U30 ( .A1(n90), .A2(n89), .ZN(Z[5]) );
  AOI22_X1 U31 ( .A1(D[5]), .A2(n7), .B1(C[5]), .B2(n5), .ZN(n89) );
  AOI22_X1 U32 ( .A1(B[5]), .A2(n21), .B1(A[5]), .B2(n9), .ZN(n90) );
  NAND2_X1 U33 ( .A1(n88), .A2(n87), .ZN(Z[4]) );
  AOI22_X1 U34 ( .A1(D[4]), .A2(n7), .B1(C[4]), .B2(n5), .ZN(n87) );
  AOI22_X1 U35 ( .A1(B[4]), .A2(n21), .B1(A[4]), .B2(n9), .ZN(n88) );
  AND2_X1 U36 ( .A1(S[0]), .A2(S[1]), .ZN(n4) );
  INV_X1 U37 ( .A(S[1]), .ZN(n23) );
  INV_X1 U38 ( .A(S[0]), .ZN(n26) );
  AOI22_X1 U39 ( .A1(B[8]), .A2(n22), .B1(A[8]), .B2(n20), .ZN(n28) );
  AOI22_X1 U40 ( .A1(D[8]), .A2(n8), .B1(C[8]), .B2(n6), .ZN(n27) );
  NAND2_X1 U41 ( .A1(n28), .A2(n27), .ZN(Z[8]) );
  AOI22_X1 U42 ( .A1(B[9]), .A2(n22), .B1(A[9]), .B2(n20), .ZN(n30) );
  AOI22_X1 U43 ( .A1(D[9]), .A2(n8), .B1(C[9]), .B2(n6), .ZN(n29) );
  NAND2_X1 U44 ( .A1(n30), .A2(n29), .ZN(Z[9]) );
  AOI22_X1 U45 ( .A1(B[10]), .A2(n22), .B1(A[10]), .B2(n20), .ZN(n32) );
  AOI22_X1 U46 ( .A1(D[10]), .A2(n8), .B1(C[10]), .B2(n6), .ZN(n31) );
  NAND2_X1 U47 ( .A1(n32), .A2(n31), .ZN(Z[10]) );
  AOI22_X1 U48 ( .A1(B[11]), .A2(n22), .B1(A[11]), .B2(n20), .ZN(n34) );
  AOI22_X1 U49 ( .A1(D[11]), .A2(n8), .B1(C[11]), .B2(n6), .ZN(n33) );
  NAND2_X1 U50 ( .A1(n34), .A2(n33), .ZN(Z[11]) );
  AOI22_X1 U51 ( .A1(B[12]), .A2(n22), .B1(A[12]), .B2(n20), .ZN(n36) );
  AOI22_X1 U52 ( .A1(D[12]), .A2(n8), .B1(C[12]), .B2(n6), .ZN(n35) );
  NAND2_X1 U53 ( .A1(n36), .A2(n35), .ZN(Z[12]) );
  AOI22_X1 U54 ( .A1(B[13]), .A2(n22), .B1(A[13]), .B2(n20), .ZN(n38) );
  AOI22_X1 U55 ( .A1(D[13]), .A2(n8), .B1(C[13]), .B2(n6), .ZN(n37) );
  NAND2_X1 U56 ( .A1(n38), .A2(n37), .ZN(Z[13]) );
  AOI22_X1 U57 ( .A1(B[14]), .A2(n22), .B1(A[14]), .B2(n20), .ZN(n40) );
  AOI22_X1 U58 ( .A1(D[14]), .A2(n8), .B1(C[14]), .B2(n6), .ZN(n39) );
  NAND2_X1 U59 ( .A1(n40), .A2(n39), .ZN(Z[14]) );
  AOI22_X1 U60 ( .A1(B[15]), .A2(n22), .B1(A[15]), .B2(n20), .ZN(n42) );
  AOI22_X1 U61 ( .A1(D[15]), .A2(n8), .B1(C[15]), .B2(n6), .ZN(n41) );
  NAND2_X1 U62 ( .A1(n42), .A2(n41), .ZN(Z[15]) );
  AOI22_X1 U63 ( .A1(B[16]), .A2(n22), .B1(A[16]), .B2(n20), .ZN(n44) );
  AOI22_X1 U64 ( .A1(D[16]), .A2(n8), .B1(C[16]), .B2(n6), .ZN(n43) );
  NAND2_X1 U65 ( .A1(n44), .A2(n43), .ZN(Z[16]) );
  AOI22_X1 U66 ( .A1(B[17]), .A2(n22), .B1(A[17]), .B2(n20), .ZN(n48) );
  AOI22_X1 U67 ( .A1(D[17]), .A2(n8), .B1(C[17]), .B2(n6), .ZN(n45) );
  NAND2_X1 U68 ( .A1(n48), .A2(n45), .ZN(Z[17]) );
  AOI22_X1 U69 ( .A1(B[18]), .A2(n22), .B1(A[18]), .B2(n20), .ZN(n50) );
  AOI22_X1 U70 ( .A1(D[18]), .A2(n8), .B1(C[18]), .B2(n6), .ZN(n49) );
  NAND2_X1 U71 ( .A1(n50), .A2(n49), .ZN(Z[18]) );
  AOI22_X1 U72 ( .A1(B[19]), .A2(n22), .B1(A[19]), .B2(n20), .ZN(n52) );
  AOI22_X1 U73 ( .A1(D[19]), .A2(n8), .B1(C[19]), .B2(n6), .ZN(n51) );
  NAND2_X1 U74 ( .A1(n52), .A2(n51), .ZN(Z[19]) );
  AOI22_X1 U75 ( .A1(B[20]), .A2(n22), .B1(A[20]), .B2(n20), .ZN(n54) );
  AOI22_X1 U76 ( .A1(D[20]), .A2(n8), .B1(C[20]), .B2(n6), .ZN(n53) );
  NAND2_X1 U77 ( .A1(n54), .A2(n53), .ZN(Z[20]) );
  AOI22_X1 U78 ( .A1(B[21]), .A2(n22), .B1(A[21]), .B2(n20), .ZN(n56) );
  AOI22_X1 U79 ( .A1(D[21]), .A2(n8), .B1(C[21]), .B2(n6), .ZN(n55) );
  NAND2_X1 U80 ( .A1(n56), .A2(n55), .ZN(Z[21]) );
  AOI22_X1 U81 ( .A1(B[22]), .A2(n22), .B1(A[22]), .B2(n20), .ZN(n58) );
  AOI22_X1 U82 ( .A1(D[22]), .A2(n8), .B1(C[22]), .B2(n6), .ZN(n57) );
  NAND2_X1 U83 ( .A1(n58), .A2(n57), .ZN(Z[22]) );
  AOI22_X1 U84 ( .A1(B[23]), .A2(n22), .B1(A[23]), .B2(n20), .ZN(n60) );
  AOI22_X1 U85 ( .A1(D[23]), .A2(n8), .B1(C[23]), .B2(n6), .ZN(n59) );
  NAND2_X1 U86 ( .A1(n60), .A2(n59), .ZN(Z[23]) );
  AOI22_X1 U87 ( .A1(B[24]), .A2(n22), .B1(A[24]), .B2(n20), .ZN(n62) );
  AOI22_X1 U88 ( .A1(D[24]), .A2(n8), .B1(C[24]), .B2(n6), .ZN(n61) );
  NAND2_X1 U89 ( .A1(n62), .A2(n61), .ZN(Z[24]) );
  AOI22_X1 U90 ( .A1(B[25]), .A2(n21), .B1(A[25]), .B2(n9), .ZN(n64) );
  AOI22_X1 U91 ( .A1(D[25]), .A2(n7), .B1(C[25]), .B2(n5), .ZN(n63) );
  NAND2_X1 U92 ( .A1(n64), .A2(n63), .ZN(Z[25]) );
  AOI22_X1 U93 ( .A1(B[26]), .A2(n21), .B1(A[26]), .B2(n9), .ZN(n66) );
  AOI22_X1 U94 ( .A1(D[26]), .A2(n7), .B1(C[26]), .B2(n5), .ZN(n65) );
  NAND2_X1 U95 ( .A1(n66), .A2(n65), .ZN(Z[26]) );
  AOI22_X1 U96 ( .A1(B[27]), .A2(n21), .B1(A[27]), .B2(n9), .ZN(n70) );
  AOI22_X1 U97 ( .A1(D[27]), .A2(n7), .B1(C[27]), .B2(n5), .ZN(n67) );
  NAND2_X1 U98 ( .A1(n70), .A2(n67), .ZN(Z[27]) );
  AOI22_X1 U99 ( .A1(B[28]), .A2(n21), .B1(A[28]), .B2(n9), .ZN(n72) );
  AOI22_X1 U100 ( .A1(D[28]), .A2(n7), .B1(C[28]), .B2(n5), .ZN(n71) );
  NAND2_X1 U101 ( .A1(n72), .A2(n71), .ZN(Z[28]) );
  AOI22_X1 U102 ( .A1(B[29]), .A2(n21), .B1(A[29]), .B2(n9), .ZN(n74) );
  AOI22_X1 U103 ( .A1(D[29]), .A2(n7), .B1(C[29]), .B2(n5), .ZN(n73) );
  NAND2_X1 U104 ( .A1(n74), .A2(n73), .ZN(Z[29]) );
  AOI22_X1 U105 ( .A1(B[30]), .A2(n21), .B1(A[30]), .B2(n9), .ZN(n76) );
  AOI22_X1 U106 ( .A1(D[30]), .A2(n7), .B1(C[30]), .B2(n5), .ZN(n75) );
  NAND2_X1 U107 ( .A1(n76), .A2(n75), .ZN(Z[30]) );
  AOI22_X1 U108 ( .A1(B[31]), .A2(n21), .B1(A[31]), .B2(n9), .ZN(n78) );
  AOI22_X1 U109 ( .A1(D[31]), .A2(n7), .B1(C[31]), .B2(n5), .ZN(n77) );
  NAND2_X1 U110 ( .A1(n78), .A2(n77), .ZN(Z[31]) );
endmodule


module Memory ( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, PC_SEL, NPC_IN, 
        NPC_ABS, NPC_REL, ALU_RES_IN, B_IN, ADD_WR_IN, DRAM_DATA_IN, 
        LOAD_TYPE_IN, STORE_TYPE_IN, PC_OUT, DRAM_R_OUT, DRAM_W_OUT, 
        DRAM_ADDR_OUT, DRAM_DATA_OUT, DATA_OUT, ALU_RES_OUT, OP_MEM, 
        ADD_WR_MEM, ADD_WR_OUT, LOAD_TYPE_OUT, STORE_TYPE_OUT );
  input [1:0] PC_SEL;
  input [31:0] NPC_IN;
  input [31:0] NPC_ABS;
  input [31:0] NPC_REL;
  input [31:0] ALU_RES_IN;
  input [31:0] B_IN;
  input [4:0] ADD_WR_IN;
  input [31:0] DRAM_DATA_IN;
  input [1:0] LOAD_TYPE_IN;
  output [31:0] PC_OUT;
  output [31:0] DRAM_ADDR_OUT;
  output [31:0] DRAM_DATA_OUT;
  output [31:0] DATA_OUT;
  output [31:0] ALU_RES_OUT;
  output [31:0] OP_MEM;
  output [4:0] ADD_WR_MEM;
  output [4:0] ADD_WR_OUT;
  output [1:0] LOAD_TYPE_OUT;
  input CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, STORE_TYPE_IN;
  output DRAM_R_OUT, DRAM_W_OUT, STORE_TYPE_OUT;
  wire   DRAM_R_IN, DRAM_W_IN, STORE_TYPE_IN;
  assign DRAM_R_OUT = DRAM_R_IN;
  assign DRAM_W_OUT = DRAM_W_IN;
  assign OP_MEM[31] = ALU_RES_IN[31];
  assign DRAM_ADDR_OUT[31] = ALU_RES_IN[31];
  assign OP_MEM[30] = ALU_RES_IN[30];
  assign DRAM_ADDR_OUT[30] = ALU_RES_IN[30];
  assign OP_MEM[29] = ALU_RES_IN[29];
  assign DRAM_ADDR_OUT[29] = ALU_RES_IN[29];
  assign OP_MEM[28] = ALU_RES_IN[28];
  assign DRAM_ADDR_OUT[28] = ALU_RES_IN[28];
  assign OP_MEM[27] = ALU_RES_IN[27];
  assign DRAM_ADDR_OUT[27] = ALU_RES_IN[27];
  assign OP_MEM[26] = ALU_RES_IN[26];
  assign DRAM_ADDR_OUT[26] = ALU_RES_IN[26];
  assign OP_MEM[25] = ALU_RES_IN[25];
  assign DRAM_ADDR_OUT[25] = ALU_RES_IN[25];
  assign OP_MEM[24] = ALU_RES_IN[24];
  assign DRAM_ADDR_OUT[24] = ALU_RES_IN[24];
  assign OP_MEM[23] = ALU_RES_IN[23];
  assign DRAM_ADDR_OUT[23] = ALU_RES_IN[23];
  assign OP_MEM[22] = ALU_RES_IN[22];
  assign DRAM_ADDR_OUT[22] = ALU_RES_IN[22];
  assign OP_MEM[21] = ALU_RES_IN[21];
  assign DRAM_ADDR_OUT[21] = ALU_RES_IN[21];
  assign OP_MEM[20] = ALU_RES_IN[20];
  assign DRAM_ADDR_OUT[20] = ALU_RES_IN[20];
  assign OP_MEM[19] = ALU_RES_IN[19];
  assign DRAM_ADDR_OUT[19] = ALU_RES_IN[19];
  assign OP_MEM[18] = ALU_RES_IN[18];
  assign DRAM_ADDR_OUT[18] = ALU_RES_IN[18];
  assign OP_MEM[17] = ALU_RES_IN[17];
  assign DRAM_ADDR_OUT[17] = ALU_RES_IN[17];
  assign OP_MEM[16] = ALU_RES_IN[16];
  assign DRAM_ADDR_OUT[16] = ALU_RES_IN[16];
  assign OP_MEM[15] = ALU_RES_IN[15];
  assign DRAM_ADDR_OUT[15] = ALU_RES_IN[15];
  assign OP_MEM[14] = ALU_RES_IN[14];
  assign DRAM_ADDR_OUT[14] = ALU_RES_IN[14];
  assign OP_MEM[13] = ALU_RES_IN[13];
  assign DRAM_ADDR_OUT[13] = ALU_RES_IN[13];
  assign OP_MEM[12] = ALU_RES_IN[12];
  assign DRAM_ADDR_OUT[12] = ALU_RES_IN[12];
  assign OP_MEM[11] = ALU_RES_IN[11];
  assign DRAM_ADDR_OUT[11] = ALU_RES_IN[11];
  assign OP_MEM[10] = ALU_RES_IN[10];
  assign DRAM_ADDR_OUT[10] = ALU_RES_IN[10];
  assign OP_MEM[9] = ALU_RES_IN[9];
  assign DRAM_ADDR_OUT[9] = ALU_RES_IN[9];
  assign OP_MEM[8] = ALU_RES_IN[8];
  assign DRAM_ADDR_OUT[8] = ALU_RES_IN[8];
  assign OP_MEM[7] = ALU_RES_IN[7];
  assign DRAM_ADDR_OUT[7] = ALU_RES_IN[7];
  assign OP_MEM[6] = ALU_RES_IN[6];
  assign DRAM_ADDR_OUT[6] = ALU_RES_IN[6];
  assign OP_MEM[5] = ALU_RES_IN[5];
  assign DRAM_ADDR_OUT[5] = ALU_RES_IN[5];
  assign OP_MEM[4] = ALU_RES_IN[4];
  assign DRAM_ADDR_OUT[4] = ALU_RES_IN[4];
  assign OP_MEM[3] = ALU_RES_IN[3];
  assign DRAM_ADDR_OUT[3] = ALU_RES_IN[3];
  assign OP_MEM[2] = ALU_RES_IN[2];
  assign DRAM_ADDR_OUT[2] = ALU_RES_IN[2];
  assign OP_MEM[1] = ALU_RES_IN[1];
  assign DRAM_ADDR_OUT[1] = ALU_RES_IN[1];
  assign OP_MEM[0] = ALU_RES_IN[0];
  assign DRAM_ADDR_OUT[0] = ALU_RES_IN[0];
  assign DRAM_DATA_OUT[31] = B_IN[31];
  assign DRAM_DATA_OUT[30] = B_IN[30];
  assign DRAM_DATA_OUT[29] = B_IN[29];
  assign DRAM_DATA_OUT[28] = B_IN[28];
  assign DRAM_DATA_OUT[27] = B_IN[27];
  assign DRAM_DATA_OUT[26] = B_IN[26];
  assign DRAM_DATA_OUT[25] = B_IN[25];
  assign DRAM_DATA_OUT[24] = B_IN[24];
  assign DRAM_DATA_OUT[23] = B_IN[23];
  assign DRAM_DATA_OUT[22] = B_IN[22];
  assign DRAM_DATA_OUT[21] = B_IN[21];
  assign DRAM_DATA_OUT[20] = B_IN[20];
  assign DRAM_DATA_OUT[19] = B_IN[19];
  assign DRAM_DATA_OUT[18] = B_IN[18];
  assign DRAM_DATA_OUT[17] = B_IN[17];
  assign DRAM_DATA_OUT[16] = B_IN[16];
  assign DRAM_DATA_OUT[15] = B_IN[15];
  assign DRAM_DATA_OUT[14] = B_IN[14];
  assign DRAM_DATA_OUT[13] = B_IN[13];
  assign DRAM_DATA_OUT[12] = B_IN[12];
  assign DRAM_DATA_OUT[11] = B_IN[11];
  assign DRAM_DATA_OUT[10] = B_IN[10];
  assign DRAM_DATA_OUT[9] = B_IN[9];
  assign DRAM_DATA_OUT[8] = B_IN[8];
  assign DRAM_DATA_OUT[7] = B_IN[7];
  assign DRAM_DATA_OUT[6] = B_IN[6];
  assign DRAM_DATA_OUT[5] = B_IN[5];
  assign DRAM_DATA_OUT[4] = B_IN[4];
  assign DRAM_DATA_OUT[3] = B_IN[3];
  assign DRAM_DATA_OUT[2] = B_IN[2];
  assign DRAM_DATA_OUT[1] = B_IN[1];
  assign DRAM_DATA_OUT[0] = B_IN[0];
  assign DATA_OUT[31] = DRAM_DATA_IN[31];
  assign DATA_OUT[30] = DRAM_DATA_IN[30];
  assign DATA_OUT[29] = DRAM_DATA_IN[29];
  assign DATA_OUT[28] = DRAM_DATA_IN[28];
  assign DATA_OUT[27] = DRAM_DATA_IN[27];
  assign DATA_OUT[26] = DRAM_DATA_IN[26];
  assign DATA_OUT[25] = DRAM_DATA_IN[25];
  assign DATA_OUT[24] = DRAM_DATA_IN[24];
  assign DATA_OUT[23] = DRAM_DATA_IN[23];
  assign DATA_OUT[22] = DRAM_DATA_IN[22];
  assign DATA_OUT[21] = DRAM_DATA_IN[21];
  assign DATA_OUT[20] = DRAM_DATA_IN[20];
  assign DATA_OUT[19] = DRAM_DATA_IN[19];
  assign DATA_OUT[18] = DRAM_DATA_IN[18];
  assign DATA_OUT[17] = DRAM_DATA_IN[17];
  assign DATA_OUT[16] = DRAM_DATA_IN[16];
  assign DATA_OUT[15] = DRAM_DATA_IN[15];
  assign DATA_OUT[14] = DRAM_DATA_IN[14];
  assign DATA_OUT[13] = DRAM_DATA_IN[13];
  assign DATA_OUT[12] = DRAM_DATA_IN[12];
  assign DATA_OUT[11] = DRAM_DATA_IN[11];
  assign DATA_OUT[10] = DRAM_DATA_IN[10];
  assign DATA_OUT[9] = DRAM_DATA_IN[9];
  assign DATA_OUT[8] = DRAM_DATA_IN[8];
  assign DATA_OUT[7] = DRAM_DATA_IN[7];
  assign DATA_OUT[6] = DRAM_DATA_IN[6];
  assign DATA_OUT[5] = DRAM_DATA_IN[5];
  assign DATA_OUT[4] = DRAM_DATA_IN[4];
  assign DATA_OUT[3] = DRAM_DATA_IN[3];
  assign DATA_OUT[2] = DRAM_DATA_IN[2];
  assign DATA_OUT[1] = DRAM_DATA_IN[1];
  assign DATA_OUT[0] = DRAM_DATA_IN[0];
  assign ADD_WR_MEM[4] = ADD_WR_IN[4];
  assign ADD_WR_MEM[3] = ADD_WR_IN[3];
  assign ADD_WR_MEM[2] = ADD_WR_IN[2];
  assign ADD_WR_MEM[1] = ADD_WR_IN[1];
  assign ADD_WR_MEM[0] = ADD_WR_IN[0];
  assign LOAD_TYPE_OUT[1] = LOAD_TYPE_IN[1];
  assign LOAD_TYPE_OUT[0] = LOAD_TYPE_IN[0];
  assign STORE_TYPE_OUT = STORE_TYPE_IN;

  regn_N5_1 reg0 ( .DIN(ADD_WR_IN), .CLK(CLK), .EN(MEM_EN_IN), .RST(RST), 
        .DOUT(ADD_WR_OUT) );
  regn_N32_1 reg1 ( .DIN(ALU_RES_IN), .CLK(CLK), .EN(MEM_EN_IN), .RST(RST), 
        .DOUT(ALU_RES_OUT) );
  mux41_NBIT32_2 PCsel ( .A(NPC_IN), .B(NPC_REL), .C(NPC_ABS), .D({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(PC_SEL), .Z(PC_OUT) );
endmodule


module ff_2 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n4, n5, n6;

  DFFR_X1 Q_reg ( .D(n4), .CK(CLK), .RN(RST), .Q(Q), .QN(n5) );
  OAI21_X1 U2 ( .B1(n5), .B2(EN), .A(n6), .ZN(n4) );
  NAND2_X1 U3 ( .A1(EN), .A2(D), .ZN(n6) );
endmodule


module mux21_NBIT32_3 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100;

  BUF_X1 U1 ( .A(n68), .Z(n1) );
  BUF_X1 U2 ( .A(n68), .Z(n2) );
  BUF_X1 U3 ( .A(n68), .Z(n3) );
  INV_X1 U4 ( .A(n100), .ZN(Z[9]) );
  AOI22_X1 U5 ( .A1(A[9]), .A2(n3), .B1(S), .B2(B[9]), .ZN(n100) );
  INV_X1 U6 ( .A(n82), .ZN(Z[21]) );
  AOI22_X1 U7 ( .A1(A[21]), .A2(n2), .B1(B[21]), .B2(S), .ZN(n82) );
  INV_X1 U8 ( .A(n83), .ZN(Z[22]) );
  AOI22_X1 U9 ( .A1(A[22]), .A2(n2), .B1(B[22]), .B2(S), .ZN(n83) );
  INV_X1 U10 ( .A(n84), .ZN(Z[23]) );
  AOI22_X1 U11 ( .A1(A[23]), .A2(n2), .B1(B[23]), .B2(S), .ZN(n84) );
  INV_X1 U12 ( .A(n77), .ZN(Z[17]) );
  AOI22_X1 U13 ( .A1(A[17]), .A2(n1), .B1(B[17]), .B2(S), .ZN(n77) );
  INV_X1 U14 ( .A(n78), .ZN(Z[18]) );
  AOI22_X1 U15 ( .A1(A[18]), .A2(n1), .B1(B[18]), .B2(S), .ZN(n78) );
  INV_X1 U16 ( .A(n79), .ZN(Z[19]) );
  AOI22_X1 U17 ( .A1(A[19]), .A2(n1), .B1(B[19]), .B2(S), .ZN(n79) );
  INV_X1 U18 ( .A(n80), .ZN(Z[1]) );
  AOI22_X1 U19 ( .A1(A[1]), .A2(n1), .B1(B[1]), .B2(S), .ZN(n80) );
  INV_X1 U20 ( .A(n73), .ZN(Z[13]) );
  AOI22_X1 U21 ( .A1(A[13]), .A2(n1), .B1(B[13]), .B2(S), .ZN(n73) );
  INV_X1 U22 ( .A(n74), .ZN(Z[14]) );
  AOI22_X1 U23 ( .A1(A[14]), .A2(n1), .B1(B[14]), .B2(S), .ZN(n74) );
  INV_X1 U24 ( .A(n75), .ZN(Z[15]) );
  AOI22_X1 U25 ( .A1(A[15]), .A2(n1), .B1(B[15]), .B2(S), .ZN(n75) );
  INV_X1 U26 ( .A(n76), .ZN(Z[16]) );
  AOI22_X1 U27 ( .A1(A[16]), .A2(n1), .B1(B[16]), .B2(S), .ZN(n76) );
  INV_X1 U28 ( .A(n69), .ZN(Z[0]) );
  AOI22_X1 U29 ( .A1(A[0]), .A2(n1), .B1(B[0]), .B2(S), .ZN(n69) );
  INV_X1 U30 ( .A(n72), .ZN(Z[12]) );
  AOI22_X1 U31 ( .A1(A[12]), .A2(n1), .B1(B[12]), .B2(S), .ZN(n72) );
  INV_X1 U32 ( .A(n97), .ZN(Z[6]) );
  AOI22_X1 U33 ( .A1(A[6]), .A2(n3), .B1(B[6]), .B2(S), .ZN(n97) );
  INV_X1 U34 ( .A(n98), .ZN(Z[7]) );
  AOI22_X1 U35 ( .A1(A[7]), .A2(n3), .B1(B[7]), .B2(S), .ZN(n98) );
  INV_X1 U36 ( .A(n99), .ZN(Z[8]) );
  AOI22_X1 U37 ( .A1(A[8]), .A2(n3), .B1(B[8]), .B2(S), .ZN(n99) );
  INV_X1 U38 ( .A(n94), .ZN(Z[3]) );
  AOI22_X1 U39 ( .A1(A[3]), .A2(n3), .B1(B[3]), .B2(S), .ZN(n94) );
  INV_X1 U40 ( .A(n95), .ZN(Z[4]) );
  AOI22_X1 U41 ( .A1(A[4]), .A2(n3), .B1(B[4]), .B2(S), .ZN(n95) );
  INV_X1 U42 ( .A(n96), .ZN(Z[5]) );
  AOI22_X1 U43 ( .A1(A[5]), .A2(n3), .B1(B[5]), .B2(S), .ZN(n96) );
  INV_X1 U44 ( .A(n89), .ZN(Z[28]) );
  AOI22_X1 U45 ( .A1(A[28]), .A2(n2), .B1(B[28]), .B2(S), .ZN(n89) );
  INV_X1 U46 ( .A(n90), .ZN(Z[29]) );
  AOI22_X1 U47 ( .A1(A[29]), .A2(n2), .B1(B[29]), .B2(S), .ZN(n90) );
  INV_X1 U48 ( .A(n91), .ZN(Z[2]) );
  AOI22_X1 U49 ( .A1(A[2]), .A2(n2), .B1(B[2]), .B2(S), .ZN(n91) );
  INV_X1 U50 ( .A(n92), .ZN(Z[30]) );
  AOI22_X1 U51 ( .A1(A[30]), .A2(n2), .B1(B[30]), .B2(S), .ZN(n92) );
  INV_X1 U52 ( .A(n86), .ZN(Z[25]) );
  AOI22_X1 U53 ( .A1(A[25]), .A2(n2), .B1(B[25]), .B2(S), .ZN(n86) );
  INV_X1 U54 ( .A(n87), .ZN(Z[26]) );
  AOI22_X1 U55 ( .A1(A[26]), .A2(n2), .B1(B[26]), .B2(S), .ZN(n87) );
  INV_X1 U56 ( .A(n88), .ZN(Z[27]) );
  AOI22_X1 U57 ( .A1(A[27]), .A2(n2), .B1(B[27]), .B2(S), .ZN(n88) );
  INV_X1 U58 ( .A(n93), .ZN(Z[31]) );
  AOI22_X1 U59 ( .A1(A[31]), .A2(n3), .B1(B[31]), .B2(S), .ZN(n93) );
  INV_X1 U60 ( .A(n81), .ZN(Z[20]) );
  AOI22_X1 U61 ( .A1(A[20]), .A2(n2), .B1(B[20]), .B2(S), .ZN(n81) );
  INV_X1 U62 ( .A(n70), .ZN(Z[10]) );
  AOI22_X1 U63 ( .A1(A[10]), .A2(n1), .B1(B[10]), .B2(S), .ZN(n70) );
  INV_X1 U64 ( .A(n85), .ZN(Z[24]) );
  AOI22_X1 U65 ( .A1(A[24]), .A2(n2), .B1(B[24]), .B2(S), .ZN(n85) );
  INV_X1 U66 ( .A(n71), .ZN(Z[11]) );
  AOI22_X1 U67 ( .A1(A[11]), .A2(n1), .B1(B[11]), .B2(S), .ZN(n71) );
  INV_X1 U68 ( .A(S), .ZN(n68) );
endmodule


module Writeback ( WB_MUX_SEL, DATA_IN, ALU_RES_IN, ADD_WR_IN, DATA_OUT, 
        ADD_WR_OUT );
  input [31:0] DATA_IN;
  input [31:0] ALU_RES_IN;
  input [4:0] ADD_WR_IN;
  output [31:0] DATA_OUT;
  output [4:0] ADD_WR_OUT;
  input WB_MUX_SEL;

  assign ADD_WR_OUT[4] = ADD_WR_IN[4];
  assign ADD_WR_OUT[3] = ADD_WR_IN[3];
  assign ADD_WR_OUT[2] = ADD_WR_IN[2];
  assign ADD_WR_OUT[1] = ADD_WR_IN[1];
  assign ADD_WR_OUT[0] = ADD_WR_IN[0];

  mux21_NBIT32_3 WBmux ( .A(ALU_RES_IN), .B(DATA_IN), .S(WB_MUX_SEL), .Z(
        DATA_OUT) );
endmodule


module HazardDetection_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n57;
  assign SUM[1] = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XNOR2_X1 U1 ( .A(A[31]), .B(n57), .ZN(SUM[31]) );
  XOR2_X1 U2 ( .A(A[30]), .B(n51), .Z(SUM[30]) );
  XOR2_X1 U3 ( .A(A[9]), .B(n31), .Z(SUM[9]) );
  XOR2_X1 U4 ( .A(A[8]), .B(n30), .Z(SUM[8]) );
  XOR2_X1 U5 ( .A(A[10]), .B(n25), .Z(SUM[10]) );
  XOR2_X1 U6 ( .A(A[11]), .B(n32), .Z(SUM[11]) );
  XOR2_X1 U7 ( .A(A[12]), .B(n33), .Z(SUM[12]) );
  XOR2_X1 U8 ( .A(A[13]), .B(n34), .Z(SUM[13]) );
  XOR2_X1 U9 ( .A(A[14]), .B(n35), .Z(SUM[14]) );
  XOR2_X1 U10 ( .A(A[15]), .B(n36), .Z(SUM[15]) );
  XOR2_X1 U11 ( .A(A[16]), .B(n37), .Z(SUM[16]) );
  XOR2_X1 U12 ( .A(A[17]), .B(n38), .Z(SUM[17]) );
  XOR2_X1 U13 ( .A(A[18]), .B(n39), .Z(SUM[18]) );
  XOR2_X1 U14 ( .A(A[19]), .B(n40), .Z(SUM[19]) );
  XOR2_X1 U15 ( .A(A[20]), .B(n41), .Z(SUM[20]) );
  XOR2_X1 U16 ( .A(A[21]), .B(n42), .Z(SUM[21]) );
  XOR2_X1 U17 ( .A(A[22]), .B(n43), .Z(SUM[22]) );
  XOR2_X1 U18 ( .A(A[23]), .B(n44), .Z(SUM[23]) );
  XOR2_X1 U19 ( .A(A[24]), .B(n45), .Z(SUM[24]) );
  XOR2_X1 U20 ( .A(A[25]), .B(n46), .Z(SUM[25]) );
  XOR2_X1 U21 ( .A(A[26]), .B(n47), .Z(SUM[26]) );
  XOR2_X1 U22 ( .A(A[27]), .B(n48), .Z(SUM[27]) );
  XOR2_X1 U23 ( .A(A[28]), .B(n49), .Z(SUM[28]) );
  XOR2_X1 U24 ( .A(A[29]), .B(n50), .Z(SUM[29]) );
  NAND2_X1 U25 ( .A1(A[30]), .A2(n51), .ZN(n57) );
  AND2_X1 U26 ( .A1(A[9]), .A2(n31), .ZN(n25) );
  AND2_X1 U27 ( .A1(A[3]), .A2(A[2]), .ZN(n26) );
  AND2_X1 U28 ( .A1(A[4]), .A2(n26), .ZN(n27) );
  AND2_X1 U29 ( .A1(A[5]), .A2(n27), .ZN(n28) );
  AND2_X1 U30 ( .A1(A[6]), .A2(n28), .ZN(n29) );
  AND2_X1 U31 ( .A1(A[7]), .A2(n29), .ZN(n30) );
  AND2_X1 U32 ( .A1(A[8]), .A2(n30), .ZN(n31) );
  AND2_X1 U33 ( .A1(A[10]), .A2(n25), .ZN(n32) );
  AND2_X1 U34 ( .A1(A[11]), .A2(n32), .ZN(n33) );
  AND2_X1 U35 ( .A1(A[12]), .A2(n33), .ZN(n34) );
  AND2_X1 U36 ( .A1(A[13]), .A2(n34), .ZN(n35) );
  AND2_X1 U37 ( .A1(A[14]), .A2(n35), .ZN(n36) );
  AND2_X1 U38 ( .A1(A[15]), .A2(n36), .ZN(n37) );
  AND2_X1 U39 ( .A1(A[16]), .A2(n37), .ZN(n38) );
  AND2_X1 U40 ( .A1(A[17]), .A2(n38), .ZN(n39) );
  AND2_X1 U41 ( .A1(A[18]), .A2(n39), .ZN(n40) );
  AND2_X1 U42 ( .A1(A[19]), .A2(n40), .ZN(n41) );
  AND2_X1 U43 ( .A1(A[20]), .A2(n41), .ZN(n42) );
  AND2_X1 U44 ( .A1(A[21]), .A2(n42), .ZN(n43) );
  AND2_X1 U45 ( .A1(A[22]), .A2(n43), .ZN(n44) );
  AND2_X1 U46 ( .A1(A[23]), .A2(n44), .ZN(n45) );
  AND2_X1 U47 ( .A1(A[24]), .A2(n45), .ZN(n46) );
  AND2_X1 U48 ( .A1(A[25]), .A2(n46), .ZN(n47) );
  AND2_X1 U49 ( .A1(A[26]), .A2(n47), .ZN(n48) );
  AND2_X1 U50 ( .A1(A[27]), .A2(n48), .ZN(n49) );
  AND2_X1 U51 ( .A1(A[28]), .A2(n49), .ZN(n50) );
  AND2_X1 U52 ( .A1(A[29]), .A2(n50), .ZN(n51) );
  INV_X1 U53 ( .A(A[2]), .ZN(SUM[2]) );
  XOR2_X1 U54 ( .A(A[3]), .B(A[2]), .Z(SUM[3]) );
  XOR2_X1 U55 ( .A(A[4]), .B(n26), .Z(SUM[4]) );
  XOR2_X1 U56 ( .A(A[5]), .B(n27), .Z(SUM[5]) );
  XOR2_X1 U57 ( .A(A[6]), .B(n28), .Z(SUM[6]) );
  XOR2_X1 U58 ( .A(A[7]), .B(n29), .Z(SUM[7]) );
endmodule


module HazardDetection ( RST, ADD_RS1, ADD_RS2, ADD_WR, DRAM_R, INS_IN, PC_IN, 
        Bubble, HDU_INS_OUT, HDU_PC_OUT, HDU_NPC_OUT );
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [4:0] ADD_WR;
  input [31:0] INS_IN;
  input [31:0] PC_IN;
  output [31:0] HDU_INS_OUT;
  output [31:0] HDU_PC_OUT;
  output [31:0] HDU_NPC_OUT;
  input RST, DRAM_R;
  output Bubble;
  wire   n1, n2, n3, n4, n5, n6, n9, n10, n12, n13, n14, n15, n16;
  assign HDU_INS_OUT[31] = INS_IN[31];
  assign HDU_INS_OUT[30] = INS_IN[30];
  assign HDU_INS_OUT[29] = INS_IN[29];
  assign HDU_INS_OUT[28] = INS_IN[28];
  assign HDU_INS_OUT[27] = INS_IN[27];
  assign HDU_INS_OUT[26] = INS_IN[26];
  assign HDU_INS_OUT[25] = INS_IN[25];
  assign HDU_INS_OUT[24] = INS_IN[24];
  assign HDU_INS_OUT[23] = INS_IN[23];
  assign HDU_INS_OUT[22] = INS_IN[22];
  assign HDU_INS_OUT[21] = INS_IN[21];
  assign HDU_INS_OUT[20] = INS_IN[20];
  assign HDU_INS_OUT[19] = INS_IN[19];
  assign HDU_INS_OUT[18] = INS_IN[18];
  assign HDU_INS_OUT[17] = INS_IN[17];
  assign HDU_INS_OUT[16] = INS_IN[16];
  assign HDU_INS_OUT[15] = INS_IN[15];
  assign HDU_INS_OUT[14] = INS_IN[14];
  assign HDU_INS_OUT[13] = INS_IN[13];
  assign HDU_INS_OUT[12] = INS_IN[12];
  assign HDU_INS_OUT[11] = INS_IN[11];
  assign HDU_INS_OUT[10] = INS_IN[10];
  assign HDU_INS_OUT[9] = INS_IN[9];
  assign HDU_INS_OUT[8] = INS_IN[8];
  assign HDU_INS_OUT[7] = INS_IN[7];
  assign HDU_INS_OUT[6] = INS_IN[6];
  assign HDU_INS_OUT[5] = INS_IN[5];
  assign HDU_INS_OUT[4] = INS_IN[4];
  assign HDU_INS_OUT[3] = INS_IN[3];
  assign HDU_INS_OUT[2] = INS_IN[2];
  assign HDU_INS_OUT[1] = INS_IN[1];
  assign HDU_INS_OUT[0] = INS_IN[0];
  assign HDU_PC_OUT[31] = PC_IN[31];
  assign HDU_PC_OUT[30] = PC_IN[30];
  assign HDU_PC_OUT[29] = PC_IN[29];
  assign HDU_PC_OUT[28] = PC_IN[28];
  assign HDU_PC_OUT[27] = PC_IN[27];
  assign HDU_PC_OUT[26] = PC_IN[26];
  assign HDU_PC_OUT[25] = PC_IN[25];
  assign HDU_PC_OUT[24] = PC_IN[24];
  assign HDU_PC_OUT[23] = PC_IN[23];
  assign HDU_PC_OUT[22] = PC_IN[22];
  assign HDU_PC_OUT[21] = PC_IN[21];
  assign HDU_PC_OUT[20] = PC_IN[20];
  assign HDU_PC_OUT[19] = PC_IN[19];
  assign HDU_PC_OUT[18] = PC_IN[18];
  assign HDU_PC_OUT[17] = PC_IN[17];
  assign HDU_PC_OUT[16] = PC_IN[16];
  assign HDU_PC_OUT[15] = PC_IN[15];
  assign HDU_PC_OUT[14] = PC_IN[14];
  assign HDU_PC_OUT[13] = PC_IN[13];
  assign HDU_PC_OUT[12] = PC_IN[12];
  assign HDU_PC_OUT[11] = PC_IN[11];
  assign HDU_PC_OUT[10] = PC_IN[10];
  assign HDU_PC_OUT[9] = PC_IN[9];
  assign HDU_PC_OUT[8] = PC_IN[8];
  assign HDU_PC_OUT[7] = PC_IN[7];
  assign HDU_PC_OUT[6] = PC_IN[6];
  assign HDU_PC_OUT[5] = PC_IN[5];
  assign HDU_PC_OUT[4] = PC_IN[4];
  assign HDU_PC_OUT[3] = PC_IN[3];
  assign HDU_PC_OUT[2] = PC_IN[2];
  assign HDU_PC_OUT[1] = PC_IN[1];
  assign HDU_PC_OUT[0] = PC_IN[0];

  HazardDetection_DW01_add_0 add_32 ( .A(PC_IN), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(HDU_NPC_OUT) );
  AND3_X1 U4 ( .A1(DRAM_R), .A2(n1), .A3(RST), .ZN(Bubble) );
  OAI33_X1 U5 ( .A1(n2), .A2(n3), .A3(n4), .B1(n5), .B2(n6), .B3(n9), .ZN(n1)
         );
  XOR2_X1 U6 ( .A(ADD_WR[4]), .B(ADD_RS2[4]), .Z(n9) );
  XOR2_X1 U8 ( .A(ADD_WR[2]), .B(ADD_RS2[2]), .Z(n6) );
  NAND3_X1 U9 ( .A1(n10), .A2(n12), .A3(n13), .ZN(n5) );
  XNOR2_X1 U11 ( .A(ADD_WR[0]), .B(ADD_RS2[0]), .ZN(n13) );
  XNOR2_X1 U12 ( .A(ADD_WR[1]), .B(ADD_RS2[1]), .ZN(n12) );
  XNOR2_X1 U13 ( .A(ADD_WR[3]), .B(ADD_RS2[3]), .ZN(n10) );
  XOR2_X1 U14 ( .A(ADD_WR[4]), .B(ADD_RS1[4]), .Z(n4) );
  XOR2_X1 U15 ( .A(ADD_WR[2]), .B(ADD_RS1[2]), .Z(n3) );
  NAND3_X1 U16 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n2) );
  XNOR2_X1 U17 ( .A(ADD_WR[0]), .B(ADD_RS1[0]), .ZN(n16) );
  XNOR2_X1 U18 ( .A(ADD_WR[1]), .B(ADD_RS1[1]), .ZN(n15) );
  XNOR2_X1 U19 ( .A(ADD_WR[3]), .B(ADD_RS1[3]), .ZN(n14) );
endmodule


module Datapath ( CLK, RST, INS_IN, DATA_IN, MUX_A_SEL, MUX_B_SEL, .ALU_OPC({
        \ALU_OPC[4] , \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), 
        ALU_OUTREG_EN, JUMP_TYPE, DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, RF_WE, 
        LOAD_TYPE_IN, STORE_TYPE_IN, WB_MUX_SEL, INS_OUT, IRAM_ADDR_OUT, 
        DRAM_ADDR_OUT, DATA_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble_out, 
        LOAD_TYPE_OUT, STORE_TYPE_OUT );
  input [31:0] INS_IN;
  input [31:0] DATA_IN;
  input [1:0] MUX_B_SEL;
  input [1:0] JUMP_TYPE;
  input [1:0] LOAD_TYPE_IN;
  output [31:0] INS_OUT;
  output [31:0] IRAM_ADDR_OUT;
  output [31:0] DRAM_ADDR_OUT;
  output [31:0] DATA_OUT;
  output [1:0] LOAD_TYPE_OUT;
  input CLK, RST, MUX_A_SEL, \ALU_OPC[4] , \ALU_OPC[3] , \ALU_OPC[2] ,
         \ALU_OPC[1] , \ALU_OPC[0] , ALU_OUTREG_EN, DRAM_R_IN, MEM_EN_IN,
         DRAM_W_IN, RF_WE, STORE_TYPE_IN, WB_MUX_SEL;
  output DRAM_R_OUT, DRAM_W_OUT, Bubble_out, STORE_TYPE_OUT;
  wire   n6, n7, n8, n9, n10, ZERO_FLAG_EX, RF_WE_WB, DRAM_R_MEM;
  wire   [4:0] ALU_OPC;
  wire   [31:0] PC_MEM_OUT;
  wire   [31:0] sig_HDU_INS_OUT;
  wire   [31:0] sig_HDU_PC_OUT;
  wire   [31:0] sig_HDU_NPC_OUT;
  wire   [31:0] PC_FETCH_OUT;
  wire   [31:0] NPC_FETCH_OUT;
  wire   [4:0] ADD_WR_WB;
  wire   [31:0] OP_WB;
  wire   [31:0] PC_DECODE_OUT;
  wire   [31:0] A_DECODE_OUT;
  wire   [31:0] B_DECODE_OUT;
  wire   [31:0] IMM_DECODE_OUT;
  wire   [4:0] ADD_RS1_HDU;
  wire   [4:0] ADD_RS2_HDU;
  wire   [4:0] ADD_WR_DECODE_OUT;
  wire   [4:0] ADD_RS1_DECODE_OUT;
  wire   [4:0] ADD_RS2_DECODE_OUT;
  wire   [4:0] ADD_WR_MEM;
  wire   [31:0] OP_MEM;
  wire   [1:0] PC_SEL_EX;
  wire   [31:0] NPC_ABS_EX;
  wire   [31:0] NPC_REL_EX;
  wire   [31:0] ALU_RES_EX;
  wire   [31:0] B_EX_OUT;
  wire   [4:0] ADD_WR_EX_OUT;
  wire   [31:0] DATA_MEM_OUT;
  wire   [31:0] ALU_RES_MEM;
  wire   [4:0] ADD_WR_MEM_OUT;

  Fetch FetchStage ( .CLK(CLK), .RST(RST), .ZERO_FLAG(ZERO_FLAG_EX), .PC_EXT(
        PC_MEM_OUT), .INS_IN(INS_IN), .Bubble_in(Bubble_out), .HDU_INS_IN(
        sig_HDU_INS_OUT), .HDU_PC_IN(sig_HDU_PC_OUT), .HDU_NPC_IN(
        sig_HDU_NPC_OUT), .PC_OUT(PC_FETCH_OUT), .ADDR_OUT(IRAM_ADDR_OUT), 
        .NPC_OUT(NPC_FETCH_OUT), .INS_OUT({n6, INS_OUT[30], n7, n8, n9, n10, 
        INS_OUT[25:0]}) );
  Decode DecodeStage ( .CLK(CLK), .RST(RST), .Bubble(Bubble_out), .RF_WE(
        RF_WE_WB), .ZERO_FLAG(ZERO_FLAG_EX), .PC_IN(PC_FETCH_OUT), .INS_IN({n6, 
        INS_OUT[30], n7, n8, n9, n10, INS_OUT[25:0]}), .ADD_WR(ADD_WR_WB), 
        .DATA_WR_IN(OP_WB), .PC_OUT(PC_DECODE_OUT), .A_OUT(A_DECODE_OUT), 
        .B_OUT(B_DECODE_OUT), .IMM_OUT(IMM_DECODE_OUT), .ADD_RS1_HDU(
        ADD_RS1_HDU), .ADD_RS2_HDU(ADD_RS2_HDU), .ADD_WR_OUT(ADD_WR_DECODE_OUT), .ADD_RS1_OUT(ADD_RS1_DECODE_OUT), .ADD_RS2_OUT(ADD_RS2_DECODE_OUT) );
  Execute ExecuteStage ( .CLK(CLK), .RST(RST), .MUX_A_SEL(MUX_A_SEL), 
        .MUX_B_SEL(MUX_B_SEL), .ALU_OPC({\ALU_OPC[4] , \ALU_OPC[3] , 
        \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), .ALU_OUTREG_EN(
        ALU_OUTREG_EN), .JUMP_TYPE(JUMP_TYPE), .PC_IN(PC_DECODE_OUT), .A_IN(
        A_DECODE_OUT), .B_IN(B_DECODE_OUT), .IMM_IN(IMM_DECODE_OUT), 
        .ADD_WR_IN(ADD_WR_DECODE_OUT), .ADD_RS1_IN(ADD_RS1_DECODE_OUT), 
        .ADD_RS2_IN(ADD_RS2_DECODE_OUT), .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_WB(
        ADD_WR_WB), .RF_WE_MEM(RF_WE), .RF_WE_WB(RF_WE_WB), .OP_MEM(OP_MEM), 
        .OP_WB(OP_WB), .PC_SEL(PC_SEL_EX), .ZERO_FLAG(ZERO_FLAG_EX), .NPC_ABS(
        NPC_ABS_EX), .NPC_REL(NPC_REL_EX), .ALU_RES(ALU_RES_EX), .B_OUT(
        B_EX_OUT), .ADD_WR_OUT(ADD_WR_EX_OUT) );
  ff_0 DRAM_R_ff ( .D(DRAM_R_IN), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(
        DRAM_R_MEM) );
  Memory MemoryStage ( .CLK(CLK), .RST(RST), .MEM_EN_IN(MEM_EN_IN), 
        .DRAM_R_IN(DRAM_R_MEM), .DRAM_W_IN(DRAM_W_IN), .PC_SEL(PC_SEL_EX), 
        .NPC_IN(NPC_FETCH_OUT), .NPC_ABS(NPC_ABS_EX), .NPC_REL(NPC_REL_EX), 
        .ALU_RES_IN(ALU_RES_EX), .B_IN(B_EX_OUT), .ADD_WR_IN(ADD_WR_EX_OUT), 
        .DRAM_DATA_IN(DATA_IN), .LOAD_TYPE_IN(LOAD_TYPE_IN), .STORE_TYPE_IN(
        STORE_TYPE_IN), .PC_OUT(PC_MEM_OUT), .DRAM_R_OUT(DRAM_R_OUT), 
        .DRAM_W_OUT(DRAM_W_OUT), .DRAM_ADDR_OUT(DRAM_ADDR_OUT), 
        .DRAM_DATA_OUT(DATA_OUT), .DATA_OUT(DATA_MEM_OUT), .ALU_RES_OUT(
        ALU_RES_MEM), .OP_MEM(OP_MEM), .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_OUT(
        ADD_WR_MEM_OUT), .LOAD_TYPE_OUT(LOAD_TYPE_OUT), .STORE_TYPE_OUT(
        STORE_TYPE_OUT) );
  ff_2 RF_WE_ff ( .D(RF_WE), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(RF_WE_WB) );
  Writeback WritebackStage ( .WB_MUX_SEL(WB_MUX_SEL), .DATA_IN(DATA_MEM_OUT), 
        .ALU_RES_IN(ALU_RES_MEM), .ADD_WR_IN(ADD_WR_MEM_OUT), .DATA_OUT(OP_WB), 
        .ADD_WR_OUT(ADD_WR_WB) );
  HazardDetection HDU ( .RST(RST), .ADD_RS1(ADD_RS1_HDU), .ADD_RS2(ADD_RS2_HDU), .ADD_WR(ADD_WR_DECODE_OUT), .DRAM_R(DRAM_R_IN), .INS_IN(INS_OUT), .PC_IN(
        PC_FETCH_OUT), .Bubble(Bubble_out), .HDU_INS_OUT(sig_HDU_INS_OUT), 
        .HDU_PC_OUT(sig_HDU_PC_OUT), .HDU_NPC_OUT(sig_HDU_NPC_OUT) );
  CLKBUF_X1 U2 ( .A(n7), .Z(INS_OUT[29]) );
  CLKBUF_X1 U3 ( .A(n8), .Z(INS_OUT[28]) );
  CLKBUF_X1 U4 ( .A(n10), .Z(INS_OUT[26]) );
  CLKBUF_X1 U5 ( .A(n6), .Z(INS_OUT[31]) );
  CLKBUF_X1 U6 ( .A(n9), .Z(INS_OUT[27]) );
endmodule


module hardwired_cu_NBIT32 ( MUX_A_SEL, MUX_B_SEL, .ALU_OPC({\ALU_OPC[4] , 
        \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), 
        ALU_OUTREG_EN, DRAM_R_IN, JUMP_TYPE, MEM_EN_IN, DRAM_W_IN, RF_WE, 
        LOAD_TYPE_IN, STORE_TYPE_IN, WB_MUX_SEL, INS_IN, Bubble, Clk, Rst );
  output [1:0] MUX_B_SEL;
  output [1:0] JUMP_TYPE;
  output [1:0] LOAD_TYPE_IN;
  input [31:0] INS_IN;
  input Bubble, Clk, Rst;
  output MUX_A_SEL, \ALU_OPC[4] , \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] ,
         \ALU_OPC[0] , ALU_OUTREG_EN, DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, RF_WE,
         STORE_TYPE_IN, WB_MUX_SEL;
  wire   INS_IN_31, INS_IN_30, INS_IN_29, INS_IN_28, INS_IN_27, INS_IN_26, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28;
  wire   [4:0] ALU_OPC;
  wire   [4:0] AluOP_E;
  assign MUX_A_SEL = 1'b0;
  assign MUX_B_SEL[1] = 1'b0;
  assign MUX_B_SEL[0] = 1'b0;
  assign ALU_OUTREG_EN = 1'b0;
  assign DRAM_R_IN = 1'b0;
  assign JUMP_TYPE[1] = 1'b0;
  assign JUMP_TYPE[0] = 1'b0;
  assign MEM_EN_IN = 1'b0;
  assign DRAM_W_IN = 1'b0;
  assign RF_WE = 1'b0;
  assign LOAD_TYPE_IN[1] = 1'b0;
  assign LOAD_TYPE_IN[0] = 1'b0;
  assign STORE_TYPE_IN = 1'b0;
  assign WB_MUX_SEL = 1'b0;
  assign INS_IN_31 = INS_IN[31];
  assign INS_IN_30 = INS_IN[30];
  assign INS_IN_29 = INS_IN[29];
  assign INS_IN_28 = INS_IN[28];
  assign INS_IN_27 = INS_IN[27];
  assign INS_IN_26 = INS_IN[26];

  DFFR_X1 \ALU_OPC_reg[4]  ( .D(AluOP_E[4]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[4]) );
  DFFR_X1 \ALU_OPC_reg[3]  ( .D(AluOP_E[3]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[3]) );
  DFFR_X1 \ALU_OPC_reg[2]  ( .D(AluOP_E[2]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[2]) );
  DFFR_X1 \ALU_OPC_reg[1]  ( .D(AluOP_E[1]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[1]) );
  NAND3_X1 U126 ( .A1(INS_IN[1]), .A2(n25), .A3(INS_IN[0]), .ZN(n65) );
  NAND3_X1 U127 ( .A1(n87), .A2(n64), .A3(n88), .ZN(n51) );
  XOR2_X1 U128 ( .A(n28), .B(INS_IN[1]), .Z(n91) );
  NAND3_X1 U129 ( .A1(n92), .A2(n27), .A3(INS_IN[0]), .ZN(n37) );
  NAND3_X1 U130 ( .A1(n10), .A2(n7), .A3(n33), .ZN(n103) );
  NAND3_X1 U131 ( .A1(n28), .A2(n27), .A3(n92), .ZN(n39) );
  NAND3_X1 U132 ( .A1(n110), .A2(n25), .A3(INS_IN[1]), .ZN(n38) );
  NAND3_X1 U133 ( .A1(n26), .A2(n27), .A3(n53), .ZN(n106) );
  NAND3_X1 U134 ( .A1(INS_IN[1]), .A2(n28), .A3(n92), .ZN(n43) );
  NAND3_X1 U135 ( .A1(n23), .A2(n21), .A3(n113), .ZN(n112) );
  DFFR_X2 \ALU_OPC_reg[0]  ( .D(AluOP_E[0]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[0]) );
  INV_X1 U17 ( .A(n77), .ZN(n11) );
  INV_X1 U18 ( .A(n79), .ZN(n4) );
  INV_X1 U19 ( .A(n59), .ZN(n14) );
  NAND2_X1 U20 ( .A1(n82), .A2(n66), .ZN(n73) );
  INV_X1 U21 ( .A(n82), .ZN(n5) );
  INV_X1 U22 ( .A(n66), .ZN(n2) );
  INV_X1 U23 ( .A(n51), .ZN(n17) );
  INV_X1 U24 ( .A(n34), .ZN(n13) );
  AOI21_X1 U25 ( .B1(n44), .B2(n45), .A(Bubble), .ZN(AluOP_E[3]) );
  AOI211_X1 U26 ( .C1(n14), .C2(n4), .A(n54), .B(n1), .ZN(n44) );
  AOI221_X1 U27 ( .B1(n46), .B2(n34), .C1(n35), .C2(n47), .A(n48), .ZN(n45) );
  OAI21_X1 U28 ( .B1(n49), .B2(n50), .A(n17), .ZN(n47) );
  AOI21_X1 U29 ( .B1(n71), .B2(n72), .A(Bubble), .ZN(AluOP_E[1]) );
  AOI221_X1 U30 ( .B1(n46), .B2(n34), .C1(n14), .C2(n73), .A(n32), .ZN(n72) );
  AOI221_X1 U31 ( .B1(n35), .B2(n76), .C1(n5), .C2(n77), .A(n67), .ZN(n71) );
  NAND4_X1 U32 ( .A1(n43), .A2(n37), .A3(n83), .A4(n84), .ZN(n76) );
  AOI21_X1 U33 ( .B1(n93), .B2(n94), .A(Bubble), .ZN(AluOP_E[0]) );
  NOR3_X1 U34 ( .A1(n95), .A2(n6), .A3(n96), .ZN(n94) );
  AOI221_X1 U35 ( .B1(n35), .B2(n104), .C1(n77), .C2(n4), .A(n1), .ZN(n93) );
  INV_X1 U36 ( .A(n68), .ZN(n6) );
  NOR3_X1 U37 ( .A1(n33), .A2(n99), .A3(n11), .ZN(n81) );
  NAND2_X1 U38 ( .A1(n52), .A2(n89), .ZN(n83) );
  NAND4_X1 U39 ( .A1(n37), .A2(n38), .A3(n39), .A4(n40), .ZN(n36) );
  AOI21_X1 U40 ( .B1(n41), .B2(n42), .A(n20), .ZN(n40) );
  INV_X1 U41 ( .A(n43), .ZN(n20) );
  OAI21_X1 U42 ( .B1(n52), .B2(n41), .A(n27), .ZN(n90) );
  NAND2_X1 U43 ( .A1(n70), .A2(n8), .ZN(n79) );
  NAND2_X1 U44 ( .A1(n70), .A2(n9), .ZN(n82) );
  OAI21_X1 U45 ( .B1(n100), .B2(n75), .A(n101), .ZN(n95) );
  NOR3_X1 U46 ( .A1(n102), .A2(n4), .A3(n46), .ZN(n100) );
  OAI21_X1 U47 ( .B1(n14), .B2(n57), .A(n73), .ZN(n101) );
  OAI21_X1 U48 ( .B1(n3), .B2(n60), .A(n103), .ZN(n102) );
  AND4_X1 U49 ( .A1(n70), .A2(n57), .A3(n10), .A4(n7), .ZN(n35) );
  NAND2_X1 U50 ( .A1(n75), .A2(n59), .ZN(n34) );
  AOI21_X1 U51 ( .B1(n55), .B2(n56), .A(Bubble), .ZN(AluOP_E[2]) );
  AOI211_X1 U52 ( .C1(n5), .C2(n12), .A(n67), .B(n54), .ZN(n55) );
  AOI221_X1 U53 ( .B1(n2), .B2(n57), .C1(n35), .C2(n16), .A(n58), .ZN(n56) );
  NOR3_X1 U54 ( .A1(n59), .A2(n33), .A3(n60), .ZN(n58) );
  INV_X1 U55 ( .A(n60), .ZN(n9) );
  NAND2_X1 U56 ( .A1(n9), .A2(n74), .ZN(n66) );
  NAND2_X1 U57 ( .A1(n89), .A2(n110), .ZN(n87) );
  NAND2_X1 U58 ( .A1(n89), .A2(n41), .ZN(n64) );
  INV_X1 U59 ( .A(n75), .ZN(n12) );
  AOI21_X1 U60 ( .B1(n29), .B2(n30), .A(Bubble), .ZN(AluOP_E[4]) );
  AOI211_X1 U61 ( .C1(n31), .C2(n9), .A(n2), .B(n32), .ZN(n30) );
  AOI22_X1 U62 ( .A1(n35), .A2(n36), .B1(n12), .B2(n4), .ZN(n29) );
  NOR2_X1 U63 ( .A1(n13), .A2(n33), .ZN(n31) );
  OAI221_X1 U64 ( .B1(n78), .B2(n79), .C1(n66), .C2(n11), .A(n80), .ZN(n67) );
  NOR3_X1 U65 ( .A1(n77), .A2(n57), .A3(n12), .ZN(n78) );
  NOR2_X1 U66 ( .A1(n48), .A2(n81), .ZN(n80) );
  AND3_X1 U67 ( .A1(n8), .A2(n74), .A3(n57), .ZN(n32) );
  AND3_X1 U68 ( .A1(n8), .A2(n74), .A3(n77), .ZN(n48) );
  INV_X1 U69 ( .A(n99), .ZN(n8) );
  INV_X1 U70 ( .A(n105), .ZN(n1) );
  AOI21_X1 U71 ( .B1(n57), .B2(n46), .A(n81), .ZN(n105) );
  INV_X1 U72 ( .A(n53), .ZN(n19) );
  INV_X1 U73 ( .A(n38), .ZN(n18) );
  AND2_X1 U74 ( .A1(n41), .A2(n25), .ZN(n92) );
  INV_X1 U75 ( .A(n50), .ZN(n26) );
  NOR3_X1 U76 ( .A1(n22), .A2(INS_IN[3]), .A3(n112), .ZN(n52) );
  NOR3_X1 U77 ( .A1(n22), .A2(n24), .A3(n112), .ZN(n41) );
  INV_X1 U78 ( .A(INS_IN[3]), .ZN(n24) );
  NOR3_X1 U79 ( .A1(INS_IN[3]), .A2(INS_IN[5]), .A3(n112), .ZN(n53) );
  NOR3_X1 U80 ( .A1(n28), .A2(INS_IN[1]), .A3(n25), .ZN(n89) );
  NOR4_X1 U81 ( .A1(INS_IN[7]), .A2(INS_IN[10]), .A3(INS_IN[9]), .A4(INS_IN[8]), .ZN(n113) );
  AOI221_X1 U82 ( .B1(n85), .B2(n52), .C1(n26), .C2(n86), .A(n51), .ZN(n84) );
  NOR2_X1 U83 ( .A1(INS_IN[2]), .A2(n91), .ZN(n85) );
  OAI21_X1 U84 ( .B1(n27), .B2(n19), .A(n90), .ZN(n86) );
  NAND4_X1 U85 ( .A1(n88), .A2(n43), .A3(n106), .A4(n107), .ZN(n104) );
  AOI221_X1 U86 ( .B1(n108), .B2(n52), .C1(n18), .C2(INS_IN[0]), .A(n62), .ZN(
        n107) );
  NOR2_X1 U87 ( .A1(INS_IN[2]), .A2(INS_IN[0]), .ZN(n108) );
  AOI22_X1 U88 ( .A1(n98), .A2(n77), .B1(n57), .B2(n99), .ZN(n97) );
  OAI21_X1 U89 ( .B1(INS_IN[1]), .B2(n50), .A(n65), .ZN(n42) );
  NAND4_X1 U90 ( .A1(n53), .A2(INS_IN[2]), .A3(INS_IN[0]), .A4(INS_IN[1]), 
        .ZN(n88) );
  NAND2_X1 U91 ( .A1(INS_IN[2]), .A2(n28), .ZN(n50) );
  INV_X1 U92 ( .A(INS_IN[1]), .ZN(n27) );
  AOI21_X1 U93 ( .B1(n52), .B2(INS_IN[1]), .A(n53), .ZN(n49) );
  NAND4_X1 U94 ( .A1(n109), .A2(n83), .A3(n87), .A4(n39), .ZN(n62) );
  NAND4_X1 U95 ( .A1(INS_IN[3]), .A2(n22), .A3(INS_IN[1]), .A4(n111), .ZN(n109) );
  NOR2_X1 U96 ( .A1(n112), .A2(n50), .ZN(n111) );
  INV_X1 U97 ( .A(INS_IN[0]), .ZN(n28) );
  NAND2_X1 U98 ( .A1(n68), .A2(n69), .ZN(n54) );
  INV_X1 U99 ( .A(INS_IN[5]), .ZN(n22) );
  AND4_X1 U100 ( .A1(n113), .A2(n21), .A3(INS_IN[3]), .A4(n114), .ZN(n110) );
  NOR2_X1 U101 ( .A1(n23), .A2(n22), .ZN(n114) );
  INV_X1 U102 ( .A(INS_IN[2]), .ZN(n25) );
  INV_X1 U103 ( .A(INS_IN[4]), .ZN(n23) );
  INV_X1 U104 ( .A(INS_IN[6]), .ZN(n21) );
  INV_X1 U105 ( .A(n61), .ZN(n16) );
  AOI211_X1 U106 ( .C1(n42), .C2(n52), .A(n62), .B(n63), .ZN(n61) );
  OAI211_X1 U107 ( .C1(n38), .C2(INS_IN[0]), .A(n37), .B(n64), .ZN(n63) );
  NOR2_X1 U108 ( .A1(INS_IN_29), .A2(n10), .ZN(n98) );
  INV_X1 U109 ( .A(INS_IN_29), .ZN(n7) );
  NAND2_X1 U110 ( .A1(INS_IN_29), .A2(n10), .ZN(n60) );
  NOR3_X1 U111 ( .A1(n3), .A2(INS_IN_30), .A3(n97), .ZN(n96) );
  AND2_X1 U112 ( .A1(INS_IN_30), .A2(n3), .ZN(n74) );
  NAND2_X1 U113 ( .A1(INS_IN_27), .A2(n15), .ZN(n59) );
  NOR2_X1 U114 ( .A1(n15), .A2(INS_IN_27), .ZN(n77) );
  NAND4_X1 U115 ( .A1(n70), .A2(n57), .A3(INS_IN_28), .A4(n7), .ZN(n69) );
  NAND4_X1 U116 ( .A1(n77), .A2(n70), .A3(INS_IN_28), .A4(n7), .ZN(n68) );
  AND3_X1 U117 ( .A1(INS_IN_28), .A2(n7), .A3(n74), .ZN(n46) );
  NAND2_X1 U118 ( .A1(INS_IN_29), .A2(INS_IN_28), .ZN(n99) );
  INV_X1 U119 ( .A(INS_IN_28), .ZN(n10) );
  NOR2_X1 U120 ( .A1(INS_IN_27), .A2(INS_IN_26), .ZN(n57) );
  NAND2_X1 U121 ( .A1(INS_IN_26), .A2(INS_IN_27), .ZN(n75) );
  INV_X1 U122 ( .A(INS_IN_26), .ZN(n15) );
  NAND2_X1 U123 ( .A1(INS_IN_31), .A2(INS_IN_30), .ZN(n33) );
  NOR2_X1 U124 ( .A1(INS_IN_31), .A2(INS_IN_30), .ZN(n70) );
  INV_X1 U125 ( .A(INS_IN_31), .ZN(n3) );
endmodule


module DLX ( Clk, Rst );
  input Clk, Rst;
  wire   DRAM_R_OUT, DRAM_W_OUT, Bubble, STORE_TYPE_OUT;
  wire   [31:0] INS_IN;
  wire   [31:0] DATA_IN;
  wire   [1:0] MUX_B_SEL;
  wire   [4:0] ALU_OPC;
  wire   [1:0] JUMP_TYPE;
  wire   [1:0] LOAD_TYPE_IN;
  wire   [31:0] INST;
  wire   [31:0] IRAM_ADDR_OUT;
  wire   [31:0] DRAM_ADDR_OUT;
  wire   [31:0] DATA_OUT;
  wire   [1:0] LOAD_TYPE_OUT;

  Datapath DP ( .CLK(Clk), .RST(Rst), .INS_IN(INS_IN), .DATA_IN(DATA_IN), 
        .MUX_A_SEL(1'b0), .MUX_B_SEL({1'b0, 1'b0}), .ALU_OPC(ALU_OPC), 
        .ALU_OUTREG_EN(1'b0), .JUMP_TYPE({1'b0, 1'b0}), .DRAM_R_IN(1'b0), 
        .MEM_EN_IN(1'b0), .DRAM_W_IN(1'b0), .RF_WE(1'b0), .LOAD_TYPE_IN({1'b0, 
        1'b0}), .STORE_TYPE_IN(1'b0), .WB_MUX_SEL(1'b0), .INS_OUT(INST), 
        .IRAM_ADDR_OUT(IRAM_ADDR_OUT), .DRAM_ADDR_OUT(DRAM_ADDR_OUT), 
        .DATA_OUT(DATA_OUT), .DRAM_R_OUT(DRAM_R_OUT), .DRAM_W_OUT(DRAM_W_OUT), 
        .Bubble_out(Bubble), .LOAD_TYPE_OUT(LOAD_TYPE_OUT), .STORE_TYPE_OUT(
        STORE_TYPE_OUT) );
  hardwired_cu_NBIT32 CU ( .ALU_OPC(ALU_OPC), .INS_IN(INST), .Bubble(Bubble), 
        .Clk(Clk), .Rst(Rst) );
  IRAM IRAM_I ( .Rst(Rst), .Addr(IRAM_ADDR_OUT), .Iout(INS_IN) );
  DRAM DRAM_I ( .Clk(Clk), .Rst(Rst), .ADDR_IN(DRAM_ADDR_OUT), .DATA_IN(
        DATA_OUT), .LOAD_TYPE(LOAD_TYPE_OUT), .STORE_TYPE(STORE_TYPE_OUT), 
        .DRAM_W(DRAM_W_OUT), .DRAM_R(DRAM_R_OUT), .DATA_OUT(DATA_IN) );
endmodule

