
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type VHDLOUT_TYPE is range 0 to 5;
type aluOp is (NOP, ADDS, ADDUS, SUBS, SUBUS, MULTS, ANDS, ORS, XORS, SLLS, 
   SRLS, SRAS, BEQZS, BNEZS, SGES, SGEUS, SGTS, SGTUS, SLES, SLTS, SLTUS, SEQS,
   NEQS, LHIS);
attribute ENUM_ENCODING of aluOp : type is 
   "00000 00001 00010 00011 00100 00101 00110 00111 01000 01001 01010 01011 01100 01101 01110 01111 10000 10001 10010 10011 10100 10101 10110 10111";
   
   -- Declarations for conversion functions.
   function integer_to_unsigned(arg, size : in INTEGER) return std_logic_vector
               ;
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
               return aluOp;
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX;

package body CONV_PACK_DLX is
   
   -- integer type to std_logic_vector function
   function integer_to_unsigned(arg, size : in INTEGER) return std_logic_vector
   is 
      variable result: std_logic_vector(size-1 downto 0);
      variable temp: INTEGER;
      -- synopsys built_in SYN_INTEGER_TO_UNSIGNED
   begin
      temp := arg;
      for i in 0 to size-1 loop
         if (temp mod 2) = 1 then
            result(i) := '1';
         else
            result(i) := '0';
         end if;
         temp := temp / 2;
      end loop;
      return result;
   end;
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
   return aluOp is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "00000" => return NOP;
         when "00001" => return ADDS;
         when "00010" => return ADDUS;
         when "00011" => return SUBS;
         when "00100" => return SUBUS;
         when "00101" => return MULTS;
         when "00110" => return ANDS;
         when "00111" => return ORS;
         when "01000" => return XORS;
         when "01001" => return SLLS;
         when "01010" => return SRLS;
         when "01011" => return SRAS;
         when "01100" => return BEQZS;
         when "01101" => return BNEZS;
         when "01110" => return SGES;
         when "01111" => return SGEUS;
         when "10000" => return SGTS;
         when "10001" => return SGTUS;
         when "10010" => return SLES;
         when "10011" => return SLTS;
         when "10100" => return SLTUS;
         when "10101" => return SEQS;
         when "10110" => return NEQS;
         when "10111" => return LHIS;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "00000";
         when ADDS => return "00001";
         when ADDUS => return "00010";
         when SUBS => return "00011";
         when SUBUS => return "00100";
         when MULTS => return "00101";
         when ANDS => return "00110";
         when ORS => return "00111";
         when XORS => return "01000";
         when SLLS => return "01001";
         when SRLS => return "01010";
         when SRAS => return "01011";
         when BEQZS => return "01100";
         when BNEZS => return "01101";
         when SGES => return "01110";
         when SGEUS => return "01111";
         when SGTS => return "10000";
         when SGTUS => return "10001";
         when SLES => return "10010";
         when SLTS => return "10011";
         when SLTUS => return "10100";
         when SEQS => return "10101";
         when NEQS => return "10110";
         when LHIS => return "10111";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "00000";
      end case;
   end;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Fetch_DW01_add_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Fetch_DW01_add_1;

architecture SYN_cla of Fetch_DW01_add_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, SUM_2_port, n36, n37,
      n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52
      , n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, 
      n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111 : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U2 : AND3_X1 port map( A1 => n38, A2 => n39, A3 => n40, ZN => n1);
   U3 : AND2_X1 port map( A1 => n40, A2 => n53, ZN => n2);
   U4 : AND2_X1 port map( A1 => n40, A2 => n66, ZN => n3);
   U5 : AND2_X1 port map( A1 => n12, A2 => n25, ZN => n23);
   U6 : NOR2_X1 port map( A1 => n15, A2 => n17, ZN => n108);
   U7 : NOR2_X1 port map( A1 => n45, A2 => n47, ZN => n49);
   U8 : NOR2_X1 port map( A1 => n45, A2 => n41, ZN => n44);
   U9 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => n15);
   U10 : NOR2_X1 port map( A1 => n99, A2 => n5, ZN => n4);
   U11 : OR2_X1 port map( A1 => n97, A2 => n98, ZN => n5);
   U12 : AND2_X1 port map( A1 => n38, A2 => n40, ZN => n6);
   U13 : AND2_X1 port map( A1 => n59, A2 => n40, ZN => n7);
   U14 : OR2_X1 port map( A1 => n98, A2 => n99, ZN => n100);
   U15 : INV_X1 port map( A => n34, ZN => n33);
   U16 : INV_X1 port map( A => n97, ZN => n101);
   U17 : AND2_X1 port map( A1 => n22, A2 => n23, ZN => n8);
   U18 : AND2_X1 port map( A1 => n107, A2 => n108, ZN => n9);
   U19 : INV_X1 port map( A => n29, ZN => n31);
   U20 : INV_X1 port map( A => n22, ZN => n24);
   U21 : INV_X1 port map( A => n25, ZN => n27);
   U22 : INV_X1 port map( A => n17, ZN => n16);
   U23 : INV_X1 port map( A => n20, ZN => n18);
   U24 : INV_X1 port map( A => n107, ZN => n109);
   U25 : INV_X1 port map( A => n80, ZN => n40);
   U26 : NOR2_X1 port map( A1 => n83, A2 => n84, ZN => n82);
   U27 : NOR2_X1 port map( A1 => n85, A2 => n86, ZN => n81);
   U28 : NAND4_X1 port map( A1 => A(16), A2 => A(17), A3 => A(18), A4 => A(19),
                           ZN => n68);
   U29 : AND2_X1 port map( A1 => n4, A2 => A(13), ZN => n94);
   U30 : NOR2_X1 port map( A1 => n111, A2 => n103, ZN => n19);
   U31 : NAND4_X1 port map( A1 => A(24), A2 => A(25), A3 => A(26), A4 => A(27),
                           ZN => n47);
   U32 : NAND4_X1 port map( A1 => A(4), A2 => A(5), A3 => n90, A4 => A(7), ZN 
                           => n103);
   U33 : NAND4_X1 port map( A1 => n107, A2 => n110, A3 => n20, A4 => A(11), ZN 
                           => n98);
   U34 : INV_X1 port map( A => n105, ZN => n110);
   U35 : NAND4_X1 port map( A1 => A(14), A2 => A(15), A3 => A(3), A4 => A(7), 
                           ZN => n83);
   U36 : NOR2_X1 port map( A1 => n41, A2 => n43, ZN => n39);
   U37 : AND3_X1 port map( A1 => A(16), A2 => A(17), A3 => n40, ZN => n10);
   U38 : AND2_X1 port map( A1 => n40, A2 => A(16), ZN => n11);
   U39 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => n55);
   U40 : NOR2_X1 port map( A1 => n60, A2 => n61, ZN => n58);
   U41 : NAND2_X1 port map( A1 => A(22), A2 => A(23), ZN => n60);
   U42 : NAND2_X1 port map( A1 => n62, A2 => A(21), ZN => n61);
   U43 : NAND2_X1 port map( A1 => n102, A2 => n28, ZN => n99);
   U44 : NAND2_X1 port map( A1 => n46, A2 => A(28), ZN => n41);
   U45 : NOR2_X1 port map( A1 => n54, A2 => n55, ZN => n53);
   U46 : NAND2_X1 port map( A1 => A(25), A2 => A(24), ZN => n54);
   U47 : AND2_X1 port map( A1 => n28, A2 => n29, ZN => n12);
   U48 : NOR2_X1 port map( A1 => n67, A2 => n68, ZN => n66);
   U49 : NAND2_X1 port map( A1 => A(21), A2 => n62, ZN => n67);
   U50 : INV_X1 port map( A => n32, ZN => n29);
   U51 : INV_X1 port map( A => n104, ZN => n20);
   U52 : NAND2_X1 port map( A1 => n72, A2 => n40, ZN => n69);
   U53 : NOR2_X1 port map( A1 => n68, A2 => n73, ZN => n72);
   U54 : INV_X1 port map( A => n26, ZN => n22);
   U55 : INV_X1 port map( A => n89, ZN => n107);
   U56 : AND2_X1 port map( A1 => n10, A2 => A(18), ZN => n76);
   U57 : AND2_X1 port map( A1 => n2, A2 => A(26), ZN => n51);
   U58 : AND2_X1 port map( A1 => n3, A2 => A(22), ZN => n64);
   U59 : NAND2_X1 port map( A1 => A(14), A2 => n94, ZN => n91);
   U60 : AND2_X1 port map( A1 => n6, A2 => A(24), ZN => n13);
   U61 : INV_X1 port map( A => n26, ZN => n90);
   U62 : INV_X1 port map( A => n30, ZN => n25);
   U63 : INV_X1 port map( A => A(24), ZN => n57);
   U64 : INV_X1 port map( A => A(16), ZN => n79);
   U65 : AND2_X1 port map( A1 => n1, A2 => A(30), ZN => n14);
   U66 : INV_X1 port map( A => n71, ZN => n70);
   U67 : INV_X1 port map( A => n93, ZN => n92);
   U68 : INV_X1 port map( A => n62, ZN => n73);
   U69 : INV_X1 port map( A => A(7), ZN => n21);
   U70 : INV_X1 port map( A => A(25), ZN => n56);
   U71 : INV_X1 port map( A => A(11), ZN => n106);
   U72 : INV_X1 port map( A => A(18), ZN => n77);
   U73 : INV_X1 port map( A => A(26), ZN => n52);
   U74 : INV_X1 port map( A => A(17), ZN => n78);
   U75 : INV_X1 port map( A => A(22), ZN => n65);
   U76 : INV_X1 port map( A => A(13), ZN => n96);
   U77 : INV_X1 port map( A => A(28), ZN => n48);
   U78 : INV_X1 port map( A => A(29), ZN => n43);
   U79 : INV_X1 port map( A => A(14), ZN => n95);
   U80 : INV_X1 port map( A => A(19), ZN => n75);
   U81 : INV_X1 port map( A => A(27), ZN => n50);
   U82 : INV_X1 port map( A => A(23), ZN => n63);
   U83 : NOR2_X1 port map( A1 => n34, A2 => n42, ZN => n28);
   U84 : INV_X1 port map( A => A(2), ZN => n42);
   U85 : XNOR2_X1 port map( A => n106, B => n9, ZN => SUM_11_port);
   U86 : XNOR2_X1 port map( A => n40, B => n79, ZN => SUM_16_port);
   U87 : XNOR2_X1 port map( A => n21, B => n8, ZN => SUM_7_port);
   U88 : INV_X1 port map( A => n74, ZN => n62);
   U89 : INV_X1 port map( A => A(20), ZN => n74);
   U90 : XNOR2_X1 port map( A => n69, B => n70, ZN => SUM_21_port);
   U91 : XNOR2_X1 port map( A => n91, B => n92, ZN => SUM_15_port);
   U92 : XNOR2_X1 port map( A => n100, B => n101, ZN => SUM_12_port);
   U93 : XNOR2_X1 port map( A => n1, B => n37, ZN => SUM_30_port);
   U94 : XNOR2_X1 port map( A => n6, B => n57, ZN => SUM_24_port);
   U95 : XNOR2_X1 port map( A => n73, B => n7, ZN => SUM_20_port);
   U96 : XNOR2_X1 port map( A => n56, B => n13, ZN => SUM_25_port);
   U97 : XNOR2_X1 port map( A => n77, B => n10, ZN => SUM_18_port);
   U98 : XNOR2_X1 port map( A => n52, B => n2, ZN => SUM_26_port);
   U99 : XNOR2_X1 port map( A => n48, B => n49, ZN => SUM_28_port);
   U100 : XNOR2_X1 port map( A => n78, B => n11, ZN => SUM_17_port);
   U101 : XNOR2_X1 port map( A => n43, B => n44, ZN => SUM_29_port);
   U102 : XNOR2_X1 port map( A => n65, B => n3, ZN => SUM_22_port);
   U103 : XNOR2_X1 port map( A => n96, B => n4, ZN => SUM_13_port);
   U104 : INV_X1 port map( A => A(6), ZN => n26);
   U105 : INV_X1 port map( A => A(4), ZN => n32);
   U106 : INV_X1 port map( A => A(8), ZN => n104);
   U107 : INV_X1 port map( A => A(9), ZN => n105);
   U108 : INV_X1 port map( A => A(5), ZN => n30);
   U109 : INV_X1 port map( A => A(30), ZN => n37);
   U110 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U111 : XNOR2_X1 port map( A => SUM_2_port, B => n33, ZN => SUM_3_port);
   U112 : XNOR2_X1 port map( A => n24, B => n23, ZN => SUM_6_port);
   U113 : XNOR2_X1 port map( A => n27, B => n12, ZN => SUM_5_port);
   U114 : XNOR2_X1 port map( A => n31, B => n28, ZN => SUM_4_port);
   U115 : XNOR2_X1 port map( A => n36, B => n14, ZN => SUM_31_port);
   U116 : INV_X1 port map( A => A(15), ZN => n93);
   U117 : INV_X1 port map( A => A(31), ZN => n36);
   U118 : XNOR2_X1 port map( A => n15, B => n16, ZN => SUM_9_port);
   U119 : XNOR2_X1 port map( A => n18, B => n19, ZN => SUM_8_port);
   U120 : INV_X1 port map( A => n47, ZN => n46);
   U121 : INV_X1 port map( A => n6, ZN => n45);
   U122 : XNOR2_X1 port map( A => n50, B => n51, ZN => SUM_27_port);
   U123 : INV_X1 port map( A => n55, ZN => n38);
   U124 : XNOR2_X1 port map( A => n63, B => n64, ZN => SUM_23_port);
   U125 : INV_X1 port map( A => A(21), ZN => n71);
   U126 : INV_X1 port map( A => n68, ZN => n59);
   U127 : XNOR2_X1 port map( A => n75, B => n76, ZN => SUM_19_port);
   U128 : NAND2_X1 port map( A1 => n81, A2 => n82, ZN => n80);
   U129 : NAND3_X1 port map( A1 => A(11), A2 => A(13), A3 => A(12), ZN => n84);
   U130 : NAND3_X1 port map( A1 => A(4), A2 => A(5), A3 => A(2), ZN => n86);
   U131 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => n85);
   U132 : NOR2_X1 port map( A1 => n104, A2 => n105, ZN => n88);
   U133 : NOR2_X1 port map( A1 => n89, A2 => n26, ZN => n87);
   U134 : INV_X1 port map( A => A(10), ZN => n89);
   U135 : XNOR2_X1 port map( A => n95, B => n94, ZN => SUM_14_port);
   U136 : INV_X1 port map( A => A(12), ZN => n97);
   U137 : INV_X1 port map( A => n103, ZN => n102);
   U138 : XNOR2_X1 port map( A => n109, B => n108, ZN => SUM_10_port);
   U139 : INV_X1 port map( A => n110, ZN => n17);
   U140 : INV_X1 port map( A => n28, ZN => n111);
   U141 : INV_X1 port map( A => A(3), ZN => n34);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute_DW01_add_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Execute_DW01_add_1;

architecture SYN_rpl of Execute_DW01_add_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_3_port, SUM_4_port, SUM_5_port, SUM_6_port, 
      SUM_7_port, SUM_8_port, SUM_9_port, SUM_10_port, SUM_11_port, SUM_12_port
      , SUM_13_port, SUM_14_port, SUM_15_port, SUM_16_port, SUM_17_port, 
      SUM_18_port, SUM_19_port, SUM_20_port, SUM_21_port, SUM_22_port, 
      SUM_23_port, SUM_24_port, SUM_25_port, SUM_26_port, SUM_27_port, 
      SUM_28_port, SUM_29_port, SUM_30_port, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n54, n55, n56, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, B(1), B(0) );
   
   U1 : XNOR2_X1 port map( A => B(31), B => n57, ZN => SUM_31_port);
   U2 : NAND2_X1 port map( A1 => B(30), A2 => n56, ZN => n57);
   U3 : INV_X1 port map( A => B(2), ZN => SUM_2_port);
   U4 : XOR2_X1 port map( A => B(3), B => B(2), Z => SUM_3_port);
   U5 : XOR2_X1 port map( A => B(4), B => n30, Z => SUM_4_port);
   U6 : XOR2_X1 port map( A => B(5), B => n31, Z => SUM_5_port);
   U7 : XOR2_X1 port map( A => B(6), B => n32, Z => SUM_6_port);
   U8 : XOR2_X1 port map( A => B(7), B => n33, Z => SUM_7_port);
   U9 : XOR2_X1 port map( A => B(8), B => n34, Z => SUM_8_port);
   U10 : XOR2_X1 port map( A => B(9), B => n35, Z => SUM_9_port);
   U11 : XOR2_X1 port map( A => B(10), B => n36, Z => SUM_10_port);
   U12 : XOR2_X1 port map( A => B(11), B => n37, Z => SUM_11_port);
   U13 : XOR2_X1 port map( A => B(12), B => n38, Z => SUM_12_port);
   U14 : XOR2_X1 port map( A => B(13), B => n39, Z => SUM_13_port);
   U15 : XOR2_X1 port map( A => B(14), B => n40, Z => SUM_14_port);
   U16 : XOR2_X1 port map( A => B(15), B => n41, Z => SUM_15_port);
   U17 : XOR2_X1 port map( A => B(16), B => n42, Z => SUM_16_port);
   U18 : XOR2_X1 port map( A => B(17), B => n43, Z => SUM_17_port);
   U19 : XOR2_X1 port map( A => B(18), B => n44, Z => SUM_18_port);
   U20 : XOR2_X1 port map( A => B(19), B => n45, Z => SUM_19_port);
   U21 : XOR2_X1 port map( A => B(20), B => n46, Z => SUM_20_port);
   U22 : XOR2_X1 port map( A => B(21), B => n47, Z => SUM_21_port);
   U23 : XOR2_X1 port map( A => B(22), B => n48, Z => SUM_22_port);
   U24 : XOR2_X1 port map( A => B(23), B => n49, Z => SUM_23_port);
   U25 : XOR2_X1 port map( A => B(24), B => n50, Z => SUM_24_port);
   U26 : XOR2_X1 port map( A => B(25), B => n51, Z => SUM_25_port);
   U27 : XOR2_X1 port map( A => B(26), B => n52, Z => SUM_26_port);
   U28 : XOR2_X1 port map( A => B(27), B => n53, Z => SUM_27_port);
   U29 : XOR2_X1 port map( A => B(28), B => n54, Z => SUM_28_port);
   U30 : XOR2_X1 port map( A => B(29), B => n55, Z => SUM_29_port);
   U31 : XOR2_X1 port map( A => B(30), B => n56, Z => SUM_30_port);
   U32 : AND2_X1 port map( A1 => B(3), A2 => B(2), ZN => n30);
   U33 : AND2_X1 port map( A1 => B(4), A2 => n30, ZN => n31);
   U34 : AND2_X1 port map( A1 => B(5), A2 => n31, ZN => n32);
   U35 : AND2_X1 port map( A1 => B(6), A2 => n32, ZN => n33);
   U36 : AND2_X1 port map( A1 => B(7), A2 => n33, ZN => n34);
   U37 : AND2_X1 port map( A1 => B(8), A2 => n34, ZN => n35);
   U38 : AND2_X1 port map( A1 => B(9), A2 => n35, ZN => n36);
   U39 : AND2_X1 port map( A1 => B(10), A2 => n36, ZN => n37);
   U40 : AND2_X1 port map( A1 => B(11), A2 => n37, ZN => n38);
   U41 : AND2_X1 port map( A1 => B(12), A2 => n38, ZN => n39);
   U42 : AND2_X1 port map( A1 => B(13), A2 => n39, ZN => n40);
   U43 : AND2_X1 port map( A1 => B(14), A2 => n40, ZN => n41);
   U44 : AND2_X1 port map( A1 => B(15), A2 => n41, ZN => n42);
   U45 : AND2_X1 port map( A1 => B(16), A2 => n42, ZN => n43);
   U46 : AND2_X1 port map( A1 => B(17), A2 => n43, ZN => n44);
   U47 : AND2_X1 port map( A1 => B(18), A2 => n44, ZN => n45);
   U48 : AND2_X1 port map( A1 => B(19), A2 => n45, ZN => n46);
   U49 : AND2_X1 port map( A1 => B(20), A2 => n46, ZN => n47);
   U50 : AND2_X1 port map( A1 => B(21), A2 => n47, ZN => n48);
   U51 : AND2_X1 port map( A1 => B(22), A2 => n48, ZN => n49);
   U52 : AND2_X1 port map( A1 => B(23), A2 => n49, ZN => n50);
   U53 : AND2_X1 port map( A1 => B(24), A2 => n50, ZN => n51);
   U54 : AND2_X1 port map( A1 => B(25), A2 => n51, ZN => n52);
   U55 : AND2_X1 port map( A1 => B(26), A2 => n52, ZN => n53);
   U56 : AND2_X1 port map( A1 => B(27), A2 => n53, ZN => n54);
   U57 : AND2_X1 port map( A1 => B(28), A2 => n54, ZN => n55);
   U58 : AND2_X1 port map( A1 => B(29), A2 => n55, ZN => n56);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Execute_DW01_add_0;

architecture SYN_rpl of Execute_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n2, n_1070 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1070, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n2, CO => carry_2_port, S
                           => SUM(1));
   U1 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U2 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n2);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity comparator_NBIT32_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end comparator_NBIT32_DW01_cmp6_0;

architecture SYN_rpl of comparator_NBIT32_DW01_cmp6_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal GT_port, GE_port, NE_port, LE_port, n3, n5, n6, n7, n8, n9, n10, n11,
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55
      , n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, 
      n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84
      , n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, 
      n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202 : std_logic;

begin
   GT <= GT_port;
   LE <= LE_port;
   GE <= GE_port;
   NE <= NE_port;
   
   U1 : INV_X1 port map( A => NE_port, ZN => EQ);
   U2 : INV_X1 port map( A => n142, ZN => n55);
   U3 : INV_X1 port map( A => n130, ZN => n7);
   U4 : INV_X1 port map( A => n118, ZN => n15);
   U5 : INV_X1 port map( A => n106, ZN => n23);
   U6 : INV_X1 port map( A => n94, ZN => n31);
   U7 : INV_X1 port map( A => n82, ZN => n39);
   U8 : INV_X1 port map( A => n139, ZN => n58);
   U9 : INV_X1 port map( A => n127, ZN => n10);
   U10 : INV_X1 port map( A => n115, ZN => n18);
   U11 : INV_X1 port map( A => n103, ZN => n26);
   U12 : INV_X1 port map( A => n91, ZN => n34);
   U13 : INV_X1 port map( A => n79, ZN => n42);
   U14 : INV_X1 port map( A => GT_port, ZN => LE_port);
   U15 : INV_X1 port map( A => n132, ZN => n61);
   U16 : INV_X1 port map( A => n141, ZN => n56);
   U17 : INV_X1 port map( A => n144, ZN => n53);
   U18 : INV_X1 port map( A => n120, ZN => n13);
   U19 : INV_X1 port map( A => n108, ZN => n21);
   U20 : INV_X1 port map( A => n96, ZN => n29);
   U21 : INV_X1 port map( A => n84, ZN => n37);
   U22 : INV_X1 port map( A => n129, ZN => n8);
   U23 : INV_X1 port map( A => n117, ZN => n16);
   U24 : INV_X1 port map( A => n105, ZN => n24);
   U25 : INV_X1 port map( A => n93, ZN => n32);
   U26 : INV_X1 port map( A => n81, ZN => n40);
   U27 : INV_X1 port map( A => n154, ZN => n47);
   U28 : INV_X1 port map( A => n68, ZN => n5);
   U29 : INV_X1 port map( A => A(30), ZN => n49);
   U30 : INV_X1 port map( A => n72, ZN => n45);
   U31 : INV_X1 port map( A => n151, ZN => n50);
   U32 : INV_X1 port map( A => B(30), ZN => n64);
   U33 : INV_X1 port map( A => n202, ZN => n3);
   U34 : INV_X1 port map( A => B(1), ZN => n63);
   U35 : INV_X1 port map( A => A(0), ZN => n6);
   U36 : INV_X1 port map( A => A(3), ZN => n51);
   U37 : INV_X1 port map( A => A(5), ZN => n54);
   U38 : INV_X1 port map( A => A(7), ZN => n59);
   U39 : INV_X1 port map( A => A(9), ZN => n62);
   U40 : INV_X1 port map( A => A(11), ZN => n11);
   U41 : INV_X1 port map( A => A(13), ZN => n14);
   U42 : INV_X1 port map( A => A(15), ZN => n19);
   U43 : INV_X1 port map( A => B(31), ZN => n65);
   U44 : INV_X1 port map( A => A(17), ZN => n22);
   U45 : INV_X1 port map( A => A(19), ZN => n27);
   U46 : INV_X1 port map( A => A(21), ZN => n30);
   U47 : INV_X1 port map( A => A(23), ZN => n35);
   U48 : INV_X1 port map( A => A(25), ZN => n38);
   U49 : INV_X1 port map( A => A(27), ZN => n43);
   U50 : INV_X1 port map( A => A(29), ZN => n46);
   U51 : INV_X1 port map( A => A(4), ZN => n52);
   U52 : INV_X1 port map( A => A(8), ZN => n60);
   U53 : INV_X1 port map( A => A(12), ZN => n12);
   U54 : INV_X1 port map( A => A(2), ZN => n48);
   U55 : INV_X1 port map( A => A(6), ZN => n57);
   U56 : INV_X1 port map( A => A(10), ZN => n9);
   U57 : INV_X1 port map( A => A(14), ZN => n17);
   U58 : INV_X1 port map( A => A(16), ZN => n20);
   U59 : INV_X1 port map( A => A(20), ZN => n28);
   U60 : INV_X1 port map( A => A(24), ZN => n36);
   U61 : INV_X1 port map( A => A(28), ZN => n44);
   U62 : INV_X1 port map( A => A(18), ZN => n25);
   U63 : INV_X1 port map( A => A(22), ZN => n33);
   U64 : INV_X1 port map( A => A(26), ZN => n41);
   U65 : INV_X1 port map( A => GE_port, ZN => LT);
   U66 : NAND2_X1 port map( A1 => LE_port, A2 => GE_port, ZN => NE_port);
   U67 : AOI21_X1 port map( B1 => n66, B2 => n5, A => n67, ZN => GE_port);
   U68 : AOI22_X1 port map( A1 => B(30), A2 => n49, B1 => n69, B2 => n70, ZN =>
                           n68);
   U69 : AOI21_X1 port map( B1 => n71, B2 => n72, A => n73, ZN => n69);
   U70 : AOI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => n71);
   U71 : AOI21_X1 port map( B1 => n77, B2 => n78, A => n79, ZN => n74);
   U72 : AOI21_X1 port map( B1 => n80, B2 => n39, A => n40, ZN => n77);
   U73 : AOI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n80);
   U74 : AOI21_X1 port map( B1 => n86, B2 => n87, A => n88, ZN => n83);
   U75 : AOI21_X1 port map( B1 => n89, B2 => n90, A => n91, ZN => n86);
   U76 : AOI21_X1 port map( B1 => n92, B2 => n31, A => n32, ZN => n89);
   U77 : AOI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n92);
   U78 : AOI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => n95);
   U79 : AOI21_X1 port map( B1 => n101, B2 => n102, A => n103, ZN => n98);
   U80 : AOI21_X1 port map( B1 => n104, B2 => n23, A => n24, ZN => n101);
   U81 : AOI21_X1 port map( B1 => n107, B2 => n108, A => n109, ZN => n104);
   U82 : AOI21_X1 port map( B1 => n110, B2 => n111, A => n112, ZN => n107);
   U83 : AOI21_X1 port map( B1 => n113, B2 => n114, A => n115, ZN => n110);
   U84 : AOI21_X1 port map( B1 => n116, B2 => n15, A => n16, ZN => n113);
   U85 : AOI21_X1 port map( B1 => n119, B2 => n120, A => n121, ZN => n116);
   U86 : AOI21_X1 port map( B1 => n122, B2 => n123, A => n124, ZN => n119);
   U87 : AOI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n122);
   U88 : AOI21_X1 port map( B1 => n128, B2 => n7, A => n8, ZN => n125);
   U89 : AOI21_X1 port map( B1 => n131, B2 => n132, A => n133, ZN => n128);
   U90 : AOI21_X1 port map( B1 => n134, B2 => n135, A => n136, ZN => n131);
   U91 : AOI21_X1 port map( B1 => n137, B2 => n138, A => n139, ZN => n134);
   U92 : AOI21_X1 port map( B1 => n140, B2 => n55, A => n56, ZN => n137);
   U93 : AOI21_X1 port map( B1 => n143, B2 => n144, A => n145, ZN => n140);
   U94 : AOI21_X1 port map( B1 => n146, B2 => n147, A => n148, ZN => n143);
   U95 : AOI21_X1 port map( B1 => n149, B2 => n150, A => n151, ZN => n146);
   U96 : AOI21_X1 port map( B1 => n152, B2 => n153, A => n47, ZN => n149);
   U97 : AOI22_X1 port map( A1 => n155, A2 => n63, B1 => A(1), B2 => n156, ZN 
                           => n152);
   U98 : OR2_X1 port map( A1 => n156, A2 => A(1), ZN => n155);
   U99 : NAND2_X1 port map( A1 => B(0), A2 => n6, ZN => n156);
   U100 : OAI21_X1 port map( B1 => n67, B2 => n157, A => n66, ZN => GT_port);
   U101 : NAND2_X1 port map( A1 => A(31), A2 => n65, ZN => n66);
   U102 : AOI22_X1 port map( A1 => A(30), A2 => n64, B1 => n158, B2 => n70, ZN 
                           => n157);
   U103 : XOR2_X1 port map( A => A(30), B => n64, Z => n70);
   U104 : AOI21_X1 port map( B1 => n159, B2 => n160, A => n45, ZN => n158);
   U105 : NAND2_X1 port map( A1 => B(29), A2 => n46, ZN => n72);
   U106 : OAI211_X1 port map( C1 => n161, C2 => n162, A => n78, B => n75, ZN =>
                           n160);
   U107 : NOR2_X1 port map( A1 => n163, A2 => n76, ZN => n75);
   U108 : AND2_X1 port map( A1 => B(28), A2 => n44, ZN => n76);
   U109 : NAND2_X1 port map( A1 => B(27), A2 => n43, ZN => n78);
   U110 : NAND2_X1 port map( A1 => n42, A2 => n164, ZN => n162);
   U111 : NOR2_X1 port map( A1 => n43, A2 => B(27), ZN => n79);
   U112 : AOI211_X1 port map( C1 => n165, C2 => n166, A => n82, B => n37, ZN =>
                           n161);
   U113 : NAND2_X1 port map( A1 => B(25), A2 => n38, ZN => n84);
   U114 : NAND2_X1 port map( A1 => n164, A2 => n81, ZN => n82);
   U115 : NAND2_X1 port map( A1 => B(26), A2 => n41, ZN => n81);
   U116 : OR2_X1 port map( A1 => n41, A2 => B(26), ZN => n164);
   U117 : OAI211_X1 port map( C1 => n167, C2 => n168, A => n90, B => n87, ZN =>
                           n166);
   U118 : NOR2_X1 port map( A1 => n169, A2 => n88, ZN => n87);
   U119 : AND2_X1 port map( A1 => B(24), A2 => n36, ZN => n88);
   U120 : NAND2_X1 port map( A1 => B(23), A2 => n35, ZN => n90);
   U121 : NAND2_X1 port map( A1 => n34, A2 => n170, ZN => n168);
   U122 : NOR2_X1 port map( A1 => n35, A2 => B(23), ZN => n91);
   U123 : AOI211_X1 port map( C1 => n171, C2 => n172, A => n94, B => n29, ZN =>
                           n167);
   U124 : NAND2_X1 port map( A1 => B(21), A2 => n30, ZN => n96);
   U125 : NAND2_X1 port map( A1 => n170, A2 => n93, ZN => n94);
   U126 : NAND2_X1 port map( A1 => B(22), A2 => n33, ZN => n93);
   U127 : OR2_X1 port map( A1 => n33, A2 => B(22), ZN => n170);
   U128 : OAI211_X1 port map( C1 => n173, C2 => n174, A => n102, B => n99, ZN 
                           => n172);
   U129 : NOR2_X1 port map( A1 => n175, A2 => n100, ZN => n99);
   U130 : AND2_X1 port map( A1 => B(20), A2 => n28, ZN => n100);
   U131 : NAND2_X1 port map( A1 => B(19), A2 => n27, ZN => n102);
   U132 : NAND2_X1 port map( A1 => n26, A2 => n176, ZN => n174);
   U133 : NOR2_X1 port map( A1 => n27, A2 => B(19), ZN => n103);
   U134 : AOI211_X1 port map( C1 => n177, C2 => n178, A => n106, B => n21, ZN 
                           => n173);
   U135 : NAND2_X1 port map( A1 => B(17), A2 => n22, ZN => n108);
   U136 : NAND2_X1 port map( A1 => n176, A2 => n105, ZN => n106);
   U137 : NAND2_X1 port map( A1 => B(18), A2 => n25, ZN => n105);
   U138 : OR2_X1 port map( A1 => n25, A2 => B(18), ZN => n176);
   U139 : OAI211_X1 port map( C1 => n179, C2 => n180, A => n114, B => n111, ZN 
                           => n178);
   U140 : NOR2_X1 port map( A1 => n181, A2 => n112, ZN => n111);
   U141 : AND2_X1 port map( A1 => B(16), A2 => n20, ZN => n112);
   U142 : NAND2_X1 port map( A1 => B(15), A2 => n19, ZN => n114);
   U143 : NAND2_X1 port map( A1 => n18, A2 => n182, ZN => n180);
   U144 : NOR2_X1 port map( A1 => n19, A2 => B(15), ZN => n115);
   U145 : AOI211_X1 port map( C1 => n183, C2 => n184, A => n118, B => n13, ZN 
                           => n179);
   U146 : NAND2_X1 port map( A1 => B(13), A2 => n14, ZN => n120);
   U147 : NAND2_X1 port map( A1 => n182, A2 => n117, ZN => n118);
   U148 : NAND2_X1 port map( A1 => B(14), A2 => n17, ZN => n117);
   U149 : OR2_X1 port map( A1 => n17, A2 => B(14), ZN => n182);
   U150 : OAI211_X1 port map( C1 => n185, C2 => n186, A => n126, B => n123, ZN 
                           => n184);
   U151 : NOR2_X1 port map( A1 => n187, A2 => n124, ZN => n123);
   U152 : AND2_X1 port map( A1 => B(12), A2 => n12, ZN => n124);
   U153 : NAND2_X1 port map( A1 => B(11), A2 => n11, ZN => n126);
   U154 : NAND2_X1 port map( A1 => n10, A2 => n188, ZN => n186);
   U155 : NOR2_X1 port map( A1 => n11, A2 => B(11), ZN => n127);
   U156 : AOI211_X1 port map( C1 => n189, C2 => n190, A => n130, B => n61, ZN 
                           => n185);
   U157 : NAND2_X1 port map( A1 => B(9), A2 => n62, ZN => n132);
   U158 : NAND2_X1 port map( A1 => n188, A2 => n129, ZN => n130);
   U159 : NAND2_X1 port map( A1 => B(10), A2 => n9, ZN => n129);
   U160 : OR2_X1 port map( A1 => n9, A2 => B(10), ZN => n188);
   U161 : OAI211_X1 port map( C1 => n191, C2 => n192, A => n138, B => n135, ZN 
                           => n190);
   U162 : NOR2_X1 port map( A1 => n193, A2 => n136, ZN => n135);
   U163 : AND2_X1 port map( A1 => B(8), A2 => n60, ZN => n136);
   U164 : NAND2_X1 port map( A1 => B(7), A2 => n59, ZN => n138);
   U165 : NAND2_X1 port map( A1 => n58, A2 => n194, ZN => n192);
   U166 : NOR2_X1 port map( A1 => n59, A2 => B(7), ZN => n139);
   U167 : AOI211_X1 port map( C1 => n195, C2 => n196, A => n142, B => n53, ZN 
                           => n191);
   U168 : NAND2_X1 port map( A1 => B(5), A2 => n54, ZN => n144);
   U169 : NAND2_X1 port map( A1 => n194, A2 => n141, ZN => n142);
   U170 : NAND2_X1 port map( A1 => B(6), A2 => n57, ZN => n141);
   U171 : OR2_X1 port map( A1 => n57, A2 => B(6), ZN => n194);
   U172 : NAND3_X1 port map( A1 => n197, A2 => n150, A3 => n147, ZN => n196);
   U173 : NOR2_X1 port map( A1 => n198, A2 => n148, ZN => n147);
   U174 : AND2_X1 port map( A1 => B(4), A2 => n52, ZN => n148);
   U175 : NAND2_X1 port map( A1 => B(3), A2 => n51, ZN => n150);
   U176 : NAND3_X1 port map( A1 => n50, A2 => n199, A3 => n200, ZN => n197);
   U177 : OAI211_X1 port map( C1 => A(1), C2 => n201, A => n3, B => n153, ZN =>
                           n200);
   U178 : AND2_X1 port map( A1 => n199, A2 => n154, ZN => n153);
   U179 : NAND2_X1 port map( A1 => B(2), A2 => n48, ZN => n154);
   U180 : AOI21_X1 port map( B1 => A(1), B2 => n201, A => n63, ZN => n202);
   U181 : NOR2_X1 port map( A1 => n6, A2 => B(0), ZN => n201);
   U182 : OR2_X1 port map( A1 => n48, A2 => B(2), ZN => n199);
   U183 : NOR2_X1 port map( A1 => n51, A2 => B(3), ZN => n151);
   U184 : NOR2_X1 port map( A1 => n198, A2 => n145, ZN => n195);
   U185 : NOR2_X1 port map( A1 => n54, A2 => B(5), ZN => n145);
   U186 : NOR2_X1 port map( A1 => n52, A2 => B(4), ZN => n198);
   U187 : NOR2_X1 port map( A1 => n193, A2 => n133, ZN => n189);
   U188 : NOR2_X1 port map( A1 => n62, A2 => B(9), ZN => n133);
   U189 : NOR2_X1 port map( A1 => n60, A2 => B(8), ZN => n193);
   U190 : NOR2_X1 port map( A1 => n187, A2 => n121, ZN => n183);
   U191 : NOR2_X1 port map( A1 => n14, A2 => B(13), ZN => n121);
   U192 : NOR2_X1 port map( A1 => n12, A2 => B(12), ZN => n187);
   U193 : NOR2_X1 port map( A1 => n181, A2 => n109, ZN => n177);
   U194 : NOR2_X1 port map( A1 => n22, A2 => B(17), ZN => n109);
   U195 : NOR2_X1 port map( A1 => n20, A2 => B(16), ZN => n181);
   U196 : NOR2_X1 port map( A1 => n175, A2 => n97, ZN => n171);
   U197 : NOR2_X1 port map( A1 => n30, A2 => B(21), ZN => n97);
   U198 : NOR2_X1 port map( A1 => n28, A2 => B(20), ZN => n175);
   U199 : NOR2_X1 port map( A1 => n169, A2 => n85, ZN => n165);
   U200 : NOR2_X1 port map( A1 => n38, A2 => B(25), ZN => n85);
   U201 : NOR2_X1 port map( A1 => n36, A2 => B(24), ZN => n169);
   U202 : NOR2_X1 port map( A1 => n163, A2 => n73, ZN => n159);
   U203 : NOR2_X1 port map( A1 => n46, A2 => B(29), ZN => n73);
   U204 : NOR2_X1 port map( A1 => n44, A2 => B(28), ZN => n163);
   U205 : NOR2_X1 port map( A1 => n65, A2 => A(31), ZN => n67);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_0_DW01_add_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end rca_bhv_numBit32_0_DW01_add_0;

architecture SYN_rpl of rca_bhv_numBit32_0_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1075 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1075, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_6_DW01_add_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end rca_bhv_numBit32_6_DW01_add_0;

architecture SYN_rpl of rca_bhv_numBit32_6_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1079 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1079, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_5_DW01_add_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end rca_bhv_numBit32_5_DW01_add_0;

architecture SYN_rpl of rca_bhv_numBit32_5_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1083 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1083, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_4_DW01_add_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end rca_bhv_numBit32_4_DW01_add_0;

architecture SYN_rpl of rca_bhv_numBit32_4_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1087 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1087, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_3_DW01_add_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end rca_bhv_numBit32_3_DW01_add_0;

architecture SYN_rpl of rca_bhv_numBit32_3_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1091 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1091, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_2_DW01_add_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end rca_bhv_numBit32_2_DW01_add_0;

architecture SYN_rpl of rca_bhv_numBit32_2_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1095 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1095, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_1_DW01_add_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end rca_bhv_numBit32_1_DW01_add_0;

architecture SYN_rpl of rca_bhv_numBit32_1_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1099 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1099, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HazardDetection_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end HazardDetection_DW01_add_0;

architecture SYN_rpl of HazardDetection_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_30_port, SUM_9_port, SUM_8_port, SUM_10_port, 
      SUM_11_port, SUM_12_port, SUM_13_port, SUM_14_port, SUM_15_port, 
      SUM_16_port, SUM_17_port, SUM_18_port, SUM_19_port, SUM_20_port, 
      SUM_21_port, SUM_22_port, SUM_23_port, SUM_24_port, SUM_25_port, 
      SUM_26_port, SUM_27_port, SUM_28_port, SUM_29_port, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49, n50, n51, SUM_3_port, SUM_4_port, 
      SUM_5_port, SUM_6_port, SUM_7_port, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U1 : XNOR2_X1 port map( A => A(31), B => n57, ZN => SUM_31_port);
   U2 : XOR2_X1 port map( A => A(30), B => n51, Z => SUM_30_port);
   U3 : XOR2_X1 port map( A => A(9), B => n31, Z => SUM_9_port);
   U4 : XOR2_X1 port map( A => A(8), B => n30, Z => SUM_8_port);
   U5 : XOR2_X1 port map( A => A(10), B => n25, Z => SUM_10_port);
   U6 : XOR2_X1 port map( A => A(11), B => n32, Z => SUM_11_port);
   U7 : XOR2_X1 port map( A => A(12), B => n33, Z => SUM_12_port);
   U8 : XOR2_X1 port map( A => A(13), B => n34, Z => SUM_13_port);
   U9 : XOR2_X1 port map( A => A(14), B => n35, Z => SUM_14_port);
   U10 : XOR2_X1 port map( A => A(15), B => n36, Z => SUM_15_port);
   U11 : XOR2_X1 port map( A => A(16), B => n37, Z => SUM_16_port);
   U12 : XOR2_X1 port map( A => A(17), B => n38, Z => SUM_17_port);
   U13 : XOR2_X1 port map( A => A(18), B => n39, Z => SUM_18_port);
   U14 : XOR2_X1 port map( A => A(19), B => n40, Z => SUM_19_port);
   U15 : XOR2_X1 port map( A => A(20), B => n41, Z => SUM_20_port);
   U16 : XOR2_X1 port map( A => A(21), B => n42, Z => SUM_21_port);
   U17 : XOR2_X1 port map( A => A(22), B => n43, Z => SUM_22_port);
   U18 : XOR2_X1 port map( A => A(23), B => n44, Z => SUM_23_port);
   U19 : XOR2_X1 port map( A => A(24), B => n45, Z => SUM_24_port);
   U20 : XOR2_X1 port map( A => A(25), B => n46, Z => SUM_25_port);
   U21 : XOR2_X1 port map( A => A(26), B => n47, Z => SUM_26_port);
   U22 : XOR2_X1 port map( A => A(27), B => n48, Z => SUM_27_port);
   U23 : XOR2_X1 port map( A => A(28), B => n49, Z => SUM_28_port);
   U24 : XOR2_X1 port map( A => A(29), B => n50, Z => SUM_29_port);
   U25 : NAND2_X1 port map( A1 => A(30), A2 => n51, ZN => n57);
   U26 : AND2_X1 port map( A1 => A(9), A2 => n31, ZN => n25);
   U27 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n26);
   U28 : AND2_X1 port map( A1 => A(4), A2 => n26, ZN => n27);
   U29 : AND2_X1 port map( A1 => A(5), A2 => n27, ZN => n28);
   U30 : AND2_X1 port map( A1 => A(6), A2 => n28, ZN => n29);
   U31 : AND2_X1 port map( A1 => A(7), A2 => n29, ZN => n30);
   U32 : AND2_X1 port map( A1 => A(8), A2 => n30, ZN => n31);
   U33 : AND2_X1 port map( A1 => A(10), A2 => n25, ZN => n32);
   U34 : AND2_X1 port map( A1 => A(11), A2 => n32, ZN => n33);
   U35 : AND2_X1 port map( A1 => A(12), A2 => n33, ZN => n34);
   U36 : AND2_X1 port map( A1 => A(13), A2 => n34, ZN => n35);
   U37 : AND2_X1 port map( A1 => A(14), A2 => n35, ZN => n36);
   U38 : AND2_X1 port map( A1 => A(15), A2 => n36, ZN => n37);
   U39 : AND2_X1 port map( A1 => A(16), A2 => n37, ZN => n38);
   U40 : AND2_X1 port map( A1 => A(17), A2 => n38, ZN => n39);
   U41 : AND2_X1 port map( A1 => A(18), A2 => n39, ZN => n40);
   U42 : AND2_X1 port map( A1 => A(19), A2 => n40, ZN => n41);
   U43 : AND2_X1 port map( A1 => A(20), A2 => n41, ZN => n42);
   U44 : AND2_X1 port map( A1 => A(21), A2 => n42, ZN => n43);
   U45 : AND2_X1 port map( A1 => A(22), A2 => n43, ZN => n44);
   U46 : AND2_X1 port map( A1 => A(23), A2 => n44, ZN => n45);
   U47 : AND2_X1 port map( A1 => A(24), A2 => n45, ZN => n46);
   U48 : AND2_X1 port map( A1 => A(25), A2 => n46, ZN => n47);
   U49 : AND2_X1 port map( A1 => A(26), A2 => n47, ZN => n48);
   U50 : AND2_X1 port map( A1 => A(27), A2 => n48, ZN => n49);
   U51 : AND2_X1 port map( A1 => A(28), A2 => n49, ZN => n50);
   U52 : AND2_X1 port map( A1 => A(29), A2 => n50, ZN => n51);
   U53 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U54 : XOR2_X1 port map( A => A(3), B => A(2), Z => SUM_3_port);
   U55 : XOR2_X1 port map( A => A(4), B => n26, Z => SUM_4_port);
   U56 : XOR2_X1 port map( A => A(5), B => n27, Z => SUM_5_port);
   U57 : XOR2_X1 port map( A => A(6), B => n28, Z => SUM_6_port);
   U58 : XOR2_X1 port map( A => A(7), B => n29, Z => SUM_7_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_15;

architecture SYN_STRUCTURAL of RCA_N4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_14;

architecture SYN_STRUCTURAL of RCA_N4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_13;

architecture SYN_STRUCTURAL of RCA_N4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_12;

architecture SYN_STRUCTURAL of RCA_N4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_11;

architecture SYN_STRUCTURAL of RCA_N4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_10;

architecture SYN_STRUCTURAL of RCA_N4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_9;

architecture SYN_STRUCTURAL of RCA_N4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_8;

architecture SYN_STRUCTURAL of RCA_N4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_7;

architecture SYN_STRUCTURAL of RCA_N4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_6;

architecture SYN_STRUCTURAL of RCA_N4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_5;

architecture SYN_STRUCTURAL of RCA_N4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_4;

architecture SYN_STRUCTURAL of RCA_N4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_3;

architecture SYN_STRUCTURAL of RCA_N4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_2;

architecture SYN_STRUCTURAL of RCA_N4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_1;

architecture SYN_STRUCTURAL of RCA_N4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_7;

architecture SYN_struct of carry_select_basic_N4_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1134, n_1135 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1134);
   RCA1 : RCA_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1135);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n11, ZN => S(1));
   U5 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n13, ZN => S(3));
   U9 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_6;

architecture SYN_struct of carry_select_basic_N4_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1136, n_1137 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1136);
   RCA1 : RCA_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1137);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n11, ZN => S(1));
   U5 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n13, ZN => S(3));
   U9 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_5;

architecture SYN_struct of carry_select_basic_N4_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1138, n_1139 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1138);
   RCA1 : RCA_N4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1139);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n11, ZN => S(1));
   U5 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n13, ZN => S(3));
   U9 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_4;

architecture SYN_struct of carry_select_basic_N4_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1140, n_1141 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1140);
   RCA1 : RCA_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1141);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n11, ZN => S(1));
   U5 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n13, ZN => S(3));
   U9 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_3;

architecture SYN_struct of carry_select_basic_N4_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1142, n_1143 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1142);
   RCA1 : RCA_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1143);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n11, ZN => S(1));
   U5 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n13, ZN => S(3));
   U9 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_2;

architecture SYN_struct of carry_select_basic_N4_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1144, n_1145 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1144);
   RCA1 : RCA_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1145);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n11, ZN => S(1));
   U5 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n13, ZN => S(3));
   U9 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_1;

architecture SYN_struct of carry_select_basic_N4_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1146, n_1147 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1146);
   RCA1 : RCA_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1147);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n11, ZN => S(1));
   U7 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U8 : INV_X1 port map( A => n12, ZN => S(2));
   U9 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_26 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_26;

architecture SYN_bhv of PGblock_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_25 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_25;

architecture SYN_bhv of PGblock_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_24 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_24;

architecture SYN_bhv of PGblock_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_23 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_23;

architecture SYN_bhv of PGblock_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_22 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_22;

architecture SYN_bhv of PGblock_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_21 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_21;

architecture SYN_bhv of PGblock_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_20 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_20;

architecture SYN_bhv of PGblock_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_19 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_19;

architecture SYN_bhv of PGblock_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_18 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_18;

architecture SYN_bhv of PGblock_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_17 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_17;

architecture SYN_bhv of PGblock_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_16 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_16;

architecture SYN_bhv of PGblock_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_15 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_15;

architecture SYN_bhv of PGblock_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_14 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_14;

architecture SYN_bhv of PGblock_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_13 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_13;

architecture SYN_bhv of PGblock_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_12 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_12;

architecture SYN_bhv of PGblock_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_11 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_11;

architecture SYN_bhv of PGblock_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_10 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_10;

architecture SYN_bhv of PGblock_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_9 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_9;

architecture SYN_bhv of PGblock_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_8 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_8;

architecture SYN_bhv of PGblock_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_7 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_7;

architecture SYN_bhv of PGblock_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_6 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_6;

architecture SYN_bhv of PGblock_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_5 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_5;

architecture SYN_bhv of PGblock_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_4 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_4;

architecture SYN_bhv of PGblock_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_3 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_3;

architecture SYN_bhv of PGblock_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_2 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_2;

architecture SYN_bhv of PGblock_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_1 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_1;

architecture SYN_bhv of PGblock_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_8 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_8;

architecture SYN_bhv of Gblock_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_7 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_7;

architecture SYN_bhv of Gblock_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_6 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_6;

architecture SYN_bhv of Gblock_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_5 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_5;

architecture SYN_bhv of Gblock_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_4 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_4;

architecture SYN_bhv of Gblock_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_3 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_3;

architecture SYN_bhv of Gblock_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_2 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_2;

architecture SYN_bhv of Gblock_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_1 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_1;

architecture SYN_bhv of Gblock_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_30 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_30;

architecture SYN_bhv of PG_net_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_29 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_29;

architecture SYN_bhv of PG_net_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_28 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_28;

architecture SYN_bhv of PG_net_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_27 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_27;

architecture SYN_bhv of PG_net_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_26 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_26;

architecture SYN_bhv of PG_net_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_25 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_25;

architecture SYN_bhv of PG_net_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_24 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_24;

architecture SYN_bhv of PG_net_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_23 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_23;

architecture SYN_bhv of PG_net_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_22 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_22;

architecture SYN_bhv of PG_net_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_21 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_21;

architecture SYN_bhv of PG_net_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_20 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_20;

architecture SYN_bhv of PG_net_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_19 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_19;

architecture SYN_bhv of PG_net_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_18 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_18;

architecture SYN_bhv of PG_net_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_17 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_17;

architecture SYN_bhv of PG_net_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_16 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_16;

architecture SYN_bhv of PG_net_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_15 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_15;

architecture SYN_bhv of PG_net_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_14 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_14;

architecture SYN_bhv of PG_net_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_13 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_13;

architecture SYN_bhv of PG_net_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_12 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_12;

architecture SYN_bhv of PG_net_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_11 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_11;

architecture SYN_bhv of PG_net_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_10 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_10;

architecture SYN_bhv of PG_net_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_9 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_9;

architecture SYN_bhv of PG_net_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_8 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_8;

architecture SYN_bhv of PG_net_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_7 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_7;

architecture SYN_bhv of PG_net_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_6 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_6;

architecture SYN_bhv of PG_net_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_5 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_5;

architecture SYN_bhv of PG_net_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_4 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_4;

architecture SYN_bhv of PG_net_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_3 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_3;

architecture SYN_bhv of PG_net_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_2 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_2;

architecture SYN_bhv of PG_net_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_1 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_1;

architecture SYN_bhv of PG_net_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_6 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end rca_bhv_numBit32_6;

architecture SYN_BEHAVIORAL of rca_bhv_numBit32_6 is

   component rca_bhv_numBit32_6_DW01_add_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   signal n_1148 : std_logic;

begin
   
   add_1_root_add_35_2 : rca_bhv_numBit32_6_DW01_add_0 port map( A(32) => A(31)
                           , A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(32) => Co, SUM(31)
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1148);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end rca_bhv_numBit32_5;

architecture SYN_BEHAVIORAL of rca_bhv_numBit32_5 is

   component rca_bhv_numBit32_5_DW01_add_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   signal n_1149 : std_logic;

begin
   
   add_1_root_add_35_2 : rca_bhv_numBit32_5_DW01_add_0 port map( A(32) => A(31)
                           , A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(32) => Co, SUM(31)
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1149);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end rca_bhv_numBit32_4;

architecture SYN_BEHAVIORAL of rca_bhv_numBit32_4 is

   component rca_bhv_numBit32_4_DW01_add_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   signal n_1150 : std_logic;

begin
   
   add_1_root_add_35_2 : rca_bhv_numBit32_4_DW01_add_0 port map( A(32) => A(31)
                           , A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(32) => Co, SUM(31)
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1150);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end rca_bhv_numBit32_3;

architecture SYN_BEHAVIORAL of rca_bhv_numBit32_3 is

   component rca_bhv_numBit32_3_DW01_add_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   signal n_1151 : std_logic;

begin
   
   add_1_root_add_35_2 : rca_bhv_numBit32_3_DW01_add_0 port map( A(32) => A(31)
                           , A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(32) => Co, SUM(31)
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1151);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end rca_bhv_numBit32_2;

architecture SYN_BEHAVIORAL of rca_bhv_numBit32_2 is

   component rca_bhv_numBit32_2_DW01_add_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   signal n_1152 : std_logic;

begin
   
   add_1_root_add_35_2 : rca_bhv_numBit32_2_DW01_add_0 port map( A(32) => A(31)
                           , A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(32) => Co, SUM(31)
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1152);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end rca_bhv_numBit32_1;

architecture SYN_BEHAVIORAL of rca_bhv_numBit32_1 is

   component rca_bhv_numBit32_1_DW01_add_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   signal n_1153 : std_logic;

begin
   
   add_1_root_add_35_2 : rca_bhv_numBit32_1_DW01_add_0 port map( A(32) => A(31)
                           , A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(32) => Co, SUM(31)
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1153);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_7 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_7;

architecture SYN_bhv of mux5to1_numBit32_7 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n91, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n160);
   U2 : BUF_X1 port map( A => n158, Z => n4);
   U3 : BUF_X1 port map( A => n158, Z => n77);
   U4 : BUF_X1 port map( A => n158, Z => n78);
   U5 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84,
                           C1 => IN5(25), C2 => n81, ZN => n146);
   U6 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84,
                           C1 => IN5(26), C2 => n81, ZN => n148);
   U7 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84,
                           C1 => IN5(27), C2 => n81, ZN => n150);
   U8 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => n84,
                           C1 => IN5(28), C2 => n81, ZN => n152);
   U9 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => n84,
                           C1 => IN5(29), C2 => n81, ZN => n154);
   U10 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => n84
                           , C1 => IN5(30), C2 => n81, ZN => n156);
   U11 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n132);
   U12 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n134);
   U13 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n136);
   U14 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n138);
   U15 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n140);
   U16 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n142);
   U17 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n144);
   U18 : BUF_X1 port map( A => n89, Z => n1);
   U19 : BUF_X1 port map( A => n89, Z => n2);
   U20 : NOR2_X1 port map( A1 => n88, A2 => n93, ZN => n158);
   U21 : INV_X1 port map( A => n94, ZN => n88);
   U22 : BUF_X1 port map( A => n89, Z => n3);
   U23 : NOR4_X1 port map( A1 => n92, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n94);
   U24 : BUF_X1 port map( A => n160, Z => n82);
   U25 : BUF_X1 port map( A => n160, Z => n83);
   U26 : BUF_X1 port map( A => n159, Z => n79);
   U27 : BUF_X1 port map( A => n159, Z => n80);
   U28 : BUF_X1 port map( A => n161, Z => n85);
   U29 : BUF_X1 port map( A => n161, Z => n86);
   U30 : BUF_X1 port map( A => n160, Z => n84);
   U31 : NOR2_X1 port map( A1 => n91, A2 => n90, ZN => n93);
   U32 : BUF_X1 port map( A => n159, Z => n81);
   U33 : BUF_X1 port map( A => n161, Z => n87);
   U34 : INV_X1 port map( A => n95, ZN => n89);
   U35 : AOI21_X1 port map( B1 => n94, B2 => n93, A => n92, ZN => n95);
   U36 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82, 
                           C1 => IN5(4), C2 => n79, ZN => n104);
   U37 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82, 
                           C1 => IN5(5), C2 => n79, ZN => n106);
   U38 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82, 
                           C1 => IN5(6), C2 => n79, ZN => n108);
   U39 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82, 
                           C1 => IN5(7), C2 => n79, ZN => n110);
   U40 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82, 
                           C1 => IN5(8), C2 => n79, ZN => n112);
   U41 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82, 
                           C1 => IN5(9), C2 => n79, ZN => n114);
   U42 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => n82
                           , C1 => IN5(10), C2 => n79, ZN => n116);
   U43 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => n82
                           , C1 => IN5(11), C2 => n79, ZN => n118);
   U44 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => n83
                           , C1 => IN5(12), C2 => n80, ZN => n120);
   U45 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => n83
                           , C1 => IN5(13), C2 => n80, ZN => n122);
   U46 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n124);
   U47 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n126);
   U48 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n128);
   U49 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n130);
   U50 : NOR3_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => n90, ZN => n161);
   U51 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n92);
   U52 : INV_X1 port map( A => SEL_in(0), ZN => n90);
   U53 : AND3_X1 port map( A1 => n90, A2 => n91, A3 => SEL_in(2), ZN => n159);
   U54 : INV_X1 port map( A => SEL_in(1), ZN => n91);
   U55 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(3));
   U56 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82, 
                           C1 => IN5(3), C2 => n79, ZN => n102);
   U57 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN 
                           => n103);
   U58 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2, 
                           ZN => n129);
   U59 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82, 
                           C1 => IN5(2), C2 => n79, ZN => n100);
   U60 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2, 
                           ZN => n131);
   U61 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2, 
                           ZN => n133);
   U62 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(4));
   U63 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN 
                           => n105);
   U64 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(5));
   U65 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN 
                           => n107);
   U66 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(6));
   U67 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN 
                           => n109);
   U68 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(7));
   U69 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN 
                           => n111);
   U70 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(8));
   U71 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN 
                           => n113);
   U72 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(9));
   U73 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN 
                           => n115);
   U74 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(10));
   U75 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n117);
   U76 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(11));
   U77 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n119);
   U78 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(12));
   U79 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2, 
                           ZN => n121);
   U80 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(13));
   U81 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2, 
                           ZN => n123);
   U82 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(14));
   U83 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n125);
   U84 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(15));
   U85 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n127);
   U86 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(16));
   U87 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(17));
   U88 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(18));
   U89 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(19));
   U90 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n135);
   U91 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(20));
   U92 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n137);
   U93 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(21));
   U94 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n139);
   U95 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(22));
   U96 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n141);
   U97 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(23));
   U98 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n143);
   U99 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Z(24));
   U100 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3,
                           ZN => n145);
   U101 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Z(25));
   U102 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3,
                           ZN => n147);
   U103 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(26));
   U104 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3,
                           ZN => n149);
   U105 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Z(27));
   U106 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3,
                           ZN => n151);
   U107 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Z(28));
   U108 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3,
                           ZN => n153);
   U110 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Z(29));
   U111 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3,
                           ZN => n155);
   U112 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => Z(30));
   U113 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3,
                           ZN => n157);
   U114 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(2));
   U115 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN
                           => n101);
   U116 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(0));
   U117 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN
                           => n97);
   U118 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(1));
   U119 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN
                           => n99);
   U120 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => Z(31));
   U121 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n163);
   U122 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => 
                           n84, C1 => IN5(31), C2 => n81, ZN => n162);
   U123 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82,
                           C1 => IN5(0), C2 => n79, ZN => n96);
   U124 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82,
                           C1 => IN5(1), C2 => n79, ZN => n98);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_6 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_6;

architecture SYN_bhv of mux5to1_numBit32_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n91, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n160);
   U2 : BUF_X1 port map( A => n158, Z => n4);
   U3 : BUF_X1 port map( A => n158, Z => n77);
   U4 : BUF_X1 port map( A => n158, Z => n78);
   U5 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => n84,
                           C1 => IN5(31), C2 => n81, ZN => n162);
   U6 : BUF_X1 port map( A => n89, Z => n1);
   U7 : BUF_X1 port map( A => n89, Z => n2);
   U8 : NOR2_X1 port map( A1 => n88, A2 => n93, ZN => n158);
   U9 : INV_X1 port map( A => n94, ZN => n88);
   U10 : BUF_X1 port map( A => n89, Z => n3);
   U11 : NOR4_X1 port map( A1 => n92, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n94);
   U12 : BUF_X1 port map( A => n160, Z => n82);
   U13 : BUF_X1 port map( A => n160, Z => n83);
   U14 : BUF_X1 port map( A => n159, Z => n79);
   U15 : BUF_X1 port map( A => n159, Z => n80);
   U16 : BUF_X1 port map( A => n161, Z => n85);
   U17 : BUF_X1 port map( A => n161, Z => n86);
   U18 : BUF_X1 port map( A => n160, Z => n84);
   U19 : NOR2_X1 port map( A1 => n91, A2 => n90, ZN => n93);
   U20 : BUF_X1 port map( A => n159, Z => n81);
   U21 : BUF_X1 port map( A => n161, Z => n87);
   U22 : INV_X1 port map( A => n95, ZN => n89);
   U23 : AOI21_X1 port map( B1 => n94, B2 => n93, A => n92, ZN => n95);
   U24 : NOR3_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => n90, ZN => n161);
   U25 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n92);
   U26 : INV_X1 port map( A => SEL_in(0), ZN => n90);
   U27 : AND3_X1 port map( A1 => n90, A2 => n91, A3 => SEL_in(2), ZN => n159);
   U28 : INV_X1 port map( A => SEL_in(1), ZN => n91);
   U29 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(5));
   U30 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82, 
                           C1 => IN5(5), C2 => n79, ZN => n106);
   U31 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN 
                           => n107);
   U32 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(6));
   U33 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN 
                           => n109);
   U34 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82, 
                           C1 => IN5(6), C2 => n79, ZN => n108);
   U35 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(7));
   U36 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN 
                           => n111);
   U37 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82, 
                           C1 => IN5(7), C2 => n79, ZN => n110);
   U38 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(8));
   U39 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN 
                           => n113);
   U40 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82, 
                           C1 => IN5(8), C2 => n79, ZN => n112);
   U41 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(9));
   U42 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN 
                           => n115);
   U43 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82, 
                           C1 => IN5(9), C2 => n79, ZN => n114);
   U44 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(10));
   U45 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n117);
   U46 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => n82
                           , C1 => IN5(10), C2 => n79, ZN => n116);
   U47 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(11));
   U48 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n119);
   U49 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => n82
                           , C1 => IN5(11), C2 => n79, ZN => n118);
   U50 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(12));
   U51 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2, 
                           ZN => n121);
   U52 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => n83
                           , C1 => IN5(12), C2 => n80, ZN => n120);
   U53 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(13));
   U54 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2, 
                           ZN => n123);
   U55 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => n83
                           , C1 => IN5(13), C2 => n80, ZN => n122);
   U56 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(14));
   U57 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n125);
   U58 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n124);
   U59 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(15));
   U60 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n127);
   U61 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n126);
   U62 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(16));
   U63 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2, 
                           ZN => n129);
   U64 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n128);
   U65 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(17));
   U66 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2, 
                           ZN => n131);
   U67 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n130);
   U68 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(18));
   U69 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2, 
                           ZN => n133);
   U70 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n132);
   U71 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(19));
   U72 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n135);
   U73 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n134);
   U74 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(20));
   U75 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n137);
   U76 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n136);
   U77 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(21));
   U78 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n139);
   U79 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n138);
   U80 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(22));
   U81 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n141);
   U82 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n140);
   U83 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(23));
   U84 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n143);
   U85 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n142);
   U86 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Z(24));
   U87 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3, 
                           ZN => n145);
   U88 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n144);
   U89 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Z(25));
   U90 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3, 
                           ZN => n147);
   U91 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84
                           , C1 => IN5(25), C2 => n81, ZN => n146);
   U92 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(26));
   U93 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3, 
                           ZN => n149);
   U94 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84
                           , C1 => IN5(26), C2 => n81, ZN => n148);
   U95 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Z(27));
   U96 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3, 
                           ZN => n151);
   U97 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84
                           , C1 => IN5(27), C2 => n81, ZN => n150);
   U98 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Z(28));
   U99 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3, 
                           ZN => n153);
   U100 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => 
                           n84, C1 => IN5(28), C2 => n81, ZN => n152);
   U101 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Z(29));
   U102 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3,
                           ZN => n155);
   U103 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => 
                           n84, C1 => IN5(29), C2 => n81, ZN => n154);
   U104 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => Z(30));
   U105 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3,
                           ZN => n157);
   U106 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => 
                           n84, C1 => IN5(30), C2 => n81, ZN => n156);
   U107 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(4));
   U108 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN
                           => n105);
   U110 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82,
                           C1 => IN5(4), C2 => n79, ZN => n104);
   U111 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(0));
   U112 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN
                           => n97);
   U113 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82,
                           C1 => IN5(0), C2 => n79, ZN => n96);
   U114 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(1));
   U115 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN
                           => n99);
   U116 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82,
                           C1 => IN5(1), C2 => n79, ZN => n98);
   U117 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(2));
   U118 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN
                           => n101);
   U119 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82,
                           C1 => IN5(2), C2 => n79, ZN => n100);
   U120 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(3));
   U121 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN
                           => n103);
   U122 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82,
                           C1 => IN5(3), C2 => n79, ZN => n102);
   U123 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => Z(31));
   U124 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n163);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_5 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_5;

architecture SYN_bhv of mux5to1_numBit32_5 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n91, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n160);
   U2 : BUF_X1 port map( A => n158, Z => n4);
   U3 : BUF_X1 port map( A => n158, Z => n77);
   U4 : BUF_X1 port map( A => n158, Z => n78);
   U5 : BUF_X1 port map( A => n89, Z => n1);
   U6 : BUF_X1 port map( A => n89, Z => n2);
   U7 : NOR2_X1 port map( A1 => n88, A2 => n93, ZN => n158);
   U8 : INV_X1 port map( A => n94, ZN => n88);
   U9 : BUF_X1 port map( A => n89, Z => n3);
   U10 : NOR4_X1 port map( A1 => n92, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n94);
   U11 : BUF_X1 port map( A => n160, Z => n82);
   U12 : BUF_X1 port map( A => n160, Z => n83);
   U13 : BUF_X1 port map( A => n159, Z => n79);
   U14 : BUF_X1 port map( A => n159, Z => n80);
   U15 : BUF_X1 port map( A => n161, Z => n85);
   U16 : BUF_X1 port map( A => n161, Z => n86);
   U17 : BUF_X1 port map( A => n160, Z => n84);
   U18 : NOR2_X1 port map( A1 => n91, A2 => n90, ZN => n93);
   U19 : BUF_X1 port map( A => n159, Z => n81);
   U20 : BUF_X1 port map( A => n161, Z => n87);
   U21 : INV_X1 port map( A => n95, ZN => n89);
   U22 : AOI21_X1 port map( B1 => n94, B2 => n93, A => n92, ZN => n95);
   U23 : NOR3_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => n90, ZN => n161);
   U24 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n92);
   U25 : INV_X1 port map( A => SEL_in(0), ZN => n90);
   U26 : AND3_X1 port map( A1 => n90, A2 => n91, A3 => SEL_in(2), ZN => n159);
   U27 : INV_X1 port map( A => SEL_in(1), ZN => n91);
   U28 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(7));
   U29 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82, 
                           C1 => IN5(7), C2 => n79, ZN => n110);
   U30 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN 
                           => n111);
   U31 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(8));
   U32 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN 
                           => n113);
   U33 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82, 
                           C1 => IN5(8), C2 => n79, ZN => n112);
   U34 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(9));
   U35 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN 
                           => n115);
   U36 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82, 
                           C1 => IN5(9), C2 => n79, ZN => n114);
   U37 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(10));
   U38 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n117);
   U39 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => n82
                           , C1 => IN5(10), C2 => n79, ZN => n116);
   U40 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(11));
   U41 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n119);
   U42 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => n82
                           , C1 => IN5(11), C2 => n79, ZN => n118);
   U43 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(12));
   U44 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2, 
                           ZN => n121);
   U45 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => n83
                           , C1 => IN5(12), C2 => n80, ZN => n120);
   U46 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(13));
   U47 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2, 
                           ZN => n123);
   U48 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => n83
                           , C1 => IN5(13), C2 => n80, ZN => n122);
   U49 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(14));
   U50 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n125);
   U51 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n124);
   U52 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(15));
   U53 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n127);
   U54 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n126);
   U55 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(16));
   U56 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2, 
                           ZN => n129);
   U57 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n128);
   U58 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(17));
   U59 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2, 
                           ZN => n131);
   U60 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n130);
   U61 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(18));
   U62 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2, 
                           ZN => n133);
   U63 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n132);
   U64 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(19));
   U65 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n135);
   U66 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n134);
   U67 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(20));
   U68 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n137);
   U69 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n136);
   U70 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(21));
   U71 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n139);
   U72 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n138);
   U73 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(22));
   U74 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n141);
   U75 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n140);
   U76 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(23));
   U77 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n143);
   U78 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n142);
   U79 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Z(24));
   U80 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3, 
                           ZN => n145);
   U81 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n144);
   U82 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Z(25));
   U83 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3, 
                           ZN => n147);
   U84 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84
                           , C1 => IN5(25), C2 => n81, ZN => n146);
   U85 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(26));
   U86 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3, 
                           ZN => n149);
   U87 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84
                           , C1 => IN5(26), C2 => n81, ZN => n148);
   U88 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Z(27));
   U89 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3, 
                           ZN => n151);
   U90 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84
                           , C1 => IN5(27), C2 => n81, ZN => n150);
   U91 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Z(28));
   U92 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3, 
                           ZN => n153);
   U93 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => n84
                           , C1 => IN5(28), C2 => n81, ZN => n152);
   U94 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Z(29));
   U95 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3, 
                           ZN => n155);
   U96 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => n84
                           , C1 => IN5(29), C2 => n81, ZN => n154);
   U97 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => Z(30));
   U98 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3, 
                           ZN => n157);
   U99 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => n84
                           , C1 => IN5(30), C2 => n81, ZN => n156);
   U100 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(6));
   U101 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN
                           => n109);
   U102 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82,
                           C1 => IN5(6), C2 => n79, ZN => n108);
   U103 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(0));
   U104 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN
                           => n97);
   U105 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82,
                           C1 => IN5(0), C2 => n79, ZN => n96);
   U106 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(1));
   U107 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN
                           => n99);
   U108 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82,
                           C1 => IN5(1), C2 => n79, ZN => n98);
   U110 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(2));
   U111 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN
                           => n101);
   U112 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82,
                           C1 => IN5(2), C2 => n79, ZN => n100);
   U113 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(3));
   U114 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN
                           => n103);
   U115 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82,
                           C1 => IN5(3), C2 => n79, ZN => n102);
   U116 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(4));
   U117 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN
                           => n105);
   U118 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82,
                           C1 => IN5(4), C2 => n79, ZN => n104);
   U119 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(5));
   U120 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN
                           => n107);
   U121 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82,
                           C1 => IN5(5), C2 => n79, ZN => n106);
   U122 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => Z(31));
   U123 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n163);
   U124 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => 
                           n84, C1 => IN5(31), C2 => n81, ZN => n162);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_4 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_4;

architecture SYN_bhv of mux5to1_numBit32_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n91, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n160);
   U2 : BUF_X1 port map( A => n158, Z => n4);
   U3 : BUF_X1 port map( A => n158, Z => n77);
   U4 : BUF_X1 port map( A => n158, Z => n78);
   U5 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => n84,
                           C1 => IN5(31), C2 => n81, ZN => n162);
   U6 : BUF_X1 port map( A => n89, Z => n1);
   U7 : BUF_X1 port map( A => n89, Z => n2);
   U8 : NOR2_X1 port map( A1 => n88, A2 => n93, ZN => n158);
   U9 : INV_X1 port map( A => n94, ZN => n88);
   U10 : BUF_X1 port map( A => n89, Z => n3);
   U11 : NOR4_X1 port map( A1 => n92, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n94);
   U12 : BUF_X1 port map( A => n160, Z => n82);
   U13 : BUF_X1 port map( A => n160, Z => n83);
   U14 : BUF_X1 port map( A => n159, Z => n79);
   U15 : BUF_X1 port map( A => n159, Z => n80);
   U16 : BUF_X1 port map( A => n161, Z => n85);
   U17 : BUF_X1 port map( A => n161, Z => n86);
   U18 : BUF_X1 port map( A => n160, Z => n84);
   U19 : NOR2_X1 port map( A1 => n91, A2 => n90, ZN => n93);
   U20 : BUF_X1 port map( A => n159, Z => n81);
   U21 : BUF_X1 port map( A => n161, Z => n87);
   U22 : INV_X1 port map( A => n95, ZN => n89);
   U23 : AOI21_X1 port map( B1 => n94, B2 => n93, A => n92, ZN => n95);
   U24 : NOR3_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => n90, ZN => n161);
   U25 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n92);
   U26 : INV_X1 port map( A => SEL_in(0), ZN => n90);
   U27 : AND3_X1 port map( A1 => n90, A2 => n91, A3 => SEL_in(2), ZN => n159);
   U28 : INV_X1 port map( A => SEL_in(1), ZN => n91);
   U29 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(9));
   U30 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82, 
                           C1 => IN5(9), C2 => n79, ZN => n114);
   U31 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN 
                           => n115);
   U32 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(10));
   U33 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n117);
   U34 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => n82
                           , C1 => IN5(10), C2 => n79, ZN => n116);
   U35 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(11));
   U36 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n119);
   U37 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => n82
                           , C1 => IN5(11), C2 => n79, ZN => n118);
   U38 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(12));
   U39 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2, 
                           ZN => n121);
   U40 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => n83
                           , C1 => IN5(12), C2 => n80, ZN => n120);
   U41 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(13));
   U42 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2, 
                           ZN => n123);
   U43 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => n83
                           , C1 => IN5(13), C2 => n80, ZN => n122);
   U44 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(14));
   U45 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n125);
   U46 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n124);
   U47 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(15));
   U48 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n127);
   U49 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n126);
   U50 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(16));
   U51 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2, 
                           ZN => n129);
   U52 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n128);
   U53 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(17));
   U54 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2, 
                           ZN => n131);
   U55 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n130);
   U56 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(18));
   U57 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2, 
                           ZN => n133);
   U58 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n132);
   U59 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(19));
   U60 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n135);
   U61 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n134);
   U62 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(20));
   U63 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n137);
   U64 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n136);
   U65 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(21));
   U66 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n139);
   U67 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n138);
   U68 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(22));
   U69 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n141);
   U70 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n140);
   U71 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(23));
   U72 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n143);
   U73 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n142);
   U74 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Z(24));
   U75 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3, 
                           ZN => n145);
   U76 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n144);
   U77 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Z(25));
   U78 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3, 
                           ZN => n147);
   U79 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84
                           , C1 => IN5(25), C2 => n81, ZN => n146);
   U80 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(26));
   U81 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3, 
                           ZN => n149);
   U82 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84
                           , C1 => IN5(26), C2 => n81, ZN => n148);
   U83 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Z(27));
   U84 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3, 
                           ZN => n151);
   U85 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84
                           , C1 => IN5(27), C2 => n81, ZN => n150);
   U86 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Z(28));
   U87 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3, 
                           ZN => n153);
   U88 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => n84
                           , C1 => IN5(28), C2 => n81, ZN => n152);
   U89 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Z(29));
   U90 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3, 
                           ZN => n155);
   U91 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => n84
                           , C1 => IN5(29), C2 => n81, ZN => n154);
   U92 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => Z(30));
   U93 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3, 
                           ZN => n157);
   U94 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => n84
                           , C1 => IN5(30), C2 => n81, ZN => n156);
   U95 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(8));
   U96 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN 
                           => n113);
   U97 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82, 
                           C1 => IN5(8), C2 => n79, ZN => n112);
   U98 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(0));
   U99 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN 
                           => n97);
   U100 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82,
                           C1 => IN5(0), C2 => n79, ZN => n96);
   U101 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(1));
   U102 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN
                           => n99);
   U103 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82,
                           C1 => IN5(1), C2 => n79, ZN => n98);
   U104 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(2));
   U105 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN
                           => n101);
   U106 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82,
                           C1 => IN5(2), C2 => n79, ZN => n100);
   U107 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(3));
   U108 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN
                           => n103);
   U110 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82,
                           C1 => IN5(3), C2 => n79, ZN => n102);
   U111 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(4));
   U112 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN
                           => n105);
   U113 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82,
                           C1 => IN5(4), C2 => n79, ZN => n104);
   U114 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(5));
   U115 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN
                           => n107);
   U116 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82,
                           C1 => IN5(5), C2 => n79, ZN => n106);
   U117 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(6));
   U118 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN
                           => n109);
   U119 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82,
                           C1 => IN5(6), C2 => n79, ZN => n108);
   U120 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(7));
   U121 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN
                           => n111);
   U122 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82,
                           C1 => IN5(7), C2 => n79, ZN => n110);
   U123 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => Z(31));
   U124 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n163);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_3 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_3;

architecture SYN_bhv of mux5to1_numBit32_3 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n90, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n160);
   U2 : BUF_X1 port map( A => n158, Z => n4);
   U3 : BUF_X1 port map( A => n158, Z => n77);
   U4 : BUF_X1 port map( A => n158, Z => n78);
   U5 : BUF_X1 port map( A => n89, Z => n1);
   U6 : BUF_X1 port map( A => n89, Z => n2);
   U7 : NOR2_X1 port map( A1 => n88, A2 => n93, ZN => n158);
   U8 : INV_X1 port map( A => n94, ZN => n88);
   U9 : BUF_X1 port map( A => n89, Z => n3);
   U10 : NOR4_X1 port map( A1 => n92, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n94);
   U11 : BUF_X1 port map( A => n160, Z => n82);
   U12 : BUF_X1 port map( A => n160, Z => n83);
   U13 : BUF_X1 port map( A => n159, Z => n79);
   U14 : BUF_X1 port map( A => n159, Z => n80);
   U15 : BUF_X1 port map( A => n161, Z => n85);
   U16 : BUF_X1 port map( A => n161, Z => n86);
   U17 : BUF_X1 port map( A => n160, Z => n84);
   U18 : NOR2_X1 port map( A1 => n90, A2 => n91, ZN => n93);
   U19 : BUF_X1 port map( A => n159, Z => n81);
   U20 : BUF_X1 port map( A => n161, Z => n87);
   U21 : INV_X1 port map( A => n95, ZN => n89);
   U22 : AOI21_X1 port map( B1 => n94, B2 => n93, A => n92, ZN => n95);
   U23 : NOR3_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => n91, ZN => n161);
   U24 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n92);
   U25 : INV_X1 port map( A => SEL_in(0), ZN => n91);
   U26 : AND3_X1 port map( A1 => n91, A2 => n90, A3 => SEL_in(2), ZN => n159);
   U27 : INV_X1 port map( A => SEL_in(1), ZN => n90);
   U28 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(11));
   U29 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => n82
                           , C1 => IN5(11), C2 => n79, ZN => n118);
   U30 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n119);
   U31 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(12));
   U32 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2, 
                           ZN => n121);
   U33 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => n83
                           , C1 => IN5(12), C2 => n80, ZN => n120);
   U34 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(13));
   U35 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2, 
                           ZN => n123);
   U36 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => n83
                           , C1 => IN5(13), C2 => n80, ZN => n122);
   U37 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(14));
   U38 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n125);
   U39 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n124);
   U40 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(15));
   U41 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n127);
   U42 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n126);
   U43 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(16));
   U44 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2, 
                           ZN => n129);
   U45 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n128);
   U46 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(17));
   U47 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2, 
                           ZN => n131);
   U48 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n130);
   U49 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(18));
   U50 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2, 
                           ZN => n133);
   U51 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n132);
   U52 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(19));
   U53 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n135);
   U54 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n134);
   U55 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(20));
   U56 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n137);
   U57 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n136);
   U58 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(21));
   U59 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n139);
   U60 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n138);
   U61 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(22));
   U62 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n141);
   U63 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n140);
   U64 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(23));
   U65 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n143);
   U66 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n142);
   U67 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Z(24));
   U68 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3, 
                           ZN => n145);
   U69 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n144);
   U70 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Z(25));
   U71 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3, 
                           ZN => n147);
   U72 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84
                           , C1 => IN5(25), C2 => n81, ZN => n146);
   U73 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(26));
   U74 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3, 
                           ZN => n149);
   U75 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84
                           , C1 => IN5(26), C2 => n81, ZN => n148);
   U76 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Z(27));
   U77 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3, 
                           ZN => n151);
   U78 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84
                           , C1 => IN5(27), C2 => n81, ZN => n150);
   U79 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Z(28));
   U80 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3, 
                           ZN => n153);
   U81 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => n84
                           , C1 => IN5(28), C2 => n81, ZN => n152);
   U82 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Z(29));
   U83 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3, 
                           ZN => n155);
   U84 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => n84
                           , C1 => IN5(29), C2 => n81, ZN => n154);
   U85 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => Z(30));
   U86 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3, 
                           ZN => n157);
   U87 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => n84
                           , C1 => IN5(30), C2 => n81, ZN => n156);
   U88 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(10));
   U89 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n117);
   U90 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => n82
                           , C1 => IN5(10), C2 => n79, ZN => n116);
   U91 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(0));
   U92 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN 
                           => n97);
   U93 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82, 
                           C1 => IN5(0), C2 => n79, ZN => n96);
   U94 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(1));
   U95 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN 
                           => n99);
   U96 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82, 
                           C1 => IN5(1), C2 => n79, ZN => n98);
   U97 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(2));
   U98 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN 
                           => n101);
   U99 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82, 
                           C1 => IN5(2), C2 => n79, ZN => n100);
   U100 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(3));
   U101 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN
                           => n103);
   U102 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82,
                           C1 => IN5(3), C2 => n79, ZN => n102);
   U103 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(4));
   U104 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN
                           => n105);
   U105 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82,
                           C1 => IN5(4), C2 => n79, ZN => n104);
   U106 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(5));
   U107 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN
                           => n107);
   U108 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82,
                           C1 => IN5(5), C2 => n79, ZN => n106);
   U110 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(6));
   U111 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN
                           => n109);
   U112 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82,
                           C1 => IN5(6), C2 => n79, ZN => n108);
   U113 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(7));
   U114 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN
                           => n111);
   U115 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82,
                           C1 => IN5(7), C2 => n79, ZN => n110);
   U116 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(8));
   U117 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN
                           => n113);
   U118 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82,
                           C1 => IN5(8), C2 => n79, ZN => n112);
   U119 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(9));
   U120 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN
                           => n115);
   U121 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82,
                           C1 => IN5(9), C2 => n79, ZN => n114);
   U122 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => Z(31));
   U123 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n163);
   U124 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => 
                           n84, C1 => IN5(31), C2 => n81, ZN => n162);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_2 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_2;

architecture SYN_bhv of mux5to1_numBit32_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n91, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n160);
   U2 : BUF_X1 port map( A => n158, Z => n4);
   U3 : BUF_X1 port map( A => n158, Z => n77);
   U4 : BUF_X1 port map( A => n158, Z => n78);
   U5 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => n84,
                           C1 => IN5(31), C2 => n81, ZN => n162);
   U6 : BUF_X1 port map( A => n89, Z => n1);
   U7 : BUF_X1 port map( A => n89, Z => n2);
   U8 : NOR2_X1 port map( A1 => n88, A2 => n93, ZN => n158);
   U9 : INV_X1 port map( A => n94, ZN => n88);
   U10 : BUF_X1 port map( A => n89, Z => n3);
   U11 : NOR4_X1 port map( A1 => n92, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n94);
   U12 : BUF_X1 port map( A => n160, Z => n82);
   U13 : BUF_X1 port map( A => n160, Z => n83);
   U14 : BUF_X1 port map( A => n159, Z => n79);
   U15 : BUF_X1 port map( A => n159, Z => n80);
   U16 : BUF_X1 port map( A => n161, Z => n85);
   U17 : BUF_X1 port map( A => n161, Z => n86);
   U18 : BUF_X1 port map( A => n160, Z => n84);
   U19 : NOR2_X1 port map( A1 => n91, A2 => n90, ZN => n93);
   U20 : BUF_X1 port map( A => n159, Z => n81);
   U21 : BUF_X1 port map( A => n161, Z => n87);
   U22 : INV_X1 port map( A => n95, ZN => n89);
   U23 : AOI21_X1 port map( B1 => n94, B2 => n93, A => n92, ZN => n95);
   U24 : NOR3_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => n90, ZN => n161);
   U25 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n92);
   U26 : INV_X1 port map( A => SEL_in(0), ZN => n90);
   U27 : AND3_X1 port map( A1 => n90, A2 => n91, A3 => SEL_in(2), ZN => n159);
   U28 : INV_X1 port map( A => SEL_in(1), ZN => n91);
   U29 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(13));
   U30 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => n83
                           , C1 => IN5(13), C2 => n80, ZN => n122);
   U31 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2, 
                           ZN => n123);
   U32 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(14));
   U33 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n125);
   U34 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n124);
   U35 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(15));
   U36 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n127);
   U37 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n126);
   U38 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(16));
   U39 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2, 
                           ZN => n129);
   U40 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n128);
   U41 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(17));
   U42 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2, 
                           ZN => n131);
   U43 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n130);
   U44 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(18));
   U45 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2, 
                           ZN => n133);
   U46 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n132);
   U47 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(19));
   U48 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n135);
   U49 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n134);
   U50 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(20));
   U51 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n137);
   U52 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n136);
   U53 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(21));
   U54 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n139);
   U55 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n138);
   U56 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(22));
   U57 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n141);
   U58 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n140);
   U59 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(23));
   U60 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n143);
   U61 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n142);
   U62 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Z(24));
   U63 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3, 
                           ZN => n145);
   U64 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n144);
   U65 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Z(25));
   U66 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3, 
                           ZN => n147);
   U67 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84
                           , C1 => IN5(25), C2 => n81, ZN => n146);
   U68 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(26));
   U69 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3, 
                           ZN => n149);
   U70 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84
                           , C1 => IN5(26), C2 => n81, ZN => n148);
   U71 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Z(27));
   U72 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3, 
                           ZN => n151);
   U73 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84
                           , C1 => IN5(27), C2 => n81, ZN => n150);
   U74 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Z(28));
   U75 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3, 
                           ZN => n153);
   U76 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => n84
                           , C1 => IN5(28), C2 => n81, ZN => n152);
   U77 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Z(29));
   U78 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3, 
                           ZN => n155);
   U79 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => n84
                           , C1 => IN5(29), C2 => n81, ZN => n154);
   U80 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => Z(30));
   U81 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3, 
                           ZN => n157);
   U82 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => n84
                           , C1 => IN5(30), C2 => n81, ZN => n156);
   U83 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(12));
   U84 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2, 
                           ZN => n121);
   U85 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => n83
                           , C1 => IN5(12), C2 => n80, ZN => n120);
   U86 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(0));
   U87 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN 
                           => n97);
   U88 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82, 
                           C1 => IN5(0), C2 => n79, ZN => n96);
   U89 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(1));
   U90 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN 
                           => n99);
   U91 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82, 
                           C1 => IN5(1), C2 => n79, ZN => n98);
   U92 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(2));
   U93 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN 
                           => n101);
   U94 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82, 
                           C1 => IN5(2), C2 => n79, ZN => n100);
   U95 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(3));
   U96 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN 
                           => n103);
   U97 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82, 
                           C1 => IN5(3), C2 => n79, ZN => n102);
   U98 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(4));
   U99 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN 
                           => n105);
   U100 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82,
                           C1 => IN5(4), C2 => n79, ZN => n104);
   U101 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(5));
   U102 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN
                           => n107);
   U103 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82,
                           C1 => IN5(5), C2 => n79, ZN => n106);
   U104 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(6));
   U105 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN
                           => n109);
   U106 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82,
                           C1 => IN5(6), C2 => n79, ZN => n108);
   U107 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(7));
   U108 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN
                           => n111);
   U110 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82,
                           C1 => IN5(7), C2 => n79, ZN => n110);
   U111 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(8));
   U112 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN
                           => n113);
   U113 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82,
                           C1 => IN5(8), C2 => n79, ZN => n112);
   U114 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(9));
   U115 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN
                           => n115);
   U116 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82,
                           C1 => IN5(9), C2 => n79, ZN => n114);
   U117 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(10));
   U118 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n117);
   U119 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => 
                           n82, C1 => IN5(10), C2 => n79, ZN => n116);
   U120 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(11));
   U121 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n119);
   U122 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => 
                           n82, C1 => IN5(11), C2 => n79, ZN => n118);
   U123 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => Z(31));
   U124 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n163);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_1 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_1;

architecture SYN_bhv of mux5to1_numBit32_1 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n91, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n160);
   U2 : BUF_X1 port map( A => n158, Z => n4);
   U3 : BUF_X1 port map( A => n158, Z => n77);
   U4 : BUF_X1 port map( A => n158, Z => n78);
   U5 : BUF_X1 port map( A => n89, Z => n1);
   U6 : BUF_X1 port map( A => n89, Z => n2);
   U7 : NOR2_X1 port map( A1 => n88, A2 => n93, ZN => n158);
   U8 : INV_X1 port map( A => n94, ZN => n88);
   U9 : BUF_X1 port map( A => n89, Z => n3);
   U10 : NOR4_X1 port map( A1 => n92, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n94);
   U11 : BUF_X1 port map( A => n160, Z => n82);
   U12 : BUF_X1 port map( A => n160, Z => n83);
   U13 : BUF_X1 port map( A => n159, Z => n79);
   U14 : BUF_X1 port map( A => n159, Z => n80);
   U15 : BUF_X1 port map( A => n161, Z => n85);
   U16 : BUF_X1 port map( A => n161, Z => n86);
   U17 : BUF_X1 port map( A => n160, Z => n84);
   U18 : NOR2_X1 port map( A1 => n91, A2 => n90, ZN => n93);
   U19 : BUF_X1 port map( A => n159, Z => n81);
   U20 : BUF_X1 port map( A => n161, Z => n87);
   U21 : INV_X1 port map( A => n95, ZN => n89);
   U22 : AOI21_X1 port map( B1 => n94, B2 => n93, A => n92, ZN => n95);
   U23 : NOR3_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => n90, ZN => n161);
   U24 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n92);
   U25 : INV_X1 port map( A => SEL_in(0), ZN => n90);
   U26 : AND3_X1 port map( A1 => n90, A2 => n91, A3 => SEL_in(2), ZN => n159);
   U27 : INV_X1 port map( A => SEL_in(1), ZN => n91);
   U28 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(15));
   U29 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n126);
   U30 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n127);
   U31 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(16));
   U32 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2, 
                           ZN => n129);
   U33 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n128);
   U34 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(17));
   U35 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2, 
                           ZN => n131);
   U36 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n130);
   U37 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(18));
   U38 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2, 
                           ZN => n133);
   U39 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n132);
   U40 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(19));
   U41 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n135);
   U42 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n134);
   U43 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(20));
   U44 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n137);
   U45 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n136);
   U46 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(21));
   U47 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n139);
   U48 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n138);
   U49 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(22));
   U50 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n141);
   U51 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n140);
   U52 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(23));
   U53 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n143);
   U54 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n142);
   U55 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Z(24));
   U56 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3, 
                           ZN => n145);
   U57 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n144);
   U58 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Z(25));
   U59 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3, 
                           ZN => n147);
   U60 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84
                           , C1 => IN5(25), C2 => n81, ZN => n146);
   U61 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(26));
   U62 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3, 
                           ZN => n149);
   U63 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84
                           , C1 => IN5(26), C2 => n81, ZN => n148);
   U64 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Z(27));
   U65 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3, 
                           ZN => n151);
   U66 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84
                           , C1 => IN5(27), C2 => n81, ZN => n150);
   U67 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Z(28));
   U68 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3, 
                           ZN => n153);
   U69 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => n84
                           , C1 => IN5(28), C2 => n81, ZN => n152);
   U70 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Z(29));
   U71 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3, 
                           ZN => n155);
   U72 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => n84
                           , C1 => IN5(29), C2 => n81, ZN => n154);
   U73 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => Z(30));
   U74 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3, 
                           ZN => n157);
   U75 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => n84
                           , C1 => IN5(30), C2 => n81, ZN => n156);
   U76 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(14));
   U77 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n125);
   U78 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n124);
   U79 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(0));
   U80 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN 
                           => n97);
   U81 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82, 
                           C1 => IN5(0), C2 => n79, ZN => n96);
   U82 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(1));
   U83 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN 
                           => n99);
   U84 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82, 
                           C1 => IN5(1), C2 => n79, ZN => n98);
   U85 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(2));
   U86 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN 
                           => n101);
   U87 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82, 
                           C1 => IN5(2), C2 => n79, ZN => n100);
   U88 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(3));
   U89 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN 
                           => n103);
   U90 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82, 
                           C1 => IN5(3), C2 => n79, ZN => n102);
   U91 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(4));
   U92 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN 
                           => n105);
   U93 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82, 
                           C1 => IN5(4), C2 => n79, ZN => n104);
   U94 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(5));
   U95 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN 
                           => n107);
   U96 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82, 
                           C1 => IN5(5), C2 => n79, ZN => n106);
   U97 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(6));
   U98 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN 
                           => n109);
   U99 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82, 
                           C1 => IN5(6), C2 => n79, ZN => n108);
   U100 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(7));
   U101 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN
                           => n111);
   U102 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82,
                           C1 => IN5(7), C2 => n79, ZN => n110);
   U103 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(8));
   U104 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN
                           => n113);
   U105 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82,
                           C1 => IN5(8), C2 => n79, ZN => n112);
   U106 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(9));
   U107 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN
                           => n115);
   U108 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82,
                           C1 => IN5(9), C2 => n79, ZN => n114);
   U110 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(10));
   U111 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n117);
   U112 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => 
                           n82, C1 => IN5(10), C2 => n79, ZN => n116);
   U113 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(11));
   U114 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n119);
   U115 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => 
                           n82, C1 => IN5(11), C2 => n79, ZN => n118);
   U116 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(12));
   U117 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2,
                           ZN => n121);
   U118 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => 
                           n83, C1 => IN5(12), C2 => n80, ZN => n120);
   U119 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(13));
   U120 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2,
                           ZN => n123);
   U121 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => 
                           n83, C1 => IN5(13), C2 => n80, ZN => n122);
   U122 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => Z(31));
   U123 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n163);
   U124 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => 
                           n84, C1 => IN5(31), C2 => n81, ZN => n162);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_4 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_4;

architecture SYN_bhv of mux41_NBIT32_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n145, Z => n73);
   U2 : BUF_X1 port map( A => n147, Z => n79);
   U3 : BUF_X1 port map( A => n144, Z => n70);
   U4 : BUF_X1 port map( A => n146, Z => n76);
   U5 : BUF_X1 port map( A => n145, Z => n72);
   U6 : BUF_X1 port map( A => n147, Z => n78);
   U7 : BUF_X1 port map( A => n144, Z => n1);
   U8 : BUF_X1 port map( A => n146, Z => n75);
   U9 : BUF_X1 port map( A => n145, Z => n74);
   U10 : BUF_X1 port map( A => n147, Z => n80);
   U11 : BUF_X1 port map( A => n144, Z => n71);
   U12 : BUF_X1 port map( A => n146, Z => n77);
   U13 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n145);
   U14 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n144);
   U15 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n147);
   U16 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n146);
   U17 : INV_X1 port map( A => S(0), ZN => n81);
   U18 : NAND2_X1 port map( A1 => n87, A2 => n86, ZN => Z(11));
   U19 : NAND2_X1 port map( A1 => n83, A2 => n82, ZN => Z(0));
   U20 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n83);
   U21 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n82);
   U22 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(4));
   U23 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN =>
                           n135);
   U24 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN =>
                           n134);
   U25 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(8));
   U26 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n143);
   U27 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n142);
   U28 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => Z(12));
   U29 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n89);
   U30 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN 
                           => n88);
   U31 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(16));
   U32 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n97);
   U33 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n96);
   U34 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(5));
   U35 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN =>
                           n137);
   U36 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN =>
                           n136);
   U37 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(1));
   U38 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN => 
                           n105);
   U39 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN =>
                           n104);
   U40 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => Z(13));
   U41 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n91);
   U42 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN 
                           => n90);
   U43 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(17));
   U44 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n99);
   U45 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n98);
   U46 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(25));
   U47 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n117);
   U48 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n116);
   U49 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(2));
   U50 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN =>
                           n127);
   U51 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN =>
                           n126);
   U52 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(6));
   U53 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n139);
   U54 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n138);
   U55 : NAND2_X1 port map( A1 => n93, A2 => n92, ZN => Z(14));
   U56 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n93);
   U57 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN 
                           => n92);
   U58 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(18));
   U59 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n101);
   U60 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n100);
   U61 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(26));
   U62 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n119);
   U63 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n118);
   U64 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(22));
   U65 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n111);
   U66 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n110);
   U67 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(21));
   U68 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n109);
   U69 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n108);
   U70 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(30));
   U71 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN 
                           => n129);
   U72 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN 
                           => n128);
   U73 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(29));
   U74 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n125);
   U75 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n124);
   U76 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(28));
   U77 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n123);
   U78 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n122);
   U79 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(3));
   U80 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN =>
                           n133);
   U81 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN =>
                           n132);
   U82 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(7));
   U83 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n141);
   U84 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n140);
   U85 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => Z(15));
   U86 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n95);
   U87 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN 
                           => n94);
   U88 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(19));
   U89 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n103);
   U90 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN 
                           => n102);
   U91 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(23));
   U92 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN 
                           => n113);
   U93 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN 
                           => n112);
   U94 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(27));
   U95 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN 
                           => n121);
   U96 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN 
                           => n120);
   U97 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(31));
   U98 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN 
                           => n131);
   U99 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN 
                           => n130);
   U100 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(24));
   U101 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN
                           => n115);
   U102 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN
                           => n114);
   U103 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(9));
   U104 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN 
                           => n149);
   U105 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN 
                           => n148);
   U106 : NAND2_X1 port map( A1 => n85, A2 => n84, ZN => Z(10));
   U107 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n85);
   U108 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN
                           => n84);
   U109 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(20));
   U110 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN
                           => n107);
   U111 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN
                           => n106);
   U112 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n87);
   U113 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN
                           => n86);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_3 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_3;

architecture SYN_bhv of mux41_NBIT32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n145, Z => n72);
   U2 : BUF_X1 port map( A => n147, Z => n78);
   U3 : BUF_X1 port map( A => n145, Z => n73);
   U4 : BUF_X1 port map( A => n147, Z => n79);
   U5 : BUF_X1 port map( A => n144, Z => n1);
   U6 : BUF_X1 port map( A => n146, Z => n75);
   U7 : BUF_X1 port map( A => n144, Z => n70);
   U8 : BUF_X1 port map( A => n146, Z => n76);
   U9 : BUF_X1 port map( A => n145, Z => n74);
   U10 : BUF_X1 port map( A => n147, Z => n80);
   U11 : BUF_X1 port map( A => n144, Z => n71);
   U12 : BUF_X1 port map( A => n146, Z => n77);
   U13 : NAND2_X1 port map( A1 => n83, A2 => n82, ZN => Z(0));
   U14 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n82);
   U15 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n83);
   U16 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(4));
   U17 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN =>
                           n134);
   U18 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN =>
                           n135);
   U19 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(8));
   U20 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n142);
   U21 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n143);
   U22 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => Z(12));
   U23 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN 
                           => n88);
   U24 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n89);
   U25 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(16));
   U26 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n96);
   U27 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n97);
   U28 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(24));
   U29 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN 
                           => n114);
   U30 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN 
                           => n115);
   U31 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(5));
   U32 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN =>
                           n136);
   U33 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN =>
                           n137);
   U34 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(1));
   U35 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN =>
                           n104);
   U36 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN => 
                           n105);
   U37 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(9));
   U38 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN =>
                           n148);
   U39 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN =>
                           n149);
   U40 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => Z(13));
   U41 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN 
                           => n90);
   U42 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n91);
   U43 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(17));
   U44 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n98);
   U45 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n99);
   U46 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(25));
   U47 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n116);
   U48 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n117);
   U49 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(2));
   U50 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN =>
                           n126);
   U51 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN =>
                           n127);
   U52 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(6));
   U53 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n138);
   U54 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n139);
   U55 : NAND2_X1 port map( A1 => n85, A2 => n84, ZN => Z(10));
   U56 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN 
                           => n84);
   U57 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n85);
   U58 : NAND2_X1 port map( A1 => n93, A2 => n92, ZN => Z(14));
   U59 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN 
                           => n92);
   U60 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n93);
   U61 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(18));
   U62 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n100);
   U63 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n101);
   U64 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(26));
   U65 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n118);
   U66 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n119);
   U67 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(22));
   U68 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n110);
   U69 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n111);
   U70 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(21));
   U71 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n108);
   U72 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n109);
   U73 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(20));
   U74 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN 
                           => n106);
   U75 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN 
                           => n107);
   U76 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(30));
   U77 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN 
                           => n128);
   U78 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN 
                           => n129);
   U79 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(29));
   U80 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n124);
   U81 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n125);
   U82 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(28));
   U83 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n122);
   U84 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n123);
   U85 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(3));
   U86 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN =>
                           n132);
   U87 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN =>
                           n133);
   U88 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(7));
   U89 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n140);
   U90 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n141);
   U91 : NAND2_X1 port map( A1 => n87, A2 => n86, ZN => Z(11));
   U92 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN 
                           => n86);
   U93 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n87);
   U94 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => Z(15));
   U95 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN 
                           => n94);
   U96 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n95);
   U97 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(19));
   U98 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN 
                           => n102);
   U99 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n103);
   U100 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(23));
   U101 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN
                           => n112);
   U102 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN
                           => n113);
   U103 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(27));
   U104 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN
                           => n120);
   U105 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN
                           => n121);
   U106 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(31));
   U107 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN
                           => n130);
   U108 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN
                           => n131);
   U109 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n145);
   U110 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n144);
   U111 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n147);
   U112 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n146);
   U113 : INV_X1 port map( A => S(0), ZN => n81);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_2 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_2;

architecture SYN_bhv of mux41_NBIT32_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n20, n21, n22, n23, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65, n66, n67, n70, n71, n72, n73, n74, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, n93, n94 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n1, Z => n20);
   U2 : BUF_X1 port map( A => n1, Z => n9);
   U3 : BUF_X1 port map( A => n3, Z => n22);
   U4 : BUF_X1 port map( A => n2, Z => n6);
   U5 : BUF_X1 port map( A => n3, Z => n21);
   U6 : BUF_X1 port map( A => n2, Z => n5);
   U7 : AND2_X1 port map( A1 => n23, A2 => n26, ZN => n1);
   U8 : BUF_X1 port map( A => n4, Z => n8);
   U9 : BUF_X1 port map( A => n4, Z => n7);
   U10 : NAND2_X1 port map( A1 => n80, A2 => n79, ZN => Z(0));
   U11 : AOI22_X1 port map( A1 => D(0), A2 => n7, B1 => C(0), B2 => n5, ZN => 
                           n79);
   U12 : AOI22_X1 port map( A1 => B(0), A2 => n21, B1 => A(0), B2 => n9, ZN => 
                           n80);
   U13 : NAND2_X1 port map( A1 => n94, A2 => n93, ZN => Z(7));
   U14 : AOI22_X1 port map( A1 => D(7), A2 => n7, B1 => C(7), B2 => n5, ZN => 
                           n93);
   U15 : AOI22_X1 port map( A1 => B(7), A2 => n21, B1 => A(7), B2 => n9, ZN => 
                           n94);
   U16 : AND2_X1 port map( A1 => S(1), A2 => n26, ZN => n2);
   U17 : AND2_X1 port map( A1 => S(0), A2 => n23, ZN => n3);
   U18 : NAND2_X1 port map( A1 => n82, A2 => n81, ZN => Z(1));
   U19 : AOI22_X1 port map( A1 => D(1), A2 => n7, B1 => C(1), B2 => n5, ZN => 
                           n81);
   U20 : AOI22_X1 port map( A1 => B(1), A2 => n21, B1 => A(1), B2 => n9, ZN => 
                           n82);
   U21 : NAND2_X1 port map( A1 => n84, A2 => n83, ZN => Z(2));
   U22 : AOI22_X1 port map( A1 => D(2), A2 => n7, B1 => C(2), B2 => n5, ZN => 
                           n83);
   U23 : AOI22_X1 port map( A1 => B(2), A2 => n21, B1 => A(2), B2 => n9, ZN => 
                           n84);
   U24 : NAND2_X1 port map( A1 => n86, A2 => n85, ZN => Z(3));
   U25 : AOI22_X1 port map( A1 => D(3), A2 => n7, B1 => C(3), B2 => n5, ZN => 
                           n85);
   U26 : AOI22_X1 port map( A1 => B(3), A2 => n21, B1 => A(3), B2 => n9, ZN => 
                           n86);
   U27 : NAND2_X1 port map( A1 => n92, A2 => n91, ZN => Z(6));
   U28 : AOI22_X1 port map( A1 => D(6), A2 => n7, B1 => C(6), B2 => n5, ZN => 
                           n91);
   U29 : AOI22_X1 port map( A1 => B(6), A2 => n21, B1 => A(6), B2 => n9, ZN => 
                           n92);
   U30 : NAND2_X1 port map( A1 => n90, A2 => n89, ZN => Z(5));
   U31 : AOI22_X1 port map( A1 => D(5), A2 => n7, B1 => C(5), B2 => n5, ZN => 
                           n89);
   U32 : AOI22_X1 port map( A1 => B(5), A2 => n21, B1 => A(5), B2 => n9, ZN => 
                           n90);
   U33 : NAND2_X1 port map( A1 => n88, A2 => n87, ZN => Z(4));
   U34 : AOI22_X1 port map( A1 => D(4), A2 => n7, B1 => C(4), B2 => n5, ZN => 
                           n87);
   U35 : AOI22_X1 port map( A1 => B(4), A2 => n21, B1 => A(4), B2 => n9, ZN => 
                           n88);
   U36 : AND2_X1 port map( A1 => S(0), A2 => S(1), ZN => n4);
   U37 : INV_X1 port map( A => S(1), ZN => n23);
   U38 : INV_X1 port map( A => S(0), ZN => n26);
   U39 : AOI22_X1 port map( A1 => B(8), A2 => n22, B1 => A(8), B2 => n20, ZN =>
                           n28);
   U40 : AOI22_X1 port map( A1 => D(8), A2 => n8, B1 => C(8), B2 => n6, ZN => 
                           n27);
   U41 : NAND2_X1 port map( A1 => n28, A2 => n27, ZN => Z(8));
   U42 : AOI22_X1 port map( A1 => B(9), A2 => n22, B1 => A(9), B2 => n20, ZN =>
                           n30);
   U43 : AOI22_X1 port map( A1 => D(9), A2 => n8, B1 => C(9), B2 => n6, ZN => 
                           n29);
   U44 : NAND2_X1 port map( A1 => n30, A2 => n29, ZN => Z(9));
   U45 : AOI22_X1 port map( A1 => B(10), A2 => n22, B1 => A(10), B2 => n20, ZN 
                           => n32);
   U46 : AOI22_X1 port map( A1 => D(10), A2 => n8, B1 => C(10), B2 => n6, ZN =>
                           n31);
   U47 : NAND2_X1 port map( A1 => n32, A2 => n31, ZN => Z(10));
   U48 : AOI22_X1 port map( A1 => B(11), A2 => n22, B1 => A(11), B2 => n20, ZN 
                           => n34);
   U49 : AOI22_X1 port map( A1 => D(11), A2 => n8, B1 => C(11), B2 => n6, ZN =>
                           n33);
   U50 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => Z(11));
   U51 : AOI22_X1 port map( A1 => B(12), A2 => n22, B1 => A(12), B2 => n20, ZN 
                           => n36);
   U52 : AOI22_X1 port map( A1 => D(12), A2 => n8, B1 => C(12), B2 => n6, ZN =>
                           n35);
   U53 : NAND2_X1 port map( A1 => n36, A2 => n35, ZN => Z(12));
   U54 : AOI22_X1 port map( A1 => B(13), A2 => n22, B1 => A(13), B2 => n20, ZN 
                           => n38);
   U55 : AOI22_X1 port map( A1 => D(13), A2 => n8, B1 => C(13), B2 => n6, ZN =>
                           n37);
   U56 : NAND2_X1 port map( A1 => n38, A2 => n37, ZN => Z(13));
   U57 : AOI22_X1 port map( A1 => B(14), A2 => n22, B1 => A(14), B2 => n20, ZN 
                           => n40);
   U58 : AOI22_X1 port map( A1 => D(14), A2 => n8, B1 => C(14), B2 => n6, ZN =>
                           n39);
   U59 : NAND2_X1 port map( A1 => n40, A2 => n39, ZN => Z(14));
   U60 : AOI22_X1 port map( A1 => B(15), A2 => n22, B1 => A(15), B2 => n20, ZN 
                           => n42);
   U61 : AOI22_X1 port map( A1 => D(15), A2 => n8, B1 => C(15), B2 => n6, ZN =>
                           n41);
   U62 : NAND2_X1 port map( A1 => n42, A2 => n41, ZN => Z(15));
   U63 : AOI22_X1 port map( A1 => B(16), A2 => n22, B1 => A(16), B2 => n20, ZN 
                           => n44);
   U64 : AOI22_X1 port map( A1 => D(16), A2 => n8, B1 => C(16), B2 => n6, ZN =>
                           n43);
   U65 : NAND2_X1 port map( A1 => n44, A2 => n43, ZN => Z(16));
   U66 : AOI22_X1 port map( A1 => B(17), A2 => n22, B1 => A(17), B2 => n20, ZN 
                           => n48);
   U67 : AOI22_X1 port map( A1 => D(17), A2 => n8, B1 => C(17), B2 => n6, ZN =>
                           n45);
   U68 : NAND2_X1 port map( A1 => n48, A2 => n45, ZN => Z(17));
   U69 : AOI22_X1 port map( A1 => B(18), A2 => n22, B1 => A(18), B2 => n20, ZN 
                           => n50);
   U70 : AOI22_X1 port map( A1 => D(18), A2 => n8, B1 => C(18), B2 => n6, ZN =>
                           n49);
   U71 : NAND2_X1 port map( A1 => n50, A2 => n49, ZN => Z(18));
   U72 : AOI22_X1 port map( A1 => B(19), A2 => n22, B1 => A(19), B2 => n20, ZN 
                           => n52);
   U73 : AOI22_X1 port map( A1 => D(19), A2 => n8, B1 => C(19), B2 => n6, ZN =>
                           n51);
   U74 : NAND2_X1 port map( A1 => n52, A2 => n51, ZN => Z(19));
   U75 : AOI22_X1 port map( A1 => B(20), A2 => n22, B1 => A(20), B2 => n20, ZN 
                           => n54);
   U76 : AOI22_X1 port map( A1 => D(20), A2 => n8, B1 => C(20), B2 => n6, ZN =>
                           n53);
   U77 : NAND2_X1 port map( A1 => n54, A2 => n53, ZN => Z(20));
   U78 : AOI22_X1 port map( A1 => B(21), A2 => n22, B1 => A(21), B2 => n20, ZN 
                           => n56);
   U79 : AOI22_X1 port map( A1 => D(21), A2 => n8, B1 => C(21), B2 => n6, ZN =>
                           n55);
   U80 : NAND2_X1 port map( A1 => n56, A2 => n55, ZN => Z(21));
   U81 : AOI22_X1 port map( A1 => B(22), A2 => n22, B1 => A(22), B2 => n20, ZN 
                           => n58);
   U82 : AOI22_X1 port map( A1 => D(22), A2 => n8, B1 => C(22), B2 => n6, ZN =>
                           n57);
   U83 : NAND2_X1 port map( A1 => n58, A2 => n57, ZN => Z(22));
   U84 : AOI22_X1 port map( A1 => B(23), A2 => n22, B1 => A(23), B2 => n20, ZN 
                           => n60);
   U85 : AOI22_X1 port map( A1 => D(23), A2 => n8, B1 => C(23), B2 => n6, ZN =>
                           n59);
   U86 : NAND2_X1 port map( A1 => n60, A2 => n59, ZN => Z(23));
   U87 : AOI22_X1 port map( A1 => B(24), A2 => n22, B1 => A(24), B2 => n20, ZN 
                           => n62);
   U88 : AOI22_X1 port map( A1 => D(24), A2 => n8, B1 => C(24), B2 => n6, ZN =>
                           n61);
   U89 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => Z(24));
   U90 : AOI22_X1 port map( A1 => B(25), A2 => n21, B1 => A(25), B2 => n9, ZN 
                           => n64);
   U91 : AOI22_X1 port map( A1 => D(25), A2 => n7, B1 => C(25), B2 => n5, ZN =>
                           n63);
   U92 : NAND2_X1 port map( A1 => n64, A2 => n63, ZN => Z(25));
   U93 : AOI22_X1 port map( A1 => B(26), A2 => n21, B1 => A(26), B2 => n9, ZN 
                           => n66);
   U94 : AOI22_X1 port map( A1 => D(26), A2 => n7, B1 => C(26), B2 => n5, ZN =>
                           n65);
   U95 : NAND2_X1 port map( A1 => n66, A2 => n65, ZN => Z(26));
   U96 : AOI22_X1 port map( A1 => B(27), A2 => n21, B1 => A(27), B2 => n9, ZN 
                           => n70);
   U97 : AOI22_X1 port map( A1 => D(27), A2 => n7, B1 => C(27), B2 => n5, ZN =>
                           n67);
   U98 : NAND2_X1 port map( A1 => n70, A2 => n67, ZN => Z(27));
   U99 : AOI22_X1 port map( A1 => B(28), A2 => n21, B1 => A(28), B2 => n9, ZN 
                           => n72);
   U100 : AOI22_X1 port map( A1 => D(28), A2 => n7, B1 => C(28), B2 => n5, ZN 
                           => n71);
   U101 : NAND2_X1 port map( A1 => n72, A2 => n71, ZN => Z(28));
   U102 : AOI22_X1 port map( A1 => B(29), A2 => n21, B1 => A(29), B2 => n9, ZN 
                           => n74);
   U103 : AOI22_X1 port map( A1 => D(29), A2 => n7, B1 => C(29), B2 => n5, ZN 
                           => n73);
   U104 : NAND2_X1 port map( A1 => n74, A2 => n73, ZN => Z(29));
   U105 : AOI22_X1 port map( A1 => B(30), A2 => n21, B1 => A(30), B2 => n9, ZN 
                           => n76);
   U106 : AOI22_X1 port map( A1 => D(30), A2 => n7, B1 => C(30), B2 => n5, ZN 
                           => n75);
   U107 : NAND2_X1 port map( A1 => n76, A2 => n75, ZN => Z(30));
   U108 : AOI22_X1 port map( A1 => B(31), A2 => n21, B1 => A(31), B2 => n9, ZN 
                           => n78);
   U109 : AOI22_X1 port map( A1 => D(31), A2 => n7, B1 => C(31), B2 => n5, ZN 
                           => n77);
   U110 : NAND2_X1 port map( A1 => n78, A2 => n77, ZN => Z(31));

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_1 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_1;

architecture SYN_bhv of mux41_NBIT32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n145, Z => n72);
   U2 : BUF_X1 port map( A => n145, Z => n73);
   U3 : BUF_X1 port map( A => n146, Z => n75);
   U4 : BUF_X1 port map( A => n146, Z => n76);
   U5 : BUF_X1 port map( A => n145, Z => n74);
   U6 : BUF_X1 port map( A => n146, Z => n77);
   U7 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n145);
   U8 : BUF_X1 port map( A => n147, Z => n78);
   U9 : BUF_X1 port map( A => n147, Z => n79);
   U10 : BUF_X1 port map( A => n144, Z => n1);
   U11 : BUF_X1 port map( A => n144, Z => n70);
   U12 : BUF_X1 port map( A => n147, Z => n80);
   U13 : BUF_X1 port map( A => n144, Z => n71);
   U14 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n146);
   U15 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n144);
   U16 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n82);
   U17 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN =>
                           n137);
   U18 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n139);
   U19 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n141);
   U20 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN =>
                           n149);
   U21 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN 
                           => n131);
   U22 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n85);
   U23 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n87);
   U24 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n91);
   U25 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n93);
   U26 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n95);
   U27 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n99);
   U28 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n101);
   U29 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n103);
   U30 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n109);
   U31 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n111);
   U32 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN 
                           => n113);
   U33 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n117);
   U34 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n119);
   U35 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN 
                           => n121);
   U36 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n125);
   U37 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN 
                           => n129);
   U38 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n147);
   U39 : INV_X1 port map( A => S(0), ZN => n81);
   U40 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN =>
                           n133);
   U41 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN =>
                           n135);
   U42 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n143);
   U43 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN => 
                           n105);
   U44 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN =>
                           n127);
   U45 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n89);
   U46 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n97);
   U47 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN 
                           => n107);
   U48 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN 
                           => n115);
   U49 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n123);
   U50 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(31));
   U51 : NAND2_X1 port map( A1 => n83, A2 => n82, ZN => Z(0));
   U52 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n83);
   U53 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN 
                           => n130);
   U54 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(3));
   U55 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN =>
                           n132);
   U56 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(4));
   U57 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN =>
                           n134);
   U58 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(5));
   U59 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN =>
                           n136);
   U60 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(6));
   U61 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n138);
   U62 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(7));
   U63 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n140);
   U64 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(8));
   U65 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n142);
   U66 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(9));
   U67 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN =>
                           n148);
   U68 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => Z(15));
   U69 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN 
                           => n94);
   U70 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(16));
   U71 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n96);
   U72 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(17));
   U73 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n98);
   U74 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(18));
   U75 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n100);
   U76 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(19));
   U77 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN 
                           => n102);
   U78 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(20));
   U79 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN 
                           => n106);
   U80 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(21));
   U81 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n108);
   U82 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(22));
   U83 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n110);
   U84 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(23));
   U85 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN 
                           => n112);
   U86 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(24));
   U87 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN 
                           => n114);
   U88 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(25));
   U89 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n116);
   U90 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(26));
   U91 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n118);
   U92 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(27));
   U93 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN 
                           => n120);
   U94 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(28));
   U95 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n122);
   U96 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(29));
   U97 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n124);
   U98 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(30));
   U99 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN 
                           => n128);
   U100 : NAND2_X1 port map( A1 => n93, A2 => n92, ZN => Z(14));
   U101 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN
                           => n92);
   U102 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(1));
   U103 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN 
                           => n104);
   U104 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(2));
   U105 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN 
                           => n126);
   U106 : NAND2_X1 port map( A1 => n85, A2 => n84, ZN => Z(10));
   U107 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN
                           => n84);
   U108 : NAND2_X1 port map( A1 => n87, A2 => n86, ZN => Z(11));
   U109 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN
                           => n86);
   U110 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => Z(12));
   U111 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN
                           => n88);
   U112 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => Z(13));
   U113 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN
                           => n90);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT5_2 is

   port( A, B : in std_logic_vector (4 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (4 downto 0));

end mux21_NBIT5_2;

architecture SYN_bhv of mux21_NBIT5_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n14, n15, n16, n17, n18 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => S, Z => n1);
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : INV_X1 port map( A => n17, ZN => Z(3));
   U4 : INV_X1 port map( A => n18, ZN => Z(4));
   U5 : INV_X1 port map( A => n15, ZN => Z(1));
   U6 : INV_X1 port map( A => n16, ZN => Z(2));
   U7 : INV_X1 port map( A => n14, ZN => Z(0));
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => n1, ZN => 
                           n17);
   U9 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => n2, B2 => B(4), ZN => 
                           n18);
   U10 : AOI22_X1 port map( A1 => A(1), A2 => n3, B1 => B(1), B2 => n1, ZN => 
                           n15);
   U11 : AOI22_X1 port map( A1 => A(0), A2 => n3, B1 => B(0), B2 => n1, ZN => 
                           n14);
   U12 : AOI22_X1 port map( A1 => A(2), A2 => n3, B1 => B(2), B2 => n1, ZN => 
                           n16);
   U13 : INV_X1 port map( A => n2, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT5_1 is

   port( A, B : in std_logic_vector (4 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (4 downto 0));

end mux21_NBIT5_1;

architecture SYN_bhv of mux21_NBIT5_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n14, n15, n16, n17, n18 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => S, Z => n1);
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : INV_X1 port map( A => n15, ZN => Z(1));
   U4 : AOI22_X1 port map( A1 => A(1), A2 => n3, B1 => B(1), B2 => n1, ZN => 
                           n15);
   U5 : INV_X1 port map( A => n16, ZN => Z(2));
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n3, B1 => B(2), B2 => n1, ZN => 
                           n16);
   U7 : INV_X1 port map( A => n17, ZN => Z(3));
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => n1, ZN => 
                           n17);
   U9 : INV_X1 port map( A => n18, ZN => Z(4));
   U10 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => n2, B2 => B(4), ZN => 
                           n18);
   U11 : INV_X1 port map( A => n14, ZN => Z(0));
   U12 : AOI22_X1 port map( A1 => A(0), A2 => n3, B1 => B(0), B2 => n1, ZN => 
                           n14);
   U13 : INV_X1 port map( A => n2, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_4 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_4;

architecture SYN_bhv of regn_N5_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n16, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n21);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n17, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n22);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n18, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n23);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n19, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n24);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n20, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n25);
   U2 : OAI21_X1 port map( B1 => n24, B2 => EN, A => n29, ZN => n19);
   U3 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n29);
   U4 : OAI21_X1 port map( B1 => n23, B2 => EN, A => n28, ZN => n18);
   U5 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n28);
   U6 : OAI21_X1 port map( B1 => n21, B2 => EN, A => n26, ZN => n16);
   U7 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n26);
   U8 : OAI21_X1 port map( B1 => n25, B2 => EN, A => n30, ZN => n20);
   U9 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n30);
   U10 : OAI21_X1 port map( B1 => n22, B2 => EN, A => n27, ZN => n17);
   U11 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n27);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_3 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_3;

architecture SYN_bhv of regn_N5_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n16, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n21);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n17, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n22);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n18, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n23);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n19, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n24);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n20, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n25);
   U2 : OAI21_X1 port map( B1 => n22, B2 => EN, A => n27, ZN => n17);
   U3 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n27);
   U4 : OAI21_X1 port map( B1 => n21, B2 => EN, A => n26, ZN => n16);
   U5 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n26);
   U6 : OAI21_X1 port map( B1 => n24, B2 => EN, A => n29, ZN => n19);
   U7 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n29);
   U8 : OAI21_X1 port map( B1 => n23, B2 => EN, A => n28, ZN => n18);
   U9 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n28);
   U10 : OAI21_X1 port map( B1 => n25, B2 => EN, A => n30, ZN => n20);
   U11 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n30);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_2 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_2;

architecture SYN_bhv of regn_N5_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n16, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n21);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n17, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n22);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n18, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n23);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n19, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n24);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n20, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n25);
   U2 : OAI21_X1 port map( B1 => n25, B2 => EN, A => n30, ZN => n20);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n30);
   U4 : OAI21_X1 port map( B1 => n24, B2 => EN, A => n29, ZN => n19);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n29);
   U6 : OAI21_X1 port map( B1 => n22, B2 => EN, A => n27, ZN => n17);
   U7 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n27);
   U8 : OAI21_X1 port map( B1 => n23, B2 => EN, A => n28, ZN => n18);
   U9 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n28);
   U10 : OAI21_X1 port map( B1 => n21, B2 => EN, A => n26, ZN => n16);
   U11 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n26);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_1 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_1;

architecture SYN_bhv of regn_N5_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n16, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n21);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n17, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n22);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n18, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n23);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n19, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n24);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n20, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n25);
   U2 : OAI21_X1 port map( B1 => n25, B2 => EN, A => n30, ZN => n20);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n30);
   U4 : OAI21_X1 port map( B1 => n24, B2 => EN, A => n29, ZN => n19);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n29);
   U6 : OAI21_X1 port map( B1 => n23, B2 => EN, A => n28, ZN => n18);
   U7 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n28);
   U8 : OAI21_X1 port map( B1 => n22, B2 => EN, A => n27, ZN => n17);
   U9 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n27);
   U10 : OAI21_X1 port map( B1 => n21, B2 => EN, A => n26, ZN => n16);
   U11 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n26);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_9 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_9;

architecture SYN_bhv of regn_N32_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U6 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U7 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U10 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U11 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U24 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U25 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U26 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U27 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U28 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U29 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U30 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U31 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U32 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U33 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U34 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U35 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U36 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U37 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U38 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U39 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U40 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U41 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U42 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U43 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U44 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U45 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U46 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U47 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U48 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U49 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U50 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U51 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U52 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U53 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U54 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U55 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U56 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U57 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U58 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U59 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U60 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U61 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U62 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U63 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U64 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U65 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U66 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);
   U67 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U68 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_8 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_8;

architecture SYN_bhv of regn_N32_8 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   DOUT_reg_30_inst : DFFR_X2 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_29_inst : DFFR_X2 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X2 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U6 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U7 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U8 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);
   U9 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U10 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U11 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U12 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U13 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U14 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U15 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U16 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U17 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U18 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U19 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U20 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U21 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U22 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U23 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U24 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U25 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U26 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U27 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U28 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U29 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U30 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U31 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U32 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U33 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U34 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U35 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U36 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U37 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U38 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U39 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U40 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U41 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U42 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U43 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U44 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U45 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U46 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U47 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U48 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U49 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U50 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U51 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U52 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U53 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U54 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U55 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U56 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U57 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U58 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U59 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U60 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U61 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U62 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U63 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U64 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U65 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U66 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_7 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_7;

architecture SYN_bhv of regn_N32_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U6 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U7 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U8 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U9 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U10 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U11 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U12 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U13 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U14 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U15 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U16 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U17 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U18 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U19 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U20 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U21 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U22 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U23 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U24 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U25 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U26 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U27 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U28 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U29 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U30 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U31 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U32 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U33 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U34 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U35 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U36 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U37 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U38 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U39 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U40 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U41 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U42 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U43 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U44 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U45 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U46 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U47 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U48 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U49 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U50 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U51 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U52 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U53 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U54 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U55 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U56 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U57 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U58 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U59 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U60 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U61 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U62 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);
   U63 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U64 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U65 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U66 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U67 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U68 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_6 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_6;

architecture SYN_bhv of regn_N32_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U6 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U7 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U8 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U9 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U10 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U11 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U12 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U13 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U14 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U15 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U16 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U17 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U18 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U19 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U20 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U21 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U22 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U23 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U24 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U25 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U26 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U27 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U28 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U29 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U30 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U31 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U32 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U33 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U34 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U35 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U36 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);
   U37 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U38 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U39 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U40 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U41 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U42 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U43 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U44 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U45 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U46 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U47 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U48 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U49 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U50 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U51 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U52 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U53 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U54 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U55 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U56 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U57 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U58 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U59 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U60 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U61 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U62 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U63 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U64 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U65 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U66 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U67 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U68 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_5 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_5;

architecture SYN_bhv of regn_N32_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_4 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_4;

architecture SYN_bhv of regn_N32_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_3 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_3;

architecture SYN_bhv of regn_N32_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_2 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_2;

architecture SYN_bhv of regn_N32_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_1 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_1;

architecture SYN_bhv of regn_N32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U4 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U6 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U7 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U8 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U9 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U10 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U11 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U12 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U13 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U14 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U15 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U16 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U17 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U18 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U19 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U20 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U21 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U22 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U23 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U24 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U25 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U26 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U27 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U28 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U29 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U30 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U31 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U32 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U33 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U34 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U35 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U36 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U37 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U38 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U39 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U40 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U41 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U42 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U43 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U44 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U45 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U46 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U47 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U48 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U49 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U50 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U51 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U52 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U53 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U54 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U55 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U56 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U57 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U58 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U59 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U60 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U61 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U62 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U63 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U64 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U65 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);
   U66 : BUF_X1 port map( A => RST, Z => n97);
   U67 : BUF_X1 port map( A => RST, Z => n98);
   U68 : BUF_X1 port map( A => RST, Z => n99);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_6 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_6;

architecture SYN_bhv of mux21_NBIT32_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104 : std_logic;

begin
   
   U1 : BUF_X2 port map( A => n2, Z => n7);
   U2 : INV_X2 port map( A => S, ZN => n3);
   U3 : CLKBUF_X1 port map( A => S, Z => n2);
   U4 : CLKBUF_X1 port map( A => S, Z => n1);
   U5 : CLKBUF_X1 port map( A => n4, Z => n8);
   U6 : CLKBUF_X1 port map( A => n1, Z => n4);
   U7 : BUF_X1 port map( A => n1, Z => n6);
   U8 : BUF_X1 port map( A => n1, Z => n5);
   U9 : INV_X1 port map( A => n95, ZN => Z(2));
   U10 : AOI22_X1 port map( A1 => A(2), A2 => n3, B1 => B(2), B2 => n5, ZN => 
                           n95);
   U11 : INV_X1 port map( A => n84, ZN => Z(1));
   U12 : AOI22_X1 port map( A1 => A(1), A2 => n3, B1 => B(1), B2 => n7, ZN => 
                           n84);
   U13 : INV_X1 port map( A => n73, ZN => Z(0));
   U14 : AOI22_X1 port map( A1 => A(0), A2 => n3, B1 => B(0), B2 => n8, ZN => 
                           n73);
   U15 : INV_X1 port map( A => n98, ZN => Z(3));
   U16 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => n5, ZN => 
                           n98);
   U17 : INV_X1 port map( A => n99, ZN => Z(4));
   U18 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => n5, ZN => 
                           n99);
   U19 : INV_X1 port map( A => n100, ZN => Z(5));
   U20 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => n4, ZN => 
                           n100);
   U21 : INV_X1 port map( A => n101, ZN => Z(6));
   U22 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => n4, ZN => 
                           n101);
   U23 : INV_X1 port map( A => n102, ZN => Z(7));
   U24 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => n4, ZN => 
                           n102);
   U25 : INV_X1 port map( A => n103, ZN => Z(8));
   U26 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => n4, ZN => 
                           n103);
   U27 : INV_X1 port map( A => n74, ZN => Z(10));
   U28 : AOI22_X1 port map( A1 => A(10), A2 => n3, B1 => B(10), B2 => n8, ZN =>
                           n74);
   U29 : INV_X1 port map( A => n75, ZN => Z(11));
   U30 : AOI22_X1 port map( A1 => A(11), A2 => n3, B1 => B(11), B2 => n8, ZN =>
                           n75);
   U31 : INV_X1 port map( A => n76, ZN => Z(12));
   U32 : AOI22_X1 port map( A1 => A(12), A2 => n3, B1 => B(12), B2 => n8, ZN =>
                           n76);
   U33 : INV_X1 port map( A => n77, ZN => Z(13));
   U34 : AOI22_X1 port map( A1 => A(13), A2 => n3, B1 => B(13), B2 => n1, ZN =>
                           n77);
   U35 : INV_X1 port map( A => n78, ZN => Z(14));
   U36 : AOI22_X1 port map( A1 => A(14), A2 => n3, B1 => B(14), B2 => n2, ZN =>
                           n78);
   U37 : INV_X1 port map( A => n79, ZN => Z(15));
   U38 : AOI22_X1 port map( A1 => A(15), A2 => n3, B1 => B(15), B2 => n2, ZN =>
                           n79);
   U39 : INV_X1 port map( A => n80, ZN => Z(16));
   U40 : AOI22_X1 port map( A1 => A(16), A2 => n3, B1 => B(16), B2 => n2, ZN =>
                           n80);
   U41 : INV_X1 port map( A => n81, ZN => Z(17));
   U42 : AOI22_X1 port map( A1 => A(17), A2 => n3, B1 => B(17), B2 => n1, ZN =>
                           n81);
   U43 : INV_X1 port map( A => n82, ZN => Z(18));
   U44 : AOI22_X1 port map( A1 => A(18), A2 => n3, B1 => B(18), B2 => n2, ZN =>
                           n82);
   U45 : INV_X1 port map( A => n83, ZN => Z(19));
   U46 : AOI22_X1 port map( A1 => A(19), A2 => n3, B1 => B(19), B2 => n1, ZN =>
                           n83);
   U47 : INV_X1 port map( A => n85, ZN => Z(20));
   U48 : AOI22_X1 port map( A1 => A(20), A2 => n3, B1 => B(20), B2 => n2, ZN =>
                           n85);
   U49 : INV_X1 port map( A => n86, ZN => Z(21));
   U50 : AOI22_X1 port map( A1 => A(21), A2 => n3, B1 => B(21), B2 => n6, ZN =>
                           n86);
   U51 : INV_X1 port map( A => n87, ZN => Z(22));
   U52 : AOI22_X1 port map( A1 => A(22), A2 => n3, B1 => B(22), B2 => n7, ZN =>
                           n87);
   U53 : INV_X1 port map( A => n88, ZN => Z(23));
   U54 : AOI22_X1 port map( A1 => A(23), A2 => n3, B1 => B(23), B2 => n7, ZN =>
                           n88);
   U55 : INV_X1 port map( A => n89, ZN => Z(24));
   U56 : AOI22_X1 port map( A1 => A(24), A2 => n3, B1 => B(24), B2 => n7, ZN =>
                           n89);
   U57 : INV_X1 port map( A => n90, ZN => Z(25));
   U58 : AOI22_X1 port map( A1 => A(25), A2 => n3, B1 => B(25), B2 => n7, ZN =>
                           n90);
   U59 : INV_X1 port map( A => n91, ZN => Z(26));
   U60 : AOI22_X1 port map( A1 => A(26), A2 => n3, B1 => B(26), B2 => n6, ZN =>
                           n91);
   U61 : INV_X1 port map( A => n92, ZN => Z(27));
   U62 : AOI22_X1 port map( A1 => A(27), A2 => n3, B1 => B(27), B2 => n6, ZN =>
                           n92);
   U63 : INV_X1 port map( A => n93, ZN => Z(28));
   U64 : AOI22_X1 port map( A1 => A(28), A2 => n3, B1 => B(28), B2 => n6, ZN =>
                           n93);
   U65 : INV_X1 port map( A => n94, ZN => Z(29));
   U66 : AOI22_X1 port map( A1 => A(29), A2 => n3, B1 => B(29), B2 => n6, ZN =>
                           n94);
   U67 : INV_X1 port map( A => n96, ZN => Z(30));
   U68 : AOI22_X1 port map( A1 => A(30), A2 => n3, B1 => B(30), B2 => n5, ZN =>
                           n96);
   U69 : INV_X1 port map( A => n97, ZN => Z(31));
   U70 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => n5, ZN =>
                           n97);
   U71 : INV_X1 port map( A => n104, ZN => Z(9));
   U72 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => n8, B2 => B(9), ZN => 
                           n104);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_5;

architecture SYN_bhv of mux21_NBIT32_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   U1 : BUF_X2 port map( A => S, Z => n3);
   U2 : INV_X2 port map( A => n3, ZN => n1);
   U3 : BUF_X1 port map( A => S, Z => n2);
   U4 : INV_X1 port map( A => n86, ZN => Z(26));
   U5 : INV_X1 port map( A => n91, ZN => Z(30));
   U6 : INV_X1 port map( A => n88, ZN => Z(28));
   U7 : INV_X1 port map( A => n92, ZN => Z(31));
   U8 : INV_X1 port map( A => n87, ZN => Z(27));
   U9 : INV_X1 port map( A => n89, ZN => Z(29));
   U10 : INV_X1 port map( A => n79, ZN => Z(1));
   U11 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => n3, ZN => 
                           n79);
   U12 : INV_X1 port map( A => n90, ZN => Z(2));
   U13 : AOI22_X1 port map( A1 => A(2), A2 => n1, B1 => B(2), B2 => n2, ZN => 
                           n90);
   U14 : INV_X1 port map( A => n93, ZN => Z(3));
   U15 : AOI22_X1 port map( A1 => A(3), A2 => n1, B1 => B(3), B2 => n2, ZN => 
                           n93);
   U16 : INV_X1 port map( A => n94, ZN => Z(4));
   U17 : AOI22_X1 port map( A1 => A(4), A2 => n1, B1 => B(4), B2 => n2, ZN => 
                           n94);
   U18 : INV_X1 port map( A => n95, ZN => Z(5));
   U19 : AOI22_X1 port map( A1 => A(5), A2 => n1, B1 => B(5), B2 => n3, ZN => 
                           n95);
   U20 : INV_X1 port map( A => n96, ZN => Z(6));
   U21 : AOI22_X1 port map( A1 => A(6), A2 => n1, B1 => B(6), B2 => n3, ZN => 
                           n96);
   U22 : INV_X1 port map( A => n97, ZN => Z(7));
   U23 : AOI22_X1 port map( A1 => A(7), A2 => n1, B1 => B(7), B2 => n3, ZN => 
                           n97);
   U24 : INV_X1 port map( A => n98, ZN => Z(8));
   U25 : AOI22_X1 port map( A1 => A(8), A2 => n1, B1 => B(8), B2 => n3, ZN => 
                           n98);
   U26 : INV_X1 port map( A => n69, ZN => Z(10));
   U27 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => n3, ZN =>
                           n69);
   U28 : INV_X1 port map( A => n70, ZN => Z(11));
   U29 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => n3, ZN =>
                           n70);
   U30 : INV_X1 port map( A => n71, ZN => Z(12));
   U31 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => n3, ZN =>
                           n71);
   U32 : INV_X1 port map( A => n72, ZN => Z(13));
   U33 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => n3, ZN =>
                           n72);
   U34 : INV_X1 port map( A => n73, ZN => Z(14));
   U35 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => n3, ZN =>
                           n73);
   U36 : INV_X1 port map( A => n74, ZN => Z(15));
   U37 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => n3, ZN =>
                           n74);
   U38 : INV_X1 port map( A => n75, ZN => Z(16));
   U39 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => n3, ZN =>
                           n75);
   U40 : INV_X1 port map( A => n76, ZN => Z(17));
   U41 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => n3, ZN =>
                           n76);
   U42 : INV_X1 port map( A => n77, ZN => Z(18));
   U43 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => n3, ZN =>
                           n77);
   U44 : INV_X1 port map( A => n78, ZN => Z(19));
   U45 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => n3, ZN =>
                           n78);
   U46 : INV_X1 port map( A => n80, ZN => Z(20));
   U47 : AOI22_X1 port map( A1 => A(20), A2 => n1, B1 => B(20), B2 => n3, ZN =>
                           n80);
   U48 : INV_X1 port map( A => n81, ZN => Z(21));
   U49 : AOI22_X1 port map( A1 => A(21), A2 => n1, B1 => B(21), B2 => n3, ZN =>
                           n81);
   U50 : INV_X1 port map( A => n82, ZN => Z(22));
   U51 : AOI22_X1 port map( A1 => A(22), A2 => n1, B1 => B(22), B2 => n3, ZN =>
                           n82);
   U52 : INV_X1 port map( A => n83, ZN => Z(23));
   U53 : AOI22_X1 port map( A1 => A(23), A2 => n1, B1 => B(23), B2 => n3, ZN =>
                           n83);
   U54 : INV_X1 port map( A => n84, ZN => Z(24));
   U55 : AOI22_X1 port map( A1 => A(24), A2 => n1, B1 => B(24), B2 => n3, ZN =>
                           n84);
   U56 : INV_X1 port map( A => n85, ZN => Z(25));
   U57 : AOI22_X1 port map( A1 => A(25), A2 => n1, B1 => B(25), B2 => n3, ZN =>
                           n85);
   U58 : INV_X1 port map( A => n99, ZN => Z(9));
   U59 : AOI22_X1 port map( A1 => A(9), A2 => n1, B1 => n3, B2 => B(9), ZN => 
                           n99);
   U60 : INV_X1 port map( A => n68, ZN => Z(0));
   U61 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => n3, ZN => 
                           n68);
   U62 : AOI22_X1 port map( A1 => A(29), A2 => n1, B1 => B(29), B2 => n3, ZN =>
                           n89);
   U63 : AOI22_X1 port map( A1 => A(30), A2 => n1, B1 => B(30), B2 => n3, ZN =>
                           n91);
   U64 : AOI22_X1 port map( A1 => A(27), A2 => n1, B1 => B(27), B2 => n3, ZN =>
                           n87);
   U65 : AOI22_X1 port map( A1 => A(28), A2 => n1, B1 => B(28), B2 => n3, ZN =>
                           n88);
   U66 : AOI22_X1 port map( A1 => A(26), A2 => n1, B1 => B(26), B2 => n3, ZN =>
                           n86);
   U67 : AOI22_X1 port map( A1 => A(31), A2 => n1, B1 => B(31), B2 => n2, ZN =>
                           n92);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_4;

architecture SYN_bhv of mux21_NBIT32_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n68, Z => n1);
   U2 : BUF_X1 port map( A => n68, Z => n2);
   U3 : BUF_X1 port map( A => n68, Z => n3);
   U4 : INV_X1 port map( A => n69, ZN => Z(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => S, ZN => n69
                           );
   U6 : INV_X1 port map( A => n81, ZN => Z(20));
   U7 : AOI22_X1 port map( A1 => A(20), A2 => n2, B1 => B(20), B2 => S, ZN => 
                           n81);
   U8 : INV_X1 port map( A => n85, ZN => Z(24));
   U9 : AOI22_X1 port map( A1 => A(24), A2 => n2, B1 => B(24), B2 => S, ZN => 
                           n85);
   U10 : INV_X1 port map( A => n97, ZN => Z(6));
   U11 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => S, ZN => 
                           n97);
   U12 : INV_X1 port map( A => n70, ZN => Z(10));
   U13 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => S, ZN => 
                           n70);
   U14 : INV_X1 port map( A => n73, ZN => Z(13));
   U15 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => S, ZN => 
                           n73);
   U16 : INV_X1 port map( A => n77, ZN => Z(17));
   U17 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => S, ZN => 
                           n77);
   U18 : INV_X1 port map( A => n89, ZN => Z(28));
   U19 : AOI22_X1 port map( A1 => A(28), A2 => n2, B1 => B(28), B2 => S, ZN => 
                           n89);
   U20 : INV_X1 port map( A => n93, ZN => Z(31));
   U21 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => S, ZN => 
                           n93);
   U22 : INV_X1 port map( A => n94, ZN => Z(3));
   U23 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => S, ZN => 
                           n94);
   U24 : INV_X1 port map( A => n98, ZN => Z(7));
   U25 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => S, ZN => 
                           n98);
   U26 : INV_X1 port map( A => n74, ZN => Z(14));
   U27 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => S, ZN => 
                           n74);
   U28 : INV_X1 port map( A => n78, ZN => Z(18));
   U29 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => S, ZN => 
                           n78);
   U30 : INV_X1 port map( A => n82, ZN => Z(21));
   U31 : AOI22_X1 port map( A1 => A(21), A2 => n2, B1 => B(21), B2 => S, ZN => 
                           n82);
   U32 : INV_X1 port map( A => n86, ZN => Z(25));
   U33 : AOI22_X1 port map( A1 => A(25), A2 => n2, B1 => B(25), B2 => S, ZN => 
                           n86);
   U34 : INV_X1 port map( A => n90, ZN => Z(29));
   U35 : AOI22_X1 port map( A1 => A(29), A2 => n2, B1 => B(29), B2 => S, ZN => 
                           n90);
   U36 : INV_X1 port map( A => n71, ZN => Z(11));
   U37 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => S, ZN => 
                           n71);
   U38 : INV_X1 port map( A => n91, ZN => Z(2));
   U39 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => S, ZN => 
                           n91);
   U40 : INV_X1 port map( A => n95, ZN => Z(4));
   U41 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => S, ZN => 
                           n95);
   U42 : INV_X1 port map( A => n99, ZN => Z(8));
   U43 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => S, ZN => 
                           n99);
   U44 : INV_X1 port map( A => n75, ZN => Z(15));
   U45 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => S, ZN => 
                           n75);
   U46 : INV_X1 port map( A => n79, ZN => Z(19));
   U47 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => S, ZN => 
                           n79);
   U48 : INV_X1 port map( A => n83, ZN => Z(22));
   U49 : AOI22_X1 port map( A1 => A(22), A2 => n2, B1 => B(22), B2 => S, ZN => 
                           n83);
   U50 : INV_X1 port map( A => n87, ZN => Z(26));
   U51 : AOI22_X1 port map( A1 => A(26), A2 => n2, B1 => B(26), B2 => S, ZN => 
                           n87);
   U52 : INV_X1 port map( A => n80, ZN => Z(1));
   U53 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => S, ZN => 
                           n80);
   U54 : INV_X1 port map( A => n96, ZN => Z(5));
   U55 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => S, ZN => 
                           n96);
   U56 : INV_X1 port map( A => n72, ZN => Z(12));
   U57 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => S, ZN => 
                           n72);
   U58 : INV_X1 port map( A => n76, ZN => Z(16));
   U59 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => S, ZN => 
                           n76);
   U60 : INV_X1 port map( A => n84, ZN => Z(23));
   U61 : AOI22_X1 port map( A1 => A(23), A2 => n2, B1 => B(23), B2 => S, ZN => 
                           n84);
   U62 : INV_X1 port map( A => n88, ZN => Z(27));
   U63 : AOI22_X1 port map( A1 => A(27), A2 => n2, B1 => B(27), B2 => S, ZN => 
                           n88);
   U64 : INV_X1 port map( A => n92, ZN => Z(30));
   U65 : AOI22_X1 port map( A1 => A(30), A2 => n2, B1 => B(30), B2 => S, ZN => 
                           n92);
   U66 : INV_X1 port map( A => n100, ZN => Z(9));
   U67 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => S, B2 => B(9), ZN => 
                           n100);
   U68 : INV_X1 port map( A => S, ZN => n68);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_3;

architecture SYN_bhv of mux21_NBIT32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n68, Z => n1);
   U2 : BUF_X1 port map( A => n68, Z => n2);
   U3 : BUF_X1 port map( A => n68, Z => n3);
   U4 : INV_X1 port map( A => n100, ZN => Z(9));
   U5 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => S, B2 => B(9), ZN => 
                           n100);
   U6 : INV_X1 port map( A => n82, ZN => Z(21));
   U7 : AOI22_X1 port map( A1 => A(21), A2 => n2, B1 => B(21), B2 => S, ZN => 
                           n82);
   U8 : INV_X1 port map( A => n83, ZN => Z(22));
   U9 : AOI22_X1 port map( A1 => A(22), A2 => n2, B1 => B(22), B2 => S, ZN => 
                           n83);
   U10 : INV_X1 port map( A => n84, ZN => Z(23));
   U11 : AOI22_X1 port map( A1 => A(23), A2 => n2, B1 => B(23), B2 => S, ZN => 
                           n84);
   U12 : INV_X1 port map( A => n77, ZN => Z(17));
   U13 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => S, ZN => 
                           n77);
   U14 : INV_X1 port map( A => n78, ZN => Z(18));
   U15 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => S, ZN => 
                           n78);
   U16 : INV_X1 port map( A => n79, ZN => Z(19));
   U17 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => S, ZN => 
                           n79);
   U18 : INV_X1 port map( A => n80, ZN => Z(1));
   U19 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => S, ZN => 
                           n80);
   U20 : INV_X1 port map( A => n73, ZN => Z(13));
   U21 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => S, ZN => 
                           n73);
   U22 : INV_X1 port map( A => n74, ZN => Z(14));
   U23 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => S, ZN => 
                           n74);
   U24 : INV_X1 port map( A => n75, ZN => Z(15));
   U25 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => S, ZN => 
                           n75);
   U26 : INV_X1 port map( A => n76, ZN => Z(16));
   U27 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => S, ZN => 
                           n76);
   U28 : INV_X1 port map( A => n69, ZN => Z(0));
   U29 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => S, ZN => 
                           n69);
   U30 : INV_X1 port map( A => n72, ZN => Z(12));
   U31 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => S, ZN => 
                           n72);
   U32 : INV_X1 port map( A => n97, ZN => Z(6));
   U33 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => S, ZN => 
                           n97);
   U34 : INV_X1 port map( A => n98, ZN => Z(7));
   U35 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => S, ZN => 
                           n98);
   U36 : INV_X1 port map( A => n99, ZN => Z(8));
   U37 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => S, ZN => 
                           n99);
   U38 : INV_X1 port map( A => n94, ZN => Z(3));
   U39 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => S, ZN => 
                           n94);
   U40 : INV_X1 port map( A => n95, ZN => Z(4));
   U41 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => S, ZN => 
                           n95);
   U42 : INV_X1 port map( A => n96, ZN => Z(5));
   U43 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => S, ZN => 
                           n96);
   U44 : INV_X1 port map( A => n89, ZN => Z(28));
   U45 : AOI22_X1 port map( A1 => A(28), A2 => n2, B1 => B(28), B2 => S, ZN => 
                           n89);
   U46 : INV_X1 port map( A => n90, ZN => Z(29));
   U47 : AOI22_X1 port map( A1 => A(29), A2 => n2, B1 => B(29), B2 => S, ZN => 
                           n90);
   U48 : INV_X1 port map( A => n91, ZN => Z(2));
   U49 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => S, ZN => 
                           n91);
   U50 : INV_X1 port map( A => n92, ZN => Z(30));
   U51 : AOI22_X1 port map( A1 => A(30), A2 => n2, B1 => B(30), B2 => S, ZN => 
                           n92);
   U52 : INV_X1 port map( A => n86, ZN => Z(25));
   U53 : AOI22_X1 port map( A1 => A(25), A2 => n2, B1 => B(25), B2 => S, ZN => 
                           n86);
   U54 : INV_X1 port map( A => n87, ZN => Z(26));
   U55 : AOI22_X1 port map( A1 => A(26), A2 => n2, B1 => B(26), B2 => S, ZN => 
                           n87);
   U56 : INV_X1 port map( A => n88, ZN => Z(27));
   U57 : AOI22_X1 port map( A1 => A(27), A2 => n2, B1 => B(27), B2 => S, ZN => 
                           n88);
   U58 : INV_X1 port map( A => n93, ZN => Z(31));
   U59 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => S, ZN => 
                           n93);
   U60 : INV_X1 port map( A => n81, ZN => Z(20));
   U61 : AOI22_X1 port map( A1 => A(20), A2 => n2, B1 => B(20), B2 => S, ZN => 
                           n81);
   U62 : INV_X1 port map( A => n70, ZN => Z(10));
   U63 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => S, ZN => 
                           n70);
   U64 : INV_X1 port map( A => n85, ZN => Z(24));
   U65 : AOI22_X1 port map( A1 => A(24), A2 => n2, B1 => B(24), B2 => S, ZN => 
                           n85);
   U66 : INV_X1 port map( A => n71, ZN => Z(11));
   U67 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => S, ZN => 
                           n71);
   U68 : INV_X1 port map( A => S, ZN => n68);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_2;

architecture SYN_bhv of mux21_NBIT32_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => n4);
   U2 : INV_X1 port map( A => n14, ZN => n5);
   U3 : BUF_X1 port map( A => n1, Z => n6);
   U4 : BUF_X1 port map( A => n3, Z => n12);
   U5 : BUF_X1 port map( A => n2, Z => n11);
   U6 : BUF_X1 port map( A => n2, Z => n9);
   U7 : BUF_X1 port map( A => n1, Z => n8);
   U8 : BUF_X1 port map( A => n2, Z => n10);
   U9 : BUF_X1 port map( A => n1, Z => n7);
   U10 : BUF_X1 port map( A => n3, Z => n14);
   U11 : BUF_X1 port map( A => n3, Z => n13);
   U12 : INV_X1 port map( A => n103, ZN => Z(31));
   U13 : AOI22_X1 port map( A1 => A(31), A2 => n4, B1 => B(31), B2 => n7, ZN =>
                           n103);
   U14 : BUF_X1 port map( A => S, Z => n3);
   U15 : BUF_X1 port map( A => S, Z => n2);
   U16 : BUF_X1 port map( A => S, Z => n1);
   U17 : INV_X1 port map( A => n79, ZN => Z(0));
   U18 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => n13, ZN => 
                           n79);
   U19 : INV_X1 port map( A => n104, ZN => Z(3));
   U20 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => B(3), B2 => n7, ZN => 
                           n104);
   U21 : INV_X1 port map( A => n105, ZN => Z(4));
   U22 : AOI22_X1 port map( A1 => A(4), A2 => n4, B1 => B(4), B2 => n7, ZN => 
                           n105);
   U23 : INV_X1 port map( A => n106, ZN => Z(5));
   U24 : AOI22_X1 port map( A1 => A(5), A2 => n5, B1 => B(5), B2 => n6, ZN => 
                           n106);
   U25 : INV_X1 port map( A => n107, ZN => Z(6));
   U26 : AOI22_X1 port map( A1 => A(6), A2 => n4, B1 => B(6), B2 => n6, ZN => 
                           n107);
   U27 : INV_X1 port map( A => n108, ZN => Z(7));
   U28 : AOI22_X1 port map( A1 => A(7), A2 => n5, B1 => B(7), B2 => n6, ZN => 
                           n108);
   U29 : INV_X1 port map( A => n109, ZN => Z(8));
   U30 : AOI22_X1 port map( A1 => A(8), A2 => n4, B1 => B(8), B2 => n6, ZN => 
                           n109);
   U31 : INV_X1 port map( A => n110, ZN => Z(9));
   U32 : AOI22_X1 port map( A1 => A(9), A2 => n5, B1 => n13, B2 => B(9), ZN => 
                           n110);
   U33 : INV_X1 port map( A => n85, ZN => Z(15));
   U34 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n12, ZN 
                           => n85);
   U35 : INV_X1 port map( A => n86, ZN => Z(16));
   U36 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => B(16), B2 => n11, ZN 
                           => n86);
   U37 : INV_X1 port map( A => n87, ZN => Z(17));
   U38 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n11, ZN 
                           => n87);
   U39 : INV_X1 port map( A => n88, ZN => Z(18));
   U40 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => B(18), B2 => n11, ZN 
                           => n88);
   U41 : INV_X1 port map( A => n89, ZN => Z(19));
   U42 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => B(19), B2 => n11, ZN 
                           => n89);
   U43 : INV_X1 port map( A => n91, ZN => Z(20));
   U44 : AOI22_X1 port map( A1 => A(20), A2 => n5, B1 => B(20), B2 => n10, ZN 
                           => n91);
   U45 : INV_X1 port map( A => n92, ZN => Z(21));
   U46 : AOI22_X1 port map( A1 => A(21), A2 => n5, B1 => B(21), B2 => n10, ZN 
                           => n92);
   U47 : INV_X1 port map( A => n93, ZN => Z(22));
   U48 : AOI22_X1 port map( A1 => A(22), A2 => n5, B1 => B(22), B2 => n9, ZN =>
                           n93);
   U49 : INV_X1 port map( A => n94, ZN => Z(23));
   U50 : AOI22_X1 port map( A1 => A(23), A2 => n5, B1 => B(23), B2 => n9, ZN =>
                           n94);
   U51 : INV_X1 port map( A => n95, ZN => Z(24));
   U52 : AOI22_X1 port map( A1 => A(24), A2 => n5, B1 => B(24), B2 => n9, ZN =>
                           n95);
   U53 : INV_X1 port map( A => n96, ZN => Z(25));
   U54 : AOI22_X1 port map( A1 => A(25), A2 => n5, B1 => B(25), B2 => n9, ZN =>
                           n96);
   U55 : INV_X1 port map( A => n97, ZN => Z(26));
   U56 : AOI22_X1 port map( A1 => A(26), A2 => n5, B1 => B(26), B2 => n8, ZN =>
                           n97);
   U57 : INV_X1 port map( A => n98, ZN => Z(27));
   U58 : AOI22_X1 port map( A1 => A(27), A2 => n5, B1 => B(27), B2 => n8, ZN =>
                           n98);
   U59 : INV_X1 port map( A => n99, ZN => Z(28));
   U60 : AOI22_X1 port map( A1 => A(28), A2 => n5, B1 => B(28), B2 => n8, ZN =>
                           n99);
   U61 : INV_X1 port map( A => n100, ZN => Z(29));
   U62 : AOI22_X1 port map( A1 => A(29), A2 => n5, B1 => B(29), B2 => n8, ZN =>
                           n100);
   U63 : INV_X1 port map( A => n102, ZN => Z(30));
   U64 : AOI22_X1 port map( A1 => A(30), A2 => n5, B1 => B(30), B2 => n10, ZN 
                           => n102);
   U65 : INV_X1 port map( A => n84, ZN => Z(14));
   U66 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n12, ZN 
                           => n84);
   U67 : INV_X1 port map( A => n90, ZN => Z(1));
   U68 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n10, ZN => 
                           n90);
   U69 : INV_X1 port map( A => n101, ZN => Z(2));
   U70 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           n101);
   U71 : INV_X1 port map( A => n80, ZN => Z(10));
   U72 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => B(10), B2 => n13, ZN 
                           => n80);
   U73 : INV_X1 port map( A => n81, ZN => Z(11));
   U74 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => B(11), B2 => n13, ZN 
                           => n81);
   U75 : INV_X1 port map( A => n82, ZN => Z(12));
   U76 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => B(12), B2 => n12, ZN 
                           => n82);
   U77 : INV_X1 port map( A => n83, ZN => Z(13));
   U78 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n12, ZN 
                           => n83);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_1;

architecture SYN_bhv of mux21_NBIT32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => n4);
   U2 : INV_X1 port map( A => n14, ZN => n5);
   U3 : BUF_X1 port map( A => n1, Z => n6);
   U4 : BUF_X1 port map( A => n3, Z => n12);
   U5 : BUF_X1 port map( A => n2, Z => n11);
   U6 : BUF_X1 port map( A => n2, Z => n9);
   U7 : BUF_X1 port map( A => n1, Z => n8);
   U8 : BUF_X1 port map( A => n2, Z => n10);
   U9 : BUF_X1 port map( A => n1, Z => n7);
   U10 : BUF_X1 port map( A => n3, Z => n14);
   U11 : BUF_X1 port map( A => n3, Z => n13);
   U12 : BUF_X1 port map( A => S, Z => n3);
   U13 : BUF_X1 port map( A => S, Z => n2);
   U14 : BUF_X1 port map( A => S, Z => n1);
   U15 : INV_X1 port map( A => n79, ZN => Z(0));
   U16 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => n13, ZN => 
                           n79);
   U17 : INV_X1 port map( A => n90, ZN => Z(1));
   U18 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n10, ZN => 
                           n90);
   U19 : INV_X1 port map( A => n101, ZN => Z(2));
   U20 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           n101);
   U21 : INV_X1 port map( A => n104, ZN => Z(3));
   U22 : AOI22_X1 port map( A1 => A(3), A2 => n4, B1 => B(3), B2 => n7, ZN => 
                           n104);
   U23 : INV_X1 port map( A => n105, ZN => Z(4));
   U24 : AOI22_X1 port map( A1 => A(4), A2 => n5, B1 => B(4), B2 => n7, ZN => 
                           n105);
   U25 : INV_X1 port map( A => n106, ZN => Z(5));
   U26 : AOI22_X1 port map( A1 => A(5), A2 => n4, B1 => B(5), B2 => n6, ZN => 
                           n106);
   U27 : INV_X1 port map( A => n107, ZN => Z(6));
   U28 : AOI22_X1 port map( A1 => A(6), A2 => n5, B1 => B(6), B2 => n6, ZN => 
                           n107);
   U29 : INV_X1 port map( A => n108, ZN => Z(7));
   U30 : AOI22_X1 port map( A1 => A(7), A2 => n4, B1 => B(7), B2 => n6, ZN => 
                           n108);
   U31 : INV_X1 port map( A => n109, ZN => Z(8));
   U32 : AOI22_X1 port map( A1 => A(8), A2 => n5, B1 => B(8), B2 => n6, ZN => 
                           n109);
   U33 : INV_X1 port map( A => n110, ZN => Z(9));
   U34 : AOI22_X1 port map( A1 => A(9), A2 => n4, B1 => n13, B2 => B(9), ZN => 
                           n110);
   U35 : INV_X1 port map( A => n80, ZN => Z(10));
   U36 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => B(10), B2 => n13, ZN 
                           => n80);
   U37 : INV_X1 port map( A => n81, ZN => Z(11));
   U38 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => B(11), B2 => n13, ZN 
                           => n81);
   U39 : INV_X1 port map( A => n82, ZN => Z(12));
   U40 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => B(12), B2 => n12, ZN 
                           => n82);
   U41 : INV_X1 port map( A => n83, ZN => Z(13));
   U42 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n12, ZN 
                           => n83);
   U43 : INV_X1 port map( A => n84, ZN => Z(14));
   U44 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n12, ZN 
                           => n84);
   U45 : INV_X1 port map( A => n85, ZN => Z(15));
   U46 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n12, ZN 
                           => n85);
   U47 : INV_X1 port map( A => n86, ZN => Z(16));
   U48 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => B(16), B2 => n11, ZN 
                           => n86);
   U49 : INV_X1 port map( A => n87, ZN => Z(17));
   U50 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n11, ZN 
                           => n87);
   U51 : INV_X1 port map( A => n88, ZN => Z(18));
   U52 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => B(18), B2 => n11, ZN 
                           => n88);
   U53 : INV_X1 port map( A => n89, ZN => Z(19));
   U54 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => B(19), B2 => n11, ZN 
                           => n89);
   U55 : INV_X1 port map( A => n91, ZN => Z(20));
   U56 : AOI22_X1 port map( A1 => A(20), A2 => n5, B1 => B(20), B2 => n10, ZN 
                           => n91);
   U57 : INV_X1 port map( A => n92, ZN => Z(21));
   U58 : AOI22_X1 port map( A1 => A(21), A2 => n5, B1 => B(21), B2 => n10, ZN 
                           => n92);
   U59 : INV_X1 port map( A => n93, ZN => Z(22));
   U60 : AOI22_X1 port map( A1 => A(22), A2 => n5, B1 => B(22), B2 => n9, ZN =>
                           n93);
   U61 : INV_X1 port map( A => n94, ZN => Z(23));
   U62 : AOI22_X1 port map( A1 => A(23), A2 => n5, B1 => B(23), B2 => n9, ZN =>
                           n94);
   U63 : INV_X1 port map( A => n95, ZN => Z(24));
   U64 : AOI22_X1 port map( A1 => A(24), A2 => n5, B1 => B(24), B2 => n9, ZN =>
                           n95);
   U65 : INV_X1 port map( A => n96, ZN => Z(25));
   U66 : AOI22_X1 port map( A1 => A(25), A2 => n5, B1 => B(25), B2 => n9, ZN =>
                           n96);
   U67 : INV_X1 port map( A => n97, ZN => Z(26));
   U68 : AOI22_X1 port map( A1 => A(26), A2 => n5, B1 => B(26), B2 => n8, ZN =>
                           n97);
   U69 : INV_X1 port map( A => n98, ZN => Z(27));
   U70 : AOI22_X1 port map( A1 => A(27), A2 => n5, B1 => B(27), B2 => n8, ZN =>
                           n98);
   U71 : INV_X1 port map( A => n99, ZN => Z(28));
   U72 : AOI22_X1 port map( A1 => A(28), A2 => n5, B1 => B(28), B2 => n8, ZN =>
                           n99);
   U73 : INV_X1 port map( A => n100, ZN => Z(29));
   U74 : AOI22_X1 port map( A1 => A(29), A2 => n5, B1 => B(29), B2 => n8, ZN =>
                           n100);
   U75 : INV_X1 port map( A => n102, ZN => Z(30));
   U76 : AOI22_X1 port map( A1 => A(30), A2 => n5, B1 => B(30), B2 => n10, ZN 
                           => n102);
   U77 : INV_X1 port map( A => n103, ZN => Z(31));
   U78 : AOI22_X1 port map( A1 => A(31), A2 => n5, B1 => B(31), B2 => n7, ZN =>
                           n103);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ff_2 is

   port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);

end ff_2;

architecture SYN_bhv of ff_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CLK, RN => RST, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => EN, A => n6, ZN => n4);
   U3 : NAND2_X1 port map( A1 => EN, A2 => D, ZN => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ff_1 is

   port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);

end ff_1;

architecture SYN_bhv of ff_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CLK, RN => RST, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => EN, A => n6, ZN => n4);
   U3 : NAND2_X1 port map( A1 => EN, A2 => D, ZN => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_0;

architecture SYN_STRUCTURAL of RCA_N4_0 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_0;

architecture SYN_struct of carry_select_basic_N4_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n6, n7, n8, n9, n5
      , n_1154, n_1155 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1154);
   RCA1 : RCA_N4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1155);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n6);
   U6 : INV_X1 port map( A => n8, ZN => S(1));
   U7 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n8);
   U8 : INV_X1 port map( A => n7, ZN => S(2));
   U9 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n7);
   U10 : INV_X1 port map( A => n9, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n9);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_0 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_0;

architecture SYN_bhv of PGblock_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n2);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_0 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_0;

architecture SYN_bhv of Gblock_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_0 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_0;

architecture SYN_bhv of PG_net_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end rca_bhv_numBit32_0;

architecture SYN_BEHAVIORAL of rca_bhv_numBit32_0 is

   component rca_bhv_numBit32_0_DW01_add_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   signal n_1156 : std_logic;

begin
   
   add_1_root_add_35_2 : rca_bhv_numBit32_0_DW01_add_0 port map( A(32) => A(31)
                           , A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(32) => Co, SUM(31)
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1156);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_0 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_0;

architecture SYN_bhv of mux5to1_numBit32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n1, n2
      , n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n90, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n8);
   U2 : BUF_X1 port map( A => n10, Z => n4);
   U3 : BUF_X1 port map( A => n10, Z => n77);
   U4 : BUF_X1 port map( A => n10, Z => n78);
   U5 : INV_X1 port map( A => SEL_in(1), ZN => n90);
   U6 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82, 
                           C1 => IN5(2), C2 => n79, ZN => n68);
   U7 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82, 
                           C1 => IN5(3), C2 => n79, ZN => n66);
   U8 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82, 
                           C1 => IN5(4), C2 => n79, ZN => n64);
   U9 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82, 
                           C1 => IN5(5), C2 => n79, ZN => n62);
   U10 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82, 
                           C1 => IN5(6), C2 => n79, ZN => n60);
   U11 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82, 
                           C1 => IN5(7), C2 => n79, ZN => n58);
   U12 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82, 
                           C1 => IN5(8), C2 => n79, ZN => n56);
   U13 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82, 
                           C1 => IN5(9), C2 => n79, ZN => n54);
   U14 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => n82
                           , C1 => IN5(10), C2 => n79, ZN => n52);
   U15 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => n82
                           , C1 => IN5(11), C2 => n79, ZN => n50);
   U16 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => n83
                           , C1 => IN5(12), C2 => n80, ZN => n48);
   U17 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => n83
                           , C1 => IN5(13), C2 => n80, ZN => n46);
   U18 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n44);
   U19 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n42);
   U20 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84
                           , C1 => IN5(25), C2 => n81, ZN => n22);
   U21 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84
                           , C1 => IN5(26), C2 => n81, ZN => n20);
   U22 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84
                           , C1 => IN5(27), C2 => n81, ZN => n18);
   U23 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => n84
                           , C1 => IN5(28), C2 => n81, ZN => n16);
   U24 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => n84
                           , C1 => IN5(29), C2 => n81, ZN => n14);
   U25 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => n84
                           , C1 => IN5(30), C2 => n81, ZN => n12);
   U26 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82, 
                           C1 => IN5(1), C2 => n79, ZN => n70);
   U27 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n40);
   U28 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n38);
   U29 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n36);
   U30 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n34);
   U31 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n32);
   U32 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n30);
   U33 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n28);
   U34 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n26);
   U35 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n24);
   U36 : BUF_X1 port map( A => n9, Z => n79);
   U37 : BUF_X1 port map( A => n9, Z => n80);
   U38 : BUF_X1 port map( A => n7, Z => n85);
   U39 : BUF_X1 port map( A => n7, Z => n86);
   U40 : BUF_X1 port map( A => n89, Z => n1);
   U41 : BUF_X1 port map( A => n89, Z => n2);
   U42 : NOR2_X1 port map( A1 => n88, A2 => n75, ZN => n10);
   U43 : INV_X1 port map( A => n74, ZN => n88);
   U44 : BUF_X1 port map( A => n89, Z => n3);
   U45 : BUF_X1 port map( A => n9, Z => n81);
   U46 : BUF_X1 port map( A => n7, Z => n87);
   U47 : NOR4_X1 port map( A1 => n76, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n74);
   U48 : NOR3_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => n91, ZN => n7);
   U49 : BUF_X1 port map( A => n8, Z => n82);
   U50 : BUF_X1 port map( A => n8, Z => n83);
   U51 : BUF_X1 port map( A => n8, Z => n84);
   U52 : NOR2_X1 port map( A1 => n90, A2 => n91, ZN => n75);
   U53 : AND3_X1 port map( A1 => n91, A2 => n90, A3 => SEL_in(2), ZN => n9);
   U54 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => Z(3));
   U55 : INV_X1 port map( A => n73, ZN => n89);
   U56 : AOI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => n73);
   U57 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN 
                           => n69);
   U58 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN 
                           => n67);
   U59 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN 
                           => n65);
   U60 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN 
                           => n63);
   U61 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN 
                           => n61);
   U62 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN 
                           => n59);
   U63 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN 
                           => n57);
   U64 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN 
                           => n55);
   U65 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN 
                           => n53);
   U66 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n51);
   U67 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n49);
   U68 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2, 
                           ZN => n47);
   U69 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2, 
                           ZN => n45);
   U70 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n43);
   U71 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n76);
   U72 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82, 
                           C1 => IN5(0), C2 => n79, ZN => n72);
   U73 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n41);
   U74 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3, 
                           ZN => n23);
   U75 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3, 
                           ZN => n21);
   U76 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3, 
                           ZN => n19);
   U77 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3, 
                           ZN => n17);
   U78 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3, 
                           ZN => n15);
   U79 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3, 
                           ZN => n13);
   U80 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3, 
                           ZN => n11);
   U81 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN 
                           => n71);
   U82 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n33);
   U83 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n31);
   U84 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n29);
   U85 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n27);
   U86 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n25);
   U87 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => Z(4));
   U88 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => Z(5));
   U89 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => Z(6));
   U90 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => Z(7));
   U91 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => Z(8));
   U92 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => Z(9));
   U93 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => Z(10));
   U94 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => Z(11));
   U95 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => Z(12));
   U96 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => Z(13));
   U97 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => Z(14));
   U98 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => Z(15));
   U99 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => Z(16));
   U100 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2,
                           ZN => n39);
   U101 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => Z(17));
   U102 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2,
                           ZN => n37);
   U103 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => Z(18));
   U104 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2,
                           ZN => n35);
   U105 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => Z(19));
   U106 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => Z(20));
   U107 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => Z(21));
   U108 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => Z(22));
   U110 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => Z(23));
   U111 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => Z(24));
   U112 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => Z(25));
   U113 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => Z(26));
   U114 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => Z(27));
   U115 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => Z(28));
   U116 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => Z(29));
   U117 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => Z(30));
   U118 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => Z(2));
   U119 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => Z(0));
   U120 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => Z(1));
   U121 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Z(31));
   U122 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n5);
   U123 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => 
                           n84, C1 => IN5(31), C2 => n81, ZN => n6);
   U124 : INV_X1 port map( A => SEL_in(0), ZN => n91);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity booth_encoder_numBit16 is

   port( B : in std_logic_vector (15 downto 0);  SEL_out : out std_logic_vector
         (23 downto 0));

end booth_encoder_numBit16;

architecture SYN_structural of booth_encoder_numBit16 is

signal X_Logic0_port : std_logic;

begin
   SEL_out <= ( B(15), B(14), B(13), B(13), B(12), B(11), B(11), B(10), B(9), 
      B(9), B(8), B(7), B(7), B(6), B(5), B(5), B(4), B(3), B(3), B(2), B(1), 
      B(1), B(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8;

architecture SYN_structural of SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   component carry_select_basic_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CSBI_1 : carry_select_basic_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) 
                           => A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), 
                           B(1) => B(1), B(0) => B(0), C_i => Ci(0), S(3) => 
                           S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CSBI_2 : carry_select_basic_N4_7 port map( A(3) => A(7), A(2) => A(6), A(1) 
                           => A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), 
                           B(1) => B(5), B(0) => B(4), C_i => Ci(1), S(3) => 
                           S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   CSBI_3 : carry_select_basic_N4_6 port map( A(3) => A(11), A(2) => A(10), 
                           A(1) => A(9), A(0) => A(8), B(3) => B(11), B(2) => 
                           B(10), B(1) => B(9), B(0) => B(8), C_i => Ci(2), 
                           S(3) => S(11), S(2) => S(10), S(1) => S(9), S(0) => 
                           S(8));
   CSBI_4 : carry_select_basic_N4_5 port map( A(3) => A(15), A(2) => A(14), 
                           A(1) => A(13), A(0) => A(12), B(3) => B(15), B(2) =>
                           B(14), B(1) => B(13), B(0) => B(12), C_i => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   CSBI_5 : carry_select_basic_N4_4 port map( A(3) => A(19), A(2) => A(18), 
                           A(1) => A(17), A(0) => A(16), B(3) => B(19), B(2) =>
                           B(18), B(1) => B(17), B(0) => B(16), C_i => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   CSBI_6 : carry_select_basic_N4_3 port map( A(3) => A(23), A(2) => A(22), 
                           A(1) => A(21), A(0) => A(20), B(3) => B(23), B(2) =>
                           B(22), B(1) => B(21), B(0) => B(20), C_i => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   CSBI_7 : carry_select_basic_N4_2 port map( A(3) => A(27), A(2) => A(26), 
                           A(1) => A(25), A(0) => A(24), B(3) => B(27), B(2) =>
                           B(26), B(1) => B(25), B(0) => B(24), C_i => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   CSBI_8 : carry_select_basic_N4_1 port map( A(3) => A(31), A(2) => A(30), 
                           A(1) => A(29), A(0) => A(28), B(3) => B(31), B(2) =>
                           B(30), B(1) => B(29), B(0) => B(28), C_i => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_generator_NBIT32_NBIT_PER_BLOCK4 is

   port( A, B : in std_logic_vector (32 downto 1);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end carry_generator_NBIT32_NBIT_PER_BLOCK4;

architecture SYN_struct of carry_generator_NBIT32_NBIT_PER_BLOCK4 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component PGblock_1
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_2
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_3
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_4
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_5
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_6
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_7
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_8
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_9
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_10
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_11
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_12
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_13
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_14
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_15
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_16
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_17
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_18
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_19
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_20
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_21
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_22
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_23
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_24
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_25
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_26
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_0
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component Gblock_1
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_2
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_3
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_4
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_5
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_6
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_7
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_8
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_0
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_net_1
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_2
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_3
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_4
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_5
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_6
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_7
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_8
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_9
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_10
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_11
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_12
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_13
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_14
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_15
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_16
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_17
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_18
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_19
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_20
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_21
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_22
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_23
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_24
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_25
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_26
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_27
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_28
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_29
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_30
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_0
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   signal Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port, G_16_16_port, G_16_15_port, G_16_13_port, 
      G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, G_13_13_port, 
      G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, G_10_10_port, 
      G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port, G_7_7_port, 
      G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port, G_3_3_port, 
      G_2_2_port, G_2_1_port, G_1_1_port, P_16_16_port, P_16_15_port, 
      P_16_13_port, P_16_9_port, P_15_15_port, P_14_14_port, P_14_13_port, 
      P_13_13_port, P_12_12_port, P_12_11_port, P_12_9_port, P_11_11_port, 
      P_10_10_port, P_10_9_port, P_9_9_port, P_8_8_port, P_8_7_port, P_8_5_port
      , P_7_7_port, P_6_6_port, P_6_5_port, P_5_5_port, P_4_4_port, P_4_3_port,
      P_3_3_port, P_2_2_port, G_32_32_port, G_32_31_port, G_32_29_port, 
      G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, G_30_29_port, 
      G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, G_28_17_port, 
      G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, G_24_24_port, 
      G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, G_22_22_port, 
      G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, G_20_17_port, 
      G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, P_32_32_port, 
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n3, n1, n2 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port );
   
   PGnetblock_2 : PG_net_0 port map( a => A(2), b => B(2), p => P_2_2_port, g 
                           => G_2_2_port);
   PGnetblock_3 : PG_net_30 port map( a => A(3), b => B(3), p => P_3_3_port, g 
                           => G_3_3_port);
   PGnetblock_4 : PG_net_29 port map( a => A(4), b => B(4), p => P_4_4_port, g 
                           => G_4_4_port);
   PGnetblock_5 : PG_net_28 port map( a => A(5), b => B(5), p => P_5_5_port, g 
                           => G_5_5_port);
   PGnetblock_6 : PG_net_27 port map( a => A(6), b => B(6), p => P_6_6_port, g 
                           => G_6_6_port);
   PGnetblock_7 : PG_net_26 port map( a => A(7), b => B(7), p => P_7_7_port, g 
                           => G_7_7_port);
   PGnetblock_8 : PG_net_25 port map( a => A(8), b => B(8), p => P_8_8_port, g 
                           => G_8_8_port);
   PGnetblock_9 : PG_net_24 port map( a => A(9), b => B(9), p => P_9_9_port, g 
                           => G_9_9_port);
   PGnetblock_10 : PG_net_23 port map( a => A(10), b => B(10), p => 
                           P_10_10_port, g => G_10_10_port);
   PGnetblock_11 : PG_net_22 port map( a => A(11), b => B(11), p => 
                           P_11_11_port, g => G_11_11_port);
   PGnetblock_12 : PG_net_21 port map( a => A(12), b => B(12), p => 
                           P_12_12_port, g => G_12_12_port);
   PGnetblock_13 : PG_net_20 port map( a => A(13), b => B(13), p => 
                           P_13_13_port, g => G_13_13_port);
   PGnetblock_14 : PG_net_19 port map( a => A(14), b => B(14), p => 
                           P_14_14_port, g => G_14_14_port);
   PGnetblock_15 : PG_net_18 port map( a => A(15), b => B(15), p => 
                           P_15_15_port, g => G_15_15_port);
   PGnetblock_16 : PG_net_17 port map( a => A(16), b => B(16), p => 
                           P_16_16_port, g => G_16_16_port);
   PGnetblock_17 : PG_net_16 port map( a => A(17), b => B(17), p => 
                           P_17_17_port, g => G_17_17_port);
   PGnetblock_18 : PG_net_15 port map( a => A(18), b => B(18), p => 
                           P_18_18_port, g => G_18_18_port);
   PGnetblock_19 : PG_net_14 port map( a => A(19), b => B(19), p => 
                           P_19_19_port, g => G_19_19_port);
   PGnetblock_20 : PG_net_13 port map( a => A(20), b => B(20), p => 
                           P_20_20_port, g => G_20_20_port);
   PGnetblock_21 : PG_net_12 port map( a => A(21), b => B(21), p => 
                           P_21_21_port, g => G_21_21_port);
   PGnetblock_22 : PG_net_11 port map( a => A(22), b => B(22), p => 
                           P_22_22_port, g => G_22_22_port);
   PGnetblock_23 : PG_net_10 port map( a => A(23), b => B(23), p => 
                           P_23_23_port, g => G_23_23_port);
   PGnetblock_24 : PG_net_9 port map( a => A(24), b => B(24), p => P_24_24_port
                           , g => G_24_24_port);
   PGnetblock_25 : PG_net_8 port map( a => A(25), b => B(25), p => P_25_25_port
                           , g => G_25_25_port);
   PGnetblock_26 : PG_net_7 port map( a => A(26), b => B(26), p => P_26_26_port
                           , g => G_26_26_port);
   PGnetblock_27 : PG_net_6 port map( a => A(27), b => B(27), p => P_27_27_port
                           , g => G_27_27_port);
   PGnetblock_28 : PG_net_5 port map( a => A(28), b => B(28), p => P_28_28_port
                           , g => G_28_28_port);
   PGnetblock_29 : PG_net_4 port map( a => A(29), b => B(29), p => P_29_29_port
                           , g => G_29_29_port);
   PGnetblock_30 : PG_net_3 port map( a => A(30), b => B(30), p => P_30_30_port
                           , g => G_30_30_port);
   PGnetblock_31 : PG_net_2 port map( a => A(31), b => B(31), p => P_31_31_port
                           , g => G_31_31_port);
   PGnetblock_32 : PG_net_1 port map( a => A(32), b => B(32), p => P_32_32_port
                           , g => G_32_32_port);
   GB_low_1_2 : Gblock_0 port map( Pik => P_2_2_port, Gik => G_2_2_port, Gk_1j 
                           => G_1_1_port, Gij => G_2_1_port);
   GB_low_2_4 : Gblock_8 port map( Pik => P_4_3_port, Gik => G_4_3_port, Gk_1j 
                           => G_2_1_port, Gij => Co_0_port);
   GB_low_3_8 : Gblock_7 port map( Pik => P_8_5_port, Gik => G_8_5_port, Gk_1j 
                           => Co_0_port, Gij => Co_1_port);
   GB_high_4_16_0 : Gblock_6 port map( Pik => P_16_9_port, Gik => G_16_9_port, 
                           Gk_1j => Co_1_port, Gij => Co_3_port);
   GB_high_4_16_1 : Gblock_5 port map( Pik => P_12_9_port, Gik => G_12_9_port, 
                           Gk_1j => Co_1_port, Gij => Co_2_port);
   GB_high_5_32_0 : Gblock_4 port map( Pik => P_32_17_port, Gik => G_32_17_port
                           , Gk_1j => Co_3_port, Gij => Co_7_port);
   GB_high_5_32_1 : Gblock_3 port map( Pik => P_28_17_port, Gik => G_28_17_port
                           , Gk_1j => Co_3_port, Gij => Co_6_port);
   GB_high_5_32_2 : Gblock_2 port map( Pik => P_24_17_port, Gik => G_24_17_port
                           , Gk_1j => Co_3_port, Gij => Co_5_port);
   GB_high_5_32_3 : Gblock_1 port map( Pik => P_20_17_port, Gik => G_20_17_port
                           , Gk_1j => Co_3_port, Gij => Co_4_port);
   PGB_low_1_4 : PGblock_0 port map( Pik => P_4_4_port, Gik => G_4_4_port, 
                           Pk_1j => P_3_3_port, Gk_1j => G_3_3_port, Pij => 
                           P_4_3_port, Gij => G_4_3_port);
   PGB_low_1_6 : PGblock_26 port map( Pik => P_6_6_port, Gik => G_6_6_port, 
                           Pk_1j => P_5_5_port, Gk_1j => G_5_5_port, Pij => 
                           P_6_5_port, Gij => G_6_5_port);
   PGB_low_1_8 : PGblock_25 port map( Pik => P_8_8_port, Gik => G_8_8_port, 
                           Pk_1j => P_7_7_port, Gk_1j => G_7_7_port, Pij => 
                           P_8_7_port, Gij => G_8_7_port);
   PGB_low_1_10 : PGblock_24 port map( Pik => P_10_10_port, Gik => G_10_10_port
                           , Pk_1j => P_9_9_port, Gk_1j => G_9_9_port, Pij => 
                           P_10_9_port, Gij => G_10_9_port);
   PGB_low_1_12 : PGblock_23 port map( Pik => P_12_12_port, Gik => G_12_12_port
                           , Pk_1j => P_11_11_port, Gk_1j => G_11_11_port, Pij 
                           => P_12_11_port, Gij => G_12_11_port);
   PGB_low_1_14 : PGblock_22 port map( Pik => P_14_14_port, Gik => G_14_14_port
                           , Pk_1j => P_13_13_port, Gk_1j => G_13_13_port, Pij 
                           => P_14_13_port, Gij => G_14_13_port);
   PGB_low_1_16 : PGblock_21 port map( Pik => P_16_16_port, Gik => G_16_16_port
                           , Pk_1j => P_15_15_port, Gk_1j => G_15_15_port, Pij 
                           => P_16_15_port, Gij => G_16_15_port);
   PGB_low_1_18 : PGblock_20 port map( Pik => P_18_18_port, Gik => G_18_18_port
                           , Pk_1j => P_17_17_port, Gk_1j => G_17_17_port, Pij 
                           => P_18_17_port, Gij => G_18_17_port);
   PGB_low_1_20 : PGblock_19 port map( Pik => P_20_20_port, Gik => G_20_20_port
                           , Pk_1j => P_19_19_port, Gk_1j => G_19_19_port, Pij 
                           => P_20_19_port, Gij => G_20_19_port);
   PGB_low_1_22 : PGblock_18 port map( Pik => P_22_22_port, Gik => G_22_22_port
                           , Pk_1j => P_21_21_port, Gk_1j => G_21_21_port, Pij 
                           => P_22_21_port, Gij => G_22_21_port);
   PGB_low_1_24 : PGblock_17 port map( Pik => P_24_24_port, Gik => G_24_24_port
                           , Pk_1j => P_23_23_port, Gk_1j => G_23_23_port, Pij 
                           => P_24_23_port, Gij => G_24_23_port);
   PGB_low_1_26 : PGblock_16 port map( Pik => P_26_26_port, Gik => G_26_26_port
                           , Pk_1j => P_25_25_port, Gk_1j => G_25_25_port, Pij 
                           => P_26_25_port, Gij => G_26_25_port);
   PGB_low_1_28 : PGblock_15 port map( Pik => P_28_28_port, Gik => G_28_28_port
                           , Pk_1j => P_27_27_port, Gk_1j => G_27_27_port, Pij 
                           => P_28_27_port, Gij => G_28_27_port);
   PGB_low_1_30 : PGblock_14 port map( Pik => P_30_30_port, Gik => G_30_30_port
                           , Pk_1j => P_29_29_port, Gk_1j => G_29_29_port, Pij 
                           => P_30_29_port, Gij => G_30_29_port);
   PGB_low_1_32 : PGblock_13 port map( Pik => P_32_32_port, Gik => G_32_32_port
                           , Pk_1j => P_31_31_port, Gk_1j => G_31_31_port, Pij 
                           => P_32_31_port, Gij => G_32_31_port);
   PGB_low_2_8 : PGblock_12 port map( Pik => P_8_7_port, Gik => G_8_7_port, 
                           Pk_1j => P_6_5_port, Gk_1j => G_6_5_port, Pij => 
                           P_8_5_port, Gij => G_8_5_port);
   PGB_low_2_12 : PGblock_11 port map( Pik => P_12_11_port, Gik => G_12_11_port
                           , Pk_1j => P_10_9_port, Gk_1j => G_10_9_port, Pij =>
                           P_12_9_port, Gij => G_12_9_port);
   PGB_low_2_16 : PGblock_10 port map( Pik => P_16_15_port, Gik => G_16_15_port
                           , Pk_1j => P_14_13_port, Gk_1j => G_14_13_port, Pij 
                           => P_16_13_port, Gij => G_16_13_port);
   PGB_low_2_20 : PGblock_9 port map( Pik => P_20_19_port, Gik => G_20_19_port,
                           Pk_1j => P_18_17_port, Gk_1j => G_18_17_port, Pij =>
                           P_20_17_port, Gij => G_20_17_port);
   PGB_low_2_24 : PGblock_8 port map( Pik => P_24_23_port, Gik => G_24_23_port,
                           Pk_1j => P_22_21_port, Gk_1j => G_22_21_port, Pij =>
                           P_24_21_port, Gij => G_24_21_port);
   PGB_low_2_28 : PGblock_7 port map( Pik => P_28_27_port, Gik => G_28_27_port,
                           Pk_1j => P_26_25_port, Gk_1j => G_26_25_port, Pij =>
                           P_28_25_port, Gij => G_28_25_port);
   PGB_low_2_32 : PGblock_6 port map( Pik => P_32_31_port, Gik => G_32_31_port,
                           Pk_1j => P_30_29_port, Gk_1j => G_30_29_port, Pij =>
                           P_32_29_port, Gij => G_32_29_port);
   PGB_low_3_16 : PGblock_5 port map( Pik => P_16_13_port, Gik => G_16_13_port,
                           Pk_1j => P_12_9_port, Gk_1j => G_12_9_port, Pij => 
                           P_16_9_port, Gij => G_16_9_port);
   PGB_low_3_24 : PGblock_4 port map( Pik => P_24_21_port, Gik => G_24_21_port,
                           Pk_1j => P_20_17_port, Gk_1j => G_20_17_port, Pij =>
                           P_24_17_port, Gij => G_24_17_port);
   PGB_low_3_32 : PGblock_3 port map( Pik => P_32_29_port, Gik => G_32_29_port,
                           Pk_1j => P_28_25_port, Gk_1j => G_28_25_port, Pij =>
                           P_32_25_port, Gij => G_32_25_port);
   PGB_high_4_32_0 : PGblock_2 port map( Pik => P_32_25_port, Gik => 
                           G_32_25_port, Pk_1j => P_24_17_port, Gk_1j => 
                           G_24_17_port, Pij => P_32_17_port, Gij => 
                           G_32_17_port);
   PGB_high_4_32_1 : PGblock_1 port map( Pik => P_28_25_port, Gik => 
                           G_28_25_port, Pk_1j => P_24_17_port, Gk_1j => 
                           G_24_17_port, Pij => P_28_17_port, Gij => 
                           G_28_17_port);
   U1 : INV_X1 port map( A => A(1), ZN => n1);
   U2 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => G_1_1_port);
   U3 : INV_X1 port map( A => B(1), ZN => n2);
   U4 : OAI21_X1 port map( B1 => A(1), B2 => B(1), A => Cin, ZN => n3);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BOOTHMUL_numBit16 is

   port( A, B : in std_logic_vector (15 downto 0);  P : out std_logic_vector 
         (31 downto 0));

end BOOTHMUL_numBit16;

architecture SYN_mixed of BOOTHMUL_numBit16 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component rca_bhv_numBit32_1
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component rca_bhv_numBit32_2
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component rca_bhv_numBit32_3
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component rca_bhv_numBit32_4
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component rca_bhv_numBit32_5
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component rca_bhv_numBit32_6
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component rca_bhv_numBit32_0
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component mux5to1_numBit32_1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux5to1_numBit32_2
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux5to1_numBit32_3
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux5to1_numBit32_4
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux5to1_numBit32_5
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux5to1_numBit32_6
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux5to1_numBit32_7
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux5to1_numBit32_0
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component booth_encoder_numBit16
      port( B : in std_logic_vector (15 downto 0);  SEL_out : out 
            std_logic_vector (23 downto 0));
   end component;
   
   signal X_Logic0_port, encoder_out_23_port, encoder_out_22_port, 
      encoder_out_21_port, encoder_out_20_port, encoder_out_19_port, 
      encoder_out_18_port, encoder_out_17_port, encoder_out_16_port, 
      encoder_out_15_port, encoder_out_14_port, encoder_out_13_port, 
      encoder_out_12_port, encoder_out_11_port, encoder_out_10_port, 
      encoder_out_9_port, encoder_out_8_port, encoder_out_7_port, 
      encoder_out_6_port, encoder_out_5_port, encoder_out_4_port, 
      encoder_out_3_port, encoder_out_2_port, encoder_out_1_port, 
      encoder_out_0_port, A_minus_31_port, A_minus_15_port, A_minus_14_port, 
      A_minus_13_port, A_minus_12_port, A_minus_11_port, A_minus_10_port, 
      A_minus_9_port, A_minus_8_port, A_minus_7_port, A_minus_6_port, 
      A_minus_5_port, A_minus_4_port, A_minus_3_port, A_minus_2_port, 
      A_minus_1_port, A_minus_0_port, sum_op_7_31_port, sum_op_7_30_port, 
      sum_op_7_29_port, sum_op_7_28_port, sum_op_7_27_port, sum_op_7_26_port, 
      sum_op_7_25_port, sum_op_7_24_port, sum_op_7_23_port, sum_op_7_22_port, 
      sum_op_7_21_port, sum_op_7_20_port, sum_op_7_19_port, sum_op_7_18_port, 
      sum_op_7_17_port, sum_op_7_16_port, sum_op_7_15_port, sum_op_7_14_port, 
      sum_op_7_13_port, sum_op_7_12_port, sum_op_7_11_port, sum_op_7_10_port, 
      sum_op_7_9_port, sum_op_7_8_port, sum_op_7_7_port, sum_op_7_6_port, 
      sum_op_7_5_port, sum_op_7_4_port, sum_op_7_3_port, sum_op_7_2_port, 
      sum_op_7_1_port, sum_op_7_0_port, sum_op_6_31_port, sum_op_6_30_port, 
      sum_op_6_29_port, sum_op_6_28_port, sum_op_6_27_port, sum_op_6_26_port, 
      sum_op_6_25_port, sum_op_6_24_port, sum_op_6_23_port, sum_op_6_22_port, 
      sum_op_6_21_port, sum_op_6_20_port, sum_op_6_19_port, sum_op_6_18_port, 
      sum_op_6_17_port, sum_op_6_16_port, sum_op_6_15_port, sum_op_6_14_port, 
      sum_op_6_13_port, sum_op_6_12_port, sum_op_6_11_port, sum_op_6_10_port, 
      sum_op_6_9_port, sum_op_6_8_port, sum_op_6_7_port, sum_op_6_6_port, 
      sum_op_6_5_port, sum_op_6_4_port, sum_op_6_3_port, sum_op_6_2_port, 
      sum_op_6_1_port, sum_op_6_0_port, sum_op_5_31_port, sum_op_5_30_port, 
      sum_op_5_29_port, sum_op_5_28_port, sum_op_5_27_port, sum_op_5_26_port, 
      sum_op_5_25_port, sum_op_5_24_port, sum_op_5_23_port, sum_op_5_22_port, 
      sum_op_5_21_port, sum_op_5_20_port, sum_op_5_19_port, sum_op_5_18_port, 
      sum_op_5_17_port, sum_op_5_16_port, sum_op_5_15_port, sum_op_5_14_port, 
      sum_op_5_13_port, sum_op_5_12_port, sum_op_5_11_port, sum_op_5_10_port, 
      sum_op_5_9_port, sum_op_5_8_port, sum_op_5_7_port, sum_op_5_6_port, 
      sum_op_5_5_port, sum_op_5_4_port, sum_op_5_3_port, sum_op_5_2_port, 
      sum_op_5_1_port, sum_op_5_0_port, sum_op_4_31_port, sum_op_4_30_port, 
      sum_op_4_29_port, sum_op_4_28_port, sum_op_4_27_port, sum_op_4_26_port, 
      sum_op_4_25_port, sum_op_4_24_port, sum_op_4_23_port, sum_op_4_22_port, 
      sum_op_4_21_port, sum_op_4_20_port, sum_op_4_19_port, sum_op_4_18_port, 
      sum_op_4_17_port, sum_op_4_16_port, sum_op_4_15_port, sum_op_4_14_port, 
      sum_op_4_13_port, sum_op_4_12_port, sum_op_4_11_port, sum_op_4_10_port, 
      sum_op_4_9_port, sum_op_4_8_port, sum_op_4_7_port, sum_op_4_6_port, 
      sum_op_4_5_port, sum_op_4_4_port, sum_op_4_3_port, sum_op_4_2_port, 
      sum_op_4_1_port, sum_op_4_0_port, sum_op_3_31_port, sum_op_3_30_port, 
      sum_op_3_29_port, sum_op_3_28_port, sum_op_3_27_port, sum_op_3_26_port, 
      sum_op_3_25_port, sum_op_3_24_port, sum_op_3_23_port, sum_op_3_22_port, 
      sum_op_3_21_port, sum_op_3_20_port, sum_op_3_19_port, sum_op_3_18_port, 
      sum_op_3_17_port, sum_op_3_16_port, sum_op_3_15_port, sum_op_3_14_port, 
      sum_op_3_13_port, sum_op_3_12_port, sum_op_3_11_port, sum_op_3_10_port, 
      sum_op_3_9_port, sum_op_3_8_port, sum_op_3_7_port, sum_op_3_6_port, 
      sum_op_3_5_port, sum_op_3_4_port, sum_op_3_3_port, sum_op_3_2_port, 
      sum_op_3_1_port, sum_op_3_0_port, sum_op_2_31_port, sum_op_2_30_port, 
      sum_op_2_29_port, sum_op_2_28_port, sum_op_2_27_port, sum_op_2_26_port, 
      sum_op_2_25_port, sum_op_2_24_port, sum_op_2_23_port, sum_op_2_22_port, 
      sum_op_2_21_port, sum_op_2_20_port, sum_op_2_19_port, sum_op_2_18_port, 
      sum_op_2_17_port, sum_op_2_16_port, sum_op_2_15_port, sum_op_2_14_port, 
      sum_op_2_13_port, sum_op_2_12_port, sum_op_2_11_port, sum_op_2_10_port, 
      sum_op_2_9_port, sum_op_2_8_port, sum_op_2_7_port, sum_op_2_6_port, 
      sum_op_2_5_port, sum_op_2_4_port, sum_op_2_3_port, sum_op_2_2_port, 
      sum_op_2_1_port, sum_op_2_0_port, sum_op_1_31_port, sum_op_1_30_port, 
      sum_op_1_29_port, sum_op_1_28_port, sum_op_1_27_port, sum_op_1_26_port, 
      sum_op_1_25_port, sum_op_1_24_port, sum_op_1_23_port, sum_op_1_22_port, 
      sum_op_1_21_port, sum_op_1_20_port, sum_op_1_19_port, sum_op_1_18_port, 
      sum_op_1_17_port, sum_op_1_16_port, sum_op_1_15_port, sum_op_1_14_port, 
      sum_op_1_13_port, sum_op_1_12_port, sum_op_1_11_port, sum_op_1_10_port, 
      sum_op_1_9_port, sum_op_1_8_port, sum_op_1_7_port, sum_op_1_6_port, 
      sum_op_1_5_port, sum_op_1_4_port, sum_op_1_3_port, sum_op_1_2_port, 
      sum_op_1_1_port, sum_op_1_0_port, sum_op_0_31_port, sum_op_0_30_port, 
      sum_op_0_29_port, sum_op_0_28_port, sum_op_0_27_port, sum_op_0_26_port, 
      sum_op_0_25_port, sum_op_0_24_port, sum_op_0_23_port, sum_op_0_22_port, 
      sum_op_0_21_port, sum_op_0_20_port, sum_op_0_19_port, sum_op_0_18_port, 
      sum_op_0_17_port, sum_op_0_16_port, sum_op_0_15_port, sum_op_0_14_port, 
      sum_op_0_13_port, sum_op_0_12_port, sum_op_0_11_port, sum_op_0_10_port, 
      sum_op_0_9_port, sum_op_0_8_port, sum_op_0_7_port, sum_op_0_6_port, 
      sum_op_0_5_port, sum_op_0_4_port, sum_op_0_3_port, sum_op_0_2_port, 
      sum_op_0_1_port, sum_op_0_0_port, rca_out_5_31_port, rca_out_5_30_port, 
      rca_out_5_29_port, rca_out_5_28_port, rca_out_5_27_port, 
      rca_out_5_26_port, rca_out_5_25_port, rca_out_5_24_port, 
      rca_out_5_23_port, rca_out_5_22_port, rca_out_5_21_port, 
      rca_out_5_20_port, rca_out_5_19_port, rca_out_5_18_port, 
      rca_out_5_17_port, rca_out_5_16_port, rca_out_5_15_port, 
      rca_out_5_14_port, rca_out_5_13_port, rca_out_5_12_port, 
      rca_out_5_11_port, rca_out_5_10_port, rca_out_5_9_port, rca_out_5_8_port,
      rca_out_5_7_port, rca_out_5_6_port, rca_out_5_5_port, rca_out_5_4_port, 
      rca_out_5_3_port, rca_out_5_2_port, rca_out_5_1_port, rca_out_5_0_port, 
      rca_out_4_31_port, rca_out_4_30_port, rca_out_4_29_port, 
      rca_out_4_28_port, rca_out_4_27_port, rca_out_4_26_port, 
      rca_out_4_25_port, rca_out_4_24_port, rca_out_4_23_port, 
      rca_out_4_22_port, rca_out_4_21_port, rca_out_4_20_port, 
      rca_out_4_19_port, rca_out_4_18_port, rca_out_4_17_port, 
      rca_out_4_16_port, rca_out_4_15_port, rca_out_4_14_port, 
      rca_out_4_13_port, rca_out_4_12_port, rca_out_4_11_port, 
      rca_out_4_10_port, rca_out_4_9_port, rca_out_4_8_port, rca_out_4_7_port, 
      rca_out_4_6_port, rca_out_4_5_port, rca_out_4_4_port, rca_out_4_3_port, 
      rca_out_4_2_port, rca_out_4_1_port, rca_out_4_0_port, rca_out_3_31_port, 
      rca_out_3_30_port, rca_out_3_29_port, rca_out_3_28_port, 
      rca_out_3_27_port, rca_out_3_26_port, rca_out_3_25_port, 
      rca_out_3_24_port, rca_out_3_23_port, rca_out_3_22_port, 
      rca_out_3_21_port, rca_out_3_20_port, rca_out_3_19_port, 
      rca_out_3_18_port, rca_out_3_17_port, rca_out_3_16_port, 
      rca_out_3_15_port, rca_out_3_14_port, rca_out_3_13_port, 
      rca_out_3_12_port, rca_out_3_11_port, rca_out_3_10_port, rca_out_3_9_port
      , rca_out_3_8_port, rca_out_3_7_port, rca_out_3_6_port, rca_out_3_5_port,
      rca_out_3_4_port, rca_out_3_3_port, rca_out_3_2_port, rca_out_3_1_port, 
      rca_out_3_0_port, rca_out_2_31_port, rca_out_2_30_port, rca_out_2_29_port
      , rca_out_2_28_port, rca_out_2_27_port, rca_out_2_26_port, 
      rca_out_2_25_port, rca_out_2_24_port, rca_out_2_23_port, 
      rca_out_2_22_port, rca_out_2_21_port, rca_out_2_20_port, 
      rca_out_2_19_port, rca_out_2_18_port, rca_out_2_17_port, 
      rca_out_2_16_port, rca_out_2_15_port, rca_out_2_14_port, 
      rca_out_2_13_port, rca_out_2_12_port, rca_out_2_11_port, 
      rca_out_2_10_port, rca_out_2_9_port, rca_out_2_8_port, rca_out_2_7_port, 
      rca_out_2_6_port, rca_out_2_5_port, rca_out_2_4_port, rca_out_2_3_port, 
      rca_out_2_2_port, rca_out_2_1_port, rca_out_2_0_port, rca_out_1_31_port, 
      rca_out_1_30_port, rca_out_1_29_port, rca_out_1_28_port, 
      rca_out_1_27_port, rca_out_1_26_port, rca_out_1_25_port, 
      rca_out_1_24_port, rca_out_1_23_port, rca_out_1_22_port, 
      rca_out_1_21_port, rca_out_1_20_port, rca_out_1_19_port, 
      rca_out_1_18_port, rca_out_1_17_port, rca_out_1_16_port, 
      rca_out_1_15_port, rca_out_1_14_port, rca_out_1_13_port, 
      rca_out_1_12_port, rca_out_1_11_port, rca_out_1_10_port, rca_out_1_9_port
      , rca_out_1_8_port, rca_out_1_7_port, rca_out_1_6_port, rca_out_1_5_port,
      rca_out_1_4_port, rca_out_1_3_port, rca_out_1_2_port, rca_out_1_1_port, 
      rca_out_1_0_port, rca_out_0_31_port, rca_out_0_30_port, rca_out_0_29_port
      , rca_out_0_28_port, rca_out_0_27_port, rca_out_0_26_port, 
      rca_out_0_25_port, rca_out_0_24_port, rca_out_0_23_port, 
      rca_out_0_22_port, rca_out_0_21_port, rca_out_0_20_port, 
      rca_out_0_19_port, rca_out_0_18_port, rca_out_0_17_port, 
      rca_out_0_16_port, rca_out_0_15_port, rca_out_0_14_port, 
      rca_out_0_13_port, rca_out_0_12_port, rca_out_0_11_port, 
      rca_out_0_10_port, rca_out_0_9_port, rca_out_0_8_port, rca_out_0_7_port, 
      rca_out_0_6_port, rca_out_0_5_port, rca_out_0_4_port, rca_out_0_3_port, 
      rca_out_0_2_port, rca_out_0_1_port, rca_out_0_0_port, add_65_carry_2_port
      , add_65_carry_3_port, add_65_carry_4_port, add_65_carry_5_port, 
      add_65_carry_6_port, add_65_carry_7_port, add_65_carry_8_port, 
      add_65_carry_9_port, add_65_carry_10_port, add_65_carry_11_port, 
      add_65_carry_12_port, add_65_carry_13_port, add_65_carry_14_port, 
      add_65_carry_15_port, add_65_A_0_port, add_65_A_1_port, add_65_A_2_port, 
      add_65_A_3_port, add_65_A_4_port, add_65_A_5_port, add_65_A_6_port, 
      add_65_A_7_port, add_65_A_8_port, add_65_A_9_port, add_65_A_10_port, 
      add_65_A_11_port, add_65_A_12_port, add_65_A_13_port, add_65_A_14_port, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164 : std_logic;

begin
   
   X_Logic0_port <= '0';
   encode : booth_encoder_numBit16 port map( B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           SEL_out(23) => encoder_out_23_port, SEL_out(22) => 
                           encoder_out_22_port, SEL_out(21) => 
                           encoder_out_21_port, SEL_out(20) => 
                           encoder_out_20_port, SEL_out(19) => 
                           encoder_out_19_port, SEL_out(18) => 
                           encoder_out_18_port, SEL_out(17) => 
                           encoder_out_17_port, SEL_out(16) => 
                           encoder_out_16_port, SEL_out(15) => 
                           encoder_out_15_port, SEL_out(14) => 
                           encoder_out_14_port, SEL_out(13) => 
                           encoder_out_13_port, SEL_out(12) => 
                           encoder_out_12_port, SEL_out(11) => 
                           encoder_out_11_port, SEL_out(10) => 
                           encoder_out_10_port, SEL_out(9) => 
                           encoder_out_9_port, SEL_out(8) => encoder_out_8_port
                           , SEL_out(7) => encoder_out_7_port, SEL_out(6) => 
                           encoder_out_6_port, SEL_out(5) => encoder_out_5_port
                           , SEL_out(4) => encoder_out_4_port, SEL_out(3) => 
                           encoder_out_3_port, SEL_out(2) => encoder_out_2_port
                           , SEL_out(1) => encoder_out_1_port, SEL_out(0) => 
                           n_1157);
   mux0_0 : mux5to1_numBit32_0 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => n48, IN2(30) => n48, 
                           IN2(29) => n49, IN2(28) => n48, IN2(27) => n48, 
                           IN2(26) => n49, IN2(25) => n48, IN2(24) => n49, 
                           IN2(23) => n48, IN2(22) => n48, IN2(21) => n48, 
                           IN2(20) => n49, IN2(19) => n48, IN2(18) => n49, 
                           IN2(17) => n48, IN2(16) => n49, IN2(15) => n48, 
                           IN2(14) => A(14), IN2(13) => A(13), IN2(12) => A(12)
                           , IN2(11) => A(11), IN2(10) => A(10), IN2(9) => A(9)
                           , IN2(8) => A(8), IN2(7) => A(7), IN2(6) => A(6), 
                           IN2(5) => A(5), IN2(4) => A(4), IN2(3) => A(3), 
                           IN2(2) => A(2), IN2(1) => A(1), IN2(0) => A(0), 
                           IN3(31) => n35, IN3(30) => n31, IN3(29) => n31, 
                           IN3(28) => n36, IN3(27) => n31, IN3(26) => n35, 
                           IN3(25) => n31, IN3(24) => n36, IN3(23) => n31, 
                           IN3(22) => n36, IN3(21) => n32, IN3(20) => n35, 
                           IN3(19) => n32, IN3(18) => n35, IN3(17) => n33, 
                           IN3(16) => n34, IN3(15) => A_minus_15_port, IN3(14) 
                           => n2, IN3(13) => n4, IN3(12) => n6, IN3(11) => n8, 
                           IN3(10) => n10, IN3(9) => n12, IN3(8) => n14, IN3(7)
                           => n16, IN3(6) => n18, IN3(5) => n20, IN3(4) => n22,
                           IN3(3) => n24, IN3(2) => n26, IN3(1) => n28, IN3(0) 
                           => A_minus_0_port, IN4(31) => n42, IN4(30) => n42, 
                           IN4(29) => n42, IN4(28) => n42, IN4(27) => n42, 
                           IN4(26) => n42, IN4(25) => n42, IN4(24) => n42, 
                           IN4(23) => n42, IN4(22) => n42, IN4(21) => n42, 
                           IN4(20) => n43, IN4(19) => n43, IN4(18) => n43, 
                           IN4(17) => n43, IN4(16) => n43, IN4(15) => A(14), 
                           IN4(14) => A(13), IN4(13) => A(12), IN4(12) => A(11)
                           , IN4(11) => A(10), IN4(10) => A(9), IN4(9) => A(8),
                           IN4(8) => A(7), IN4(7) => A(6), IN4(6) => A(5), 
                           IN4(5) => A(4), IN4(4) => A(3), IN4(3) => A(2), 
                           IN4(2) => A(1), IN4(1) => A(0), IN4(0) => 
                           X_Logic0_port, IN5(31) => n41, IN5(30) => n41, 
                           IN5(29) => n41, IN5(28) => n41, IN5(27) => n41, 
                           IN5(26) => n41, IN5(25) => n40, IN5(24) => n40, 
                           IN5(23) => n39, IN5(22) => n40, IN5(21) => n38, 
                           IN5(20) => n39, IN5(19) => n38, IN5(18) => n38, 
                           IN5(17) => n39, IN5(16) => A_minus_15_port, IN5(15) 
                           => n2, IN5(14) => n4, IN5(13) => n6, IN5(12) => n8, 
                           IN5(11) => n10, IN5(10) => n12, IN5(9) => n14, 
                           IN5(8) => n16, IN5(7) => n18, IN5(6) => n20, IN5(5) 
                           => n22, IN5(4) => n24, IN5(3) => n26, IN5(2) => n28,
                           IN5(1) => A_minus_0_port, IN5(0) => X_Logic0_port, 
                           SEL_in(2) => encoder_out_2_port, SEL_in(1) => 
                           encoder_out_1_port, SEL_in(0) => encoder_out_0_port,
                           Z(31) => sum_op_0_31_port, Z(30) => sum_op_0_30_port
                           , Z(29) => sum_op_0_29_port, Z(28) => 
                           sum_op_0_28_port, Z(27) => sum_op_0_27_port, Z(26) 
                           => sum_op_0_26_port, Z(25) => sum_op_0_25_port, 
                           Z(24) => sum_op_0_24_port, Z(23) => sum_op_0_23_port
                           , Z(22) => sum_op_0_22_port, Z(21) => 
                           sum_op_0_21_port, Z(20) => sum_op_0_20_port, Z(19) 
                           => sum_op_0_19_port, Z(18) => sum_op_0_18_port, 
                           Z(17) => sum_op_0_17_port, Z(16) => sum_op_0_16_port
                           , Z(15) => sum_op_0_15_port, Z(14) => 
                           sum_op_0_14_port, Z(13) => sum_op_0_13_port, Z(12) 
                           => sum_op_0_12_port, Z(11) => sum_op_0_11_port, 
                           Z(10) => sum_op_0_10_port, Z(9) => sum_op_0_9_port, 
                           Z(8) => sum_op_0_8_port, Z(7) => sum_op_0_7_port, 
                           Z(6) => sum_op_0_6_port, Z(5) => sum_op_0_5_port, 
                           Z(4) => sum_op_0_4_port, Z(3) => sum_op_0_3_port, 
                           Z(2) => sum_op_0_2_port, Z(1) => sum_op_0_1_port, 
                           Z(0) => sum_op_0_0_port);
   mux_i_1 : mux5to1_numBit32_7 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => n52, IN2(30) => n51, 
                           IN2(29) => n51, IN2(28) => n51, IN2(27) => n51, 
                           IN2(26) => n51, IN2(25) => n50, IN2(24) => n50, 
                           IN2(23) => n50, IN2(22) => n50, IN2(21) => n50, 
                           IN2(20) => n49, IN2(19) => n49, IN2(18) => n49, 
                           IN2(17) => n49, IN2(16) => A(14), IN2(15) => A(13), 
                           IN2(14) => A(12), IN2(13) => A(11), IN2(12) => A(10)
                           , IN2(11) => A(9), IN2(10) => A(8), IN2(9) => A(7), 
                           IN2(8) => A(6), IN2(7) => A(5), IN2(6) => A(4), 
                           IN2(5) => A(3), IN2(4) => A(2), IN2(3) => A(1), 
                           IN2(2) => A(0), IN2(1) => X_Logic0_port, IN2(0) => 
                           X_Logic0_port, IN3(31) => n31, IN3(30) => n36, 
                           IN3(29) => n31, IN3(28) => n35, IN3(27) => n31, 
                           IN3(26) => n35, IN3(25) => n32, IN3(24) => n36, 
                           IN3(23) => n32, IN3(22) => n35, IN3(21) => n33, 
                           IN3(20) => n34, IN3(19) => n33, IN3(18) => n34, 
                           IN3(17) => A_minus_15_port, IN3(16) => n2, IN3(15) 
                           => n4, IN3(14) => n6, IN3(13) => n8, IN3(12) => n10,
                           IN3(11) => n12, IN3(10) => n14, IN3(9) => n16, 
                           IN3(8) => n18, IN3(7) => n20, IN3(6) => n22, IN3(5) 
                           => n24, IN3(4) => n26, IN3(3) => n28, IN3(2) => 
                           A_minus_0_port, IN3(1) => X_Logic0_port, IN3(0) => 
                           X_Logic0_port, IN4(31) => n47, IN4(30) => n47, 
                           IN4(29) => n47, IN4(28) => n47, IN4(27) => n46, 
                           IN4(26) => n47, IN4(25) => n47, IN4(24) => n47, 
                           IN4(23) => n46, IN4(22) => n46, IN4(21) => n46, 
                           IN4(20) => n46, IN4(19) => n46, IN4(18) => n42, 
                           IN4(17) => A(14), IN4(16) => A(13), IN4(15) => A(12)
                           , IN4(14) => A(11), IN4(13) => A(10), IN4(12) => 
                           A(9), IN4(11) => A(8), IN4(10) => A(7), IN4(9) => 
                           A(6), IN4(8) => A(5), IN4(7) => A(4), IN4(6) => A(3)
                           , IN4(5) => A(2), IN4(4) => A(1), IN4(3) => A(0), 
                           IN4(2) => X_Logic0_port, IN4(1) => X_Logic0_port, 
                           IN4(0) => X_Logic0_port, IN5(31) => n41, IN5(30) => 
                           n41, IN5(29) => n40, IN5(28) => n40, IN5(27) => n40,
                           IN5(26) => n40, IN5(25) => n40, IN5(24) => n41, 
                           IN5(23) => n37, IN5(22) => n39, IN5(21) => n37, 
                           IN5(20) => n39, IN5(19) => n37, IN5(18) => 
                           A_minus_15_port, IN5(17) => n2, IN5(16) => n4, 
                           IN5(15) => n6, IN5(14) => n8, IN5(13) => n10, 
                           IN5(12) => n12, IN5(11) => n14, IN5(10) => n16, 
                           IN5(9) => n18, IN5(8) => n20, IN5(7) => n22, IN5(6) 
                           => n24, IN5(5) => n26, IN5(4) => n28, IN5(3) => 
                           A_minus_0_port, IN5(2) => X_Logic0_port, IN5(1) => 
                           X_Logic0_port, IN5(0) => X_Logic0_port, SEL_in(2) =>
                           encoder_out_5_port, SEL_in(1) => encoder_out_4_port,
                           SEL_in(0) => encoder_out_3_port, Z(31) => 
                           sum_op_1_31_port, Z(30) => sum_op_1_30_port, Z(29) 
                           => sum_op_1_29_port, Z(28) => sum_op_1_28_port, 
                           Z(27) => sum_op_1_27_port, Z(26) => sum_op_1_26_port
                           , Z(25) => sum_op_1_25_port, Z(24) => 
                           sum_op_1_24_port, Z(23) => sum_op_1_23_port, Z(22) 
                           => sum_op_1_22_port, Z(21) => sum_op_1_21_port, 
                           Z(20) => sum_op_1_20_port, Z(19) => sum_op_1_19_port
                           , Z(18) => sum_op_1_18_port, Z(17) => 
                           sum_op_1_17_port, Z(16) => sum_op_1_16_port, Z(15) 
                           => sum_op_1_15_port, Z(14) => sum_op_1_14_port, 
                           Z(13) => sum_op_1_13_port, Z(12) => sum_op_1_12_port
                           , Z(11) => sum_op_1_11_port, Z(10) => 
                           sum_op_1_10_port, Z(9) => sum_op_1_9_port, Z(8) => 
                           sum_op_1_8_port, Z(7) => sum_op_1_7_port, Z(6) => 
                           sum_op_1_6_port, Z(5) => sum_op_1_5_port, Z(4) => 
                           sum_op_1_4_port, Z(3) => sum_op_1_3_port, Z(2) => 
                           sum_op_1_2_port, Z(1) => sum_op_1_1_port, Z(0) => 
                           sum_op_1_0_port);
   mux_i_2 : mux5to1_numBit32_6 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => A(15), IN2(30) => A(15), 
                           IN2(29) => A(15), IN2(28) => A(15), IN2(27) => A(15)
                           , IN2(26) => A(15), IN2(25) => n48, IN2(24) => A(15)
                           , IN2(23) => A(15), IN2(22) => n53, IN2(21) => n53, 
                           IN2(20) => n53, IN2(19) => n53, IN2(18) => A(14), 
                           IN2(17) => A(13), IN2(16) => A(12), IN2(15) => A(11)
                           , IN2(14) => A(10), IN2(13) => A(9), IN2(12) => A(8)
                           , IN2(11) => A(7), IN2(10) => A(6), IN2(9) => A(5), 
                           IN2(8) => A(4), IN2(7) => A(3), IN2(6) => A(2), 
                           IN2(5) => A(1), IN2(4) => A(0), IN2(3) => 
                           X_Logic0_port, IN2(2) => X_Logic0_port, IN2(1) => 
                           X_Logic0_port, IN2(0) => X_Logic0_port, IN3(31) => 
                           n31, IN3(30) => n36, IN3(29) => n31, IN3(28) => n36,
                           IN3(27) => n32, IN3(26) => n36, IN3(25) => n32, 
                           IN3(24) => n36, IN3(23) => n33, IN3(22) => n34, 
                           IN3(21) => n33, IN3(20) => n34, IN3(19) => 
                           A_minus_15_port, IN3(18) => n2, IN3(17) => n4, 
                           IN3(16) => n6, IN3(15) => n8, IN3(14) => n10, 
                           IN3(13) => n12, IN3(12) => n14, IN3(11) => n16, 
                           IN3(10) => n18, IN3(9) => n20, IN3(8) => n22, IN3(7)
                           => n24, IN3(6) => n26, IN3(5) => n28, IN3(4) => 
                           A_minus_0_port, IN3(3) => X_Logic0_port, IN3(2) => 
                           X_Logic0_port, IN3(1) => X_Logic0_port, IN3(0) => 
                           X_Logic0_port, IN4(31) => n46, IN4(30) => n46, 
                           IN4(29) => n46, IN4(28) => n46, IN4(27) => n46, 
                           IN4(26) => n47, IN4(25) => n46, IN4(24) => n47, 
                           IN4(23) => n45, IN4(22) => n47, IN4(21) => n47, 
                           IN4(20) => n47, IN4(19) => A(14), IN4(18) => A(13), 
                           IN4(17) => A(12), IN4(16) => A(11), IN4(15) => A(10)
                           , IN4(14) => A(9), IN4(13) => A(8), IN4(12) => A(7),
                           IN4(11) => A(6), IN4(10) => A(5), IN4(9) => A(4), 
                           IN4(8) => A(3), IN4(7) => A(2), IN4(6) => A(1), 
                           IN4(5) => A(0), IN4(4) => X_Logic0_port, IN4(3) => 
                           X_Logic0_port, IN4(2) => X_Logic0_port, IN4(1) => 
                           X_Logic0_port, IN4(0) => X_Logic0_port, IN5(31) => 
                           n41, IN5(30) => n41, IN5(29) => n40, IN5(28) => n40,
                           IN5(27) => n39, IN5(26) => n39, IN5(25) => n38, 
                           IN5(24) => n38, IN5(23) => n37, IN5(22) => n37, 
                           IN5(21) => n38, IN5(20) => A_minus_15_port, IN5(19) 
                           => n2, IN5(18) => n4, IN5(17) => n6, IN5(16) => n8, 
                           IN5(15) => n10, IN5(14) => n12, IN5(13) => n14, 
                           IN5(12) => n16, IN5(11) => n18, IN5(10) => n20, 
                           IN5(9) => n22, IN5(8) => n24, IN5(7) => n26, IN5(6) 
                           => n28, IN5(5) => A_minus_0_port, IN5(4) => 
                           X_Logic0_port, IN5(3) => X_Logic0_port, IN5(2) => 
                           X_Logic0_port, IN5(1) => X_Logic0_port, IN5(0) => 
                           X_Logic0_port, SEL_in(2) => encoder_out_8_port, 
                           SEL_in(1) => encoder_out_7_port, SEL_in(0) => 
                           encoder_out_6_port, Z(31) => sum_op_2_31_port, Z(30)
                           => sum_op_2_30_port, Z(29) => sum_op_2_29_port, 
                           Z(28) => sum_op_2_28_port, Z(27) => sum_op_2_27_port
                           , Z(26) => sum_op_2_26_port, Z(25) => 
                           sum_op_2_25_port, Z(24) => sum_op_2_24_port, Z(23) 
                           => sum_op_2_23_port, Z(22) => sum_op_2_22_port, 
                           Z(21) => sum_op_2_21_port, Z(20) => sum_op_2_20_port
                           , Z(19) => sum_op_2_19_port, Z(18) => 
                           sum_op_2_18_port, Z(17) => sum_op_2_17_port, Z(16) 
                           => sum_op_2_16_port, Z(15) => sum_op_2_15_port, 
                           Z(14) => sum_op_2_14_port, Z(13) => sum_op_2_13_port
                           , Z(12) => sum_op_2_12_port, Z(11) => 
                           sum_op_2_11_port, Z(10) => sum_op_2_10_port, Z(9) =>
                           sum_op_2_9_port, Z(8) => sum_op_2_8_port, Z(7) => 
                           sum_op_2_7_port, Z(6) => sum_op_2_6_port, Z(5) => 
                           sum_op_2_5_port, Z(4) => sum_op_2_4_port, Z(3) => 
                           sum_op_2_3_port, Z(2) => sum_op_2_2_port, Z(1) => 
                           sum_op_2_1_port, Z(0) => sum_op_2_0_port);
   mux_i_3 : mux5to1_numBit32_5 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => n52, IN2(30) => n52, 
                           IN2(29) => n50, IN2(28) => n53, IN2(27) => n53, 
                           IN2(26) => n53, IN2(25) => n53, IN2(24) => n53, 
                           IN2(23) => n53, IN2(22) => n53, IN2(21) => n53, 
                           IN2(20) => A(14), IN2(19) => A(13), IN2(18) => A(12)
                           , IN2(17) => A(11), IN2(16) => A(10), IN2(15) => 
                           A(9), IN2(14) => A(8), IN2(13) => A(7), IN2(12) => 
                           A(6), IN2(11) => A(5), IN2(10) => A(4), IN2(9) => 
                           A(3), IN2(8) => A(2), IN2(7) => A(1), IN2(6) => A(0)
                           , IN2(5) => X_Logic0_port, IN2(4) => X_Logic0_port, 
                           IN2(3) => X_Logic0_port, IN2(2) => X_Logic0_port, 
                           IN2(1) => X_Logic0_port, IN2(0) => X_Logic0_port, 
                           IN3(31) => n31, IN3(30) => n35, IN3(29) => n32, 
                           IN3(28) => n35, IN3(27) => n32, IN3(26) => n36, 
                           IN3(25) => n33, IN3(24) => n34, IN3(23) => n33, 
                           IN3(22) => n34, IN3(21) => A_minus_15_port, IN3(20) 
                           => n2, IN3(19) => n4, IN3(18) => n6, IN3(17) => n8, 
                           IN3(16) => n10, IN3(15) => n12, IN3(14) => n14, 
                           IN3(13) => n16, IN3(12) => n18, IN3(11) => n20, 
                           IN3(10) => n22, IN3(9) => n24, IN3(8) => n26, IN3(7)
                           => n28, IN3(6) => A_minus_0_port, IN3(5) => 
                           X_Logic0_port, IN3(4) => X_Logic0_port, IN3(3) => 
                           X_Logic0_port, IN3(2) => X_Logic0_port, IN3(1) => 
                           X_Logic0_port, IN3(0) => X_Logic0_port, IN4(31) => 
                           n45, IN4(30) => n45, IN4(29) => n45, IN4(28) => n45,
                           IN4(27) => n45, IN4(26) => n45, IN4(25) => n45, 
                           IN4(24) => n45, IN4(23) => n45, IN4(22) => n45, 
                           IN4(21) => A(14), IN4(20) => A(13), IN4(19) => A(12)
                           , IN4(18) => A(11), IN4(17) => A(10), IN4(16) => 
                           A(9), IN4(15) => A(8), IN4(14) => A(7), IN4(13) => 
                           A(6), IN4(12) => A(5), IN4(11) => A(4), IN4(10) => 
                           A(3), IN4(9) => A(2), IN4(8) => A(1), IN4(7) => A(0)
                           , IN4(6) => X_Logic0_port, IN4(5) => X_Logic0_port, 
                           IN4(4) => X_Logic0_port, IN4(3) => X_Logic0_port, 
                           IN4(2) => X_Logic0_port, IN4(1) => X_Logic0_port, 
                           IN4(0) => X_Logic0_port, IN5(31) => n40, IN5(30) => 
                           n40, IN5(29) => n39, IN5(28) => n39, IN5(27) => n37,
                           IN5(26) => n38, IN5(25) => n38, IN5(24) => n37, 
                           IN5(23) => n38, IN5(22) => A_minus_15_port, IN5(21) 
                           => n2, IN5(20) => n4, IN5(19) => n6, IN5(18) => n8, 
                           IN5(17) => n10, IN5(16) => n12, IN5(15) => n14, 
                           IN5(14) => n16, IN5(13) => n18, IN5(12) => n20, 
                           IN5(11) => n22, IN5(10) => n24, IN5(9) => n26, 
                           IN5(8) => n28, IN5(7) => A_minus_0_port, IN5(6) => 
                           X_Logic0_port, IN5(5) => X_Logic0_port, IN5(4) => 
                           X_Logic0_port, IN5(3) => X_Logic0_port, IN5(2) => 
                           X_Logic0_port, IN5(1) => X_Logic0_port, IN5(0) => 
                           X_Logic0_port, SEL_in(2) => encoder_out_11_port, 
                           SEL_in(1) => encoder_out_10_port, SEL_in(0) => 
                           encoder_out_9_port, Z(31) => sum_op_3_31_port, Z(30)
                           => sum_op_3_30_port, Z(29) => sum_op_3_29_port, 
                           Z(28) => sum_op_3_28_port, Z(27) => sum_op_3_27_port
                           , Z(26) => sum_op_3_26_port, Z(25) => 
                           sum_op_3_25_port, Z(24) => sum_op_3_24_port, Z(23) 
                           => sum_op_3_23_port, Z(22) => sum_op_3_22_port, 
                           Z(21) => sum_op_3_21_port, Z(20) => sum_op_3_20_port
                           , Z(19) => sum_op_3_19_port, Z(18) => 
                           sum_op_3_18_port, Z(17) => sum_op_3_17_port, Z(16) 
                           => sum_op_3_16_port, Z(15) => sum_op_3_15_port, 
                           Z(14) => sum_op_3_14_port, Z(13) => sum_op_3_13_port
                           , Z(12) => sum_op_3_12_port, Z(11) => 
                           sum_op_3_11_port, Z(10) => sum_op_3_10_port, Z(9) =>
                           sum_op_3_9_port, Z(8) => sum_op_3_8_port, Z(7) => 
                           sum_op_3_7_port, Z(6) => sum_op_3_6_port, Z(5) => 
                           sum_op_3_5_port, Z(4) => sum_op_3_4_port, Z(3) => 
                           sum_op_3_3_port, Z(2) => sum_op_3_2_port, Z(1) => 
                           sum_op_3_1_port, Z(0) => sum_op_3_0_port);
   mux_i_4 : mux5to1_numBit32_4 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => n52, IN2(30) => n52, 
                           IN2(29) => n52, IN2(28) => n52, IN2(27) => n52, 
                           IN2(26) => n52, IN2(25) => n52, IN2(24) => n52, 
                           IN2(23) => n52, IN2(22) => A(14), IN2(21) => A(13), 
                           IN2(20) => A(12), IN2(19) => A(11), IN2(18) => A(10)
                           , IN2(17) => A(9), IN2(16) => A(8), IN2(15) => A(7),
                           IN2(14) => A(6), IN2(13) => A(5), IN2(12) => A(4), 
                           IN2(11) => A(3), IN2(10) => A(2), IN2(9) => A(1), 
                           IN2(8) => A(0), IN2(7) => X_Logic0_port, IN2(6) => 
                           X_Logic0_port, IN2(5) => X_Logic0_port, IN2(4) => 
                           X_Logic0_port, IN2(3) => X_Logic0_port, IN2(2) => 
                           X_Logic0_port, IN2(1) => X_Logic0_port, IN2(0) => 
                           X_Logic0_port, IN3(31) => n31, IN3(30) => n36, 
                           IN3(29) => n32, IN3(28) => n36, IN3(27) => n33, 
                           IN3(26) => n34, IN3(25) => n33, IN3(24) => n34, 
                           IN3(23) => A_minus_15_port, IN3(22) => n2, IN3(21) 
                           => n4, IN3(20) => n6, IN3(19) => n8, IN3(18) => n10,
                           IN3(17) => n12, IN3(16) => n14, IN3(15) => n16, 
                           IN3(14) => n18, IN3(13) => n20, IN3(12) => n22, 
                           IN3(11) => n24, IN3(10) => n26, IN3(9) => n28, 
                           IN3(8) => A_minus_0_port, IN3(7) => X_Logic0_port, 
                           IN3(6) => X_Logic0_port, IN3(5) => X_Logic0_port, 
                           IN3(4) => X_Logic0_port, IN3(3) => X_Logic0_port, 
                           IN3(2) => X_Logic0_port, IN3(1) => X_Logic0_port, 
                           IN3(0) => X_Logic0_port, IN4(31) => n44, IN4(30) => 
                           n44, IN4(29) => n44, IN4(28) => n44, IN4(27) => n44,
                           IN4(26) => n44, IN4(25) => n44, IN4(24) => n44, 
                           IN4(23) => A(14), IN4(22) => A(13), IN4(21) => A(12)
                           , IN4(20) => A(11), IN4(19) => A(10), IN4(18) => 
                           A(9), IN4(17) => A(8), IN4(16) => A(7), IN4(15) => 
                           A(6), IN4(14) => A(5), IN4(13) => A(4), IN4(12) => 
                           A(3), IN4(11) => A(2), IN4(10) => A(1), IN4(9) => 
                           A(0), IN4(8) => X_Logic0_port, IN4(7) => 
                           X_Logic0_port, IN4(6) => X_Logic0_port, IN4(5) => 
                           X_Logic0_port, IN4(4) => X_Logic0_port, IN4(3) => 
                           X_Logic0_port, IN4(2) => X_Logic0_port, IN4(1) => 
                           X_Logic0_port, IN4(0) => X_Logic0_port, IN5(31) => 
                           n39, IN5(30) => n39, IN5(29) => n38, IN5(28) => n41,
                           IN5(27) => n37, IN5(26) => n38, IN5(25) => n39, 
                           IN5(24) => A_minus_15_port, IN5(23) => n2, IN5(22) 
                           => n4, IN5(21) => n6, IN5(20) => n8, IN5(19) => n10,
                           IN5(18) => n12, IN5(17) => n14, IN5(16) => n16, 
                           IN5(15) => n18, IN5(14) => n20, IN5(13) => n22, 
                           IN5(12) => n24, IN5(11) => n26, IN5(10) => n28, 
                           IN5(9) => A_minus_0_port, IN5(8) => X_Logic0_port, 
                           IN5(7) => X_Logic0_port, IN5(6) => X_Logic0_port, 
                           IN5(5) => X_Logic0_port, IN5(4) => X_Logic0_port, 
                           IN5(3) => X_Logic0_port, IN5(2) => X_Logic0_port, 
                           IN5(1) => X_Logic0_port, IN5(0) => X_Logic0_port, 
                           SEL_in(2) => encoder_out_14_port, SEL_in(1) => 
                           encoder_out_13_port, SEL_in(0) => 
                           encoder_out_12_port, Z(31) => sum_op_4_31_port, 
                           Z(30) => sum_op_4_30_port, Z(29) => sum_op_4_29_port
                           , Z(28) => sum_op_4_28_port, Z(27) => 
                           sum_op_4_27_port, Z(26) => sum_op_4_26_port, Z(25) 
                           => sum_op_4_25_port, Z(24) => sum_op_4_24_port, 
                           Z(23) => sum_op_4_23_port, Z(22) => sum_op_4_22_port
                           , Z(21) => sum_op_4_21_port, Z(20) => 
                           sum_op_4_20_port, Z(19) => sum_op_4_19_port, Z(18) 
                           => sum_op_4_18_port, Z(17) => sum_op_4_17_port, 
                           Z(16) => sum_op_4_16_port, Z(15) => sum_op_4_15_port
                           , Z(14) => sum_op_4_14_port, Z(13) => 
                           sum_op_4_13_port, Z(12) => sum_op_4_12_port, Z(11) 
                           => sum_op_4_11_port, Z(10) => sum_op_4_10_port, Z(9)
                           => sum_op_4_9_port, Z(8) => sum_op_4_8_port, Z(7) =>
                           sum_op_4_7_port, Z(6) => sum_op_4_6_port, Z(5) => 
                           sum_op_4_5_port, Z(4) => sum_op_4_4_port, Z(3) => 
                           sum_op_4_3_port, Z(2) => sum_op_4_2_port, Z(1) => 
                           sum_op_4_1_port, Z(0) => sum_op_4_0_port);
   mux_i_5 : mux5to1_numBit32_3 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => n51, IN2(30) => n51, 
                           IN2(29) => n51, IN2(28) => n51, IN2(27) => n51, 
                           IN2(26) => n51, IN2(25) => n51, IN2(24) => A(14), 
                           IN2(23) => A(13), IN2(22) => A(12), IN2(21) => A(11)
                           , IN2(20) => A(10), IN2(19) => A(9), IN2(18) => A(8)
                           , IN2(17) => A(7), IN2(16) => A(6), IN2(15) => A(5),
                           IN2(14) => A(4), IN2(13) => A(3), IN2(12) => A(2), 
                           IN2(11) => A(1), IN2(10) => A(0), IN2(9) => 
                           X_Logic0_port, IN2(8) => X_Logic0_port, IN2(7) => 
                           X_Logic0_port, IN2(6) => X_Logic0_port, IN2(5) => 
                           X_Logic0_port, IN2(4) => X_Logic0_port, IN2(3) => 
                           X_Logic0_port, IN2(2) => X_Logic0_port, IN2(1) => 
                           X_Logic0_port, IN2(0) => X_Logic0_port, IN3(31) => 
                           n32, IN3(30) => n35, IN3(29) => n32, IN3(28) => n35,
                           IN3(27) => n33, IN3(26) => n34, IN3(25) => 
                           A_minus_15_port, IN3(24) => n2, IN3(23) => n4, 
                           IN3(22) => n6, IN3(21) => n8, IN3(20) => n10, 
                           IN3(19) => n12, IN3(18) => n14, IN3(17) => n16, 
                           IN3(16) => n18, IN3(15) => n20, IN3(14) => n22, 
                           IN3(13) => n24, IN3(12) => n26, IN3(11) => n28, 
                           IN3(10) => A_minus_0_port, IN3(9) => X_Logic0_port, 
                           IN3(8) => X_Logic0_port, IN3(7) => X_Logic0_port, 
                           IN3(6) => X_Logic0_port, IN3(5) => X_Logic0_port, 
                           IN3(4) => X_Logic0_port, IN3(3) => X_Logic0_port, 
                           IN3(2) => X_Logic0_port, IN3(1) => X_Logic0_port, 
                           IN3(0) => X_Logic0_port, IN4(31) => n43, IN4(30) => 
                           n43, IN4(29) => n44, IN4(28) => n44, IN4(27) => n44,
                           IN4(26) => n44, IN4(25) => A(14), IN4(24) => A(13), 
                           IN4(23) => A(12), IN4(22) => A(11), IN4(21) => A(10)
                           , IN4(20) => A(9), IN4(19) => A(8), IN4(18) => A(7),
                           IN4(17) => A(6), IN4(16) => A(5), IN4(15) => A(4), 
                           IN4(14) => A(3), IN4(13) => A(2), IN4(12) => A(1), 
                           IN4(11) => A(0), IN4(10) => X_Logic0_port, IN4(9) =>
                           X_Logic0_port, IN4(8) => X_Logic0_port, IN4(7) => 
                           X_Logic0_port, IN4(6) => X_Logic0_port, IN4(5) => 
                           X_Logic0_port, IN4(4) => X_Logic0_port, IN4(3) => 
                           X_Logic0_port, IN4(2) => X_Logic0_port, IN4(1) => 
                           X_Logic0_port, IN4(0) => X_Logic0_port, IN5(31) => 
                           n40, IN5(30) => n39, IN5(29) => n37, IN5(28) => n38,
                           IN5(27) => n37, IN5(26) => A_minus_15_port, IN5(25) 
                           => n2, IN5(24) => n4, IN5(23) => n6, IN5(22) => n8, 
                           IN5(21) => n10, IN5(20) => n12, IN5(19) => n14, 
                           IN5(18) => n16, IN5(17) => n18, IN5(16) => n20, 
                           IN5(15) => n22, IN5(14) => n24, IN5(13) => n26, 
                           IN5(12) => n28, IN5(11) => A_minus_0_port, IN5(10) 
                           => X_Logic0_port, IN5(9) => X_Logic0_port, IN5(8) =>
                           X_Logic0_port, IN5(7) => X_Logic0_port, IN5(6) => 
                           X_Logic0_port, IN5(5) => X_Logic0_port, IN5(4) => 
                           X_Logic0_port, IN5(3) => X_Logic0_port, IN5(2) => 
                           X_Logic0_port, IN5(1) => X_Logic0_port, IN5(0) => 
                           X_Logic0_port, SEL_in(2) => encoder_out_17_port, 
                           SEL_in(1) => encoder_out_16_port, SEL_in(0) => 
                           encoder_out_15_port, Z(31) => sum_op_5_31_port, 
                           Z(30) => sum_op_5_30_port, Z(29) => sum_op_5_29_port
                           , Z(28) => sum_op_5_28_port, Z(27) => 
                           sum_op_5_27_port, Z(26) => sum_op_5_26_port, Z(25) 
                           => sum_op_5_25_port, Z(24) => sum_op_5_24_port, 
                           Z(23) => sum_op_5_23_port, Z(22) => sum_op_5_22_port
                           , Z(21) => sum_op_5_21_port, Z(20) => 
                           sum_op_5_20_port, Z(19) => sum_op_5_19_port, Z(18) 
                           => sum_op_5_18_port, Z(17) => sum_op_5_17_port, 
                           Z(16) => sum_op_5_16_port, Z(15) => sum_op_5_15_port
                           , Z(14) => sum_op_5_14_port, Z(13) => 
                           sum_op_5_13_port, Z(12) => sum_op_5_12_port, Z(11) 
                           => sum_op_5_11_port, Z(10) => sum_op_5_10_port, Z(9)
                           => sum_op_5_9_port, Z(8) => sum_op_5_8_port, Z(7) =>
                           sum_op_5_7_port, Z(6) => sum_op_5_6_port, Z(5) => 
                           sum_op_5_5_port, Z(4) => sum_op_5_4_port, Z(3) => 
                           sum_op_5_3_port, Z(2) => sum_op_5_2_port, Z(1) => 
                           sum_op_5_1_port, Z(0) => sum_op_5_0_port);
   mux_i_6 : mux5to1_numBit32_2 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => n50, IN2(30) => n50, 
                           IN2(29) => n50, IN2(28) => n50, IN2(27) => n50, 
                           IN2(26) => A(14), IN2(25) => A(13), IN2(24) => A(12)
                           , IN2(23) => A(11), IN2(22) => A(10), IN2(21) => 
                           A(9), IN2(20) => A(8), IN2(19) => A(7), IN2(18) => 
                           A(6), IN2(17) => A(5), IN2(16) => A(4), IN2(15) => 
                           A(3), IN2(14) => A(2), IN2(13) => A(1), IN2(12) => 
                           A(0), IN2(11) => X_Logic0_port, IN2(10) => 
                           X_Logic0_port, IN2(9) => X_Logic0_port, IN2(8) => 
                           X_Logic0_port, IN2(7) => X_Logic0_port, IN2(6) => 
                           X_Logic0_port, IN2(5) => X_Logic0_port, IN2(4) => 
                           X_Logic0_port, IN2(3) => X_Logic0_port, IN2(2) => 
                           X_Logic0_port, IN2(1) => X_Logic0_port, IN2(0) => 
                           X_Logic0_port, IN3(31) => n32, IN3(30) => n35, 
                           IN3(29) => n33, IN3(28) => n34, IN3(27) => 
                           A_minus_15_port, IN3(26) => n2, IN3(25) => n4, 
                           IN3(24) => n6, IN3(23) => n8, IN3(22) => n10, 
                           IN3(21) => n12, IN3(20) => n14, IN3(19) => n16, 
                           IN3(18) => n18, IN3(17) => n20, IN3(16) => n22, 
                           IN3(15) => n24, IN3(14) => n26, IN3(13) => n28, 
                           IN3(12) => A_minus_0_port, IN3(11) => X_Logic0_port,
                           IN3(10) => X_Logic0_port, IN3(9) => X_Logic0_port, 
                           IN3(8) => X_Logic0_port, IN3(7) => X_Logic0_port, 
                           IN3(6) => X_Logic0_port, IN3(5) => X_Logic0_port, 
                           IN3(4) => X_Logic0_port, IN3(3) => X_Logic0_port, 
                           IN3(2) => X_Logic0_port, IN3(1) => X_Logic0_port, 
                           IN3(0) => X_Logic0_port, IN4(31) => n43, IN4(30) => 
                           n43, IN4(29) => n43, IN4(28) => n43, IN4(27) => 
                           A(14), IN4(26) => A(13), IN4(25) => A(12), IN4(24) 
                           => A(11), IN4(23) => A(10), IN4(22) => A(9), IN4(21)
                           => A(8), IN4(20) => A(7), IN4(19) => A(6), IN4(18) 
                           => A(5), IN4(17) => A(4), IN4(16) => A(3), IN4(15) 
                           => A(2), IN4(14) => A(1), IN4(13) => A(0), IN4(12) 
                           => X_Logic0_port, IN4(11) => X_Logic0_port, IN4(10) 
                           => X_Logic0_port, IN4(9) => X_Logic0_port, IN4(8) =>
                           X_Logic0_port, IN4(7) => X_Logic0_port, IN4(6) => 
                           X_Logic0_port, IN4(5) => X_Logic0_port, IN4(4) => 
                           X_Logic0_port, IN4(3) => X_Logic0_port, IN4(2) => 
                           X_Logic0_port, IN4(1) => X_Logic0_port, IN4(0) => 
                           X_Logic0_port, IN5(31) => n37, IN5(30) => n38, 
                           IN5(29) => n37, IN5(28) => A_minus_15_port, IN5(27) 
                           => n2, IN5(26) => n4, IN5(25) => n6, IN5(24) => n8, 
                           IN5(23) => n10, IN5(22) => n12, IN5(21) => n14, 
                           IN5(20) => n16, IN5(19) => n18, IN5(18) => n20, 
                           IN5(17) => n22, IN5(16) => n24, IN5(15) => n26, 
                           IN5(14) => n28, IN5(13) => A_minus_0_port, IN5(12) 
                           => X_Logic0_port, IN5(11) => X_Logic0_port, IN5(10) 
                           => X_Logic0_port, IN5(9) => X_Logic0_port, IN5(8) =>
                           X_Logic0_port, IN5(7) => X_Logic0_port, IN5(6) => 
                           X_Logic0_port, IN5(5) => X_Logic0_port, IN5(4) => 
                           X_Logic0_port, IN5(3) => X_Logic0_port, IN5(2) => 
                           X_Logic0_port, IN5(1) => X_Logic0_port, IN5(0) => 
                           X_Logic0_port, SEL_in(2) => encoder_out_20_port, 
                           SEL_in(1) => encoder_out_19_port, SEL_in(0) => 
                           encoder_out_18_port, Z(31) => sum_op_6_31_port, 
                           Z(30) => sum_op_6_30_port, Z(29) => sum_op_6_29_port
                           , Z(28) => sum_op_6_28_port, Z(27) => 
                           sum_op_6_27_port, Z(26) => sum_op_6_26_port, Z(25) 
                           => sum_op_6_25_port, Z(24) => sum_op_6_24_port, 
                           Z(23) => sum_op_6_23_port, Z(22) => sum_op_6_22_port
                           , Z(21) => sum_op_6_21_port, Z(20) => 
                           sum_op_6_20_port, Z(19) => sum_op_6_19_port, Z(18) 
                           => sum_op_6_18_port, Z(17) => sum_op_6_17_port, 
                           Z(16) => sum_op_6_16_port, Z(15) => sum_op_6_15_port
                           , Z(14) => sum_op_6_14_port, Z(13) => 
                           sum_op_6_13_port, Z(12) => sum_op_6_12_port, Z(11) 
                           => sum_op_6_11_port, Z(10) => sum_op_6_10_port, Z(9)
                           => sum_op_6_9_port, Z(8) => sum_op_6_8_port, Z(7) =>
                           sum_op_6_7_port, Z(6) => sum_op_6_6_port, Z(5) => 
                           sum_op_6_5_port, Z(4) => sum_op_6_4_port, Z(3) => 
                           sum_op_6_3_port, Z(2) => sum_op_6_2_port, Z(1) => 
                           sum_op_6_1_port, Z(0) => sum_op_6_0_port);
   mux_i_7 : mux5to1_numBit32_1 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => n49, IN2(30) => n49, 
                           IN2(29) => n50, IN2(28) => A(14), IN2(27) => A(13), 
                           IN2(26) => A(12), IN2(25) => A(11), IN2(24) => A(10)
                           , IN2(23) => A(9), IN2(22) => A(8), IN2(21) => A(7),
                           IN2(20) => A(6), IN2(19) => A(5), IN2(18) => A(4), 
                           IN2(17) => A(3), IN2(16) => A(2), IN2(15) => A(1), 
                           IN2(14) => A(0), IN2(13) => X_Logic0_port, IN2(12) 
                           => X_Logic0_port, IN2(11) => X_Logic0_port, IN2(10) 
                           => X_Logic0_port, IN2(9) => X_Logic0_port, IN2(8) =>
                           X_Logic0_port, IN2(7) => X_Logic0_port, IN2(6) => 
                           X_Logic0_port, IN2(5) => X_Logic0_port, IN2(4) => 
                           X_Logic0_port, IN2(3) => X_Logic0_port, IN2(2) => 
                           X_Logic0_port, IN2(1) => X_Logic0_port, IN2(0) => 
                           X_Logic0_port, IN3(31) => n33, IN3(30) => n34, 
                           IN3(29) => A_minus_15_port, IN3(28) => n2, IN3(27) 
                           => n4, IN3(26) => n6, IN3(25) => n8, IN3(24) => n10,
                           IN3(23) => n12, IN3(22) => n14, IN3(21) => n16, 
                           IN3(20) => n18, IN3(19) => n20, IN3(18) => n22, 
                           IN3(17) => n24, IN3(16) => n26, IN3(15) => n28, 
                           IN3(14) => A_minus_0_port, IN3(13) => X_Logic0_port,
                           IN3(12) => X_Logic0_port, IN3(11) => X_Logic0_port, 
                           IN3(10) => X_Logic0_port, IN3(9) => X_Logic0_port, 
                           IN3(8) => X_Logic0_port, IN3(7) => X_Logic0_port, 
                           IN3(6) => X_Logic0_port, IN3(5) => X_Logic0_port, 
                           IN3(4) => X_Logic0_port, IN3(3) => X_Logic0_port, 
                           IN3(2) => X_Logic0_port, IN3(1) => X_Logic0_port, 
                           IN3(0) => X_Logic0_port, IN4(31) => n43, IN4(30) => 
                           n45, IN4(29) => A(14), IN4(28) => A(13), IN4(27) => 
                           A(12), IN4(26) => A(11), IN4(25) => A(10), IN4(24) 
                           => A(9), IN4(23) => A(8), IN4(22) => A(7), IN4(21) 
                           => A(6), IN4(20) => A(5), IN4(19) => A(4), IN4(18) 
                           => A(3), IN4(17) => A(2), IN4(16) => A(1), IN4(15) 
                           => A(0), IN4(14) => X_Logic0_port, IN4(13) => 
                           X_Logic0_port, IN4(12) => X_Logic0_port, IN4(11) => 
                           X_Logic0_port, IN4(10) => X_Logic0_port, IN4(9) => 
                           X_Logic0_port, IN4(8) => X_Logic0_port, IN4(7) => 
                           X_Logic0_port, IN4(6) => X_Logic0_port, IN4(5) => 
                           X_Logic0_port, IN4(4) => X_Logic0_port, IN4(3) => 
                           X_Logic0_port, IN4(2) => X_Logic0_port, IN4(1) => 
                           X_Logic0_port, IN4(0) => X_Logic0_port, IN5(31) => 
                           n37, IN5(30) => A_minus_15_port, IN5(29) => n2, 
                           IN5(28) => n4, IN5(27) => n6, IN5(26) => n8, IN5(25)
                           => n10, IN5(24) => n12, IN5(23) => n14, IN5(22) => 
                           n16, IN5(21) => n18, IN5(20) => n20, IN5(19) => n22,
                           IN5(18) => n24, IN5(17) => n26, IN5(16) => n28, 
                           IN5(15) => A_minus_0_port, IN5(14) => X_Logic0_port,
                           IN5(13) => X_Logic0_port, IN5(12) => X_Logic0_port, 
                           IN5(11) => X_Logic0_port, IN5(10) => X_Logic0_port, 
                           IN5(9) => X_Logic0_port, IN5(8) => X_Logic0_port, 
                           IN5(7) => X_Logic0_port, IN5(6) => X_Logic0_port, 
                           IN5(5) => X_Logic0_port, IN5(4) => X_Logic0_port, 
                           IN5(3) => X_Logic0_port, IN5(2) => X_Logic0_port, 
                           IN5(1) => X_Logic0_port, IN5(0) => X_Logic0_port, 
                           SEL_in(2) => encoder_out_23_port, SEL_in(1) => 
                           encoder_out_22_port, SEL_in(0) => 
                           encoder_out_21_port, Z(31) => sum_op_7_31_port, 
                           Z(30) => sum_op_7_30_port, Z(29) => sum_op_7_29_port
                           , Z(28) => sum_op_7_28_port, Z(27) => 
                           sum_op_7_27_port, Z(26) => sum_op_7_26_port, Z(25) 
                           => sum_op_7_25_port, Z(24) => sum_op_7_24_port, 
                           Z(23) => sum_op_7_23_port, Z(22) => sum_op_7_22_port
                           , Z(21) => sum_op_7_21_port, Z(20) => 
                           sum_op_7_20_port, Z(19) => sum_op_7_19_port, Z(18) 
                           => sum_op_7_18_port, Z(17) => sum_op_7_17_port, 
                           Z(16) => sum_op_7_16_port, Z(15) => sum_op_7_15_port
                           , Z(14) => sum_op_7_14_port, Z(13) => 
                           sum_op_7_13_port, Z(12) => sum_op_7_12_port, Z(11) 
                           => sum_op_7_11_port, Z(10) => sum_op_7_10_port, Z(9)
                           => sum_op_7_9_port, Z(8) => sum_op_7_8_port, Z(7) =>
                           sum_op_7_7_port, Z(6) => sum_op_7_6_port, Z(5) => 
                           sum_op_7_5_port, Z(4) => sum_op_7_4_port, Z(3) => 
                           sum_op_7_3_port, Z(2) => sum_op_7_2_port, Z(1) => 
                           sum_op_7_1_port, Z(0) => sum_op_7_0_port);
   rca0_0 : rca_bhv_numBit32_0 port map( A(31) => sum_op_0_31_port, A(30) => 
                           sum_op_0_30_port, A(29) => sum_op_0_29_port, A(28) 
                           => sum_op_0_28_port, A(27) => sum_op_0_27_port, 
                           A(26) => sum_op_0_26_port, A(25) => sum_op_0_25_port
                           , A(24) => sum_op_0_24_port, A(23) => 
                           sum_op_0_23_port, A(22) => sum_op_0_22_port, A(21) 
                           => sum_op_0_21_port, A(20) => sum_op_0_20_port, 
                           A(19) => sum_op_0_19_port, A(18) => sum_op_0_18_port
                           , A(17) => sum_op_0_17_port, A(16) => 
                           sum_op_0_16_port, A(15) => sum_op_0_15_port, A(14) 
                           => sum_op_0_14_port, A(13) => sum_op_0_13_port, 
                           A(12) => sum_op_0_12_port, A(11) => sum_op_0_11_port
                           , A(10) => sum_op_0_10_port, A(9) => sum_op_0_9_port
                           , A(8) => sum_op_0_8_port, A(7) => sum_op_0_7_port, 
                           A(6) => sum_op_0_6_port, A(5) => sum_op_0_5_port, 
                           A(4) => sum_op_0_4_port, A(3) => sum_op_0_3_port, 
                           A(2) => sum_op_0_2_port, A(1) => sum_op_0_1_port, 
                           A(0) => sum_op_0_0_port, B(31) => sum_op_1_31_port, 
                           B(30) => sum_op_1_30_port, B(29) => sum_op_1_29_port
                           , B(28) => sum_op_1_28_port, B(27) => 
                           sum_op_1_27_port, B(26) => sum_op_1_26_port, B(25) 
                           => sum_op_1_25_port, B(24) => sum_op_1_24_port, 
                           B(23) => sum_op_1_23_port, B(22) => sum_op_1_22_port
                           , B(21) => sum_op_1_21_port, B(20) => 
                           sum_op_1_20_port, B(19) => sum_op_1_19_port, B(18) 
                           => sum_op_1_18_port, B(17) => sum_op_1_17_port, 
                           B(16) => sum_op_1_16_port, B(15) => sum_op_1_15_port
                           , B(14) => sum_op_1_14_port, B(13) => 
                           sum_op_1_13_port, B(12) => sum_op_1_12_port, B(11) 
                           => sum_op_1_11_port, B(10) => sum_op_1_10_port, B(9)
                           => sum_op_1_9_port, B(8) => sum_op_1_8_port, B(7) =>
                           sum_op_1_7_port, B(6) => sum_op_1_6_port, B(5) => 
                           sum_op_1_5_port, B(4) => sum_op_1_4_port, B(3) => 
                           sum_op_1_3_port, B(2) => sum_op_1_2_port, B(1) => 
                           sum_op_1_1_port, B(0) => sum_op_1_0_port, Ci => 
                           X_Logic0_port, S(31) => rca_out_0_31_port, S(30) => 
                           rca_out_0_30_port, S(29) => rca_out_0_29_port, S(28)
                           => rca_out_0_28_port, S(27) => rca_out_0_27_port, 
                           S(26) => rca_out_0_26_port, S(25) => 
                           rca_out_0_25_port, S(24) => rca_out_0_24_port, S(23)
                           => rca_out_0_23_port, S(22) => rca_out_0_22_port, 
                           S(21) => rca_out_0_21_port, S(20) => 
                           rca_out_0_20_port, S(19) => rca_out_0_19_port, S(18)
                           => rca_out_0_18_port, S(17) => rca_out_0_17_port, 
                           S(16) => rca_out_0_16_port, S(15) => 
                           rca_out_0_15_port, S(14) => rca_out_0_14_port, S(13)
                           => rca_out_0_13_port, S(12) => rca_out_0_12_port, 
                           S(11) => rca_out_0_11_port, S(10) => 
                           rca_out_0_10_port, S(9) => rca_out_0_9_port, S(8) =>
                           rca_out_0_8_port, S(7) => rca_out_0_7_port, S(6) => 
                           rca_out_0_6_port, S(5) => rca_out_0_5_port, S(4) => 
                           rca_out_0_4_port, S(3) => rca_out_0_3_port, S(2) => 
                           rca_out_0_2_port, S(1) => rca_out_0_1_port, S(0) => 
                           rca_out_0_0_port, Co => n_1158);
   rca_i_1 : rca_bhv_numBit32_6 port map( A(31) => rca_out_0_31_port, A(30) => 
                           rca_out_0_30_port, A(29) => rca_out_0_29_port, A(28)
                           => rca_out_0_28_port, A(27) => rca_out_0_27_port, 
                           A(26) => rca_out_0_26_port, A(25) => 
                           rca_out_0_25_port, A(24) => rca_out_0_24_port, A(23)
                           => rca_out_0_23_port, A(22) => rca_out_0_22_port, 
                           A(21) => rca_out_0_21_port, A(20) => 
                           rca_out_0_20_port, A(19) => rca_out_0_19_port, A(18)
                           => rca_out_0_18_port, A(17) => rca_out_0_17_port, 
                           A(16) => rca_out_0_16_port, A(15) => 
                           rca_out_0_15_port, A(14) => rca_out_0_14_port, A(13)
                           => rca_out_0_13_port, A(12) => rca_out_0_12_port, 
                           A(11) => rca_out_0_11_port, A(10) => 
                           rca_out_0_10_port, A(9) => rca_out_0_9_port, A(8) =>
                           rca_out_0_8_port, A(7) => rca_out_0_7_port, A(6) => 
                           rca_out_0_6_port, A(5) => rca_out_0_5_port, A(4) => 
                           rca_out_0_4_port, A(3) => rca_out_0_3_port, A(2) => 
                           rca_out_0_2_port, A(1) => rca_out_0_1_port, A(0) => 
                           rca_out_0_0_port, B(31) => sum_op_2_31_port, B(30) 
                           => sum_op_2_30_port, B(29) => sum_op_2_29_port, 
                           B(28) => sum_op_2_28_port, B(27) => sum_op_2_27_port
                           , B(26) => sum_op_2_26_port, B(25) => 
                           sum_op_2_25_port, B(24) => sum_op_2_24_port, B(23) 
                           => sum_op_2_23_port, B(22) => sum_op_2_22_port, 
                           B(21) => sum_op_2_21_port, B(20) => sum_op_2_20_port
                           , B(19) => sum_op_2_19_port, B(18) => 
                           sum_op_2_18_port, B(17) => sum_op_2_17_port, B(16) 
                           => sum_op_2_16_port, B(15) => sum_op_2_15_port, 
                           B(14) => sum_op_2_14_port, B(13) => sum_op_2_13_port
                           , B(12) => sum_op_2_12_port, B(11) => 
                           sum_op_2_11_port, B(10) => sum_op_2_10_port, B(9) =>
                           sum_op_2_9_port, B(8) => sum_op_2_8_port, B(7) => 
                           sum_op_2_7_port, B(6) => sum_op_2_6_port, B(5) => 
                           sum_op_2_5_port, B(4) => sum_op_2_4_port, B(3) => 
                           sum_op_2_3_port, B(2) => sum_op_2_2_port, B(1) => 
                           sum_op_2_1_port, B(0) => sum_op_2_0_port, Ci => 
                           X_Logic0_port, S(31) => rca_out_1_31_port, S(30) => 
                           rca_out_1_30_port, S(29) => rca_out_1_29_port, S(28)
                           => rca_out_1_28_port, S(27) => rca_out_1_27_port, 
                           S(26) => rca_out_1_26_port, S(25) => 
                           rca_out_1_25_port, S(24) => rca_out_1_24_port, S(23)
                           => rca_out_1_23_port, S(22) => rca_out_1_22_port, 
                           S(21) => rca_out_1_21_port, S(20) => 
                           rca_out_1_20_port, S(19) => rca_out_1_19_port, S(18)
                           => rca_out_1_18_port, S(17) => rca_out_1_17_port, 
                           S(16) => rca_out_1_16_port, S(15) => 
                           rca_out_1_15_port, S(14) => rca_out_1_14_port, S(13)
                           => rca_out_1_13_port, S(12) => rca_out_1_12_port, 
                           S(11) => rca_out_1_11_port, S(10) => 
                           rca_out_1_10_port, S(9) => rca_out_1_9_port, S(8) =>
                           rca_out_1_8_port, S(7) => rca_out_1_7_port, S(6) => 
                           rca_out_1_6_port, S(5) => rca_out_1_5_port, S(4) => 
                           rca_out_1_4_port, S(3) => rca_out_1_3_port, S(2) => 
                           rca_out_1_2_port, S(1) => rca_out_1_1_port, S(0) => 
                           rca_out_1_0_port, Co => n_1159);
   rca_i_2 : rca_bhv_numBit32_5 port map( A(31) => rca_out_1_31_port, A(30) => 
                           rca_out_1_30_port, A(29) => rca_out_1_29_port, A(28)
                           => rca_out_1_28_port, A(27) => rca_out_1_27_port, 
                           A(26) => rca_out_1_26_port, A(25) => 
                           rca_out_1_25_port, A(24) => rca_out_1_24_port, A(23)
                           => rca_out_1_23_port, A(22) => rca_out_1_22_port, 
                           A(21) => rca_out_1_21_port, A(20) => 
                           rca_out_1_20_port, A(19) => rca_out_1_19_port, A(18)
                           => rca_out_1_18_port, A(17) => rca_out_1_17_port, 
                           A(16) => rca_out_1_16_port, A(15) => 
                           rca_out_1_15_port, A(14) => rca_out_1_14_port, A(13)
                           => rca_out_1_13_port, A(12) => rca_out_1_12_port, 
                           A(11) => rca_out_1_11_port, A(10) => 
                           rca_out_1_10_port, A(9) => rca_out_1_9_port, A(8) =>
                           rca_out_1_8_port, A(7) => rca_out_1_7_port, A(6) => 
                           rca_out_1_6_port, A(5) => rca_out_1_5_port, A(4) => 
                           rca_out_1_4_port, A(3) => rca_out_1_3_port, A(2) => 
                           rca_out_1_2_port, A(1) => rca_out_1_1_port, A(0) => 
                           rca_out_1_0_port, B(31) => sum_op_3_31_port, B(30) 
                           => sum_op_3_30_port, B(29) => sum_op_3_29_port, 
                           B(28) => sum_op_3_28_port, B(27) => sum_op_3_27_port
                           , B(26) => sum_op_3_26_port, B(25) => 
                           sum_op_3_25_port, B(24) => sum_op_3_24_port, B(23) 
                           => sum_op_3_23_port, B(22) => sum_op_3_22_port, 
                           B(21) => sum_op_3_21_port, B(20) => sum_op_3_20_port
                           , B(19) => sum_op_3_19_port, B(18) => 
                           sum_op_3_18_port, B(17) => sum_op_3_17_port, B(16) 
                           => sum_op_3_16_port, B(15) => sum_op_3_15_port, 
                           B(14) => sum_op_3_14_port, B(13) => sum_op_3_13_port
                           , B(12) => sum_op_3_12_port, B(11) => 
                           sum_op_3_11_port, B(10) => sum_op_3_10_port, B(9) =>
                           sum_op_3_9_port, B(8) => sum_op_3_8_port, B(7) => 
                           sum_op_3_7_port, B(6) => sum_op_3_6_port, B(5) => 
                           sum_op_3_5_port, B(4) => sum_op_3_4_port, B(3) => 
                           sum_op_3_3_port, B(2) => sum_op_3_2_port, B(1) => 
                           sum_op_3_1_port, B(0) => sum_op_3_0_port, Ci => 
                           X_Logic0_port, S(31) => rca_out_2_31_port, S(30) => 
                           rca_out_2_30_port, S(29) => rca_out_2_29_port, S(28)
                           => rca_out_2_28_port, S(27) => rca_out_2_27_port, 
                           S(26) => rca_out_2_26_port, S(25) => 
                           rca_out_2_25_port, S(24) => rca_out_2_24_port, S(23)
                           => rca_out_2_23_port, S(22) => rca_out_2_22_port, 
                           S(21) => rca_out_2_21_port, S(20) => 
                           rca_out_2_20_port, S(19) => rca_out_2_19_port, S(18)
                           => rca_out_2_18_port, S(17) => rca_out_2_17_port, 
                           S(16) => rca_out_2_16_port, S(15) => 
                           rca_out_2_15_port, S(14) => rca_out_2_14_port, S(13)
                           => rca_out_2_13_port, S(12) => rca_out_2_12_port, 
                           S(11) => rca_out_2_11_port, S(10) => 
                           rca_out_2_10_port, S(9) => rca_out_2_9_port, S(8) =>
                           rca_out_2_8_port, S(7) => rca_out_2_7_port, S(6) => 
                           rca_out_2_6_port, S(5) => rca_out_2_5_port, S(4) => 
                           rca_out_2_4_port, S(3) => rca_out_2_3_port, S(2) => 
                           rca_out_2_2_port, S(1) => rca_out_2_1_port, S(0) => 
                           rca_out_2_0_port, Co => n_1160);
   rca_i_3 : rca_bhv_numBit32_4 port map( A(31) => rca_out_2_31_port, A(30) => 
                           rca_out_2_30_port, A(29) => rca_out_2_29_port, A(28)
                           => rca_out_2_28_port, A(27) => rca_out_2_27_port, 
                           A(26) => rca_out_2_26_port, A(25) => 
                           rca_out_2_25_port, A(24) => rca_out_2_24_port, A(23)
                           => rca_out_2_23_port, A(22) => rca_out_2_22_port, 
                           A(21) => rca_out_2_21_port, A(20) => 
                           rca_out_2_20_port, A(19) => rca_out_2_19_port, A(18)
                           => rca_out_2_18_port, A(17) => rca_out_2_17_port, 
                           A(16) => rca_out_2_16_port, A(15) => 
                           rca_out_2_15_port, A(14) => rca_out_2_14_port, A(13)
                           => rca_out_2_13_port, A(12) => rca_out_2_12_port, 
                           A(11) => rca_out_2_11_port, A(10) => 
                           rca_out_2_10_port, A(9) => rca_out_2_9_port, A(8) =>
                           rca_out_2_8_port, A(7) => rca_out_2_7_port, A(6) => 
                           rca_out_2_6_port, A(5) => rca_out_2_5_port, A(4) => 
                           rca_out_2_4_port, A(3) => rca_out_2_3_port, A(2) => 
                           rca_out_2_2_port, A(1) => rca_out_2_1_port, A(0) => 
                           rca_out_2_0_port, B(31) => sum_op_4_31_port, B(30) 
                           => sum_op_4_30_port, B(29) => sum_op_4_29_port, 
                           B(28) => sum_op_4_28_port, B(27) => sum_op_4_27_port
                           , B(26) => sum_op_4_26_port, B(25) => 
                           sum_op_4_25_port, B(24) => sum_op_4_24_port, B(23) 
                           => sum_op_4_23_port, B(22) => sum_op_4_22_port, 
                           B(21) => sum_op_4_21_port, B(20) => sum_op_4_20_port
                           , B(19) => sum_op_4_19_port, B(18) => 
                           sum_op_4_18_port, B(17) => sum_op_4_17_port, B(16) 
                           => sum_op_4_16_port, B(15) => sum_op_4_15_port, 
                           B(14) => sum_op_4_14_port, B(13) => sum_op_4_13_port
                           , B(12) => sum_op_4_12_port, B(11) => 
                           sum_op_4_11_port, B(10) => sum_op_4_10_port, B(9) =>
                           sum_op_4_9_port, B(8) => sum_op_4_8_port, B(7) => 
                           sum_op_4_7_port, B(6) => sum_op_4_6_port, B(5) => 
                           sum_op_4_5_port, B(4) => sum_op_4_4_port, B(3) => 
                           sum_op_4_3_port, B(2) => sum_op_4_2_port, B(1) => 
                           sum_op_4_1_port, B(0) => sum_op_4_0_port, Ci => 
                           X_Logic0_port, S(31) => rca_out_3_31_port, S(30) => 
                           rca_out_3_30_port, S(29) => rca_out_3_29_port, S(28)
                           => rca_out_3_28_port, S(27) => rca_out_3_27_port, 
                           S(26) => rca_out_3_26_port, S(25) => 
                           rca_out_3_25_port, S(24) => rca_out_3_24_port, S(23)
                           => rca_out_3_23_port, S(22) => rca_out_3_22_port, 
                           S(21) => rca_out_3_21_port, S(20) => 
                           rca_out_3_20_port, S(19) => rca_out_3_19_port, S(18)
                           => rca_out_3_18_port, S(17) => rca_out_3_17_port, 
                           S(16) => rca_out_3_16_port, S(15) => 
                           rca_out_3_15_port, S(14) => rca_out_3_14_port, S(13)
                           => rca_out_3_13_port, S(12) => rca_out_3_12_port, 
                           S(11) => rca_out_3_11_port, S(10) => 
                           rca_out_3_10_port, S(9) => rca_out_3_9_port, S(8) =>
                           rca_out_3_8_port, S(7) => rca_out_3_7_port, S(6) => 
                           rca_out_3_6_port, S(5) => rca_out_3_5_port, S(4) => 
                           rca_out_3_4_port, S(3) => rca_out_3_3_port, S(2) => 
                           rca_out_3_2_port, S(1) => rca_out_3_1_port, S(0) => 
                           rca_out_3_0_port, Co => n_1161);
   rca_i_4 : rca_bhv_numBit32_3 port map( A(31) => rca_out_3_31_port, A(30) => 
                           rca_out_3_30_port, A(29) => rca_out_3_29_port, A(28)
                           => rca_out_3_28_port, A(27) => rca_out_3_27_port, 
                           A(26) => rca_out_3_26_port, A(25) => 
                           rca_out_3_25_port, A(24) => rca_out_3_24_port, A(23)
                           => rca_out_3_23_port, A(22) => rca_out_3_22_port, 
                           A(21) => rca_out_3_21_port, A(20) => 
                           rca_out_3_20_port, A(19) => rca_out_3_19_port, A(18)
                           => rca_out_3_18_port, A(17) => rca_out_3_17_port, 
                           A(16) => rca_out_3_16_port, A(15) => 
                           rca_out_3_15_port, A(14) => rca_out_3_14_port, A(13)
                           => rca_out_3_13_port, A(12) => rca_out_3_12_port, 
                           A(11) => rca_out_3_11_port, A(10) => 
                           rca_out_3_10_port, A(9) => rca_out_3_9_port, A(8) =>
                           rca_out_3_8_port, A(7) => rca_out_3_7_port, A(6) => 
                           rca_out_3_6_port, A(5) => rca_out_3_5_port, A(4) => 
                           rca_out_3_4_port, A(3) => rca_out_3_3_port, A(2) => 
                           rca_out_3_2_port, A(1) => rca_out_3_1_port, A(0) => 
                           rca_out_3_0_port, B(31) => sum_op_5_31_port, B(30) 
                           => sum_op_5_30_port, B(29) => sum_op_5_29_port, 
                           B(28) => sum_op_5_28_port, B(27) => sum_op_5_27_port
                           , B(26) => sum_op_5_26_port, B(25) => 
                           sum_op_5_25_port, B(24) => sum_op_5_24_port, B(23) 
                           => sum_op_5_23_port, B(22) => sum_op_5_22_port, 
                           B(21) => sum_op_5_21_port, B(20) => sum_op_5_20_port
                           , B(19) => sum_op_5_19_port, B(18) => 
                           sum_op_5_18_port, B(17) => sum_op_5_17_port, B(16) 
                           => sum_op_5_16_port, B(15) => sum_op_5_15_port, 
                           B(14) => sum_op_5_14_port, B(13) => sum_op_5_13_port
                           , B(12) => sum_op_5_12_port, B(11) => 
                           sum_op_5_11_port, B(10) => sum_op_5_10_port, B(9) =>
                           sum_op_5_9_port, B(8) => sum_op_5_8_port, B(7) => 
                           sum_op_5_7_port, B(6) => sum_op_5_6_port, B(5) => 
                           sum_op_5_5_port, B(4) => sum_op_5_4_port, B(3) => 
                           sum_op_5_3_port, B(2) => sum_op_5_2_port, B(1) => 
                           sum_op_5_1_port, B(0) => sum_op_5_0_port, Ci => 
                           X_Logic0_port, S(31) => rca_out_4_31_port, S(30) => 
                           rca_out_4_30_port, S(29) => rca_out_4_29_port, S(28)
                           => rca_out_4_28_port, S(27) => rca_out_4_27_port, 
                           S(26) => rca_out_4_26_port, S(25) => 
                           rca_out_4_25_port, S(24) => rca_out_4_24_port, S(23)
                           => rca_out_4_23_port, S(22) => rca_out_4_22_port, 
                           S(21) => rca_out_4_21_port, S(20) => 
                           rca_out_4_20_port, S(19) => rca_out_4_19_port, S(18)
                           => rca_out_4_18_port, S(17) => rca_out_4_17_port, 
                           S(16) => rca_out_4_16_port, S(15) => 
                           rca_out_4_15_port, S(14) => rca_out_4_14_port, S(13)
                           => rca_out_4_13_port, S(12) => rca_out_4_12_port, 
                           S(11) => rca_out_4_11_port, S(10) => 
                           rca_out_4_10_port, S(9) => rca_out_4_9_port, S(8) =>
                           rca_out_4_8_port, S(7) => rca_out_4_7_port, S(6) => 
                           rca_out_4_6_port, S(5) => rca_out_4_5_port, S(4) => 
                           rca_out_4_4_port, S(3) => rca_out_4_3_port, S(2) => 
                           rca_out_4_2_port, S(1) => rca_out_4_1_port, S(0) => 
                           rca_out_4_0_port, Co => n_1162);
   rca_i_5 : rca_bhv_numBit32_2 port map( A(31) => rca_out_4_31_port, A(30) => 
                           rca_out_4_30_port, A(29) => rca_out_4_29_port, A(28)
                           => rca_out_4_28_port, A(27) => rca_out_4_27_port, 
                           A(26) => rca_out_4_26_port, A(25) => 
                           rca_out_4_25_port, A(24) => rca_out_4_24_port, A(23)
                           => rca_out_4_23_port, A(22) => rca_out_4_22_port, 
                           A(21) => rca_out_4_21_port, A(20) => 
                           rca_out_4_20_port, A(19) => rca_out_4_19_port, A(18)
                           => rca_out_4_18_port, A(17) => rca_out_4_17_port, 
                           A(16) => rca_out_4_16_port, A(15) => 
                           rca_out_4_15_port, A(14) => rca_out_4_14_port, A(13)
                           => rca_out_4_13_port, A(12) => rca_out_4_12_port, 
                           A(11) => rca_out_4_11_port, A(10) => 
                           rca_out_4_10_port, A(9) => rca_out_4_9_port, A(8) =>
                           rca_out_4_8_port, A(7) => rca_out_4_7_port, A(6) => 
                           rca_out_4_6_port, A(5) => rca_out_4_5_port, A(4) => 
                           rca_out_4_4_port, A(3) => rca_out_4_3_port, A(2) => 
                           rca_out_4_2_port, A(1) => rca_out_4_1_port, A(0) => 
                           rca_out_4_0_port, B(31) => sum_op_6_31_port, B(30) 
                           => sum_op_6_30_port, B(29) => sum_op_6_29_port, 
                           B(28) => sum_op_6_28_port, B(27) => sum_op_6_27_port
                           , B(26) => sum_op_6_26_port, B(25) => 
                           sum_op_6_25_port, B(24) => sum_op_6_24_port, B(23) 
                           => sum_op_6_23_port, B(22) => sum_op_6_22_port, 
                           B(21) => sum_op_6_21_port, B(20) => sum_op_6_20_port
                           , B(19) => sum_op_6_19_port, B(18) => 
                           sum_op_6_18_port, B(17) => sum_op_6_17_port, B(16) 
                           => sum_op_6_16_port, B(15) => sum_op_6_15_port, 
                           B(14) => sum_op_6_14_port, B(13) => sum_op_6_13_port
                           , B(12) => sum_op_6_12_port, B(11) => 
                           sum_op_6_11_port, B(10) => sum_op_6_10_port, B(9) =>
                           sum_op_6_9_port, B(8) => sum_op_6_8_port, B(7) => 
                           sum_op_6_7_port, B(6) => sum_op_6_6_port, B(5) => 
                           sum_op_6_5_port, B(4) => sum_op_6_4_port, B(3) => 
                           sum_op_6_3_port, B(2) => sum_op_6_2_port, B(1) => 
                           sum_op_6_1_port, B(0) => sum_op_6_0_port, Ci => 
                           X_Logic0_port, S(31) => rca_out_5_31_port, S(30) => 
                           rca_out_5_30_port, S(29) => rca_out_5_29_port, S(28)
                           => rca_out_5_28_port, S(27) => rca_out_5_27_port, 
                           S(26) => rca_out_5_26_port, S(25) => 
                           rca_out_5_25_port, S(24) => rca_out_5_24_port, S(23)
                           => rca_out_5_23_port, S(22) => rca_out_5_22_port, 
                           S(21) => rca_out_5_21_port, S(20) => 
                           rca_out_5_20_port, S(19) => rca_out_5_19_port, S(18)
                           => rca_out_5_18_port, S(17) => rca_out_5_17_port, 
                           S(16) => rca_out_5_16_port, S(15) => 
                           rca_out_5_15_port, S(14) => rca_out_5_14_port, S(13)
                           => rca_out_5_13_port, S(12) => rca_out_5_12_port, 
                           S(11) => rca_out_5_11_port, S(10) => 
                           rca_out_5_10_port, S(9) => rca_out_5_9_port, S(8) =>
                           rca_out_5_8_port, S(7) => rca_out_5_7_port, S(6) => 
                           rca_out_5_6_port, S(5) => rca_out_5_5_port, S(4) => 
                           rca_out_5_4_port, S(3) => rca_out_5_3_port, S(2) => 
                           rca_out_5_2_port, S(1) => rca_out_5_1_port, S(0) => 
                           rca_out_5_0_port, Co => n_1163);
   rca_i_6 : rca_bhv_numBit32_1 port map( A(31) => rca_out_5_31_port, A(30) => 
                           rca_out_5_30_port, A(29) => rca_out_5_29_port, A(28)
                           => rca_out_5_28_port, A(27) => rca_out_5_27_port, 
                           A(26) => rca_out_5_26_port, A(25) => 
                           rca_out_5_25_port, A(24) => rca_out_5_24_port, A(23)
                           => rca_out_5_23_port, A(22) => rca_out_5_22_port, 
                           A(21) => rca_out_5_21_port, A(20) => 
                           rca_out_5_20_port, A(19) => rca_out_5_19_port, A(18)
                           => rca_out_5_18_port, A(17) => rca_out_5_17_port, 
                           A(16) => rca_out_5_16_port, A(15) => 
                           rca_out_5_15_port, A(14) => rca_out_5_14_port, A(13)
                           => rca_out_5_13_port, A(12) => rca_out_5_12_port, 
                           A(11) => rca_out_5_11_port, A(10) => 
                           rca_out_5_10_port, A(9) => rca_out_5_9_port, A(8) =>
                           rca_out_5_8_port, A(7) => rca_out_5_7_port, A(6) => 
                           rca_out_5_6_port, A(5) => rca_out_5_5_port, A(4) => 
                           rca_out_5_4_port, A(3) => rca_out_5_3_port, A(2) => 
                           rca_out_5_2_port, A(1) => rca_out_5_1_port, A(0) => 
                           rca_out_5_0_port, B(31) => sum_op_7_31_port, B(30) 
                           => sum_op_7_30_port, B(29) => sum_op_7_29_port, 
                           B(28) => sum_op_7_28_port, B(27) => sum_op_7_27_port
                           , B(26) => sum_op_7_26_port, B(25) => 
                           sum_op_7_25_port, B(24) => sum_op_7_24_port, B(23) 
                           => sum_op_7_23_port, B(22) => sum_op_7_22_port, 
                           B(21) => sum_op_7_21_port, B(20) => sum_op_7_20_port
                           , B(19) => sum_op_7_19_port, B(18) => 
                           sum_op_7_18_port, B(17) => sum_op_7_17_port, B(16) 
                           => sum_op_7_16_port, B(15) => sum_op_7_15_port, 
                           B(14) => sum_op_7_14_port, B(13) => sum_op_7_13_port
                           , B(12) => sum_op_7_12_port, B(11) => 
                           sum_op_7_11_port, B(10) => sum_op_7_10_port, B(9) =>
                           sum_op_7_9_port, B(8) => sum_op_7_8_port, B(7) => 
                           sum_op_7_7_port, B(6) => sum_op_7_6_port, B(5) => 
                           sum_op_7_5_port, B(4) => sum_op_7_4_port, B(3) => 
                           sum_op_7_3_port, B(2) => sum_op_7_2_port, B(1) => 
                           sum_op_7_1_port, B(0) => sum_op_7_0_port, Ci => 
                           X_Logic0_port, S(31) => P(31), S(30) => P(30), S(29)
                           => P(29), S(28) => P(28), S(27) => P(27), S(26) => 
                           P(26), S(25) => P(25), S(24) => P(24), S(23) => 
                           P(23), S(22) => P(22), S(21) => P(21), S(20) => 
                           P(20), S(19) => P(19), S(18) => P(18), S(17) => 
                           P(17), S(16) => P(16), S(15) => P(15), S(14) => 
                           P(14), S(13) => P(13), S(12) => P(12), S(11) => 
                           P(11), S(10) => P(10), S(9) => P(9), S(8) => P(8), 
                           S(7) => P(7), S(6) => P(6), S(5) => P(5), S(4) => 
                           P(4), S(3) => P(3), S(2) => P(2), S(1) => P(1), S(0)
                           => P(0), Co => n_1164);
   add_65_U1_1_1 : HA_X1 port map( A => add_65_A_1_port, B => add_65_A_0_port, 
                           CO => add_65_carry_2_port, S => A_minus_1_port);
   add_65_U1_1_2 : HA_X1 port map( A => add_65_A_2_port, B => 
                           add_65_carry_2_port, CO => add_65_carry_3_port, S =>
                           A_minus_2_port);
   add_65_U1_1_3 : HA_X1 port map( A => add_65_A_3_port, B => 
                           add_65_carry_3_port, CO => add_65_carry_4_port, S =>
                           A_minus_3_port);
   add_65_U1_1_4 : HA_X1 port map( A => add_65_A_4_port, B => 
                           add_65_carry_4_port, CO => add_65_carry_5_port, S =>
                           A_minus_4_port);
   add_65_U1_1_5 : HA_X1 port map( A => add_65_A_5_port, B => 
                           add_65_carry_5_port, CO => add_65_carry_6_port, S =>
                           A_minus_5_port);
   add_65_U1_1_6 : HA_X1 port map( A => add_65_A_6_port, B => 
                           add_65_carry_6_port, CO => add_65_carry_7_port, S =>
                           A_minus_6_port);
   add_65_U1_1_7 : HA_X1 port map( A => add_65_A_7_port, B => 
                           add_65_carry_7_port, CO => add_65_carry_8_port, S =>
                           A_minus_7_port);
   add_65_U1_1_8 : HA_X1 port map( A => add_65_A_8_port, B => 
                           add_65_carry_8_port, CO => add_65_carry_9_port, S =>
                           A_minus_8_port);
   add_65_U1_1_9 : HA_X1 port map( A => add_65_A_9_port, B => 
                           add_65_carry_9_port, CO => add_65_carry_10_port, S 
                           => A_minus_9_port);
   add_65_U1_1_10 : HA_X1 port map( A => add_65_A_10_port, B => 
                           add_65_carry_10_port, CO => add_65_carry_11_port, S 
                           => A_minus_10_port);
   add_65_U1_1_11 : HA_X1 port map( A => add_65_A_11_port, B => 
                           add_65_carry_11_port, CO => add_65_carry_12_port, S 
                           => A_minus_11_port);
   add_65_U1_1_12 : HA_X1 port map( A => add_65_A_12_port, B => 
                           add_65_carry_12_port, CO => add_65_carry_13_port, S 
                           => A_minus_12_port);
   add_65_U1_1_13 : HA_X1 port map( A => add_65_A_13_port, B => 
                           add_65_carry_13_port, CO => add_65_carry_14_port, S 
                           => A_minus_13_port);
   add_65_U1_1_14 : HA_X1 port map( A => add_65_A_14_port, B => 
                           add_65_carry_14_port, CO => add_65_carry_15_port, S 
                           => A_minus_14_port);
   U3 : INV_X1 port map( A => A_minus_14_port, ZN => n1);
   U4 : INV_X1 port map( A => n1, ZN => n2);
   U5 : INV_X1 port map( A => A_minus_13_port, ZN => n3);
   U6 : INV_X1 port map( A => n3, ZN => n4);
   U7 : INV_X1 port map( A => A_minus_12_port, ZN => n5);
   U8 : INV_X1 port map( A => n5, ZN => n6);
   U9 : INV_X1 port map( A => A_minus_11_port, ZN => n7);
   U10 : INV_X1 port map( A => n7, ZN => n8);
   U11 : INV_X1 port map( A => A_minus_10_port, ZN => n9);
   U12 : INV_X1 port map( A => n9, ZN => n10);
   U13 : INV_X1 port map( A => A_minus_9_port, ZN => n11);
   U14 : INV_X1 port map( A => n11, ZN => n12);
   U15 : INV_X1 port map( A => A_minus_8_port, ZN => n13);
   U16 : INV_X1 port map( A => n13, ZN => n14);
   U17 : INV_X1 port map( A => A_minus_7_port, ZN => n15);
   U18 : INV_X1 port map( A => n15, ZN => n16);
   U19 : INV_X1 port map( A => A_minus_6_port, ZN => n17);
   U20 : INV_X1 port map( A => n17, ZN => n18);
   U21 : INV_X1 port map( A => A_minus_5_port, ZN => n19);
   U22 : INV_X1 port map( A => n19, ZN => n20);
   U23 : INV_X1 port map( A => A_minus_4_port, ZN => n21);
   U24 : INV_X1 port map( A => n21, ZN => n22);
   U25 : INV_X1 port map( A => A_minus_3_port, ZN => n23);
   U26 : INV_X1 port map( A => n23, ZN => n24);
   U27 : INV_X1 port map( A => A_minus_2_port, ZN => n25);
   U28 : INV_X1 port map( A => n25, ZN => n26);
   U29 : INV_X1 port map( A => A_minus_1_port, ZN => n27);
   U30 : INV_X1 port map( A => n27, ZN => n28);
   U31 : BUF_X1 port map( A => n30, Z => n40);
   U32 : BUF_X1 port map( A => n30, Z => n39);
   U33 : BUF_X1 port map( A => n30, Z => n37);
   U34 : BUF_X1 port map( A => n30, Z => n38);
   U35 : BUF_X1 port map( A => n29, Z => n36);
   U36 : BUF_X1 port map( A => n29, Z => n31);
   U37 : BUF_X1 port map( A => n29, Z => n33);
   U38 : BUF_X1 port map( A => n29, Z => n35);
   U39 : BUF_X1 port map( A => n29, Z => n32);
   U40 : BUF_X1 port map( A => n29, Z => n34);
   U41 : BUF_X1 port map( A => n30, Z => n41);
   U42 : BUF_X1 port map( A => A_minus_31_port, Z => n29);
   U43 : BUF_X1 port map( A => A_minus_31_port, Z => n30);
   U44 : INV_X1 port map( A => n54, ZN => n42);
   U45 : INV_X1 port map( A => n54, ZN => n43);
   U46 : INV_X1 port map( A => n54, ZN => n47);
   U47 : INV_X1 port map( A => n54, ZN => n46);
   U48 : INV_X1 port map( A => n54, ZN => n44);
   U49 : INV_X1 port map( A => n54, ZN => n45);
   U50 : INV_X1 port map( A => n54, ZN => n48);
   U51 : INV_X1 port map( A => n54, ZN => n53);
   U52 : INV_X1 port map( A => n54, ZN => n52);
   U53 : INV_X1 port map( A => n54, ZN => n51);
   U54 : INV_X1 port map( A => n54, ZN => n50);
   U55 : INV_X1 port map( A => n54, ZN => n49);
   U56 : INV_X1 port map( A => add_65_A_0_port, ZN => A_minus_0_port);
   U57 : INV_X1 port map( A => A(0), ZN => add_65_A_0_port);
   U58 : INV_X1 port map( A => A(14), ZN => add_65_A_14_port);
   U59 : INV_X1 port map( A => A(1), ZN => add_65_A_1_port);
   U60 : INV_X1 port map( A => A(2), ZN => add_65_A_2_port);
   U61 : INV_X1 port map( A => A(3), ZN => add_65_A_3_port);
   U62 : INV_X1 port map( A => A(4), ZN => add_65_A_4_port);
   U63 : INV_X1 port map( A => A(5), ZN => add_65_A_5_port);
   U64 : INV_X1 port map( A => A(6), ZN => add_65_A_6_port);
   U65 : INV_X1 port map( A => A(7), ZN => add_65_A_7_port);
   U66 : INV_X1 port map( A => A(8), ZN => add_65_A_8_port);
   U67 : INV_X1 port map( A => A(9), ZN => add_65_A_9_port);
   U68 : INV_X1 port map( A => A(10), ZN => add_65_A_10_port);
   U69 : INV_X1 port map( A => A(11), ZN => add_65_A_11_port);
   U70 : INV_X1 port map( A => A(12), ZN => add_65_A_12_port);
   U71 : INV_X1 port map( A => A(13), ZN => add_65_A_13_port);
   U72 : XOR2_X2 port map( A => add_65_carry_15_port, B => n54, Z => 
                           A_minus_15_port);
   U73 : INV_X1 port map( A => A(15), ZN => n54);
   U74 : NOR2_X1 port map( A1 => add_65_carry_15_port, A2 => A(15), ZN => 
                           A_minus_31_port);
   encoder_out_0_port <= '0';

end SYN_mixed;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity P4Adder_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (31 downto 0);  Cout : out std_logic);

end P4Adder_NBIT32;

architecture SYN_struct of P4Adder_NBIT32 is

   component SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component carry_generator_NBIT32_NBIT_PER_BLOCK4
      port( A, B : in std_logic_vector (32 downto 1);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal Csum_7_port, Csum_6_port, Csum_5_port, Csum_4_port, Csum_3_port, 
      Csum_2_port, Csum_1_port : std_logic;

begin
   
   Carrygen0 : carry_generator_NBIT32_NBIT_PER_BLOCK4 port map( A(32) => A(31),
                           A(31) => A(30), A(30) => A(29), A(29) => A(28), 
                           A(28) => A(27), A(27) => A(26), A(26) => A(25), 
                           A(25) => A(24), A(24) => A(23), A(23) => A(22), 
                           A(22) => A(21), A(21) => A(20), A(20) => A(19), 
                           A(19) => A(18), A(18) => A(17), A(17) => A(16), 
                           A(16) => A(15), A(15) => A(14), A(14) => A(13), 
                           A(13) => A(12), A(12) => A(11), A(11) => A(10), 
                           A(10) => A(9), A(9) => A(8), A(8) => A(7), A(7) => 
                           A(6), A(6) => A(5), A(5) => A(4), A(4) => A(3), A(3)
                           => A(2), A(2) => A(1), A(1) => A(0), B(32) => B(31),
                           B(31) => B(30), B(30) => B(29), B(29) => B(28), 
                           B(28) => B(27), B(27) => B(26), B(26) => B(25), 
                           B(25) => B(24), B(24) => B(23), B(23) => B(22), 
                           B(22) => B(21), B(21) => B(20), B(20) => B(19), 
                           B(19) => B(18), B(18) => B(17), B(17) => B(16), 
                           B(16) => B(15), B(15) => B(14), B(14) => B(13), 
                           B(13) => B(12), B(12) => B(11), B(11) => B(10), 
                           B(10) => B(9), B(9) => B(8), B(8) => B(7), B(7) => 
                           B(6), B(6) => B(5), B(5) => B(4), B(4) => B(3), B(3)
                           => B(2), B(2) => B(1), B(1) => B(0), Cin => Cin, 
                           Co(7) => Cout, Co(6) => Csum_7_port, Co(5) => 
                           Csum_6_port, Co(4) => Csum_5_port, Co(3) => 
                           Csum_4_port, Co(2) => Csum_3_port, Co(1) => 
                           Csum_2_port, Co(0) => Csum_1_port);
   Sumgen0 : SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), Ci(7) => 
                           Csum_7_port, Ci(6) => Csum_6_port, Ci(5) => 
                           Csum_5_port, Ci(4) => Csum_4_port, Ci(3) => 
                           Csum_3_port, Ci(2) => Csum_2_port, Ci(1) => 
                           Csum_1_port, Ci(0) => Cin, S(31) => S(31), S(30) => 
                           S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           S(21), S(20) => S(20), S(19) => S(19), S(18) => 
                           S(18), S(17) => S(17), S(16) => S(16), S(15) => 
                           S(15), S(14) => S(14), S(13) => S(13), S(12) => 
                           S(12), S(11) => S(11), S(10) => S(10), S(9) => S(9),
                           S(8) => S(8), S(7) => S(7), S(6) => S(6), S(5) => 
                           S(5), S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1)
                           => S(1), S(0) => S(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity shifter_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  LOGIC_ARITH, LEFT_RIGHT : 
         in std_logic;  RES : out std_logic_vector (31 downto 0));

end shifter_NBIT32;

architecture SYN_bhv of shifter_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X4
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X2
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, 
      n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
      n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, 
      n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, 
      n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n1, n2, n3, n4, n5, n6, 
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n266, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649 : std_logic;

begin
   
   U264 : AOI21_X2 port map( B1 => A(31), B2 => B(18), A => n483, ZN => n282);
   U267 : OAI21_X2 port map( B1 => n613, B2 => n629, A => n486, ZN => n285);
   U269 : AOI21_X2 port map( B1 => A(31), B2 => n39, A => n487, ZN => n288);
   U388 : AOI221_X2 port map( B1 => n31, B2 => A(18), C1 => n21, C2 => A(17), A
                           => n568, ZN => n196);
   U428 : NOR2_X2 port map( A1 => n639, A2 => n39, ZN => n165);
   U461 : NOR2_X2 port map( A1 => n643, A2 => n39, ZN => n199);
   U637 : NAND3_X1 port map( A1 => n227, A2 => n647, A3 => n228, ZN => n226);
   U638 : NAND3_X1 port map( A1 => n227, A2 => n647, A3 => B(4), ZN => n428);
   U639 : NAND3_X1 port map( A1 => n445, A2 => n199, A3 => LEFT_RIGHT, ZN => 
                           n240);
   U641 : NAND3_X1 port map( A1 => n489, A2 => n629, A3 => n579, ZN => n255);
   U642 : NAND3_X1 port map( A1 => n267, A2 => n199, A3 => n445, ZN => n138);
   U2 : NOR4_X1 port map( A1 => B(20), A2 => B(21), A3 => B(19), A4 => n594, ZN
                           => n484);
   U3 : NOR2_X2 port map( A1 => n640, A2 => B(3), ZN => n262);
   U4 : NOR2_X2 port map( A1 => n490, A2 => B(11), ZN => n283);
   U5 : NAND3_X1 port map( A1 => n445, A2 => n35, A3 => LEFT_RIGHT, ZN => n269)
                           ;
   U6 : INV_X1 port map( A => n167, ZN => n636);
   U7 : NOR2_X1 port map( A1 => n637, A2 => B(4), ZN => n167);
   U8 : INV_X1 port map( A => n169, ZN => n645);
   U9 : INV_X1 port map( A => n165, ZN => n638);
   U10 : INV_X1 port map( A => n199, ZN => n642);
   U11 : INV_X1 port map( A => n32, ZN => n28);
   U12 : INV_X1 port map( A => n32, ZN => n26);
   U13 : INV_X1 port map( A => n32, ZN => n27);
   U14 : INV_X1 port map( A => n22, ZN => n14);
   U15 : INV_X1 port map( A => n22, ZN => n15);
   U16 : INV_X1 port map( A => n21, ZN => n16);
   U17 : INV_X1 port map( A => n505, ZN => n644);
   U18 : INV_X1 port map( A => n31, ZN => n29);
   U19 : INV_X1 port map( A => n493, ZN => n641);
   U20 : NOR2_X1 port map( A1 => n646, A2 => n39, ZN => n169);
   U21 : NAND2_X1 port map( A1 => n488, A2 => n454, ZN => n161);
   U22 : INV_X1 port map( A => n42, ZN => n39);
   U23 : OAI222_X1 port map( A1 => n79, A2 => n645, B1 => n63, B2 => n636, C1 
                           => n91, C2 => n638, ZN => n371);
   U24 : OAI222_X1 port map( A1 => n82, A2 => n645, B1 => n62, B2 => n636, C1 
                           => n95, C2 => n638, ZN => n360);
   U25 : OAI222_X1 port map( A1 => n85, A2 => n645, B1 => n73, B2 => n636, C1 
                           => n99, C2 => n638, ZN => n349);
   U26 : OAI222_X1 port map( A1 => n87, A2 => n645, B1 => n76, B2 => n636, C1 
                           => n104, C2 => n638, ZN => n338);
   U27 : NOR2_X1 port map( A1 => n41, A2 => n643, ZN => n493);
   U28 : OAI22_X1 port map( A1 => n116, A2 => n643, B1 => n127, B2 => n639, ZN 
                           => n383);
   U29 : INV_X1 port map( A => n454, ZN => n637);
   U30 : AOI21_X1 port map( B1 => n135, B2 => n2, A => n519, ZN => n286);
   U31 : AOI21_X1 port map( B1 => n130, B2 => n3, A => n519, ZN => n312);
   U32 : BUF_X1 port map( A => n138, Z => n34);
   U33 : BUF_X1 port map( A => n138, Z => n33);
   U34 : NOR2_X1 port map( A1 => n383, A2 => n359, ZN => n197);
   U35 : NOR2_X1 port map( A1 => n119, A2 => n359, ZN => n181);
   U36 : BUF_X1 port map( A => n138, Z => n35);
   U37 : NAND2_X1 port map( A1 => n488, A2 => n5, ZN => n505);
   U38 : INV_X1 port map( A => n182, ZN => n119);
   U39 : INV_X1 port map( A => n238, ZN => n107);
   U40 : INV_X1 port map( A => n214, ZN => n56);
   U41 : INV_X1 port map( A => n202, ZN => n50);
   U42 : INV_X1 port map( A => n188, ZN => n48);
   U43 : NOR2_X1 port map( A1 => n613, A2 => n148, ZN => n150);
   U44 : OAI21_X2 port map( B1 => n612, B2 => n633, A => n481, ZN => n279);
   U45 : NOR2_X1 port map( A1 => n640, A2 => n647, ZN => n454);
   U46 : NAND2_X1 port map( A1 => n484, A2 => n631, ZN => n281);
   U47 : AOI222_X1 port map( A1 => n370, A2 => n262, B1 => n320, B2 => n260, C1
                           => n185, C2 => n3, ZN => n238);
   U48 : INV_X1 port map( A => n356, ZN => n643);
   U49 : AOI222_X1 port map( A1 => n168, A2 => n262, B1 => n355, B2 => n260, C1
                           => n170, C2 => n3, ZN => n471);
   U50 : AOI222_X1 port map( A1 => n402, A2 => n262, B1 => n403, B2 => n260, C1
                           => n464, C2 => n2, ZN => n461);
   U51 : NAND2_X1 port map( A1 => n488, A2 => n262, ZN => n157);
   U52 : NAND2_X1 port map( A1 => n488, A2 => n260, ZN => n158);
   U53 : OAI222_X1 port map( A1 => n374, A2 => n639, B1 => n646, B2 => n375, C1
                           => n376, C2 => n643, ZN => n172);
   U54 : OAI222_X1 port map( A1 => n132, A2 => n639, B1 => n362, B2 => n646, C1
                           => n363, C2 => n643, ZN => n139);
   U55 : OAI222_X1 port map( A1 => n614, A2 => n639, B1 => n293, B2 => n646, C1
                           => n405, C2 => n643, ZN => n348);
   U56 : OAI222_X1 port map( A1 => n616, A2 => n639, B1 => n46, B2 => n646, C1 
                           => n387, C2 => n643, ZN => n337);
   U57 : AOI221_X1 port map( B1 => n130, B2 => n262, C1 => n355, C2 => n2, A =>
                           n359, ZN => n159);
   U58 : AOI221_X1 port map( B1 => n135, B2 => n262, C1 => n403, C2 => n3, A =>
                           n359, ZN => n347);
   U59 : OAI221_X1 port map( B1 => n106, B2 => n639, C1 => n90, C2 => n643, A 
                           => n607, ZN => n480);
   U60 : AOI22_X1 port map( A1 => n454, A2 => n320, B1 => n260, B2 => n370, ZN 
                           => n607);
   U61 : AOI222_X1 port map( A1 => n169, A2 => n185, B1 => n493, B2 => n320, C1
                           => n167, C2 => n370, ZN => n550);
   U62 : OAI222_X1 port map( A1 => n62, A2 => n645, B1 => n363, B2 => n636, C1 
                           => n82, C2 => n638, ZN => n418);
   U63 : OAI222_X1 port map( A1 => n73, A2 => n645, B1 => n405, B2 => n636, C1 
                           => n85, C2 => n638, ZN => n404);
   U64 : OAI222_X1 port map( A1 => n76, A2 => n645, B1 => n387, B2 => n636, C1 
                           => n87, C2 => n638, ZN => n386);
   U65 : INV_X1 port map( A => n260, ZN => n646);
   U66 : NOR2_X1 port map( A1 => n648, A2 => B(4), ZN => n488);
   U67 : INV_X1 port map( A => n262, ZN => n639);
   U68 : INV_X1 port map( A => n332, ZN => n628);
   U69 : OAI222_X1 port map( A1 => n133, A2 => n14, B1 => n29, B2 => n615, C1 
                           => n1, C2 => n103, ZN => n602);
   U70 : OAI221_X1 port map( B1 => n363, B2 => n639, C1 => n62, C2 => n643, A 
                           => n522, ZN => n314);
   U71 : AOI22_X1 port map( A1 => n454, A2 => n58, B1 => n260, B2 => n420, ZN 
                           => n522);
   U72 : OAI221_X1 port map( B1 => n405, B2 => n639, C1 => n73, C2 => n643, A 
                           => n509, ZN => n290);
   U73 : AOI22_X1 port map( A1 => n454, A2 => n52, B1 => n260, B2 => n407, ZN 
                           => n509);
   U74 : OAI221_X1 port map( B1 => n387, B2 => n639, C1 => n76, C2 => n643, A 
                           => n496, ZN => n271);
   U75 : AOI22_X1 port map( A1 => n454, A2 => n390, B1 => n260, B2 => n389, ZN 
                           => n496);
   U76 : OAI21_X1 port map( B1 => n613, B2 => n631, A => n486, ZN => n253);
   U77 : NOR2_X1 port map( A1 => n613, A2 => n647, ZN => n359);
   U78 : NOR2_X1 port map( A1 => n613, A2 => n2, ZN => n519);
   U79 : AOI221_X1 port map( B1 => n219, B2 => n199, C1 => n223, C2 => n39, A 
                           => n224, ZN => n222);
   U80 : OAI222_X1 port map( A1 => n638, A2 => n71, B1 => n636, B2 => n93, C1 
                           => n645, C2 => n81, ZN => n224);
   U81 : AOI221_X1 port map( B1 => n207, B2 => n199, C1 => n211, C2 => n39, A 
                           => n212, ZN => n210);
   U82 : OAI222_X1 port map( A1 => n638, A2 => n68, B1 => n636, B2 => n97, C1 
                           => n645, C2 => n84, ZN => n212);
   U83 : AOI221_X1 port map( B1 => n193, B2 => n199, C1 => n115, C2 => n39, A 
                           => n200, ZN => n198);
   U84 : OAI222_X1 port map( A1 => n638, A2 => n75, B1 => n636, B2 => n101, C1 
                           => n645, C2 => n196, ZN => n200);
   U85 : OAI22_X1 port map( A1 => n8, A2 => n131, B1 => n1, B2 => n266, ZN => 
                           n533);
   U86 : OAI221_X1 port map( B1 => n618, B2 => n642, C1 => n238, C2 => n41, A 
                           => n239, ZN => n229);
   U87 : AOI222_X1 port map( A1 => n165, A2 => n178, B1 => n167, B2 => n186, C1
                           => n169, C2 => n184, ZN => n239);
   U88 : OAI221_X1 port map( B1 => n65, B2 => n642, C1 => n182, C2 => n41, A =>
                           n183, ZN => n173);
   U89 : AOI222_X1 port map( A1 => n165, A2 => n184, B1 => n167, B2 => n185, C1
                           => n169, C2 => n186, ZN => n183);
   U90 : OAI221_X1 port map( B1 => n71, B2 => n642, C1 => n163, C2 => n42, A =>
                           n164, ZN => n141);
   U91 : AOI222_X1 port map( A1 => n165, A2 => n166, B1 => n167, B2 => n168, C1
                           => n169, C2 => n170, ZN => n164);
   U92 : OAI221_X1 port map( B1 => n68, B2 => n642, C1 => n344, C2 => n42, A =>
                           n581, ZN => n572);
   U93 : AOI222_X1 port map( A1 => n165, A2 => n516, B1 => n167, B2 => n402, C1
                           => n169, C2 => n464, ZN => n581);
   U94 : OAI221_X1 port map( B1 => n93, B2 => n638, C1 => n81, C2 => n642, A =>
                           n534, ZN => n526);
   U95 : AOI222_X1 port map( A1 => n169, A2 => n168, B1 => n493, B2 => n129, C1
                           => n167, C2 => n355, ZN => n534);
   U96 : OAI221_X1 port map( B1 => n97, B2 => n638, C1 => n84, C2 => n642, A =>
                           n520, ZN => n511);
   U97 : AOI222_X1 port map( A1 => n169, A2 => n402, B1 => n493, B2 => n134, C1
                           => n167, C2 => n403, ZN => n520);
   U98 : OAI221_X1 port map( B1 => n101, B2 => n638, C1 => n196, C2 => n642, A 
                           => n507, ZN => n498);
   U99 : AOI222_X1 port map( A1 => n169, A2 => n453, B1 => n493, B2 => n382, C1
                           => n167, C2 => n506, ZN => n507);
   U100 : NOR2_X1 port map( A1 => n613, A2 => n8, ZN => n382);
   U101 : OAI221_X1 port map( B1 => n127, B2 => n161, C1 => n116, C2 => n158, A
                           => n162, ZN => n503);
   U102 : OAI221_X1 port map( B1 => n237, B2 => n160, C1 => n90, C2 => n161, A 
                           => n162, ZN => n235);
   U103 : OAI221_X1 port map( B1 => n110, B2 => n160, C1 => n93, C2 => n161, A 
                           => n162, ZN => n220);
   U104 : OAI221_X1 port map( B1 => n113, B2 => n160, C1 => n97, C2 => n161, A 
                           => n162, ZN => n208);
   U105 : OAI221_X1 port map( B1 => n197, B2 => n160, C1 => n101, C2 => n161, A
                           => n162, ZN => n194);
   U106 : OAI221_X1 port map( B1 => n181, B2 => n160, C1 => n106, C2 => n161, A
                           => n162, ZN => n179);
   U107 : OAI221_X1 port map( B1 => n159, B2 => n160, C1 => n109, C2 => n161, A
                           => n162, ZN => n155);
   U108 : OAI221_X1 port map( B1 => n347, B2 => n160, C1 => n112, C2 => n161, A
                           => n162, ZN => n577);
   U109 : OAI221_X1 port map( B1 => n336, B2 => n160, C1 => n116, C2 => n161, A
                           => n162, ZN => n560);
   U110 : OAI221_X1 port map( B1 => n323, B2 => n160, C1 => n118, C2 => n161, A
                           => n162, ZN => n548);
   U111 : INV_X1 port map( A => n370, ZN => n118);
   U112 : OAI221_X1 port map( B1 => n312, B2 => n160, C1 => n121, C2 => n161, A
                           => n162, ZN => n531);
   U113 : INV_X1 port map( A => n355, ZN => n121);
   U114 : OAI221_X1 port map( B1 => n286, B2 => n160, C1 => n124, C2 => n161, A
                           => n162, ZN => n517);
   U115 : INV_X1 port map( A => n403, ZN => n124);
   U116 : AND2_X1 port map( A1 => n491, A2 => n633, ZN => n276);
   U117 : AOI22_X1 port map( A1 => n480, A2 => n39, B1 => n43, B2 => n64, ZN =>
                           n587);
   U118 : INV_X1 port map( A => n601, ZN => n64);
   U119 : AOI221_X1 port map( B1 => n4, B2 => n602, C1 => n454, C2 => n184, A 
                           => n603, ZN => n601);
   U120 : OAI22_X1 port map( A1 => n618, A2 => n639, B1 => n65, B2 => n646, ZN 
                           => n603);
   U121 : AOI22_X1 port map( A1 => n420, A2 => n2, B1 => n58, B2 => n262, ZN =>
                           n214);
   U122 : AOI22_X1 port map( A1 => n407, A2 => n5, B1 => n52, B2 => n262, ZN =>
                           n202);
   U123 : AOI22_X1 port map( A1 => n389, A2 => n3, B1 => n390, B2 => n262, ZN 
                           => n188);
   U124 : AOI22_X1 port map( A1 => n168, A2 => n3, B1 => n355, B2 => n262, ZN 
                           => n413);
   U125 : AOI22_X1 port map( A1 => n402, A2 => n5, B1 => n403, B2 => n262, ZN 
                           => n396);
   U126 : AOI22_X1 port map( A1 => n452, A2 => n4, B1 => n453, B2 => n262, ZN 
                           => n449);
   U127 : AOI22_X1 port map( A1 => n370, A2 => n4, B1 => n320, B2 => n262, ZN 
                           => n182);
   U128 : AOI22_X1 port map( A1 => n355, A2 => n2, B1 => n129, B2 => n262, ZN 
                           => n163);
   U129 : AOI22_X1 port map( A1 => n403, A2 => n4, B1 => n134, B2 => n262, ZN 
                           => n344);
   U130 : AOI21_X1 port map( B1 => n148, B2 => n232, A => n150, ZN => n231);
   U131 : OAI21_X1 port map( B1 => n233, B2 => n152, A => n153, ZN => n232);
   U132 : AOI211_X1 port map( C1 => n644, C2 => n234, A => n235, B => n236, ZN 
                           => n233);
   U133 : OAI22_X1 port map( A1 => n65, A2 => n157, B1 => n78, B2 => n158, ZN 
                           => n236);
   U134 : AOI21_X1 port map( B1 => n148, B2 => n217, A => n150, ZN => n216);
   U135 : OAI21_X1 port map( B1 => n218, B2 => n152, A => n153, ZN => n217);
   U136 : AOI211_X1 port map( C1 => n644, C2 => n219, A => n220, B => n221, ZN 
                           => n218);
   U137 : OAI22_X1 port map( A1 => n71, A2 => n157, B1 => n81, B2 => n158, ZN 
                           => n221);
   U138 : AOI21_X1 port map( B1 => n148, B2 => n205, A => n150, ZN => n204);
   U139 : OAI21_X1 port map( B1 => n206, B2 => n152, A => n153, ZN => n205);
   U140 : AOI211_X1 port map( C1 => n644, C2 => n207, A => n208, B => n209, ZN 
                           => n206);
   U141 : OAI22_X1 port map( A1 => n68, A2 => n157, B1 => n84, B2 => n158, ZN 
                           => n209);
   U142 : AOI21_X1 port map( B1 => n148, B2 => n191, A => n150, ZN => n190);
   U143 : OAI21_X1 port map( B1 => n192, B2 => n152, A => n153, ZN => n191);
   U144 : AOI211_X1 port map( C1 => n644, C2 => n193, A => n194, B => n195, ZN 
                           => n192);
   U145 : OAI22_X1 port map( A1 => n75, A2 => n157, B1 => n196, B2 => n158, ZN 
                           => n195);
   U146 : AOI21_X1 port map( B1 => n148, B2 => n176, A => n150, ZN => n175);
   U147 : OAI21_X1 port map( B1 => n177, B2 => n152, A => n153, ZN => n176);
   U148 : AOI211_X1 port map( C1 => n644, C2 => n178, A => n179, B => n180, ZN 
                           => n177);
   U149 : OAI22_X1 port map( A1 => n78, A2 => n157, B1 => n90, B2 => n158, ZN 
                           => n180);
   U150 : AOI21_X1 port map( B1 => n148, B2 => n149, A => n150, ZN => n145);
   U151 : OAI21_X1 port map( B1 => n151, B2 => n152, A => n153, ZN => n149);
   U152 : AOI211_X1 port map( C1 => n644, C2 => n154, A => n155, B => n156, ZN 
                           => n151);
   U153 : OAI22_X1 port map( A1 => n81, A2 => n157, B1 => n93, B2 => n158, ZN 
                           => n156);
   U154 : AOI21_X1 port map( B1 => n148, B2 => n575, A => n150, ZN => n574);
   U155 : OAI21_X1 port map( B1 => n576, B2 => n152, A => n153, ZN => n575);
   U156 : AOI211_X1 port map( C1 => n644, C2 => n305, A => n577, B => n578, ZN 
                           => n576);
   U157 : OAI22_X1 port map( A1 => n84, A2 => n157, B1 => n97, B2 => n158, ZN 
                           => n578);
   U158 : AOI21_X1 port map( B1 => n148, B2 => n558, A => n150, ZN => n557);
   U159 : OAI21_X1 port map( B1 => n559, B2 => n152, A => n153, ZN => n558);
   U160 : AOI211_X1 port map( C1 => n644, C2 => n261, A => n560, B => n561, ZN 
                           => n559);
   U161 : OAI22_X1 port map( A1 => n196, A2 => n157, B1 => n101, B2 => n158, ZN
                           => n561);
   U162 : AOI21_X1 port map( B1 => n148, B2 => n546, A => n150, ZN => n545);
   U163 : OAI21_X1 port map( B1 => n547, B2 => n152, A => n153, ZN => n546);
   U164 : AOI211_X1 port map( C1 => n644, C2 => n184, A => n548, B => n549, ZN 
                           => n547);
   U165 : OAI22_X1 port map( A1 => n90, A2 => n157, B1 => n106, B2 => n158, ZN 
                           => n549);
   U166 : AOI21_X1 port map( B1 => n148, B2 => n529, A => n150, ZN => n528);
   U167 : OAI21_X1 port map( B1 => n530, B2 => n152, A => n153, ZN => n529);
   U168 : AOI211_X1 port map( C1 => n644, C2 => n166, A => n531, B => n532, ZN 
                           => n530);
   U169 : OAI22_X1 port map( A1 => n93, A2 => n157, B1 => n109, B2 => n158, ZN 
                           => n532);
   U170 : AOI21_X1 port map( B1 => n148, B2 => n514, A => n150, ZN => n513);
   U171 : OAI21_X1 port map( B1 => n515, B2 => n152, A => n153, ZN => n514);
   U172 : AOI211_X1 port map( C1 => n644, C2 => n516, A => n517, B => n518, ZN 
                           => n515);
   U173 : OAI22_X1 port map( A1 => n97, A2 => n157, B1 => n112, B2 => n158, ZN 
                           => n518);
   U174 : AOI21_X1 port map( B1 => n283, B2 => n415, A => n285, ZN => n414);
   U175 : OAI21_X1 port map( B1 => n110, B2 => n287, A => n288, ZN => n415);
   U176 : AOI21_X1 port map( B1 => n283, B2 => n398, A => n285, ZN => n397);
   U177 : OAI21_X1 port map( B1 => n113, B2 => n287, A => n288, ZN => n398);
   U178 : AOI21_X1 port map( B1 => n283, B2 => n385, A => n285, ZN => n384);
   U179 : OAI21_X1 port map( B1 => n197, B2 => n287, A => n288, ZN => n385);
   U180 : AOI21_X1 port map( B1 => n283, B2 => n369, A => n285, ZN => n368);
   U181 : OAI21_X1 port map( B1 => n181, B2 => n287, A => n288, ZN => n369);
   U182 : AOI21_X1 port map( B1 => n283, B2 => n335, A => n285, ZN => n334);
   U183 : OAI21_X1 port map( B1 => n336, B2 => n287, A => n288, ZN => n335);
   U184 : OAI211_X1 port map( C1 => n127, C2 => n646, A => n401, B => n449, ZN 
                           => n257);
   U185 : AOI21_X1 port map( B1 => n320, B2 => n4, A => n519, ZN => n323);
   U186 : AOI21_X1 port map( B1 => n506, B2 => n5, A => n519, ZN => n336);
   U187 : NAND2_X1 port map( A1 => n484, A2 => n633, ZN => n249);
   U188 : OAI21_X1 port map( B1 => n417, B2 => n637, A => n471, ZN => n440);
   U189 : OAI21_X1 port map( B1 => n400, B2 => n637, A => n461, ZN => n302);
   U190 : NOR2_X1 port map( A1 => n613, A2 => n484, ZN => n483);
   U191 : OAI21_X1 port map( B1 => n412, B2 => n637, A => n471, ZN => n434);
   U192 : OAI21_X1 port map( B1 => n395, B2 => n637, A => n461, ZN => n297);
   U193 : OAI21_X1 port map( B1 => n412, B2 => n646, A => n413, ZN => n223);
   U194 : OAI21_X1 port map( B1 => n395, B2 => n646, A => n396, ZN => n211);
   U195 : OAI21_X1 port map( B1 => n333, B2 => n647, A => n449, ZN => n246);
   U196 : OAI21_X1 port map( B1 => n482, B2 => n281, A => n282, ZN => n479);
   U197 : AOI21_X1 port map( B1 => n283, B2 => n485, A => n285, ZN => n482);
   U198 : OAI21_X1 port map( B1 => n89, B2 => n287, A => n288, ZN => n485);
   U199 : INV_X1 port map( A => n480, ZN => n89);
   U200 : OAI21_X1 port map( B1 => n472, B2 => n281, A => n282, ZN => n470);
   U201 : AOI21_X1 port map( B1 => n283, B2 => n473, A => n285, ZN => n472);
   U202 : OAI21_X1 port map( B1 => n94, B2 => n287, A => n288, ZN => n473);
   U203 : INV_X1 port map( A => n440, ZN => n94);
   U204 : OAI21_X1 port map( B1 => n462, B2 => n281, A => n282, ZN => n460);
   U205 : AOI21_X1 port map( B1 => n283, B2 => n463, A => n285, ZN => n462);
   U206 : OAI21_X1 port map( B1 => n98, B2 => n287, A => n288, ZN => n463);
   U207 : INV_X1 port map( A => n302, ZN => n98);
   U208 : OAI21_X1 port map( B1 => n450, B2 => n281, A => n282, ZN => n448);
   U209 : AOI21_X1 port map( B1 => n283, B2 => n451, A => n285, ZN => n450);
   U210 : OAI21_X1 port map( B1 => n102, B2 => n287, A => n288, ZN => n451);
   U211 : INV_X1 port map( A => n257, ZN => n102);
   U212 : OAI21_X1 port map( B1 => n425, B2 => n281, A => n282, ZN => n424);
   U213 : AOI21_X1 port map( B1 => n283, B2 => n426, A => n285, ZN => n425);
   U214 : OAI21_X1 port map( B1 => n237, B2 => n287, A => n288, ZN => n426);
   U215 : OAI21_X1 port map( B1 => n357, B2 => n281, A => n282, ZN => n354);
   U216 : AOI21_X1 port map( B1 => n283, B2 => n358, A => n285, ZN => n357);
   U217 : OAI21_X1 port map( B1 => n159, B2 => n287, A => n288, ZN => n358);
   U218 : OAI21_X1 port map( B1 => n345, B2 => n281, A => n282, ZN => n343);
   U219 : AOI21_X1 port map( B1 => n283, B2 => n346, A => n285, ZN => n345);
   U220 : OAI21_X1 port map( B1 => n347, B2 => n287, A => n288, ZN => n346);
   U221 : OAI21_X1 port map( B1 => n321, B2 => n281, A => n282, ZN => n319);
   U222 : AOI21_X1 port map( B1 => n283, B2 => n322, A => n285, ZN => n321);
   U223 : OAI21_X1 port map( B1 => n323, B2 => n287, A => n288, ZN => n322);
   U224 : OAI21_X1 port map( B1 => n310, B2 => n281, A => n282, ZN => n309);
   U225 : AOI21_X1 port map( B1 => n283, B2 => n311, A => n285, ZN => n310);
   U226 : OAI21_X1 port map( B1 => n312, B2 => n287, A => n288, ZN => n311);
   U227 : OAI21_X1 port map( B1 => n280, B2 => n281, A => n282, ZN => n277);
   U228 : AOI21_X1 port map( B1 => n283, B2 => n284, A => n285, ZN => n280);
   U229 : OAI21_X1 port map( B1 => n286, B2 => n287, A => n288, ZN => n284);
   U230 : AOI22_X1 port map( A1 => n246, A2 => n39, B1 => n43, B2 => n247, ZN 
                           => n245);
   U231 : AOI22_X1 port map( A1 => n434, A2 => n39, B1 => n42, B2 => n435, ZN 
                           => n433);
   U232 : AOI22_X1 port map( A1 => n297, A2 => n39, B1 => n42, B2 => n298, ZN 
                           => n296);
   U233 : INV_X1 port map( A => n452, ZN => n101);
   U234 : INV_X1 port map( A => n464, ZN => n97);
   U235 : INV_X1 port map( A => n170, ZN => n93);
   U236 : INV_X1 port map( A => n186, ZN => n90);
   U237 : INV_X1 port map( A => n516, ZN => n84);
   U238 : INV_X1 port map( A => n166, ZN => n81);
   U239 : NOR2_X1 port map( A1 => n266, A2 => n8, ZN => n580);
   U240 : AOI21_X1 port map( B1 => n251, B2 => n438, A => n253, ZN => n437);
   U241 : OAI21_X1 port map( B1 => n439, B2 => n255, A => n256, ZN => n438);
   U242 : AOI22_X1 port map( A1 => n435, A2 => n40, B1 => B(4), B2 => n440, ZN 
                           => n439);
   U243 : AOI21_X1 port map( B1 => n251, B2 => n300, A => n253, ZN => n299);
   U244 : OAI21_X1 port map( B1 => n301, B2 => n255, A => n256, ZN => n300);
   U245 : AOI22_X1 port map( A1 => n298, A2 => n40, B1 => B(4), B2 => n302, ZN 
                           => n301);
   U246 : AOI21_X1 port map( B1 => n251, B2 => n252, A => n253, ZN => n248);
   U247 : OAI21_X1 port map( B1 => n254, B2 => n255, A => n256, ZN => n252);
   U248 : AOI22_X1 port map( A1 => n247, A2 => n40, B1 => B(4), B2 => n257, ZN 
                           => n254);
   U249 : BUF_X1 port map( A => n356, Z => n2);
   U250 : BUF_X1 port map( A => n356, Z => n3);
   U251 : INV_X1 port map( A => n293, ZN => n52);
   U252 : INV_X1 port map( A => n184, ZN => n78);
   U253 : INV_X1 port map( A => n506, ZN => n127);
   U254 : INV_X1 port map( A => n185, ZN => n106);
   U255 : INV_X1 port map( A => n412, ZN => n129);
   U256 : INV_X1 port map( A => n395, ZN => n134);
   U257 : INV_X1 port map( A => n390, ZN => n46);
   U258 : BUF_X1 port map( A => n356, Z => n4);
   U259 : BUF_X1 port map( A => n356, Z => n5);
   U260 : INV_X1 port map( A => n453, ZN => n116);
   U261 : INV_X1 port map( A => n154, ZN => n71);
   U262 : INV_X1 port map( A => n305, ZN => n68);
   U263 : INV_X1 port map( A => n178, ZN => n65);
   U265 : INV_X1 port map( A => n168, ZN => n109);
   U266 : INV_X1 port map( A => n402, ZN => n112);
   U268 : INV_X1 port map( A => n261, ZN => n75);
   U270 : INV_X1 port map( A => n419, ZN => n82);
   U271 : INV_X1 port map( A => n406, ZN => n85);
   U272 : INV_X1 port map( A => n388, ZN => n87);
   U273 : BUF_X1 port map( A => n44, Z => n42);
   U274 : INV_X1 port map( A => n362, ZN => n58);
   U275 : INV_X1 port map( A => n474, ZN => n62);
   U276 : INV_X1 port map( A => n465, ZN => n73);
   U277 : INV_X1 port map( A => n455, ZN => n76);
   U278 : INV_X1 port map( A => n267, ZN => n8);
   U279 : BUF_X1 port map( A => n44, Z => n43);
   U280 : BUF_X1 port map( A => n44, Z => n40);
   U281 : INV_X1 port map( A => n417, ZN => n130);
   U282 : INV_X1 port map( A => n400, ZN => n135);
   U283 : BUF_X1 port map( A => n44, Z => n41);
   U284 : INV_X1 port map( A => n373, ZN => n79);
   U285 : INV_X1 port map( A => n420, ZN => n132);
   U286 : INV_X1 port map( A => n407, ZN => n614);
   U287 : INV_X1 port map( A => n389, ZN => n616);
   U288 : INV_X1 port map( A => n429, ZN => n63);
   U289 : INV_X1 port map( A => n372, ZN => n91);
   U290 : INV_X1 port map( A => n361, ZN => n95);
   U291 : INV_X1 port map( A => n350, ZN => n99);
   U292 : INV_X1 port map( A => n339, ZN => n104);
   U293 : AND2_X1 port map( A1 => n238, A2 => n401, ZN => n237);
   U294 : INV_X1 port map( A => n234, ZN => n618);
   U295 : INV_X1 port map( A => n416, ZN => n110);
   U296 : OAI211_X1 port map( C1 => n417, C2 => n646, A => n401, B => n413, ZN 
                           => n416);
   U297 : INV_X1 port map( A => n399, ZN => n113);
   U298 : OAI211_X1 port map( C1 => n400, C2 => n646, A => n401, B => n396, ZN 
                           => n399);
   U299 : INV_X1 port map( A => n381, ZN => n115);
   U300 : AOI21_X1 port map( B1 => n260, B2 => n382, A => n383, ZN => n381);
   U301 : OR4_X1 port map( A1 => B(21), A2 => B(20), A3 => B(19), A4 => B(18), 
                           ZN => n598);
   U302 : OAI22_X1 port map( A1 => n88, A2 => n1, B1 => n86, B2 => n8, ZN => 
                           n568);
   U303 : AOI222_X1 port map( A1 => n11, A2 => A(1), B1 => A(0), B2 => n18, C1 
                           => n7, C2 => A(2), ZN => n293);
   U304 : AOI221_X1 port map( B1 => n31, B2 => A(6), C1 => n20, C2 => A(7), A 
                           => n525, ZN => n363);
   U305 : OAI22_X1 port map( A1 => n623, A2 => n1, B1 => n624, B2 => n8, ZN => 
                           n525);
   U306 : AOI221_X1 port map( B1 => n30, B2 => A(7), C1 => n20, C2 => A(8), A 
                           => n570, ZN => n405);
   U307 : OAI22_X1 port map( A1 => n624, A2 => n1, B1 => n66, B2 => n8, ZN => 
                           n570);
   U308 : AOI221_X1 port map( B1 => n31, B2 => A(8), C1 => n21, C2 => A(9), A 
                           => n552, ZN => n387);
   U309 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n74, B2 => n8, ZN => 
                           n552);
   U310 : AOI221_X1 port map( B1 => n30, B2 => A(5), C1 => n20, C2 => A(6), A 
                           => n541, ZN => n376);
   U311 : OAI22_X1 port map( A1 => n622, A2 => n1, B1 => n623, B2 => n8, ZN => 
                           n541);
   U312 : OAI221_X1 port map( B1 => n29, B2 => n613, C1 => n17, C2 => n266, A 
                           => n609, ZN => n320);
   U313 : AOI22_X1 port map( A1 => A(29), A2 => n10, B1 => A(28), B2 => n267, 
                           ZN => n609);
   U314 : OAI221_X1 port map( B1 => n27, B2 => n128, C1 => n15, C2 => n126, A 
                           => n535, ZN => n355);
   U315 : AOI22_X1 port map( A1 => A(26), A2 => n11, B1 => A(25), B2 => n6, ZN 
                           => n535);
   U316 : OAI221_X1 port map( B1 => n28, B2 => n131, C1 => n16, C2 => n128, A 
                           => n585, ZN => n403);
   U317 : AOI22_X1 port map( A1 => A(27), A2 => n9, B1 => A(26), B2 => n267, ZN
                           => n585);
   U318 : OR3_X1 port map( A1 => B(22), A2 => B(24), A3 => B(23), ZN => n594);
   U319 : NAND3_X1 port map( A1 => n489, A2 => n629, A3 => n600, ZN => n152);
   U320 : NOR3_X1 port map( A1 => B(12), A2 => B(14), A3 => B(13), ZN => n600);
   U321 : NAND3_X1 port map( A1 => n592, A2 => n632, A3 => n599, ZN => n146);
   U322 : INV_X1 port map( A => B(22), ZN => n632);
   U323 : NOR3_X1 port map( A1 => B(23), A2 => B(25), A3 => B(24), ZN => n599);
   U324 : NAND2_X1 port map( A1 => A(31), A2 => n648, ZN => n162);
   U325 : OAI221_X1 port map( B1 => n29, B2 => n86, C1 => n17, C2 => n83, A => 
                           n606, ZN => n184);
   U326 : AOI22_X1 port map( A1 => A(13), A2 => n10, B1 => A(12), B2 => n267, 
                           ZN => n606);
   U327 : OAI221_X1 port map( B1 => n29, B2 => n126, C1 => n17, C2 => n123, A 
                           => n608, ZN => n370);
   U328 : AOI22_X1 port map( A1 => A(25), A2 => n10, B1 => A(24), B2 => n267, 
                           ZN => n608);
   U329 : NAND2_X1 port map( A1 => n488, A2 => n489, ZN => n287);
   U330 : OAI221_X1 port map( B1 => n27, B2 => n117, C1 => n15, C2 => n114, A 
                           => n536, ZN => n168);
   U331 : AOI22_X1 port map( A1 => A(22), A2 => n9, B1 => A(21), B2 => n7, ZN 
                           => n536);
   U332 : OAI221_X1 port map( B1 => n28, B2 => n120, C1 => n16, C2 => n117, A 
                           => n583, ZN => n402);
   U333 : AOI22_X1 port map( A1 => A(23), A2 => n9, B1 => A(22), B2 => n267, ZN
                           => n583);
   U334 : AOI221_X1 port map( B1 => A(1), B2 => n32, C1 => A(2), C2 => n18, A 
                           => n540, ZN => n374);
   U335 : OAI22_X1 port map( A1 => n615, A2 => n1, B1 => n617, B2 => n8, ZN => 
                           n540);
   U336 : NAND2_X1 port map( A1 => A(31), A2 => n152, ZN => n153);
   U337 : NAND2_X1 port map( A1 => A(31), A2 => n146, ZN => n147);
   U338 : NOR2_X2 port map( A1 => n612, A2 => n591, ZN => n144);
   U339 : OAI221_X1 port map( B1 => n28, B2 => n266, C1 => n16, C2 => n131, A 
                           => n564, ZN => n506);
   U340 : AOI22_X1 port map( A1 => A(28), A2 => n9, B1 => A(27), B2 => n7, ZN 
                           => n564);
   U341 : OAI221_X1 port map( B1 => n28, B2 => n123, C1 => n16, C2 => n120, A 
                           => n565, ZN => n453);
   U342 : AOI22_X1 port map( A1 => A(24), A2 => n9, B1 => A(23), B2 => n7, ZN 
                           => n565);
   U343 : NOR2_X2 port map( A1 => n647, A2 => B(2), ZN => n260);
   U344 : OAI221_X1 port map( B1 => n26, B2 => n114, C1 => n14, C2 => n111, A 
                           => n611, ZN => n185);
   U345 : AOI22_X1 port map( A1 => A(21), A2 => n11, B1 => A(20), B2 => n6, ZN 
                           => n611);
   U346 : AOI222_X1 port map( A1 => n429, A2 => n5, B1 => n620, B2 => n262, C1 
                           => n227, C2 => B(3), ZN => n327);
   U347 : INV_X1 port map( A => n376, ZN => n620);
   U348 : OAI221_X1 port map( B1 => n26, B2 => n77, C1 => n15, C2 => n74, A => 
                           n444, ZN => n154);
   U349 : AOI22_X1 port map( A1 => A(10), A2 => n11, B1 => A(9), B2 => n6, ZN 
                           => n444);
   U350 : OAI221_X1 port map( B1 => n29, B2 => n80, C1 => n16, C2 => n77, A => 
                           n586, ZN => n305);
   U351 : AOI22_X1 port map( A1 => A(11), A2 => n10, B1 => A(10), B2 => n267, 
                           ZN => n586);
   U352 : OAI221_X1 port map( B1 => n28, B2 => n83, C1 => n16, C2 => n80, A => 
                           n567, ZN => n261);
   U353 : AOI22_X1 port map( A1 => A(12), A2 => n9, B1 => A(11), B2 => n7, ZN 
                           => n567);
   U354 : OAI221_X1 port map( B1 => n26, B2 => n623, C1 => n14, C2 => n622, A 
                           => n443, ZN => n219);
   U355 : AOI22_X1 port map( A1 => A(6), A2 => n11, B1 => A(5), B2 => n7, ZN =>
                           n443);
   U356 : OAI221_X1 port map( B1 => n26, B2 => n624, C1 => n14, C2 => n623, A 
                           => n306, ZN => n207);
   U357 : AOI22_X1 port map( A1 => A(7), A2 => n11, B1 => A(6), B2 => n6, ZN =>
                           n306);
   U358 : OAI221_X1 port map( B1 => n27, B2 => n66, C1 => n15, C2 => n624, A =>
                           n265, ZN => n193);
   U359 : AOI22_X1 port map( A1 => A(8), A2 => n10, B1 => A(7), B2 => n6, ZN =>
                           n265);
   U360 : OAI221_X1 port map( B1 => n29, B2 => n100, C1 => n17, C2 => n96, A =>
                           n610, ZN => n186);
   U361 : AOI22_X1 port map( A1 => A(17), A2 => n10, B1 => A(16), B2 => n267, 
                           ZN => n610);
   U362 : OAI221_X1 port map( B1 => n29, B2 => n74, C1 => n17, C2 => n66, A => 
                           n604, ZN => n178);
   U363 : AOI22_X1 port map( A1 => A(9), A2 => n10, B1 => A(8), B2 => n267, ZN 
                           => n604);
   U364 : OAI221_X1 port map( B1 => n27, B2 => n88, C1 => n15, C2 => n86, A => 
                           n537, ZN => n166);
   U365 : AOI22_X1 port map( A1 => A(14), A2 => n11, B1 => A(13), B2 => n7, ZN 
                           => n537);
   U366 : OAI221_X1 port map( B1 => n28, B2 => n92, C1 => n16, C2 => n88, A => 
                           n584, ZN => n516);
   U367 : AOI22_X1 port map( A1 => A(15), A2 => n9, B1 => A(14), B2 => n7, ZN 
                           => n584);
   U368 : OAI221_X1 port map( B1 => n27, B2 => n80, C1 => n15, C2 => n83, A => 
                           n494, ZN => n373);
   U369 : AOI22_X1 port map( A1 => A(15), A2 => n9, B1 => A(16), B2 => n6, ZN 
                           => n494);
   U370 : OAI221_X1 port map( B1 => n27, B2 => n133, C1 => n15, C2 => n615, A 
                           => n523, ZN => n420);
   U371 : AOI22_X1 port map( A1 => A(4), A2 => n10, B1 => A(5), B2 => n7, ZN =>
                           n523);
   U372 : OAI221_X1 port map( B1 => n28, B2 => n615, C1 => n16, C2 => n617, A 
                           => n571, ZN => n407);
   U373 : AOI22_X1 port map( A1 => A(5), A2 => n9, B1 => A(6), B2 => n7, ZN => 
                           n571);
   U374 : OAI221_X1 port map( B1 => n28, B2 => n617, C1 => n16, C2 => n619, A 
                           => n554, ZN => n389);
   U375 : AOI22_X1 port map( A1 => A(6), A2 => n9, B1 => A(7), B2 => n7, ZN => 
                           n554);
   U376 : OAI221_X1 port map( B1 => n49, B2 => n29, C1 => n103, C2 => n14, A =>
                           n553, ZN => n390);
   U377 : AOI22_X1 port map( A1 => A(2), A2 => n9, B1 => A(3), B2 => n7, ZN => 
                           n553);
   U378 : OAI221_X1 port map( B1 => n28, B2 => n624, C1 => n16, C2 => n66, A =>
                           n542, ZN => n429);
   U379 : AOI22_X1 port map( A1 => A(11), A2 => n9, B1 => A(12), B2 => n7, ZN 
                           => n542);
   U380 : OAI221_X1 port map( B1 => n28, B2 => n111, C1 => n16, C2 => n108, A 
                           => n566, ZN => n452);
   U381 : AOI22_X1 port map( A1 => A(20), A2 => n9, B1 => A(19), B2 => n7, ZN 
                           => n566);
   U382 : OAI221_X1 port map( B1 => n28, B2 => n105, C1 => n16, C2 => n100, A 
                           => n538, ZN => n170);
   U383 : AOI22_X1 port map( A1 => A(18), A2 => n9, B1 => A(17), B2 => n7, ZN 
                           => n538);
   U384 : OAI221_X1 port map( B1 => n28, B2 => n108, C1 => n16, C2 => n105, A 
                           => n582, ZN => n464);
   U385 : AOI22_X1 port map( A1 => A(19), A2 => n10, B1 => A(18), B2 => n7, ZN 
                           => n582);
   U386 : INV_X1 port map( A => A(31), ZN => n613);
   U387 : AOI22_X1 port map( A1 => n267, A2 => A(1), B1 => n11, B2 => A(0), ZN 
                           => n362);
   U389 : NAND2_X1 port map( A1 => B(4), A2 => n579, ZN => n160);
   U390 : OAI222_X1 port map( A1 => n79, A2 => n636, B1 => n326, B2 => n642, C1
                           => n91, C2 => n645, ZN => n325);
   U391 : AOI222_X1 port map( A1 => A(27), A2 => n10, B1 => A(25), B2 => n30, 
                           C1 => A(26), C2 => n18, ZN => n326);
   U392 : AOI222_X1 port map( A1 => A(28), A2 => n10, B1 => A(26), B2 => n30, 
                           C1 => A(27), C2 => n19, ZN => n316);
   U393 : AOI222_X1 port map( A1 => A(29), A2 => n11, B1 => A(27), B2 => n32, 
                           C1 => A(28), C2 => n18, ZN => n292);
   U394 : AOI222_X1 port map( A1 => A(30), A2 => n11, B1 => A(28), B2 => n30, 
                           C1 => A(29), C2 => n22, ZN => n273);
   U395 : AOI21_X1 port map( B1 => A(31), B2 => B(11), A => n487, ZN => n256);
   U396 : AOI21_X1 port map( B1 => A(31), B2 => B(25), A => n483, ZN => n250);
   U397 : OAI222_X1 port map( A1 => n171, A2 => n36, B1 => n55, B2 => n626, C1 
                           => n623, C2 => n33, ZN => RES(8));
   U398 : INV_X1 port map( A => n172, ZN => n55);
   U399 : AOI221_X1 port map( B1 => n140, B2 => n173, C1 => n142, C2 => n174, A
                           => n144, ZN => n171);
   U400 : OAI21_X1 port map( B1 => n175, B2 => n146, A => n147, ZN => n174);
   U401 : OAI222_X1 port map( A1 => n187, A2 => n36, B1 => n188, B2 => n626, C1
                           => n622, C2 => n33, ZN => RES(7));
   U402 : AOI221_X1 port map( B1 => n140, B2 => n61, C1 => n142, C2 => n189, A 
                           => n144, ZN => n187);
   U403 : INV_X1 port map( A => n198, ZN => n61);
   U404 : OAI21_X1 port map( B1 => n190, B2 => n146, A => n147, ZN => n189);
   U405 : OAI222_X1 port map( A1 => n136, A2 => n36, B1 => n59, B2 => n626, C1 
                           => n624, C2 => n33, ZN => RES(9));
   U406 : INV_X1 port map( A => n139, ZN => n59);
   U407 : AOI221_X1 port map( B1 => n140, B2 => n141, C1 => n142, C2 => n143, A
                           => n144, ZN => n136);
   U408 : OAI21_X1 port map( B1 => n145, B2 => n146, A => n147, ZN => n143);
   U409 : OAI222_X1 port map( A1 => n539, A2 => n36, B1 => n327, B2 => n626, C1
                           => n77, C2 => n35, ZN => RES(12));
   U410 : AOI221_X1 port map( B1 => n140, B2 => n543, C1 => n142, C2 => n544, A
                           => n144, ZN => n539);
   U411 : OAI21_X1 port map( B1 => n545, B2 => n146, A => n147, ZN => n544);
   U412 : OAI221_X1 port map( B1 => n90, B2 => n638, C1 => n78, C2 => n642, A 
                           => n550, ZN => n543);
   U413 : OAI222_X1 port map( A1 => n521, A2 => n36, B1 => n57, B2 => n626, C1 
                           => n80, C2 => n35, ZN => RES(13));
   U414 : INV_X1 port map( A => n314, ZN => n57);
   U415 : AOI221_X1 port map( B1 => n140, B2 => n526, C1 => n142, C2 => n527, A
                           => n144, ZN => n521);
   U416 : OAI21_X1 port map( B1 => n528, B2 => n146, A => n147, ZN => n527);
   U417 : OAI222_X1 port map( A1 => n508, A2 => n36, B1 => n51, B2 => n626, C1 
                           => n83, C2 => n35, ZN => RES(14));
   U418 : INV_X1 port map( A => n290, ZN => n51);
   U419 : AOI221_X1 port map( B1 => n140, B2 => n511, C1 => n142, C2 => n512, A
                           => n144, ZN => n508);
   U420 : OAI21_X1 port map( B1 => n513, B2 => n146, A => n147, ZN => n512);
   U421 : OAI222_X1 port map( A1 => n551, A2 => n36, B1 => n45, B2 => n626, C1 
                           => n74, C2 => n35, ZN => RES(11));
   U422 : INV_X1 port map( A => n337, ZN => n45);
   U423 : AOI221_X1 port map( B1 => n140, B2 => n555, C1 => n142, C2 => n556, A
                           => n144, ZN => n551);
   U424 : OAI21_X1 port map( B1 => n557, B2 => n146, A => n147, ZN => n556);
   U425 : OAI222_X1 port map( A1 => n495, A2 => n36, B1 => n47, B2 => n626, C1 
                           => n86, C2 => n35, ZN => RES(15));
   U426 : INV_X1 port map( A => n271, ZN => n47);
   U427 : AOI221_X1 port map( B1 => n140, B2 => n498, C1 => n142, C2 => n499, A
                           => n144, ZN => n495);
   U429 : OAI21_X1 port map( B1 => n500, B2 => n146, A => n147, ZN => n499);
   U430 : OAI222_X1 port map( A1 => n569, A2 => n36, B1 => n53, B2 => n626, C1 
                           => n66, C2 => n35, ZN => RES(10));
   U431 : INV_X1 port map( A => n348, ZN => n53);
   U432 : AOI221_X1 port map( B1 => n140, B2 => n572, C1 => n142, C2 => n573, A
                           => n144, ZN => n569);
   U433 : OAI21_X1 port map( B1 => n574, B2 => n146, A => n147, ZN => n573);
   U434 : OAI222_X1 port map( A1 => n201, A2 => n36, B1 => n202, B2 => n626, C1
                           => n621, C2 => n33, ZN => RES(6));
   U435 : AOI221_X1 port map( B1 => n140, B2 => n67, C1 => n142, C2 => n203, A 
                           => n144, ZN => n201);
   U436 : INV_X1 port map( A => n210, ZN => n67);
   U437 : OAI21_X1 port map( B1 => n204, B2 => n146, A => n147, ZN => n203);
   U438 : OAI222_X1 port map( A1 => n213, A2 => n36, B1 => n214, B2 => n626, C1
                           => n619, C2 => n33, ZN => RES(5));
   U439 : AOI221_X1 port map( B1 => n140, B2 => n70, C1 => n142, C2 => n215, A 
                           => n144, ZN => n213);
   U440 : INV_X1 port map( A => n222, ZN => n70);
   U441 : OAI21_X1 port map( B1 => n216, B2 => n146, A => n147, ZN => n215);
   U442 : OAI221_X1 port map( B1 => n27, B2 => n83, C1 => n15, C2 => n86, A => 
                           n476, ZN => n419);
   U443 : AOI22_X1 port map( A1 => A(16), A2 => n11, B1 => A(17), B2 => n6, ZN 
                           => n476);
   U444 : OAI221_X1 port map( B1 => n27, B2 => n86, C1 => n15, C2 => n88, A => 
                           n467, ZN => n406);
   U445 : AOI22_X1 port map( A1 => A(17), A2 => n9, B1 => A(18), B2 => n7, ZN 
                           => n467);
   U446 : OAI221_X1 port map( B1 => n27, B2 => n88, C1 => n15, C2 => n92, A => 
                           n457, ZN => n388);
   U447 : AOI22_X1 port map( A1 => A(18), A2 => n10, B1 => A(19), B2 => n6, ZN 
                           => n457);
   U448 : OAI221_X1 port map( B1 => n26, B2 => n92, C1 => n14, C2 => n96, A => 
                           n430, ZN => n372);
   U449 : AOI22_X1 port map( A1 => A(19), A2 => n11, B1 => A(20), B2 => n6, ZN 
                           => n430);
   U450 : OAI221_X1 port map( B1 => n29, B2 => n622, C1 => n17, C2 => n621, A 
                           => n605, ZN => n234);
   U451 : AOI22_X1 port map( A1 => A(5), A2 => n10, B1 => A(4), B2 => n267, ZN 
                           => n605);
   U452 : OAI221_X1 port map( B1 => n258, B2 => n643, C1 => n196, C2 => n637, A
                           => n259, ZN => n247);
   U453 : AOI22_X1 port map( A1 => n260, A2 => n261, B1 => n262, B2 => n193, ZN
                           => n259);
   U454 : AOI222_X1 port map( A1 => A(4), A2 => n11, B1 => A(6), B2 => n31, C1 
                           => A(5), C2 => n19, ZN => n258);
   U455 : OAI221_X1 port map( B1 => n303, B2 => n643, C1 => n84, C2 => n637, A 
                           => n304, ZN => n298);
   U456 : AOI22_X1 port map( A1 => n260, A2 => n305, B1 => n262, B2 => n207, ZN
                           => n304);
   U457 : AOI222_X1 port map( A1 => A(3), A2 => n10, B1 => A(5), B2 => n32, C1 
                           => A(4), C2 => n19, ZN => n303);
   U458 : OAI221_X1 port map( B1 => n441, B2 => n643, C1 => n81, C2 => n637, A 
                           => n442, ZN => n435);
   U459 : AOI22_X1 port map( A1 => n260, A2 => n154, B1 => n262, B2 => n219, ZN
                           => n442);
   U460 : AOI222_X1 port map( A1 => A(2), A2 => n10, B1 => A(4), B2 => n30, C1 
                           => A(3), C2 => n20, ZN => n441);
   U462 : INV_X1 port map( A => n228, ZN => n626);
   U463 : OAI221_X1 port map( B1 => n27, B2 => n66, C1 => n15, C2 => n74, A => 
                           n524, ZN => n474);
   U464 : AOI22_X1 port map( A1 => A(12), A2 => n11, B1 => A(13), B2 => n7, ZN 
                           => n524);
   U465 : OAI221_X1 port map( B1 => n27, B2 => n74, C1 => n15, C2 => n77, A => 
                           n510, ZN => n465);
   U466 : AOI22_X1 port map( A1 => A(13), A2 => n9, B1 => A(14), B2 => n6, ZN 
                           => n510);
   U467 : OAI221_X1 port map( B1 => n27, B2 => n77, C1 => n15, C2 => n80, A => 
                           n497, ZN => n455);
   U468 : AOI22_X1 port map( A1 => A(14), A2 => n10, B1 => A(15), B2 => n7, ZN 
                           => n497);
   U469 : OAI221_X1 port map( B1 => n26, B2 => n96, C1 => n14, C2 => n100, A =>
                           n421, ZN => n361);
   U470 : AOI22_X1 port map( A1 => A(20), A2 => n11, B1 => A(21), B2 => n6, ZN 
                           => n421);
   U471 : OAI221_X1 port map( B1 => n26, B2 => n100, C1 => n14, C2 => n105, A 
                           => n408, ZN => n350);
   U472 : AOI22_X1 port map( A1 => A(21), A2 => n11, B1 => A(22), B2 => n6, ZN 
                           => n408);
   U473 : OAI221_X1 port map( B1 => n26, B2 => n105, C1 => n14, C2 => n108, A 
                           => n391, ZN => n339);
   U474 : AOI22_X1 port map( A1 => A(22), A2 => n9, B1 => A(23), B2 => n6, ZN 
                           => n391);
   U475 : OAI221_X1 port map( B1 => n26, B2 => n108, C1 => n14, C2 => n111, A 
                           => n377, ZN => n324);
   U476 : AOI22_X1 port map( A1 => A(23), A2 => n9, B1 => A(24), B2 => n6, ZN 
                           => n377);
   U477 : OAI221_X1 port map( B1 => n26, B2 => n111, C1 => n14, C2 => n114, A 
                           => n364, ZN => n313);
   U478 : AOI22_X1 port map( A1 => A(24), A2 => n10, B1 => A(25), B2 => n6, ZN 
                           => n364);
   U479 : OAI221_X1 port map( B1 => n26, B2 => n114, C1 => n14, C2 => n117, A 
                           => n351, ZN => n289);
   U480 : AOI22_X1 port map( A1 => A(25), A2 => n11, B1 => A(26), B2 => n6, ZN 
                           => n351);
   U481 : OAI221_X1 port map( B1 => n26, B2 => n117, C1 => n14, C2 => n120, A 
                           => n340, ZN => n270);
   U482 : AOI22_X1 port map( A1 => A(26), A2 => n10, B1 => A(27), B2 => n6, ZN 
                           => n340);
   U483 : AOI22_X1 port map( A1 => n640, A2 => n506, B1 => B(2), B2 => n382, ZN
                           => n333);
   U484 : AOI21_X1 port map( B1 => n22, B2 => A(31), A => n533, ZN => n412);
   U485 : AOI21_X1 port map( B1 => n11, B2 => A(31), A => n580, ZN => n395);
   U486 : AOI21_X1 port map( B1 => B(1), B2 => A(31), A => n533, ZN => n417);
   U487 : AOI21_X1 port map( B1 => n8, B2 => A(31), A => n580, ZN => n400);
   U488 : NOR2_X1 port map( A1 => n490, A2 => B(18), ZN => n251);
   U489 : OAI22_X1 port map( A1 => B(2), A2 => n374, B1 => n640, B2 => n375, ZN
                           => n227);
   U490 : OAI221_X1 port map( B1 => n196, B2 => n638, C1 => n75, C2 => n642, A 
                           => n562, ZN => n555);
   U491 : AOI221_X1 port map( B1 => n169, B2 => n452, C1 => n167, C2 => n453, A
                           => n563, ZN => n562);
   U492 : NOR3_X1 port map( A1 => n41, A2 => B(3), A3 => n333, ZN => n563);
   U493 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n267);
   U494 : AOI21_X1 port map( B1 => n634, B2 => n590, A => n144, ZN => n481);
   U495 : INV_X1 port map( A => n592, ZN => n634);
   U496 : NAND2_X1 port map( A1 => A(31), A2 => n490, ZN => n486);
   U497 : OAI221_X1 port map( B1 => n225, B2 => n36, C1 => n617, C2 => n33, A 
                           => n226, ZN => RES(4));
   U498 : AOI221_X1 port map( B1 => n140, B2 => n229, C1 => n142, C2 => n230, A
                           => n144, ZN => n225);
   U499 : OAI21_X1 port map( B1 => n231, B2 => n146, A => n147, ZN => n230);
   U500 : NAND2_X1 port map( A1 => n454, A2 => A(31), ZN => n401);
   U501 : NOR2_X1 port map( A1 => B(2), A2 => B(3), ZN => n356);
   U502 : AOI21_X1 port map( B1 => n148, B2 => n501, A => n150, ZN => n500);
   U503 : OAI21_X1 port map( B1 => n502, B2 => n152, A => n153, ZN => n501);
   U504 : AOI211_X1 port map( C1 => B(4), C2 => A(31), A => n503, B => n504, ZN
                           => n502);
   U505 : OAI22_X1 port map( A1 => n196, A2 => n505, B1 => n101, B2 => n157, ZN
                           => n504);
   U506 : INV_X1 port map( A => A(10), ZN => n66);
   U507 : OAI21_X1 port map( B1 => n489, B2 => n613, A => n162, ZN => n487);
   U508 : NOR3_X1 port map( A1 => n332, A2 => B(3), A3 => n333, ZN => n331);
   U509 : INV_X1 port map( A => B(3), ZN => n647);
   U510 : INV_X1 port map( A => A(11), ZN => n74);
   U511 : INV_X1 port map( A => A(15), ZN => n86);
   U512 : INV_X1 port map( A => A(9), ZN => n624);
   U513 : INV_X1 port map( A => A(16), ZN => n88);
   U514 : BUF_X1 port map( A => n137, Z => n36);
   U515 : BUF_X1 port map( A => n137, Z => n37);
   U516 : NAND2_X1 port map( A1 => A(0), A2 => n6, ZN => n375);
   U517 : INV_X1 port map( A => A(23), ZN => n114);
   U518 : INV_X1 port map( A => A(19), ZN => n100);
   U519 : INV_X1 port map( A => A(24), ZN => n117);
   U520 : INV_X1 port map( A => A(20), ZN => n105);
   U521 : INV_X1 port map( A => A(21), ZN => n108);
   U522 : INV_X1 port map( A => A(22), ZN => n111);
   U523 : INV_X1 port map( A => A(8), ZN => n623);
   U524 : INV_X1 port map( A => A(12), ZN => n77);
   U525 : INV_X1 port map( A => A(13), ZN => n80);
   U526 : INV_X1 port map( A => A(14), ZN => n83);
   U527 : INV_X1 port map( A => A(30), ZN => n266);
   U528 : INV_X1 port map( A => A(3), ZN => n615);
   U529 : OR4_X1 port map( A1 => B(13), A2 => B(14), A3 => B(12), A4 => n596, 
                           ZN => n490);
   U530 : OR3_X1 port map( A1 => B(15), A2 => B(17), A3 => B(16), ZN => n596);
   U531 : INV_X1 port map( A => B(2), ZN => n640);
   U532 : INV_X1 port map( A => A(17), ZN => n92);
   U533 : INV_X1 port map( A => A(7), ZN => n622);
   U534 : INV_X1 port map( A => A(18), ZN => n96);
   U535 : INV_X1 port map( A => A(25), ZN => n120);
   U536 : AND3_X1 port map( A1 => n579, A2 => n591, A3 => n597, ZN => n445);
   U537 : NOR3_X1 port map( A1 => n152, A2 => n146, A3 => n630, ZN => n597);
   U538 : INV_X1 port map( A => n148, ZN => n630);
   U539 : INV_X1 port map( A => A(4), ZN => n617);
   U540 : INV_X1 port map( A => n590, ZN => n612);
   U541 : INV_X1 port map( A => A(27), ZN => n126);
   U542 : INV_X1 port map( A => A(26), ZN => n123);
   U543 : INV_X1 port map( A => A(6), ZN => n621);
   U544 : INV_X1 port map( A => A(5), ZN => n619);
   U545 : INV_X1 port map( A => A(28), ZN => n128);
   U546 : INV_X1 port map( A => A(29), ZN => n131);
   U547 : INV_X1 port map( A => B(25), ZN => n633);
   U548 : INV_X1 port map( A => A(2), ZN => n133);
   U549 : AND2_X1 port map( A1 => n140, A2 => n199, ZN => n278);
   U550 : INV_X1 port map( A => A(1), ZN => n103);
   U551 : INV_X1 port map( A => n579, ZN => n648);
   U552 : INV_X1 port map( A => A(0), ZN => n49);
   U553 : OR2_X1 port map( A1 => n625, A2 => B(1), ZN => n1);
   U554 : NAND2_X1 port map( A1 => n140, A2 => n40, ZN => n332);
   U555 : INV_X1 port map( A => n436, ZN => n627);
   U556 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n263);
   U557 : NAND2_X1 port map( A1 => B(1), A2 => n625, ZN => n264);
   U558 : INV_X1 port map( A => B(11), ZN => n629);
   U559 : INV_X1 port map( A => B(18), ZN => n631);
   U560 : AND2_X1 port map( A1 => n142, A2 => n592, ZN => n491);
   U561 : BUF_X1 port map( A => n137, Z => n38);
   U562 : INV_X1 port map( A => B(0), ZN => n625);
   U563 : INV_X1 port map( A => B(4), ZN => n44);
   U564 : NOR2_X2 port map( A1 => n635, A2 => LOGIC_ARITH, ZN => n142);
   U565 : INV_X1 port map( A => n591, ZN => n635);
   U566 : NOR3_X1 port map( A1 => B(9), A2 => B(8), A3 => B(10), ZN => n489);
   U567 : NOR3_X1 port map( A1 => B(7), A2 => B(6), A3 => B(5), ZN => n579);
   U568 : NOR3_X1 port map( A1 => B(28), A2 => B(27), A3 => B(26), ZN => n592);
   U569 : OAI222_X1 port map( A1 => n468, A2 => n269, B1 => n469, B2 => n37, C1
                           => n92, C2 => n34, ZN => RES(17));
   U570 : AOI221_X1 port map( B1 => n165, B2 => n474, C1 => n199, C2 => n419, A
                           => n475, ZN => n468);
   U571 : AOI221_X1 port map( B1 => n276, B2 => n470, C1 => n628, C2 => n434, A
                           => n279, ZN => n469);
   U572 : OAI222_X1 port map( A1 => n132, A2 => n636, B1 => n362, B2 => n641, 
                           C1 => n363, C2 => n645, ZN => n475);
   U573 : OAI222_X1 port map( A1 => n458, A2 => n269, B1 => n459, B2 => n38, C1
                           => n96, C2 => n34, ZN => RES(18));
   U574 : AOI221_X1 port map( B1 => n165, B2 => n465, C1 => n199, C2 => n406, A
                           => n466, ZN => n458);
   U575 : AOI221_X1 port map( B1 => n276, B2 => n460, C1 => n628, C2 => n297, A
                           => n279, ZN => n459);
   U576 : OAI222_X1 port map( A1 => n614, A2 => n636, B1 => n293, B2 => n641, 
                           C1 => n405, C2 => n645, ZN => n466);
   U577 : OAI222_X1 port map( A1 => n446, A2 => n269, B1 => n447, B2 => n37, C1
                           => n100, C2 => n34, ZN => RES(19));
   U578 : AOI221_X1 port map( B1 => n165, B2 => n455, C1 => n199, C2 => n388, A
                           => n456, ZN => n446);
   U579 : AOI221_X1 port map( B1 => n276, B2 => n448, C1 => n628, C2 => n246, A
                           => n279, ZN => n447);
   U580 : OAI222_X1 port map( A1 => n616, A2 => n636, B1 => n46, B2 => n641, C1
                           => n387, C2 => n645, ZN => n456);
   U581 : OAI222_X1 port map( A1 => n422, A2 => n269, B1 => n423, B2 => n37, C1
                           => n105, C2 => n34, ZN => RES(20));
   U582 : AOI221_X1 port map( B1 => n165, B2 => n373, C1 => n199, C2 => n372, A
                           => n427, ZN => n422);
   U583 : AOI221_X1 port map( B1 => n276, B2 => n424, C1 => n628, C2 => n107, A
                           => n279, ZN => n423);
   U584 : OAI221_X1 port map( B1 => n376, B2 => n636, C1 => n63, C2 => n645, A 
                           => n428, ZN => n427);
   U585 : OAI222_X1 port map( A1 => n409, A2 => n269, B1 => n410, B2 => n37, C1
                           => n108, C2 => n34, ZN => RES(21));
   U586 : AOI221_X1 port map( B1 => n276, B2 => n411, C1 => n628, C2 => n223, A
                           => n279, ZN => n410);
   U587 : AOI221_X1 port map( B1 => n199, B2 => n361, C1 => B(4), C2 => n56, A 
                           => n418, ZN => n409);
   U588 : OAI21_X1 port map( B1 => n414, B2 => n281, A => n282, ZN => n411);
   U589 : OAI222_X1 port map( A1 => n392, A2 => n269, B1 => n393, B2 => n37, C1
                           => n111, C2 => n34, ZN => RES(22));
   U590 : AOI221_X1 port map( B1 => n276, B2 => n394, C1 => n628, C2 => n211, A
                           => n279, ZN => n393);
   U591 : AOI221_X1 port map( B1 => n199, B2 => n350, C1 => B(4), C2 => n50, A 
                           => n404, ZN => n392);
   U592 : OAI21_X1 port map( B1 => n397, B2 => n281, A => n282, ZN => n394);
   U593 : OAI222_X1 port map( A1 => n378, A2 => n269, B1 => n379, B2 => n37, C1
                           => n114, C2 => n34, ZN => RES(23));
   U594 : AOI221_X1 port map( B1 => n276, B2 => n380, C1 => n628, C2 => n115, A
                           => n279, ZN => n379);
   U595 : AOI221_X1 port map( B1 => n199, B2 => n339, C1 => B(4), C2 => n48, A 
                           => n386, ZN => n378);
   U596 : OAI21_X1 port map( B1 => n384, B2 => n281, A => n282, ZN => n380);
   U597 : OAI222_X1 port map( A1 => n365, A2 => n269, B1 => n366, B2 => n37, C1
                           => n117, C2 => n34, ZN => RES(24));
   U598 : AOI221_X1 port map( B1 => n276, B2 => n367, C1 => n628, C2 => n119, A
                           => n279, ZN => n366);
   U599 : AOI221_X1 port map( B1 => n199, B2 => n324, C1 => n39, C2 => n172, A 
                           => n371, ZN => n365);
   U600 : OAI21_X1 port map( B1 => n368, B2 => n281, A => n282, ZN => n367);
   U601 : OAI222_X1 port map( A1 => n352, A2 => n269, B1 => n353, B2 => n37, C1
                           => n120, C2 => n34, ZN => RES(25));
   U602 : AOI221_X1 port map( B1 => n276, B2 => n354, C1 => n628, C2 => n122, A
                           => n279, ZN => n353);
   U603 : AOI221_X1 port map( B1 => n199, B2 => n313, C1 => n39, C2 => n139, A 
                           => n360, ZN => n352);
   U604 : INV_X1 port map( A => n163, ZN => n122);
   U605 : OAI222_X1 port map( A1 => n477, A2 => n269, B1 => n478, B2 => n38, C1
                           => n88, C2 => n35, ZN => RES(16));
   U606 : AOI221_X1 port map( B1 => n165, B2 => n429, C1 => n199, C2 => n373, A
                           => n492, ZN => n477);
   U607 : AOI221_X1 port map( B1 => n276, B2 => n479, C1 => n628, C2 => n480, A
                           => n279, ZN => n478);
   U608 : OAI222_X1 port map( A1 => n374, A2 => n636, B1 => n375, B2 => n641, 
                           C1 => n376, C2 => n645, ZN => n492);
   U609 : OAI222_X1 port map( A1 => n341, A2 => n269, B1 => n342, B2 => n37, C1
                           => n123, C2 => n34, ZN => RES(26));
   U610 : AOI221_X1 port map( B1 => n276, B2 => n343, C1 => n628, C2 => n125, A
                           => n279, ZN => n342);
   U611 : AOI221_X1 port map( B1 => n199, B2 => n289, C1 => n39, C2 => n348, A 
                           => n349, ZN => n341);
   U612 : INV_X1 port map( A => n344, ZN => n125);
   U613 : OAI222_X1 port map( A1 => n328, A2 => n269, B1 => n329, B2 => n37, C1
                           => n126, C2 => n34, ZN => RES(27));
   U614 : AOI211_X1 port map( C1 => n276, C2 => n330, A => n279, B => n331, ZN 
                           => n329);
   U615 : AOI221_X1 port map( B1 => n199, B2 => n270, C1 => n39, C2 => n337, A 
                           => n338, ZN => n328);
   U616 : OAI21_X1 port map( B1 => n334, B2 => n281, A => n282, ZN => n330);
   U617 : OAI222_X1 port map( A1 => n317, A2 => n269, B1 => n318, B2 => n37, C1
                           => n128, C2 => n34, ZN => RES(28));
   U618 : AOI221_X1 port map( B1 => n165, B2 => n324, C1 => n39, C2 => n54, A 
                           => n325, ZN => n317);
   U619 : AOI221_X1 port map( B1 => n276, B2 => n319, C1 => n278, C2 => n320, A
                           => n279, ZN => n318);
   U620 : INV_X1 port map( A => n327, ZN => n54);
   U621 : OAI222_X1 port map( A1 => n307, A2 => n269, B1 => n308, B2 => n37, C1
                           => n131, C2 => n33, ZN => RES(29));
   U622 : AOI221_X1 port map( B1 => n165, B2 => n313, C1 => n39, C2 => n314, A 
                           => n315, ZN => n307);
   U623 : AOI221_X1 port map( B1 => n276, B2 => n309, C1 => n278, C2 => n129, A
                           => n279, ZN => n308);
   U624 : OAI222_X1 port map( A1 => n82, A2 => n636, B1 => n316, B2 => n642, C1
                           => n95, C2 => n645, ZN => n315);
   U625 : OAI222_X1 port map( A1 => n274, A2 => n269, B1 => n275, B2 => n38, C1
                           => n266, C2 => n33, ZN => RES(30));
   U626 : AOI221_X1 port map( B1 => n165, B2 => n289, C1 => n39, C2 => n290, A 
                           => n291, ZN => n274);
   U627 : AOI221_X1 port map( B1 => n276, B2 => n277, C1 => n278, C2 => n134, A
                           => n279, ZN => n275);
   U628 : OAI222_X1 port map( A1 => n85, A2 => n636, B1 => n292, B2 => n642, C1
                           => n99, C2 => n645, ZN => n291);
   U629 : OAI221_X1 port map( B1 => n293, B2 => n240, C1 => n133, C2 => n33, A 
                           => n294, ZN => RES(2));
   U630 : AOI221_X1 port map( B1 => n242, B2 => n295, C1 => n627, C2 => n69, A 
                           => n244, ZN => n294);
   U631 : INV_X1 port map( A => n296, ZN => n69);
   U632 : OAI21_X1 port map( B1 => n299, B2 => n249, A => n250, ZN => n295);
   U633 : OAI221_X1 port map( B1 => n362, B2 => n240, C1 => n103, C2 => n33, A 
                           => n431, ZN => RES(1));
   U634 : AOI221_X1 port map( B1 => n242, B2 => n432, C1 => n627, C2 => n72, A 
                           => n244, ZN => n431);
   U635 : INV_X1 port map( A => n433, ZN => n72);
   U636 : OAI21_X1 port map( B1 => n437, B2 => n249, A => n250, ZN => n432);
   U640 : OAI221_X1 port map( B1 => n46, B2 => n240, C1 => n615, C2 => n33, A 
                           => n241, ZN => RES(3));
   U643 : AOI221_X1 port map( B1 => n242, B2 => n243, C1 => n627, C2 => n60, A 
                           => n244, ZN => n241);
   U644 : INV_X1 port map( A => n245, ZN => n60);
   U645 : OAI21_X1 port map( B1 => n248, B2 => n249, A => n250, ZN => n243);
   U646 : NOR2_X1 port map( A1 => B(29), A2 => B(30), ZN => n591);
   U647 : AND2_X1 port map( A1 => LOGIC_ARITH, A2 => n445, ZN => n140);
   U648 : NOR2_X1 port map( A1 => n613, A2 => LOGIC_ARITH, ZN => n590);
   U649 : OAI221_X1 port map( B1 => n587, B2 => n436, C1 => n49, C2 => n33, A 
                           => n588, ZN => RES(0));
   U650 : NOR2_X1 port map( A1 => n269, A2 => n39, ZN => n228);
   U651 : AOI21_X1 port map( B1 => n242, B2 => n589, A => n244, ZN => n588);
   U652 : OAI21_X1 port map( B1 => n593, B2 => n249, A => n250, ZN => n589);
   U653 : AOI21_X1 port map( B1 => n251, B2 => n595, A => n253, ZN => n593);
   U654 : OAI21_X1 port map( B1 => n587, B2 => n255, A => n256, ZN => n595);
   U655 : AND2_X1 port map( A1 => n491, A2 => n649, ZN => n242);
   U656 : NAND2_X1 port map( A1 => n35, A2 => n649, ZN => n137);
   U657 : NAND2_X1 port map( A1 => n140, A2 => n649, ZN => n436);
   U658 : NOR2_X1 port map( A1 => n481, A2 => LEFT_RIGHT, ZN => n244);
   U659 : INV_X1 port map( A => LEFT_RIGHT, ZN => n649);
   U660 : OAI222_X1 port map( A1 => n268, A2 => n269, B1 => LEFT_RIGHT, B2 => 
                           n612, C1 => n613, C2 => n34, ZN => RES(31));
   U661 : AOI221_X1 port map( B1 => n165, B2 => n270, C1 => n39, C2 => n271, A 
                           => n272, ZN => n268);
   U662 : OAI222_X1 port map( A1 => n87, A2 => n636, B1 => n273, B2 => n642, C1
                           => n104, C2 => n645, ZN => n272);
   U663 : NOR4_X4 port map( A1 => B(16), A2 => B(17), A3 => B(15), A4 => n598, 
                           ZN => n148);
   U664 : INV_X1 port map( A => n8, ZN => n6);
   U665 : INV_X1 port map( A => n8, ZN => n7);
   U666 : INV_X1 port map( A => n1, ZN => n9);
   U667 : INV_X1 port map( A => n1, ZN => n10);
   U668 : INV_X1 port map( A => n1, ZN => n11);
   U669 : CLKBUF_X1 port map( A => n264, Z => n12);
   U670 : CLKBUF_X1 port map( A => n264, Z => n13);
   U671 : INV_X1 port map( A => n19, ZN => n17);
   U672 : INV_X1 port map( A => n12, ZN => n18);
   U673 : INV_X1 port map( A => n12, ZN => n19);
   U674 : INV_X1 port map( A => n264, ZN => n20);
   U675 : INV_X1 port map( A => n13, ZN => n21);
   U676 : INV_X1 port map( A => n13, ZN => n22);
   U677 : CLKBUF_X1 port map( A => n263, Z => n23);
   U678 : CLKBUF_X1 port map( A => n263, Z => n24);
   U679 : CLKBUF_X1 port map( A => n263, Z => n25);
   U680 : INV_X1 port map( A => n23, ZN => n30);
   U681 : INV_X1 port map( A => n24, ZN => n31);
   U682 : INV_X1 port map( A => n25, ZN => n32);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity comparator_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  OPSel : in std_logic_vector
         (0 to 2);  RES : out std_logic_vector (31 downto 0));

end comparator_NBIT32;

architecture SYN_bhv of comparator_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component comparator_NBIT32_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   signal X_Logic0_port, N26, N27, N28, N29, N30, N31, n10, n15, n16, n17, n18,
      n19, n20, RES_0_port, n2, n3, n4 : std_logic;

begin
   RES <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, RES_0_port 
      );
   
   X_Logic0_port <= '0';
   n10 <= '0';
   r57 : comparator_NBIT32_DW01_cmp6_0 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), TC => n10, LT => N30, GT => N28,
                           EQ => N26, LE => N31, GE => N29, NE => N27);
   U3 : INV_X1 port map( A => n15, ZN => RES_0_port);
   U4 : AOI21_X1 port map( B1 => n16, B2 => n4, A => n17, ZN => n15);
   U5 : INV_X1 port map( A => OPSel(2), ZN => n3);
   U6 : OAI22_X1 port map( A1 => n19, A2 => n2, B1 => OPSel(1), B2 => n20, ZN 
                           => n16);
   U7 : INV_X1 port map( A => OPSel(1), ZN => n2);
   U8 : AOI22_X1 port map( A1 => N28, A2 => n3, B1 => N29, B2 => OPSel(2), ZN 
                           => n19);
   U9 : AOI22_X1 port map( A1 => N26, A2 => n3, B1 => N27, B2 => OPSel(2), ZN 
                           => n20);
   U10 : NOR3_X1 port map( A1 => n4, A2 => OPSel(1), A3 => n18, ZN => n17);
   U11 : AOI22_X1 port map( A1 => N30, A2 => n3, B1 => OPSel(2), B2 => N31, ZN 
                           => n18);
   U12 : INV_X1 port map( A => OPSel(0), ZN => n4);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_NBIT32 is

   port( OP1, OP2 : in std_logic_vector (31 downto 0);  ALU_OPC : in 
         std_logic_vector (0 to 4);  ALU_RES : out std_logic_vector (31 downto 
         0));

end ALU_NBIT32;

architecture SYN_struct of ALU_NBIT32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux21_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux41_NBIT32_1
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component BOOTHMUL_numBit16
      port( A, B : in std_logic_vector (15 downto 0);  P : out std_logic_vector
            (31 downto 0));
   end component;
   
   component P4Adder_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component shifter_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  LOGIC_ARITH, LEFT_RIGHT 
            : in std_logic;  RES : out std_logic_vector (31 downto 0));
   end component;
   
   component comparator_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  OPSel : in 
            std_logic_vector (0 to 2);  RES : out std_logic_vector (31 downto 
            0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, select_type_sig_1_port, select_type_sig_0_port, 
      select_zero_sig, A_CMP_31_port, A_CMP_30_port, A_CMP_29_port, 
      A_CMP_28_port, A_CMP_27_port, A_CMP_26_port, A_CMP_25_port, A_CMP_24_port
      , A_CMP_23_port, A_CMP_22_port, A_CMP_21_port, A_CMP_20_port, 
      A_CMP_19_port, A_CMP_18_port, A_CMP_17_port, A_CMP_16_port, A_CMP_15_port
      , A_CMP_14_port, A_CMP_13_port, A_CMP_12_port, A_CMP_11_port, 
      A_CMP_10_port, A_CMP_9_port, A_CMP_8_port, A_CMP_7_port, A_CMP_6_port, 
      A_CMP_5_port, A_CMP_4_port, A_CMP_3_port, A_CMP_2_port, A_CMP_1_port, 
      A_CMP_0_port, B_CMP_31_port, B_CMP_30_port, B_CMP_29_port, B_CMP_28_port,
      B_CMP_27_port, B_CMP_26_port, B_CMP_25_port, B_CMP_24_port, B_CMP_23_port
      , B_CMP_22_port, B_CMP_21_port, B_CMP_20_port, B_CMP_19_port, 
      B_CMP_18_port, B_CMP_17_port, B_CMP_16_port, B_CMP_15_port, B_CMP_14_port
      , B_CMP_13_port, B_CMP_12_port, B_CMP_11_port, B_CMP_10_port, 
      B_CMP_9_port, B_CMP_8_port, B_CMP_7_port, B_CMP_6_port, B_CMP_5_port, 
      B_CMP_4_port, B_CMP_3_port, B_CMP_2_port, B_CMP_1_port, B_CMP_0_port, 
      A_SHF_31_port, A_SHF_30_port, A_SHF_29_port, A_SHF_28_port, A_SHF_27_port
      , A_SHF_26_port, A_SHF_25_port, A_SHF_24_port, A_SHF_23_port, 
      A_SHF_22_port, A_SHF_21_port, A_SHF_20_port, A_SHF_19_port, A_SHF_18_port
      , A_SHF_17_port, A_SHF_16_port, A_SHF_15_port, A_SHF_14_port, 
      A_SHF_13_port, A_SHF_12_port, A_SHF_11_port, A_SHF_10_port, A_SHF_9_port,
      A_SHF_8_port, A_SHF_7_port, A_SHF_6_port, A_SHF_5_port, A_SHF_4_port, 
      A_SHF_3_port, A_SHF_2_port, A_SHF_1_port, A_SHF_0_port, B_SHF_31_port, 
      B_SHF_30_port, B_SHF_29_port, B_SHF_28_port, B_SHF_27_port, B_SHF_26_port
      , B_SHF_25_port, B_SHF_24_port, B_SHF_23_port, B_SHF_22_port, 
      B_SHF_21_port, B_SHF_20_port, B_SHF_19_port, B_SHF_18_port, B_SHF_17_port
      , B_SHF_16_port, B_SHF_15_port, B_SHF_14_port, B_SHF_13_port, 
      B_SHF_12_port, B_SHF_11_port, B_SHF_10_port, B_SHF_9_port, B_SHF_8_port, 
      B_SHF_7_port, B_SHF_6_port, B_SHF_5_port, B_SHF_4_port, B_SHF_3_port, 
      B_SHF_2_port, B_SHF_1_port, B_SHF_0_port, A_ADD_31_port, A_ADD_30_port, 
      A_ADD_29_port, A_ADD_28_port, A_ADD_27_port, A_ADD_26_port, A_ADD_25_port
      , A_ADD_24_port, A_ADD_23_port, A_ADD_22_port, A_ADD_21_port, 
      A_ADD_20_port, A_ADD_19_port, A_ADD_18_port, A_ADD_17_port, A_ADD_16_port
      , A_ADD_15_port, A_ADD_14_port, A_ADD_13_port, A_ADD_12_port, 
      A_ADD_11_port, A_ADD_10_port, A_ADD_9_port, A_ADD_8_port, A_ADD_7_port, 
      A_ADD_6_port, A_ADD_5_port, A_ADD_4_port, A_ADD_3_port, A_ADD_2_port, 
      A_ADD_1_port, A_ADD_0_port, B_ADD_31_port, B_ADD_30_port, B_ADD_29_port, 
      B_ADD_28_port, B_ADD_27_port, B_ADD_26_port, B_ADD_25_port, B_ADD_24_port
      , B_ADD_23_port, B_ADD_22_port, B_ADD_21_port, B_ADD_20_port, 
      B_ADD_19_port, B_ADD_18_port, B_ADD_17_port, B_ADD_16_port, B_ADD_15_port
      , B_ADD_14_port, B_ADD_13_port, B_ADD_12_port, B_ADD_11_port, 
      B_ADD_10_port, B_ADD_9_port, B_ADD_8_port, B_ADD_7_port, B_ADD_6_port, 
      B_ADD_5_port, B_ADD_4_port, B_ADD_3_port, B_ADD_2_port, B_ADD_1_port, 
      B_ADD_0_port, A_MUL_15_port, A_MUL_14_port, A_MUL_13_port, A_MUL_12_port,
      A_MUL_11_port, A_MUL_10_port, A_MUL_9_port, A_MUL_8_port, A_MUL_7_port, 
      A_MUL_6_port, A_MUL_5_port, A_MUL_4_port, A_MUL_3_port, A_MUL_2_port, 
      A_MUL_1_port, A_MUL_0_port, B_MUL_15_port, B_MUL_14_port, B_MUL_13_port, 
      B_MUL_12_port, B_MUL_11_port, B_MUL_10_port, B_MUL_9_port, B_MUL_8_port, 
      B_MUL_7_port, B_MUL_6_port, B_MUL_5_port, B_MUL_4_port, B_MUL_3_port, 
      B_MUL_2_port, B_MUL_1_port, B_MUL_0_port, LOGIC_ARITH, LEFT_RIGHT, 
      OPSel_1_port, OPSel_0_port, ADD_SUB, LOGIC_RES_31_port, LOGIC_RES_30_port
      , LOGIC_RES_29_port, LOGIC_RES_28_port, LOGIC_RES_27_port, 
      LOGIC_RES_26_port, LOGIC_RES_25_port, LOGIC_RES_24_port, 
      LOGIC_RES_23_port, LOGIC_RES_22_port, LOGIC_RES_21_port, 
      LOGIC_RES_20_port, LOGIC_RES_19_port, LOGIC_RES_18_port, 
      LOGIC_RES_17_port, LOGIC_RES_16_port, LOGIC_RES_15_port, 
      LOGIC_RES_14_port, LOGIC_RES_13_port, LOGIC_RES_12_port, 
      LOGIC_RES_11_port, LOGIC_RES_10_port, LOGIC_RES_9_port, LOGIC_RES_8_port,
      LOGIC_RES_7_port, LOGIC_RES_6_port, LOGIC_RES_5_port, LOGIC_RES_4_port, 
      LOGIC_RES_3_port, LOGIC_RES_2_port, LOGIC_RES_1_port, LOGIC_RES_0_port, 
      COMP_RES_31_port, COMP_RES_30_port, COMP_RES_29_port, COMP_RES_28_port, 
      COMP_RES_27_port, COMP_RES_26_port, COMP_RES_25_port, COMP_RES_24_port, 
      COMP_RES_23_port, COMP_RES_22_port, COMP_RES_21_port, COMP_RES_20_port, 
      COMP_RES_19_port, COMP_RES_18_port, COMP_RES_17_port, COMP_RES_16_port, 
      COMP_RES_15_port, COMP_RES_14_port, COMP_RES_13_port, COMP_RES_12_port, 
      COMP_RES_11_port, COMP_RES_10_port, COMP_RES_9_port, COMP_RES_8_port, 
      COMP_RES_7_port, COMP_RES_6_port, COMP_RES_5_port, COMP_RES_4_port, 
      COMP_RES_3_port, COMP_RES_2_port, COMP_RES_1_port, COMP_RES_0_port, 
      SHIFT_RES_31_port, SHIFT_RES_30_port, SHIFT_RES_29_port, 
      SHIFT_RES_28_port, SHIFT_RES_27_port, SHIFT_RES_26_port, 
      SHIFT_RES_25_port, SHIFT_RES_24_port, SHIFT_RES_23_port, 
      SHIFT_RES_22_port, SHIFT_RES_21_port, SHIFT_RES_20_port, 
      SHIFT_RES_19_port, SHIFT_RES_18_port, SHIFT_RES_17_port, 
      SHIFT_RES_16_port, SHIFT_RES_15_port, SHIFT_RES_14_port, 
      SHIFT_RES_13_port, SHIFT_RES_12_port, SHIFT_RES_11_port, 
      SHIFT_RES_10_port, SHIFT_RES_9_port, SHIFT_RES_8_port, SHIFT_RES_7_port, 
      SHIFT_RES_6_port, SHIFT_RES_5_port, SHIFT_RES_4_port, SHIFT_RES_3_port, 
      SHIFT_RES_2_port, SHIFT_RES_1_port, SHIFT_RES_0_port, ADD_SUB_RES_31_port
      , ADD_SUB_RES_30_port, ADD_SUB_RES_29_port, ADD_SUB_RES_28_port, 
      ADD_SUB_RES_27_port, ADD_SUB_RES_26_port, ADD_SUB_RES_25_port, 
      ADD_SUB_RES_24_port, ADD_SUB_RES_23_port, ADD_SUB_RES_22_port, 
      ADD_SUB_RES_21_port, ADD_SUB_RES_20_port, ADD_SUB_RES_19_port, 
      ADD_SUB_RES_18_port, ADD_SUB_RES_17_port, ADD_SUB_RES_16_port, 
      ADD_SUB_RES_15_port, ADD_SUB_RES_14_port, ADD_SUB_RES_13_port, 
      ADD_SUB_RES_12_port, ADD_SUB_RES_11_port, ADD_SUB_RES_10_port, 
      ADD_SUB_RES_9_port, ADD_SUB_RES_8_port, ADD_SUB_RES_7_port, 
      ADD_SUB_RES_6_port, ADD_SUB_RES_5_port, ADD_SUB_RES_4_port, 
      ADD_SUB_RES_3_port, ADD_SUB_RES_2_port, ADD_SUB_RES_1_port, 
      ADD_SUB_RES_0_port, MUL_RES_31_port, MUL_RES_30_port, MUL_RES_29_port, 
      MUL_RES_28_port, MUL_RES_27_port, MUL_RES_26_port, MUL_RES_25_port, 
      MUL_RES_24_port, MUL_RES_23_port, MUL_RES_22_port, MUL_RES_21_port, 
      MUL_RES_20_port, MUL_RES_19_port, MUL_RES_18_port, MUL_RES_17_port, 
      MUL_RES_16_port, MUL_RES_15_port, MUL_RES_14_port, MUL_RES_13_port, 
      MUL_RES_12_port, MUL_RES_11_port, MUL_RES_10_port, MUL_RES_9_port, 
      MUL_RES_8_port, MUL_RES_7_port, MUL_RES_6_port, MUL_RES_5_port, 
      MUL_RES_4_port, MUL_RES_3_port, MUL_RES_2_port, MUL_RES_1_port, 
      MUL_RES_0_port, sig_intraMux_31_port, sig_intraMux_30_port, 
      sig_intraMux_29_port, sig_intraMux_28_port, sig_intraMux_27_port, 
      sig_intraMux_26_port, sig_intraMux_25_port, sig_intraMux_24_port, 
      sig_intraMux_23_port, sig_intraMux_22_port, sig_intraMux_21_port, 
      sig_intraMux_20_port, sig_intraMux_19_port, sig_intraMux_18_port, 
      sig_intraMux_17_port, sig_intraMux_16_port, sig_intraMux_15_port, 
      sig_intraMux_14_port, sig_intraMux_13_port, sig_intraMux_12_port, 
      sig_intraMux_11_port, sig_intraMux_10_port, sig_intraMux_9_port, 
      sig_intraMux_8_port, sig_intraMux_7_port, sig_intraMux_6_port, 
      sig_intraMux_5_port, sig_intraMux_4_port, sig_intraMux_3_port, 
      sig_intraMux_2_port, sig_intraMux_1_port, sig_intraMux_0_port, 
      sig_ALU_RES_31_port, sig_ALU_RES_30_port, sig_ALU_RES_29_port, 
      sig_ALU_RES_28_port, sig_ALU_RES_27_port, sig_ALU_RES_26_port, 
      sig_ALU_RES_25_port, sig_ALU_RES_24_port, sig_ALU_RES_23_port, 
      sig_ALU_RES_22_port, sig_ALU_RES_21_port, sig_ALU_RES_20_port, 
      sig_ALU_RES_19_port, sig_ALU_RES_18_port, sig_ALU_RES_17_port, 
      sig_ALU_RES_16_port, sig_ALU_RES_15_port, sig_ALU_RES_14_port, 
      sig_ALU_RES_13_port, sig_ALU_RES_12_port, sig_ALU_RES_11_port, 
      sig_ALU_RES_10_port, sig_ALU_RES_9_port, sig_ALU_RES_8_port, 
      sig_ALU_RES_7_port, sig_ALU_RES_6_port, sig_ALU_RES_5_port, 
      sig_ALU_RES_4_port, sig_ALU_RES_3_port, sig_ALU_RES_2_port, 
      sig_ALU_RES_1_port, sig_ALU_RES_0_port, n78, n79, n80, n81, n82, n83, n84
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n85, n86, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n_1165, n_1166, n_1167, 
      n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, 
      n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, 
      n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, 
      n_1195, n_1196 : std_logic;

begin
   
   X_Logic0_port <= '0';
   U227 : OAI22_X2 port map( A1 => n195, A2 => n39, B1 => n45, B2 => n72, ZN =>
                           A_SHF_31_port);
   U257 : NOR2_X2 port map( A1 => n86, A2 => n30, ZN => A_MUL_9_port);
   U258 : NOR2_X2 port map( A1 => n85, A2 => n30, ZN => A_MUL_8_port);
   U259 : NOR2_X2 port map( A1 => n77, A2 => n30, ZN => A_MUL_7_port);
   U260 : NOR2_X2 port map( A1 => n76, A2 => n30, ZN => A_MUL_6_port);
   U261 : NOR2_X2 port map( A1 => n75, A2 => n29, ZN => A_MUL_5_port);
   U262 : NOR2_X2 port map( A1 => n74, A2 => n29, ZN => A_MUL_4_port);
   U263 : NOR2_X2 port map( A1 => n73, A2 => n29, ZN => A_MUL_3_port);
   U264 : NOR2_X2 port map( A1 => n70, A2 => n29, ZN => A_MUL_2_port);
   U265 : NOR2_X2 port map( A1 => n59, A2 => n29, ZN => A_MUL_1_port);
   U267 : NOR2_X2 port map( A1 => n53, A2 => n29, ZN => A_MUL_14_port);
   U268 : NOR2_X2 port map( A1 => n52, A2 => n29, ZN => A_MUL_13_port);
   U269 : NOR2_X2 port map( A1 => n51, A2 => n29, ZN => A_MUL_12_port);
   U270 : NOR2_X2 port map( A1 => n50, A2 => n29, ZN => A_MUL_11_port);
   U271 : NOR2_X2 port map( A1 => n49, A2 => n29, ZN => A_MUL_10_port);
   U272 : NOR2_X2 port map( A1 => n48, A2 => n29, ZN => A_MUL_0_port);
   U427 : NAND3_X1 port map( A1 => n212, A2 => n211, A3 => n80, ZN => n79);
   U428 : NAND3_X1 port map( A1 => n47, A2 => n41, A3 => n38, ZN => 
                           select_type_sig_1_port);
   U429 : NAND3_X1 port map( A1 => n84, A2 => n7, A3 => n38, ZN => 
                           select_type_sig_0_port);
   U430 : NAND3_X1 port map( A1 => ALU_OPC(1), A2 => n212, A3 => n156, ZN => 
                           n84);
   U431 : NAND3_X1 port map( A1 => ALU_OPC(4), A2 => ALU_OPC(1), A3 => n156, ZN
                           => n158);
   U432 : NAND3_X1 port map( A1 => ALU_OPC(0), A2 => ALU_OPC(3), A3 => n162, ZN
                           => n82);
   U434 : NAND3_X1 port map( A1 => n211, A2 => n209, A3 => ALU_OPC(0), ZN => 
                           n164);
   U436 : NAND3_X1 port map( A1 => n209, A2 => n204, A3 => n211, ZN => n170);
   Comp : comparator_NBIT32 port map( A(31) => A_CMP_31_port, A(30) => 
                           A_CMP_30_port, A(29) => A_CMP_29_port, A(28) => 
                           A_CMP_28_port, A(27) => A_CMP_27_port, A(26) => 
                           A_CMP_26_port, A(25) => A_CMP_25_port, A(24) => 
                           A_CMP_24_port, A(23) => A_CMP_23_port, A(22) => 
                           A_CMP_22_port, A(21) => A_CMP_21_port, A(20) => 
                           A_CMP_20_port, A(19) => A_CMP_19_port, A(18) => 
                           A_CMP_18_port, A(17) => A_CMP_17_port, A(16) => 
                           A_CMP_16_port, A(15) => A_CMP_15_port, A(14) => 
                           A_CMP_14_port, A(13) => A_CMP_13_port, A(12) => 
                           A_CMP_12_port, A(11) => A_CMP_11_port, A(10) => 
                           A_CMP_10_port, A(9) => A_CMP_9_port, A(8) => 
                           A_CMP_8_port, A(7) => A_CMP_7_port, A(6) => 
                           A_CMP_6_port, A(5) => A_CMP_5_port, A(4) => 
                           A_CMP_4_port, A(3) => A_CMP_3_port, A(2) => 
                           A_CMP_2_port, A(1) => A_CMP_1_port, A(0) => 
                           A_CMP_0_port, B(31) => B_CMP_31_port, B(30) => 
                           B_CMP_30_port, B(29) => B_CMP_29_port, B(28) => 
                           B_CMP_28_port, B(27) => B_CMP_27_port, B(26) => 
                           B_CMP_26_port, B(25) => B_CMP_25_port, B(24) => 
                           B_CMP_24_port, B(23) => B_CMP_23_port, B(22) => 
                           B_CMP_22_port, B(21) => B_CMP_21_port, B(20) => 
                           B_CMP_20_port, B(19) => B_CMP_19_port, B(18) => 
                           B_CMP_18_port, B(17) => B_CMP_17_port, B(16) => 
                           B_CMP_16_port, B(15) => B_CMP_15_port, B(14) => 
                           B_CMP_14_port, B(13) => B_CMP_13_port, B(12) => 
                           B_CMP_12_port, B(11) => B_CMP_11_port, B(10) => 
                           B_CMP_10_port, B(9) => B_CMP_9_port, B(8) => 
                           B_CMP_8_port, B(7) => B_CMP_7_port, B(6) => 
                           B_CMP_6_port, B(5) => B_CMP_5_port, B(4) => 
                           B_CMP_4_port, B(3) => B_CMP_3_port, B(2) => 
                           B_CMP_2_port, B(1) => B_CMP_1_port, B(0) => 
                           B_CMP_0_port, OPSel(0) => n206, OPSel(1) => 
                           OPSel_1_port, OPSel(2) => OPSel_0_port, RES(31) => 
                           n_1165, RES(30) => n_1166, RES(29) => n_1167, 
                           RES(28) => n_1168, RES(27) => n_1169, RES(26) => 
                           n_1170, RES(25) => n_1171, RES(24) => n_1172, 
                           RES(23) => n_1173, RES(22) => n_1174, RES(21) => 
                           n_1175, RES(20) => n_1176, RES(19) => n_1177, 
                           RES(18) => n_1178, RES(17) => n_1179, RES(16) => 
                           n_1180, RES(15) => n_1181, RES(14) => n_1182, 
                           RES(13) => n_1183, RES(12) => n_1184, RES(11) => 
                           n_1185, RES(10) => n_1186, RES(9) => n_1187, RES(8) 
                           => n_1188, RES(7) => n_1189, RES(6) => n_1190, 
                           RES(5) => n_1191, RES(4) => n_1192, RES(3) => n_1193
                           , RES(2) => n_1194, RES(1) => n_1195, RES(0) => 
                           COMP_RES_0_port);
   Shift : shifter_NBIT32 port map( A(31) => A_SHF_31_port, A(30) => 
                           A_SHF_30_port, A(29) => A_SHF_29_port, A(28) => 
                           A_SHF_28_port, A(27) => A_SHF_27_port, A(26) => 
                           A_SHF_26_port, A(25) => A_SHF_25_port, A(24) => 
                           A_SHF_24_port, A(23) => A_SHF_23_port, A(22) => 
                           A_SHF_22_port, A(21) => A_SHF_21_port, A(20) => 
                           A_SHF_20_port, A(19) => A_SHF_19_port, A(18) => 
                           A_SHF_18_port, A(17) => A_SHF_17_port, A(16) => 
                           A_SHF_16_port, A(15) => A_SHF_15_port, A(14) => 
                           A_SHF_14_port, A(13) => A_SHF_13_port, A(12) => 
                           A_SHF_12_port, A(11) => A_SHF_11_port, A(10) => 
                           A_SHF_10_port, A(9) => A_SHF_9_port, A(8) => 
                           A_SHF_8_port, A(7) => A_SHF_7_port, A(6) => 
                           A_SHF_6_port, A(5) => A_SHF_5_port, A(4) => 
                           A_SHF_4_port, A(3) => A_SHF_3_port, A(2) => 
                           A_SHF_2_port, A(1) => A_SHF_1_port, A(0) => 
                           A_SHF_0_port, B(31) => B_SHF_31_port, B(30) => 
                           B_SHF_30_port, B(29) => B_SHF_29_port, B(28) => 
                           B_SHF_28_port, B(27) => B_SHF_27_port, B(26) => 
                           B_SHF_26_port, B(25) => B_SHF_25_port, B(24) => 
                           B_SHF_24_port, B(23) => B_SHF_23_port, B(22) => 
                           B_SHF_22_port, B(21) => B_SHF_21_port, B(20) => 
                           B_SHF_20_port, B(19) => B_SHF_19_port, B(18) => 
                           B_SHF_18_port, B(17) => B_SHF_17_port, B(16) => 
                           B_SHF_16_port, B(15) => B_SHF_15_port, B(14) => 
                           B_SHF_14_port, B(13) => B_SHF_13_port, B(12) => 
                           B_SHF_12_port, B(11) => B_SHF_11_port, B(10) => 
                           B_SHF_10_port, B(9) => B_SHF_9_port, B(8) => 
                           B_SHF_8_port, B(7) => B_SHF_7_port, B(6) => 
                           B_SHF_6_port, B(5) => B_SHF_5_port, B(4) => 
                           B_SHF_4_port, B(3) => B_SHF_3_port, B(2) => 
                           B_SHF_2_port, B(1) => B_SHF_1_port, B(0) => 
                           B_SHF_0_port, LOGIC_ARITH => LOGIC_ARITH, LEFT_RIGHT
                           => LEFT_RIGHT, RES(31) => SHIFT_RES_31_port, RES(30)
                           => SHIFT_RES_30_port, RES(29) => SHIFT_RES_29_port, 
                           RES(28) => SHIFT_RES_28_port, RES(27) => 
                           SHIFT_RES_27_port, RES(26) => SHIFT_RES_26_port, 
                           RES(25) => SHIFT_RES_25_port, RES(24) => 
                           SHIFT_RES_24_port, RES(23) => SHIFT_RES_23_port, 
                           RES(22) => SHIFT_RES_22_port, RES(21) => 
                           SHIFT_RES_21_port, RES(20) => SHIFT_RES_20_port, 
                           RES(19) => SHIFT_RES_19_port, RES(18) => 
                           SHIFT_RES_18_port, RES(17) => SHIFT_RES_17_port, 
                           RES(16) => SHIFT_RES_16_port, RES(15) => 
                           SHIFT_RES_15_port, RES(14) => SHIFT_RES_14_port, 
                           RES(13) => SHIFT_RES_13_port, RES(12) => 
                           SHIFT_RES_12_port, RES(11) => SHIFT_RES_11_port, 
                           RES(10) => SHIFT_RES_10_port, RES(9) => 
                           SHIFT_RES_9_port, RES(8) => SHIFT_RES_8_port, RES(7)
                           => SHIFT_RES_7_port, RES(6) => SHIFT_RES_6_port, 
                           RES(5) => SHIFT_RES_5_port, RES(4) => 
                           SHIFT_RES_4_port, RES(3) => SHIFT_RES_3_port, RES(2)
                           => SHIFT_RES_2_port, RES(1) => SHIFT_RES_1_port, 
                           RES(0) => SHIFT_RES_0_port);
   Add_Sub_unit : P4Adder_NBIT32 port map( A(31) => A_ADD_31_port, A(30) => 
                           A_ADD_30_port, A(29) => A_ADD_29_port, A(28) => 
                           A_ADD_28_port, A(27) => A_ADD_27_port, A(26) => 
                           A_ADD_26_port, A(25) => A_ADD_25_port, A(24) => 
                           A_ADD_24_port, A(23) => A_ADD_23_port, A(22) => 
                           A_ADD_22_port, A(21) => A_ADD_21_port, A(20) => 
                           A_ADD_20_port, A(19) => A_ADD_19_port, A(18) => 
                           A_ADD_18_port, A(17) => A_ADD_17_port, A(16) => 
                           A_ADD_16_port, A(15) => A_ADD_15_port, A(14) => 
                           A_ADD_14_port, A(13) => A_ADD_13_port, A(12) => 
                           A_ADD_12_port, A(11) => A_ADD_11_port, A(10) => 
                           A_ADD_10_port, A(9) => A_ADD_9_port, A(8) => 
                           A_ADD_8_port, A(7) => A_ADD_7_port, A(6) => 
                           A_ADD_6_port, A(5) => A_ADD_5_port, A(4) => 
                           A_ADD_4_port, A(3) => A_ADD_3_port, A(2) => 
                           A_ADD_2_port, A(1) => A_ADD_1_port, A(0) => 
                           A_ADD_0_port, B(31) => B_ADD_31_port, B(30) => 
                           B_ADD_30_port, B(29) => B_ADD_29_port, B(28) => 
                           B_ADD_28_port, B(27) => B_ADD_27_port, B(26) => 
                           B_ADD_26_port, B(25) => B_ADD_25_port, B(24) => 
                           B_ADD_24_port, B(23) => B_ADD_23_port, B(22) => 
                           B_ADD_22_port, B(21) => B_ADD_21_port, B(20) => 
                           B_ADD_20_port, B(19) => B_ADD_19_port, B(18) => 
                           B_ADD_18_port, B(17) => B_ADD_17_port, B(16) => 
                           B_ADD_16_port, B(15) => B_ADD_15_port, B(14) => 
                           B_ADD_14_port, B(13) => B_ADD_13_port, B(12) => 
                           B_ADD_12_port, B(11) => B_ADD_11_port, B(10) => 
                           B_ADD_10_port, B(9) => B_ADD_9_port, B(8) => 
                           B_ADD_8_port, B(7) => B_ADD_7_port, B(6) => 
                           B_ADD_6_port, B(5) => B_ADD_5_port, B(4) => 
                           B_ADD_4_port, B(3) => B_ADD_3_port, B(2) => 
                           B_ADD_2_port, B(1) => B_ADD_1_port, B(0) => 
                           B_ADD_0_port, Cin => ADD_SUB, S(31) => 
                           ADD_SUB_RES_31_port, S(30) => ADD_SUB_RES_30_port, 
                           S(29) => ADD_SUB_RES_29_port, S(28) => 
                           ADD_SUB_RES_28_port, S(27) => ADD_SUB_RES_27_port, 
                           S(26) => ADD_SUB_RES_26_port, S(25) => 
                           ADD_SUB_RES_25_port, S(24) => ADD_SUB_RES_24_port, 
                           S(23) => ADD_SUB_RES_23_port, S(22) => 
                           ADD_SUB_RES_22_port, S(21) => ADD_SUB_RES_21_port, 
                           S(20) => ADD_SUB_RES_20_port, S(19) => 
                           ADD_SUB_RES_19_port, S(18) => ADD_SUB_RES_18_port, 
                           S(17) => ADD_SUB_RES_17_port, S(16) => 
                           ADD_SUB_RES_16_port, S(15) => ADD_SUB_RES_15_port, 
                           S(14) => ADD_SUB_RES_14_port, S(13) => 
                           ADD_SUB_RES_13_port, S(12) => ADD_SUB_RES_12_port, 
                           S(11) => ADD_SUB_RES_11_port, S(10) => 
                           ADD_SUB_RES_10_port, S(9) => ADD_SUB_RES_9_port, 
                           S(8) => ADD_SUB_RES_8_port, S(7) => 
                           ADD_SUB_RES_7_port, S(6) => ADD_SUB_RES_6_port, S(5)
                           => ADD_SUB_RES_5_port, S(4) => ADD_SUB_RES_4_port, 
                           S(3) => ADD_SUB_RES_3_port, S(2) => 
                           ADD_SUB_RES_2_port, S(1) => ADD_SUB_RES_1_port, S(0)
                           => ADD_SUB_RES_0_port, Cout => n_1196);
   Booth_mul : BOOTHMUL_numBit16 port map( A(15) => A_MUL_15_port, A(14) => 
                           A_MUL_14_port, A(13) => A_MUL_13_port, A(12) => 
                           A_MUL_12_port, A(11) => A_MUL_11_port, A(10) => 
                           A_MUL_10_port, A(9) => A_MUL_9_port, A(8) => 
                           A_MUL_8_port, A(7) => A_MUL_7_port, A(6) => 
                           A_MUL_6_port, A(5) => A_MUL_5_port, A(4) => 
                           A_MUL_4_port, A(3) => A_MUL_3_port, A(2) => 
                           A_MUL_2_port, A(1) => A_MUL_1_port, A(0) => 
                           A_MUL_0_port, B(15) => B_MUL_15_port, B(14) => 
                           B_MUL_14_port, B(13) => B_MUL_13_port, B(12) => 
                           B_MUL_12_port, B(11) => B_MUL_11_port, B(10) => 
                           B_MUL_10_port, B(9) => B_MUL_9_port, B(8) => 
                           B_MUL_8_port, B(7) => B_MUL_7_port, B(6) => 
                           B_MUL_6_port, B(5) => B_MUL_5_port, B(4) => 
                           B_MUL_4_port, B(3) => B_MUL_3_port, B(2) => 
                           B_MUL_2_port, B(1) => B_MUL_1_port, B(0) => 
                           B_MUL_0_port, P(31) => MUL_RES_31_port, P(30) => 
                           MUL_RES_30_port, P(29) => MUL_RES_29_port, P(28) => 
                           MUL_RES_28_port, P(27) => MUL_RES_27_port, P(26) => 
                           MUL_RES_26_port, P(25) => MUL_RES_25_port, P(24) => 
                           MUL_RES_24_port, P(23) => MUL_RES_23_port, P(22) => 
                           MUL_RES_22_port, P(21) => MUL_RES_21_port, P(20) => 
                           MUL_RES_20_port, P(19) => MUL_RES_19_port, P(18) => 
                           MUL_RES_18_port, P(17) => MUL_RES_17_port, P(16) => 
                           MUL_RES_16_port, P(15) => MUL_RES_15_port, P(14) => 
                           MUL_RES_14_port, P(13) => MUL_RES_13_port, P(12) => 
                           MUL_RES_12_port, P(11) => MUL_RES_11_port, P(10) => 
                           MUL_RES_10_port, P(9) => MUL_RES_9_port, P(8) => 
                           MUL_RES_8_port, P(7) => MUL_RES_7_port, P(6) => 
                           MUL_RES_6_port, P(5) => MUL_RES_5_port, P(4) => 
                           MUL_RES_4_port, P(3) => MUL_RES_3_port, P(2) => 
                           MUL_RES_2_port, P(1) => MUL_RES_1_port, P(0) => 
                           MUL_RES_0_port);
   Res_mux : mux41_NBIT32_1 port map( A(31) => ADD_SUB_RES_31_port, A(30) => 
                           ADD_SUB_RES_30_port, A(29) => ADD_SUB_RES_29_port, 
                           A(28) => ADD_SUB_RES_28_port, A(27) => 
                           ADD_SUB_RES_27_port, A(26) => ADD_SUB_RES_26_port, 
                           A(25) => ADD_SUB_RES_25_port, A(24) => 
                           ADD_SUB_RES_24_port, A(23) => ADD_SUB_RES_23_port, 
                           A(22) => ADD_SUB_RES_22_port, A(21) => 
                           ADD_SUB_RES_21_port, A(20) => ADD_SUB_RES_20_port, 
                           A(19) => ADD_SUB_RES_19_port, A(18) => 
                           ADD_SUB_RES_18_port, A(17) => ADD_SUB_RES_17_port, 
                           A(16) => ADD_SUB_RES_16_port, A(15) => 
                           ADD_SUB_RES_15_port, A(14) => ADD_SUB_RES_14_port, 
                           A(13) => ADD_SUB_RES_13_port, A(12) => 
                           ADD_SUB_RES_12_port, A(11) => ADD_SUB_RES_11_port, 
                           A(10) => ADD_SUB_RES_10_port, A(9) => 
                           ADD_SUB_RES_9_port, A(8) => ADD_SUB_RES_8_port, A(7)
                           => ADD_SUB_RES_7_port, A(6) => ADD_SUB_RES_6_port, 
                           A(5) => ADD_SUB_RES_5_port, A(4) => 
                           ADD_SUB_RES_4_port, A(3) => ADD_SUB_RES_3_port, A(2)
                           => ADD_SUB_RES_2_port, A(1) => ADD_SUB_RES_1_port, 
                           A(0) => ADD_SUB_RES_0_port, B(31) => 
                           LOGIC_RES_31_port, B(30) => LOGIC_RES_30_port, B(29)
                           => LOGIC_RES_29_port, B(28) => LOGIC_RES_28_port, 
                           B(27) => LOGIC_RES_27_port, B(26) => 
                           LOGIC_RES_26_port, B(25) => LOGIC_RES_25_port, B(24)
                           => LOGIC_RES_24_port, B(23) => LOGIC_RES_23_port, 
                           B(22) => LOGIC_RES_22_port, B(21) => 
                           LOGIC_RES_21_port, B(20) => LOGIC_RES_20_port, B(19)
                           => LOGIC_RES_19_port, B(18) => LOGIC_RES_18_port, 
                           B(17) => LOGIC_RES_17_port, B(16) => 
                           LOGIC_RES_16_port, B(15) => LOGIC_RES_15_port, B(14)
                           => LOGIC_RES_14_port, B(13) => LOGIC_RES_13_port, 
                           B(12) => LOGIC_RES_12_port, B(11) => 
                           LOGIC_RES_11_port, B(10) => LOGIC_RES_10_port, B(9) 
                           => LOGIC_RES_9_port, B(8) => LOGIC_RES_8_port, B(7) 
                           => LOGIC_RES_7_port, B(6) => LOGIC_RES_6_port, B(5) 
                           => LOGIC_RES_5_port, B(4) => LOGIC_RES_4_port, B(3) 
                           => LOGIC_RES_3_port, B(2) => LOGIC_RES_2_port, B(1) 
                           => LOGIC_RES_1_port, B(0) => LOGIC_RES_0_port, C(31)
                           => SHIFT_RES_31_port, C(30) => SHIFT_RES_30_port, 
                           C(29) => SHIFT_RES_29_port, C(28) => 
                           SHIFT_RES_28_port, C(27) => SHIFT_RES_27_port, C(26)
                           => SHIFT_RES_26_port, C(25) => SHIFT_RES_25_port, 
                           C(24) => SHIFT_RES_24_port, C(23) => 
                           SHIFT_RES_23_port, C(22) => SHIFT_RES_22_port, C(21)
                           => SHIFT_RES_21_port, C(20) => SHIFT_RES_20_port, 
                           C(19) => SHIFT_RES_19_port, C(18) => 
                           SHIFT_RES_18_port, C(17) => SHIFT_RES_17_port, C(16)
                           => SHIFT_RES_16_port, C(15) => SHIFT_RES_15_port, 
                           C(14) => SHIFT_RES_14_port, C(13) => 
                           SHIFT_RES_13_port, C(12) => SHIFT_RES_12_port, C(11)
                           => SHIFT_RES_11_port, C(10) => SHIFT_RES_10_port, 
                           C(9) => SHIFT_RES_9_port, C(8) => SHIFT_RES_8_port, 
                           C(7) => SHIFT_RES_7_port, C(6) => SHIFT_RES_6_port, 
                           C(5) => SHIFT_RES_5_port, C(4) => SHIFT_RES_4_port, 
                           C(3) => SHIFT_RES_3_port, C(2) => SHIFT_RES_2_port, 
                           C(1) => SHIFT_RES_1_port, C(0) => SHIFT_RES_0_port, 
                           D(31) => COMP_RES_31_port, D(30) => COMP_RES_30_port
                           , D(29) => COMP_RES_29_port, D(28) => 
                           COMP_RES_28_port, D(27) => COMP_RES_27_port, D(26) 
                           => COMP_RES_26_port, D(25) => COMP_RES_25_port, 
                           D(24) => COMP_RES_24_port, D(23) => COMP_RES_23_port
                           , D(22) => COMP_RES_22_port, D(21) => 
                           COMP_RES_21_port, D(20) => COMP_RES_20_port, D(19) 
                           => COMP_RES_19_port, D(18) => COMP_RES_18_port, 
                           D(17) => COMP_RES_17_port, D(16) => COMP_RES_16_port
                           , D(15) => COMP_RES_15_port, D(14) => 
                           COMP_RES_14_port, D(13) => COMP_RES_13_port, D(12) 
                           => COMP_RES_12_port, D(11) => COMP_RES_11_port, 
                           D(10) => COMP_RES_10_port, D(9) => COMP_RES_9_port, 
                           D(8) => COMP_RES_8_port, D(7) => COMP_RES_7_port, 
                           D(6) => COMP_RES_6_port, D(5) => COMP_RES_5_port, 
                           D(4) => COMP_RES_4_port, D(3) => COMP_RES_3_port, 
                           D(2) => COMP_RES_2_port, D(1) => COMP_RES_1_port, 
                           D(0) => COMP_RES_0_port, S(1) => 
                           select_type_sig_1_port, S(0) => 
                           select_type_sig_0_port, Z(31) => 
                           sig_intraMux_31_port, Z(30) => sig_intraMux_30_port,
                           Z(29) => sig_intraMux_29_port, Z(28) => 
                           sig_intraMux_28_port, Z(27) => sig_intraMux_27_port,
                           Z(26) => sig_intraMux_26_port, Z(25) => 
                           sig_intraMux_25_port, Z(24) => sig_intraMux_24_port,
                           Z(23) => sig_intraMux_23_port, Z(22) => 
                           sig_intraMux_22_port, Z(21) => sig_intraMux_21_port,
                           Z(20) => sig_intraMux_20_port, Z(19) => 
                           sig_intraMux_19_port, Z(18) => sig_intraMux_18_port,
                           Z(17) => sig_intraMux_17_port, Z(16) => 
                           sig_intraMux_16_port, Z(15) => sig_intraMux_15_port,
                           Z(14) => sig_intraMux_14_port, Z(13) => 
                           sig_intraMux_13_port, Z(12) => sig_intraMux_12_port,
                           Z(11) => sig_intraMux_11_port, Z(10) => 
                           sig_intraMux_10_port, Z(9) => sig_intraMux_9_port, 
                           Z(8) => sig_intraMux_8_port, Z(7) => 
                           sig_intraMux_7_port, Z(6) => sig_intraMux_6_port, 
                           Z(5) => sig_intraMux_5_port, Z(4) => 
                           sig_intraMux_4_port, Z(3) => sig_intraMux_3_port, 
                           Z(2) => sig_intraMux_2_port, Z(1) => 
                           sig_intraMux_1_port, Z(0) => sig_intraMux_0_port);
   Mul_mux : mux21_NBIT32_2 port map( A(31) => sig_intraMux_31_port, A(30) => 
                           sig_intraMux_30_port, A(29) => sig_intraMux_29_port,
                           A(28) => sig_intraMux_28_port, A(27) => 
                           sig_intraMux_27_port, A(26) => sig_intraMux_26_port,
                           A(25) => sig_intraMux_25_port, A(24) => 
                           sig_intraMux_24_port, A(23) => sig_intraMux_23_port,
                           A(22) => sig_intraMux_22_port, A(21) => 
                           sig_intraMux_21_port, A(20) => sig_intraMux_20_port,
                           A(19) => sig_intraMux_19_port, A(18) => 
                           sig_intraMux_18_port, A(17) => sig_intraMux_17_port,
                           A(16) => sig_intraMux_16_port, A(15) => 
                           sig_intraMux_15_port, A(14) => sig_intraMux_14_port,
                           A(13) => sig_intraMux_13_port, A(12) => 
                           sig_intraMux_12_port, A(11) => sig_intraMux_11_port,
                           A(10) => sig_intraMux_10_port, A(9) => 
                           sig_intraMux_9_port, A(8) => sig_intraMux_8_port, 
                           A(7) => sig_intraMux_7_port, A(6) => 
                           sig_intraMux_6_port, A(5) => sig_intraMux_5_port, 
                           A(4) => sig_intraMux_4_port, A(3) => 
                           sig_intraMux_3_port, A(2) => sig_intraMux_2_port, 
                           A(1) => sig_intraMux_1_port, A(0) => 
                           sig_intraMux_0_port, B(31) => MUL_RES_31_port, B(30)
                           => MUL_RES_30_port, B(29) => MUL_RES_29_port, B(28) 
                           => MUL_RES_28_port, B(27) => MUL_RES_27_port, B(26) 
                           => MUL_RES_26_port, B(25) => MUL_RES_25_port, B(24) 
                           => MUL_RES_24_port, B(23) => MUL_RES_23_port, B(22) 
                           => MUL_RES_22_port, B(21) => MUL_RES_21_port, B(20) 
                           => MUL_RES_20_port, B(19) => MUL_RES_19_port, B(18) 
                           => MUL_RES_18_port, B(17) => MUL_RES_17_port, B(16) 
                           => MUL_RES_16_port, B(15) => MUL_RES_15_port, B(14) 
                           => MUL_RES_14_port, B(13) => MUL_RES_13_port, B(12) 
                           => MUL_RES_12_port, B(11) => MUL_RES_11_port, B(10) 
                           => MUL_RES_10_port, B(9) => MUL_RES_9_port, B(8) => 
                           MUL_RES_8_port, B(7) => MUL_RES_7_port, B(6) => 
                           MUL_RES_6_port, B(5) => MUL_RES_5_port, B(4) => 
                           MUL_RES_4_port, B(3) => MUL_RES_3_port, B(2) => 
                           MUL_RES_2_port, B(1) => MUL_RES_1_port, B(0) => 
                           MUL_RES_0_port, S => n1, Z(31) => 
                           sig_ALU_RES_31_port, Z(30) => sig_ALU_RES_30_port, 
                           Z(29) => sig_ALU_RES_29_port, Z(28) => 
                           sig_ALU_RES_28_port, Z(27) => sig_ALU_RES_27_port, 
                           Z(26) => sig_ALU_RES_26_port, Z(25) => 
                           sig_ALU_RES_25_port, Z(24) => sig_ALU_RES_24_port, 
                           Z(23) => sig_ALU_RES_23_port, Z(22) => 
                           sig_ALU_RES_22_port, Z(21) => sig_ALU_RES_21_port, 
                           Z(20) => sig_ALU_RES_20_port, Z(19) => 
                           sig_ALU_RES_19_port, Z(18) => sig_ALU_RES_18_port, 
                           Z(17) => sig_ALU_RES_17_port, Z(16) => 
                           sig_ALU_RES_16_port, Z(15) => sig_ALU_RES_15_port, 
                           Z(14) => sig_ALU_RES_14_port, Z(13) => 
                           sig_ALU_RES_13_port, Z(12) => sig_ALU_RES_12_port, 
                           Z(11) => sig_ALU_RES_11_port, Z(10) => 
                           sig_ALU_RES_10_port, Z(9) => sig_ALU_RES_9_port, 
                           Z(8) => sig_ALU_RES_8_port, Z(7) => 
                           sig_ALU_RES_7_port, Z(6) => sig_ALU_RES_6_port, Z(5)
                           => sig_ALU_RES_5_port, Z(4) => sig_ALU_RES_4_port, 
                           Z(3) => sig_ALU_RES_3_port, Z(2) => 
                           sig_ALU_RES_2_port, Z(1) => sig_ALU_RES_1_port, Z(0)
                           => sig_ALU_RES_0_port);
   Zeros_mux : mux21_NBIT32_1 port map( A(31) => sig_ALU_RES_31_port, A(30) => 
                           sig_ALU_RES_30_port, A(29) => sig_ALU_RES_29_port, 
                           A(28) => sig_ALU_RES_28_port, A(27) => 
                           sig_ALU_RES_27_port, A(26) => sig_ALU_RES_26_port, 
                           A(25) => sig_ALU_RES_25_port, A(24) => 
                           sig_ALU_RES_24_port, A(23) => sig_ALU_RES_23_port, 
                           A(22) => sig_ALU_RES_22_port, A(21) => 
                           sig_ALU_RES_21_port, A(20) => sig_ALU_RES_20_port, 
                           A(19) => sig_ALU_RES_19_port, A(18) => 
                           sig_ALU_RES_18_port, A(17) => sig_ALU_RES_17_port, 
                           A(16) => sig_ALU_RES_16_port, A(15) => 
                           sig_ALU_RES_15_port, A(14) => sig_ALU_RES_14_port, 
                           A(13) => sig_ALU_RES_13_port, A(12) => 
                           sig_ALU_RES_12_port, A(11) => sig_ALU_RES_11_port, 
                           A(10) => sig_ALU_RES_10_port, A(9) => 
                           sig_ALU_RES_9_port, A(8) => sig_ALU_RES_8_port, A(7)
                           => sig_ALU_RES_7_port, A(6) => sig_ALU_RES_6_port, 
                           A(5) => sig_ALU_RES_5_port, A(4) => 
                           sig_ALU_RES_4_port, A(3) => sig_ALU_RES_3_port, A(2)
                           => sig_ALU_RES_2_port, A(1) => sig_ALU_RES_1_port, 
                           A(0) => sig_ALU_RES_0_port, B(31) => X_Logic0_port, 
                           B(30) => X_Logic0_port, B(29) => X_Logic0_port, 
                           B(28) => X_Logic0_port, B(27) => X_Logic0_port, 
                           B(26) => X_Logic0_port, B(25) => X_Logic0_port, 
                           B(24) => X_Logic0_port, B(23) => X_Logic0_port, 
                           B(22) => X_Logic0_port, B(21) => X_Logic0_port, 
                           B(20) => X_Logic0_port, B(19) => X_Logic0_port, 
                           B(18) => X_Logic0_port, B(17) => X_Logic0_port, 
                           B(16) => X_Logic0_port, B(15) => X_Logic0_port, 
                           B(14) => X_Logic0_port, B(13) => X_Logic0_port, 
                           B(12) => X_Logic0_port, B(11) => X_Logic0_port, 
                           B(10) => X_Logic0_port, B(9) => X_Logic0_port, B(8) 
                           => X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, S => select_zero_sig, Z(31) => 
                           ALU_RES(31), Z(30) => ALU_RES(30), Z(29) => 
                           ALU_RES(29), Z(28) => ALU_RES(28), Z(27) => 
                           ALU_RES(27), Z(26) => ALU_RES(26), Z(25) => 
                           ALU_RES(25), Z(24) => ALU_RES(24), Z(23) => 
                           ALU_RES(23), Z(22) => ALU_RES(22), Z(21) => 
                           ALU_RES(21), Z(20) => ALU_RES(20), Z(19) => 
                           ALU_RES(19), Z(18) => ALU_RES(18), Z(17) => 
                           ALU_RES(17), Z(16) => ALU_RES(16), Z(15) => 
                           ALU_RES(15), Z(14) => ALU_RES(14), Z(13) => 
                           ALU_RES(13), Z(12) => ALU_RES(12), Z(11) => 
                           ALU_RES(11), Z(10) => ALU_RES(10), Z(9) => 
                           ALU_RES(9), Z(8) => ALU_RES(8), Z(7) => ALU_RES(7), 
                           Z(6) => ALU_RES(6), Z(5) => ALU_RES(5), Z(4) => 
                           ALU_RES(4), Z(3) => ALU_RES(3), Z(2) => ALU_RES(2), 
                           Z(1) => ALU_RES(1), Z(0) => ALU_RES(0));
   U3 : OAI22_X1 port map( A1 => n198, A2 => n39, B1 => n44, B2 => n75, ZN => 
                           A_SHF_5_port);
   U4 : OAI22_X1 port map( A1 => n199, A2 => n39, B1 => n44, B2 => n76, ZN => 
                           A_SHF_6_port);
   U5 : OAI22_X1 port map( A1 => n189, A2 => n40, B1 => n45, B2 => n66, ZN => 
                           A_SHF_26_port);
   U6 : OAI22_X1 port map( A1 => n190, A2 => n40, B1 => n45, B2 => n67, ZN => 
                           A_SHF_27_port);
   U7 : AND3_X1 port map( A1 => ALU_OPC(4), A2 => ALU_OPC(2), A3 => n163, ZN =>
                           n1);
   U8 : OR2_X1 port map( A1 => n211, A2 => n205, ZN => n2);
   U9 : OR2_X1 port map( A1 => n170, A2 => ALU_OPC(4), ZN => n3);
   U10 : INV_X1 port map( A => n4, ZN => ADD_SUB);
   U11 : NOR2_X1 port map( A1 => n210, A2 => n3, ZN => n5);
   U12 : NOR2_X1 port map( A1 => n212, A2 => n2, ZN => n6);
   U13 : NOR2_X1 port map( A1 => n5, A2 => n6, ZN => n4);
   U14 : BUF_X1 port map( A => n168, Z => n17);
   U15 : BUF_X1 port map( A => n168, Z => n18);
   U16 : BUF_X1 port map( A => n168, Z => n19);
   U17 : OAI22_X1 port map( A1 => n179, A2 => n41, B1 => n46, B2 => n56, ZN => 
                           A_SHF_17_port);
   U18 : OAI22_X1 port map( A1 => n200, A2 => n39, B1 => n44, B2 => n77, ZN => 
                           A_SHF_7_port);
   U19 : OAI22_X1 port map( A1 => n180, A2 => n41, B1 => n46, B2 => n57, ZN => 
                           A_SHF_18_port);
   U20 : OAI22_X1 port map( A1 => n188, A2 => n40, B1 => n45, B2 => n65, ZN => 
                           A_SHF_25_port);
   U21 : OAI22_X1 port map( A1 => n191, A2 => n40, B1 => n45, B2 => n68, ZN => 
                           A_SHF_28_port);
   U22 : OAI22_X1 port map( A1 => n197, A2 => n40, B1 => n45, B2 => n74, ZN => 
                           A_SHF_4_port);
   U23 : NOR2_X1 port map( A1 => n42, A2 => n196, ZN => B_SHF_3_port);
   U24 : OAI22_X1 port map( A1 => n201, A2 => n39, B1 => n44, B2 => n85, ZN => 
                           A_SHF_8_port);
   U25 : OAI22_X1 port map( A1 => n193, A2 => n39, B1 => n45, B2 => n70, ZN => 
                           A_SHF_2_port);
   U26 : OAI22_X1 port map( A1 => n186, A2 => n40, B1 => n45, B2 => n63, ZN => 
                           A_SHF_23_port);
   U27 : OAI22_X1 port map( A1 => n187, A2 => n40, B1 => n45, B2 => n64, ZN => 
                           A_SHF_24_port);
   U28 : OAI22_X1 port map( A1 => n181, A2 => n40, B1 => n46, B2 => n58, ZN => 
                           A_SHF_19_port);
   U29 : OAI22_X1 port map( A1 => n183, A2 => n40, B1 => n46, B2 => n60, ZN => 
                           A_SHF_20_port);
   U30 : OAI22_X1 port map( A1 => n184, A2 => n40, B1 => n46, B2 => n61, ZN => 
                           A_SHF_21_port);
   U31 : OAI22_X1 port map( A1 => n185, A2 => n40, B1 => n46, B2 => n62, ZN => 
                           A_SHF_22_port);
   U32 : OAI22_X1 port map( A1 => n174, A2 => n41, B1 => n47, B2 => n51, ZN => 
                           A_SHF_12_port);
   U33 : OAI22_X1 port map( A1 => n175, A2 => n41, B1 => n46, B2 => n52, ZN => 
                           A_SHF_13_port);
   U34 : OAI22_X1 port map( A1 => n176, A2 => n41, B1 => n46, B2 => n53, ZN => 
                           A_SHF_14_port);
   U35 : NOR2_X1 port map( A1 => n196, A2 => n30, ZN => B_MUL_3_port);
   U36 : NOR2_X1 port map( A1 => n198, A2 => n30, ZN => B_MUL_5_port);
   U37 : NOR2_X1 port map( A1 => n200, A2 => n30, ZN => B_MUL_7_port);
   U38 : NOR2_X1 port map( A1 => n202, A2 => n30, ZN => B_MUL_9_port);
   U39 : NOR2_X1 port map( A1 => n182, A2 => n30, ZN => B_MUL_1_port);
   U40 : NOR2_X1 port map( A1 => n173, A2 => n30, ZN => B_MUL_11_port);
   U41 : NOR2_X1 port map( A1 => n175, A2 => n30, ZN => B_MUL_13_port);
   U42 : NOR2_X1 port map( A1 => n42, A2 => n202, ZN => B_SHF_9_port);
   U43 : NOR2_X1 port map( A1 => n42, A2 => n201, ZN => B_SHF_8_port);
   U44 : NOR2_X1 port map( A1 => n44, A2 => n172, ZN => B_SHF_10_port);
   U45 : OAI22_X1 port map( A1 => n182, A2 => n40, B1 => n46, B2 => n59, ZN => 
                           A_SHF_1_port);
   U46 : NOR2_X1 port map( A1 => n42, A2 => n193, ZN => B_SHF_2_port);
   U47 : OAI22_X1 port map( A1 => n202, A2 => n39, B1 => n44, B2 => n86, ZN => 
                           A_SHF_9_port);
   U48 : OAI22_X1 port map( A1 => n171, A2 => n39, B1 => n46, B2 => n48, ZN => 
                           A_SHF_0_port);
   U49 : NOR2_X1 port map( A1 => n42, A2 => n200, ZN => B_SHF_7_port);
   U50 : NOR2_X1 port map( A1 => n42, A2 => n199, ZN => B_SHF_6_port);
   U51 : NOR2_X1 port map( A1 => n42, A2 => n198, ZN => B_SHF_5_port);
   U52 : OAI22_X1 port map( A1 => n173, A2 => n41, B1 => n47, B2 => n50, ZN => 
                           A_SHF_11_port);
   U53 : OAI22_X1 port map( A1 => n177, A2 => n41, B1 => n46, B2 => n54, ZN => 
                           A_SHF_15_port);
   U54 : OAI22_X1 port map( A1 => n192, A2 => n39, B1 => n45, B2 => n69, ZN => 
                           A_SHF_29_port);
   U55 : OAI22_X1 port map( A1 => n178, A2 => n41, B1 => n46, B2 => n55, ZN => 
                           A_SHF_16_port);
   U56 : OAI22_X1 port map( A1 => n196, A2 => n39, B1 => n45, B2 => n73, ZN => 
                           A_SHF_3_port);
   U57 : NOR2_X1 port map( A1 => n17, A2 => n48, ZN => A_ADD_0_port);
   U58 : NOR2_X1 port map( A1 => n19, A2 => n74, ZN => A_ADD_4_port);
   U59 : NOR2_X1 port map( A1 => n19, A2 => n85, ZN => A_ADD_8_port);
   U60 : NOR2_X1 port map( A1 => n19, A2 => n75, ZN => A_ADD_5_port);
   U61 : NOR2_X1 port map( A1 => n19, A2 => n86, ZN => A_ADD_9_port);
   U62 : NOR2_X1 port map( A1 => n19, A2 => n76, ZN => A_ADD_6_port);
   U63 : NOR2_X1 port map( A1 => n19, A2 => n73, ZN => A_ADD_3_port);
   U64 : NOR2_X1 port map( A1 => n19, A2 => n77, ZN => A_ADD_7_port);
   U65 : NOR2_X1 port map( A1 => n19, A2 => n72, ZN => A_ADD_31_port);
   U66 : NOR2_X1 port map( A1 => n17, A2 => n51, ZN => A_ADD_12_port);
   U67 : NOR2_X1 port map( A1 => n17, A2 => n55, ZN => A_ADD_16_port);
   U68 : NOR2_X1 port map( A1 => n18, A2 => n64, ZN => A_ADD_24_port);
   U69 : NOR2_X1 port map( A1 => n17, A2 => n59, ZN => A_ADD_1_port);
   U70 : NOR2_X1 port map( A1 => n17, A2 => n52, ZN => A_ADD_13_port);
   U71 : NOR2_X1 port map( A1 => n17, A2 => n56, ZN => A_ADD_17_port);
   U72 : NOR2_X1 port map( A1 => n18, A2 => n65, ZN => A_ADD_25_port);
   U73 : NOR2_X1 port map( A1 => n18, A2 => n70, ZN => A_ADD_2_port);
   U74 : NOR2_X1 port map( A1 => n17, A2 => n49, ZN => A_ADD_10_port);
   U75 : NOR2_X1 port map( A1 => n17, A2 => n53, ZN => A_ADD_14_port);
   U76 : NOR2_X1 port map( A1 => n17, A2 => n57, ZN => A_ADD_18_port);
   U77 : NOR2_X1 port map( A1 => n18, A2 => n66, ZN => A_ADD_26_port);
   U78 : NOR2_X1 port map( A1 => n18, A2 => n62, ZN => A_ADD_22_port);
   U79 : NOR2_X1 port map( A1 => n18, A2 => n61, ZN => A_ADD_21_port);
   U80 : NOR2_X1 port map( A1 => n18, A2 => n60, ZN => A_ADD_20_port);
   U81 : NOR2_X1 port map( A1 => n18, A2 => n71, ZN => A_ADD_30_port);
   U82 : NOR2_X1 port map( A1 => n18, A2 => n69, ZN => A_ADD_29_port);
   U83 : NOR2_X1 port map( A1 => n18, A2 => n68, ZN => A_ADD_28_port);
   U84 : NOR2_X1 port map( A1 => n17, A2 => n50, ZN => A_ADD_11_port);
   U85 : NOR2_X1 port map( A1 => n17, A2 => n54, ZN => A_ADD_15_port);
   U86 : NOR2_X1 port map( A1 => n17, A2 => n58, ZN => A_ADD_19_port);
   U87 : NOR2_X1 port map( A1 => n18, A2 => n63, ZN => A_ADD_23_port);
   U88 : NOR2_X1 port map( A1 => n18, A2 => n67, ZN => A_ADD_27_port);
   U89 : NOR2_X1 port map( A1 => n43, A2 => n182, ZN => B_SHF_1_port);
   U90 : NOR2_X1 port map( A1 => n42, A2 => n191, ZN => B_SHF_28_port);
   U91 : NOR2_X1 port map( A1 => n42, A2 => n190, ZN => B_SHF_27_port);
   U92 : NOR2_X1 port map( A1 => n43, A2 => n189, ZN => B_SHF_26_port);
   U93 : OAI22_X1 port map( A1 => n172, A2 => n41, B1 => n47, B2 => n49, ZN => 
                           A_SHF_10_port);
   U94 : NOR2_X1 port map( A1 => n44, A2 => n173, ZN => B_SHF_11_port);
   U95 : NOR2_X1 port map( A1 => n177, A2 => n30, ZN => B_MUL_15_port);
   U96 : OAI22_X1 port map( A1 => n194, A2 => n39, B1 => n45, B2 => n71, ZN => 
                           A_SHF_30_port);
   U97 : NOR2_X1 port map( A1 => n43, A2 => n180, ZN => B_SHF_18_port);
   U98 : NOR2_X1 port map( A1 => n42, A2 => n192, ZN => B_SHF_29_port);
   U99 : NOR2_X1 port map( A1 => n42, A2 => n194, ZN => B_SHF_30_port);
   U100 : BUF_X1 port map( A => n208, Z => n11);
   U101 : BUF_X1 port map( A => n208, Z => n12);
   U102 : BUF_X1 port map( A => n208, Z => n13);
   U103 : BUF_X1 port map( A => n208, Z => n15);
   U104 : BUF_X1 port map( A => n208, Z => n14);
   U105 : NOR2_X1 port map( A1 => n43, A2 => n188, ZN => B_SHF_25_port);
   U106 : NOR2_X1 port map( A1 => n44, A2 => n171, ZN => B_SHF_0_port);
   U107 : NOR2_X1 port map( A1 => n43, A2 => n178, ZN => B_SHF_16_port);
   U108 : NOR2_X1 port map( A1 => n43, A2 => n179, ZN => B_SHF_17_port);
   U109 : NOR2_X1 port map( A1 => n44, A2 => n177, ZN => B_SHF_15_port);
   U110 : NOR2_X1 port map( A1 => n54, A2 => n29, ZN => A_MUL_15_port);
   U111 : NOR2_X1 port map( A1 => n193, A2 => n30, ZN => B_MUL_2_port);
   U112 : NOR2_X1 port map( A1 => n197, A2 => n29, ZN => B_MUL_4_port);
   U113 : NOR2_X1 port map( A1 => n199, A2 => n30, ZN => B_MUL_6_port);
   U114 : NOR2_X1 port map( A1 => n201, A2 => n29, ZN => B_MUL_8_port);
   U115 : NOR2_X1 port map( A1 => n171, A2 => n30, ZN => B_MUL_0_port);
   U116 : NOR2_X1 port map( A1 => n172, A2 => n30, ZN => B_MUL_10_port);
   U117 : NOR2_X1 port map( A1 => n174, A2 => n30, ZN => B_MUL_12_port);
   U118 : NOR2_X1 port map( A1 => n176, A2 => n30, ZN => B_MUL_14_port);
   U119 : BUF_X1 port map( A => n4, Z => n9);
   U120 : BUF_X1 port map( A => n4, Z => n8);
   U121 : OAI21_X1 port map( B1 => n47, B2 => n197, A => n41, ZN => 
                           B_SHF_4_port);
   U122 : BUF_X1 port map( A => n4, Z => n10);
   U123 : NOR2_X1 port map( A1 => n43, A2 => n187, ZN => B_SHF_24_port);
   U124 : NOR2_X1 port map( A1 => n43, A2 => n186, ZN => B_SHF_23_port);
   U125 : NOR2_X1 port map( A1 => n43, A2 => n185, ZN => B_SHF_22_port);
   U126 : NOR2_X1 port map( A1 => n34, A2 => n71, ZN => A_CMP_30_port);
   U127 : OAI22_X1 port map( A1 => n99, A2 => n198, B1 => n100, B2 => n75, ZN 
                           => LOGIC_RES_5_port);
   U128 : OAI22_X1 port map( A1 => n97, A2 => n199, B1 => n98, B2 => n76, ZN =>
                           LOGIC_RES_6_port);
   U129 : OAI22_X1 port map( A1 => n95, A2 => n200, B1 => n96, B2 => n77, ZN =>
                           LOGIC_RES_7_port);
   U130 : OAI22_X1 port map( A1 => n90, A2 => n202, B1 => n91, B2 => n86, ZN =>
                           LOGIC_RES_9_port);
   U131 : OAI22_X1 port map( A1 => n105, A2 => n195, B1 => n106, B2 => n72, ZN 
                           => LOGIC_RES_31_port);
   U132 : NOR2_X1 port map( A1 => n33, A2 => n59, ZN => A_CMP_1_port);
   U133 : OAI22_X1 port map( A1 => n151, A2 => n172, B1 => n152, B2 => n49, ZN 
                           => LOGIC_RES_10_port);
   U134 : OAI22_X1 port map( A1 => n149, A2 => n173, B1 => n150, B2 => n50, ZN 
                           => LOGIC_RES_11_port);
   U135 : OAI22_X1 port map( A1 => n145, A2 => n175, B1 => n146, B2 => n52, ZN 
                           => LOGIC_RES_13_port);
   U136 : OAI22_X1 port map( A1 => n143, A2 => n176, B1 => n144, B2 => n53, ZN 
                           => LOGIC_RES_14_port);
   U137 : OAI22_X1 port map( A1 => n141, A2 => n177, B1 => n142, B2 => n54, ZN 
                           => LOGIC_RES_15_port);
   U138 : OAI22_X1 port map( A1 => n137, A2 => n179, B1 => n138, B2 => n56, ZN 
                           => LOGIC_RES_17_port);
   U139 : OAI22_X1 port map( A1 => n135, A2 => n180, B1 => n136, B2 => n57, ZN 
                           => LOGIC_RES_18_port);
   U140 : OAI22_X1 port map( A1 => n133, A2 => n181, B1 => n134, B2 => n58, ZN 
                           => LOGIC_RES_19_port);
   U141 : OAI22_X1 port map( A1 => n127, A2 => n184, B1 => n128, B2 => n61, ZN 
                           => LOGIC_RES_21_port);
   U142 : OAI22_X1 port map( A1 => n125, A2 => n185, B1 => n126, B2 => n62, ZN 
                           => LOGIC_RES_22_port);
   U143 : OAI22_X1 port map( A1 => n123, A2 => n186, B1 => n124, B2 => n63, ZN 
                           => LOGIC_RES_23_port);
   U144 : OAI22_X1 port map( A1 => n119, A2 => n188, B1 => n120, B2 => n65, ZN 
                           => LOGIC_RES_25_port);
   U145 : OAI22_X1 port map( A1 => n117, A2 => n189, B1 => n118, B2 => n66, ZN 
                           => LOGIC_RES_26_port);
   U146 : OAI22_X1 port map( A1 => n115, A2 => n190, B1 => n116, B2 => n67, ZN 
                           => LOGIC_RES_27_port);
   U147 : OAI22_X1 port map( A1 => n111, A2 => n192, B1 => n112, B2 => n69, ZN 
                           => LOGIC_RES_29_port);
   U148 : OAI22_X1 port map( A1 => n107, A2 => n194, B1 => n108, B2 => n71, ZN 
                           => LOGIC_RES_30_port);
   U149 : NOR2_X1 port map( A1 => n43, A2 => n181, ZN => B_SHF_19_port);
   U150 : NOR2_X1 port map( A1 => n43, A2 => n184, ZN => B_SHF_21_port);
   U151 : NOR2_X1 port map( A1 => n44, A2 => n175, ZN => B_SHF_13_port);
   U152 : NOR2_X1 port map( A1 => n43, A2 => n183, ZN => B_SHF_20_port);
   U153 : NOR2_X1 port map( A1 => n44, A2 => n176, ZN => B_SHF_14_port);
   U154 : NOR2_X1 port map( A1 => n44, A2 => n174, ZN => B_SHF_12_port);
   U155 : NOR2_X1 port map( A1 => n38, A2 => n200, ZN => B_CMP_7_port);
   U156 : NOR2_X1 port map( A1 => n38, A2 => n202, ZN => B_CMP_9_port);
   U157 : AOI21_X1 port map( B1 => n13, B2 => n198, A => n25, ZN => n100);
   U158 : AOI21_X1 port map( B1 => n13, B2 => n199, A => n25, ZN => n98);
   U159 : AOI21_X1 port map( B1 => n13, B2 => n201, A => n25, ZN => n94);
   U160 : AOI21_X1 port map( B1 => n15, B2 => n182, A => n27, ZN => n132);
   U161 : AOI21_X1 port map( B1 => n14, B2 => n193, A => n26, ZN => n110);
   U162 : AOI21_X1 port map( B1 => n14, B2 => n196, A => n26, ZN => n104);
   U163 : AOI21_X1 port map( B1 => n14, B2 => n197, A => n26, ZN => n102);
   U164 : AOI21_X1 port map( B1 => n14, B2 => n200, A => n26, ZN => n96);
   U165 : AOI21_X1 port map( B1 => n14, B2 => n202, A => n26, ZN => n91);
   U166 : AOI21_X1 port map( B1 => n15, B2 => n176, A => n27, ZN => n144);
   U167 : AOI21_X1 port map( B1 => n15, B2 => n177, A => n27, ZN => n142);
   U168 : AOI21_X1 port map( B1 => n15, B2 => n178, A => n27, ZN => n140);
   U169 : AOI21_X1 port map( B1 => n15, B2 => n179, A => n27, ZN => n138);
   U170 : AOI21_X1 port map( B1 => n15, B2 => n180, A => n27, ZN => n136);
   U171 : AOI21_X1 port map( B1 => n15, B2 => n181, A => n27, ZN => n134);
   U172 : AOI21_X1 port map( B1 => n15, B2 => n183, A => n27, ZN => n130);
   U173 : AOI21_X1 port map( B1 => n15, B2 => n184, A => n27, ZN => n128);
   U174 : AOI21_X1 port map( B1 => n15, B2 => n185, A => n27, ZN => n126);
   U175 : AOI21_X1 port map( B1 => n15, B2 => n186, A => n27, ZN => n124);
   U176 : AOI21_X1 port map( B1 => n15, B2 => n187, A => n26, ZN => n122);
   U177 : AOI21_X1 port map( B1 => n14, B2 => n188, A => n26, ZN => n120);
   U178 : AOI21_X1 port map( B1 => n14, B2 => n189, A => n26, ZN => n118);
   U179 : AOI21_X1 port map( B1 => n14, B2 => n190, A => n26, ZN => n116);
   U180 : AOI21_X1 port map( B1 => n14, B2 => n191, A => n26, ZN => n114);
   U181 : AOI21_X1 port map( B1 => n14, B2 => n192, A => n26, ZN => n112);
   U182 : AOI21_X1 port map( B1 => n14, B2 => n194, A => n26, ZN => n108);
   U183 : AOI21_X1 port map( B1 => n14, B2 => n195, A => n26, ZN => n106);
   U184 : AOI21_X1 port map( B1 => n16, B2 => n172, A => n28, ZN => n152);
   U185 : AOI21_X1 port map( B1 => n16, B2 => n173, A => n28, ZN => n150);
   U186 : AOI21_X1 port map( B1 => n16, B2 => n174, A => n27, ZN => n148);
   U187 : AOI21_X1 port map( B1 => n16, B2 => n175, A => n27, ZN => n146);
   U188 : NOR2_X1 port map( A1 => n38, A2 => n201, ZN => B_CMP_8_port);
   U189 : NOR2_X1 port map( A1 => n38, A2 => n199, ZN => B_CMP_6_port);
   U190 : NOR2_X1 port map( A1 => n37, A2 => n194, ZN => B_CMP_30_port);
   U191 : NOR2_X1 port map( A1 => n35, A2 => n171, ZN => B_CMP_0_port);
   U192 : NOR2_X1 port map( A1 => n37, A2 => n196, ZN => B_CMP_3_port);
   U193 : NOR2_X1 port map( A1 => n37, A2 => n198, ZN => B_CMP_5_port);
   U194 : NOR2_X1 port map( A1 => n35, A2 => n173, ZN => B_CMP_11_port);
   U195 : NOR2_X1 port map( A1 => n36, A2 => n175, ZN => B_CMP_13_port);
   U196 : NOR2_X1 port map( A1 => n36, A2 => n177, ZN => B_CMP_15_port);
   U197 : NOR2_X1 port map( A1 => n36, A2 => n179, ZN => B_CMP_17_port);
   U198 : NOR2_X1 port map( A1 => n36, A2 => n181, ZN => B_CMP_19_port);
   U199 : NOR2_X1 port map( A1 => n36, A2 => n184, ZN => B_CMP_21_port);
   U200 : NOR2_X1 port map( A1 => n36, A2 => n186, ZN => B_CMP_23_port);
   U201 : NOR2_X1 port map( A1 => n37, A2 => n188, ZN => B_CMP_25_port);
   U202 : NOR2_X1 port map( A1 => n37, A2 => n190, ZN => B_CMP_27_port);
   U203 : NOR2_X1 port map( A1 => n37, A2 => n192, ZN => B_CMP_29_port);
   U204 : NOR2_X1 port map( A1 => n35, A2 => n72, ZN => A_CMP_31_port);
   U205 : NOR2_X1 port map( A1 => n37, A2 => n197, ZN => B_CMP_4_port);
   U206 : NOR2_X1 port map( A1 => n35, A2 => n174, ZN => B_CMP_12_port);
   U207 : NOR2_X1 port map( A1 => n36, A2 => n178, ZN => B_CMP_16_port);
   U208 : NOR2_X1 port map( A1 => n36, A2 => n183, ZN => B_CMP_20_port);
   U209 : NOR2_X1 port map( A1 => n37, A2 => n187, ZN => B_CMP_24_port);
   U210 : NOR2_X1 port map( A1 => n37, A2 => n191, ZN => B_CMP_28_port);
   U211 : NOR2_X1 port map( A1 => n37, A2 => n193, ZN => B_CMP_2_port);
   U212 : NOR2_X1 port map( A1 => n35, A2 => n172, ZN => B_CMP_10_port);
   U213 : NOR2_X1 port map( A1 => n36, A2 => n176, ZN => B_CMP_14_port);
   U214 : NOR2_X1 port map( A1 => n36, A2 => n180, ZN => B_CMP_18_port);
   U215 : NOR2_X1 port map( A1 => n36, A2 => n185, ZN => B_CMP_22_port);
   U216 : NOR2_X1 port map( A1 => n37, A2 => n189, ZN => B_CMP_26_port);
   U217 : AND2_X1 port map( A1 => n22, A2 => n10, ZN => n168);
   U218 : NOR2_X1 port map( A1 => n42, A2 => n195, ZN => B_SHF_31_port);
   U219 : NOR2_X1 port map( A1 => n36, A2 => n182, ZN => B_CMP_1_port);
   U220 : NOR2_X1 port map( A1 => n33, A2 => n48, ZN => A_CMP_0_port);
   U221 : NOR2_X1 port map( A1 => n35, A2 => n73, ZN => A_CMP_3_port);
   U222 : NOR2_X1 port map( A1 => n35, A2 => n75, ZN => A_CMP_5_port);
   U223 : NOR2_X1 port map( A1 => n35, A2 => n77, ZN => A_CMP_7_port);
   U224 : NOR2_X1 port map( A1 => n35, A2 => n86, ZN => A_CMP_9_port);
   U225 : NOR2_X1 port map( A1 => n33, A2 => n50, ZN => A_CMP_11_port);
   U226 : NOR2_X1 port map( A1 => n33, A2 => n52, ZN => A_CMP_13_port);
   U228 : NOR2_X1 port map( A1 => n33, A2 => n54, ZN => A_CMP_15_port);
   U229 : NOR2_X1 port map( A1 => n37, A2 => n195, ZN => B_CMP_31_port);
   U230 : NOR2_X1 port map( A1 => n33, A2 => n56, ZN => A_CMP_17_port);
   U231 : NOR2_X1 port map( A1 => n33, A2 => n58, ZN => A_CMP_19_port);
   U232 : NOR2_X1 port map( A1 => n34, A2 => n61, ZN => A_CMP_21_port);
   U233 : NOR2_X1 port map( A1 => n34, A2 => n63, ZN => A_CMP_23_port);
   U234 : NOR2_X1 port map( A1 => n34, A2 => n65, ZN => A_CMP_25_port);
   U235 : NOR2_X1 port map( A1 => n34, A2 => n67, ZN => A_CMP_27_port);
   U236 : NOR2_X1 port map( A1 => n34, A2 => n69, ZN => A_CMP_29_port);
   U237 : NOR2_X1 port map( A1 => n35, A2 => n74, ZN => A_CMP_4_port);
   U238 : NOR2_X1 port map( A1 => n35, A2 => n85, ZN => A_CMP_8_port);
   U239 : NOR2_X1 port map( A1 => n33, A2 => n51, ZN => A_CMP_12_port);
   U240 : NOR2_X1 port map( A1 => n34, A2 => n70, ZN => A_CMP_2_port);
   U241 : NOR2_X1 port map( A1 => n35, A2 => n76, ZN => A_CMP_6_port);
   U242 : NOR2_X1 port map( A1 => n33, A2 => n49, ZN => A_CMP_10_port);
   U243 : NOR2_X1 port map( A1 => n33, A2 => n53, ZN => A_CMP_14_port);
   U244 : NOR2_X1 port map( A1 => n33, A2 => n55, ZN => A_CMP_16_port);
   U245 : NOR2_X1 port map( A1 => n34, A2 => n60, ZN => A_CMP_20_port);
   U246 : NOR2_X1 port map( A1 => n34, A2 => n64, ZN => A_CMP_24_port);
   U247 : NOR2_X1 port map( A1 => n34, A2 => n68, ZN => A_CMP_28_port);
   U248 : NOR2_X1 port map( A1 => n33, A2 => n57, ZN => A_CMP_18_port);
   U249 : NOR2_X1 port map( A1 => n34, A2 => n62, ZN => A_CMP_22_port);
   U250 : NOR2_X1 port map( A1 => n34, A2 => n66, ZN => A_CMP_26_port);
   U251 : OAI22_X1 port map( A1 => OP2(0), A2 => n10, B1 => n171, B2 => n22, ZN
                           => B_ADD_0_port);
   U252 : OAI22_X1 port map( A1 => OP2(4), A2 => n8, B1 => n197, B2 => n20, ZN 
                           => B_ADD_4_port);
   U253 : OAI22_X1 port map( A1 => OP2(8), A2 => n8, B1 => n201, B2 => n20, ZN 
                           => B_ADD_8_port);
   U254 : OAI22_X1 port map( A1 => OP2(12), A2 => n10, B1 => n174, B2 => n22, 
                           ZN => B_ADD_12_port);
   U255 : OAI22_X1 port map( A1 => OP2(16), A2 => n10, B1 => n178, B2 => n22, 
                           ZN => B_ADD_16_port);
   U256 : OAI22_X1 port map( A1 => OP2(24), A2 => n9, B1 => n187, B2 => n21, ZN
                           => B_ADD_24_port);
   U266 : OAI22_X1 port map( A1 => OP2(5), A2 => n8, B1 => n198, B2 => n20, ZN 
                           => B_ADD_5_port);
   U273 : OAI22_X1 port map( A1 => OP2(1), A2 => n9, B1 => n182, B2 => n21, ZN 
                           => B_ADD_1_port);
   U274 : OAI22_X1 port map( A1 => OP2(9), A2 => n8, B1 => n202, B2 => n20, ZN 
                           => B_ADD_9_port);
   U275 : OAI22_X1 port map( A1 => OP2(13), A2 => n10, B1 => n175, B2 => n22, 
                           ZN => B_ADD_13_port);
   U276 : OAI22_X1 port map( A1 => OP2(17), A2 => n9, B1 => n179, B2 => n21, ZN
                           => B_ADD_17_port);
   U277 : OAI22_X1 port map( A1 => OP2(25), A2 => n9, B1 => n188, B2 => n21, ZN
                           => B_ADD_25_port);
   U278 : OAI22_X1 port map( A1 => OP2(2), A2 => n8, B1 => n193, B2 => n20, ZN 
                           => B_ADD_2_port);
   U279 : OAI22_X1 port map( A1 => OP2(6), A2 => n8, B1 => n199, B2 => n20, ZN 
                           => B_ADD_6_port);
   U280 : OAI22_X1 port map( A1 => OP2(10), A2 => n10, B1 => n172, B2 => n22, 
                           ZN => B_ADD_10_port);
   U281 : OAI22_X1 port map( A1 => OP2(14), A2 => n10, B1 => n176, B2 => n22, 
                           ZN => B_ADD_14_port);
   U282 : OAI22_X1 port map( A1 => OP2(18), A2 => n9, B1 => n180, B2 => n21, ZN
                           => B_ADD_18_port);
   U283 : OAI22_X1 port map( A1 => OP2(26), A2 => n9, B1 => n189, B2 => n21, ZN
                           => B_ADD_26_port);
   U284 : OAI22_X1 port map( A1 => OP2(22), A2 => n9, B1 => n185, B2 => n21, ZN
                           => B_ADD_22_port);
   U285 : OAI22_X1 port map( A1 => OP2(21), A2 => n9, B1 => n184, B2 => n21, ZN
                           => B_ADD_21_port);
   U286 : OAI22_X1 port map( A1 => OP2(20), A2 => n9, B1 => n183, B2 => n21, ZN
                           => B_ADD_20_port);
   U287 : OAI22_X1 port map( A1 => OP2(30), A2 => n8, B1 => n194, B2 => n20, ZN
                           => B_ADD_30_port);
   U288 : OAI22_X1 port map( A1 => OP2(29), A2 => n8, B1 => n192, B2 => n20, ZN
                           => B_ADD_29_port);
   U289 : OAI22_X1 port map( A1 => OP2(28), A2 => n8, B1 => n191, B2 => n20, ZN
                           => B_ADD_28_port);
   U290 : OAI22_X1 port map( A1 => OP2(3), A2 => n8, B1 => n196, B2 => n20, ZN 
                           => B_ADD_3_port);
   U291 : OAI22_X1 port map( A1 => OP2(7), A2 => n8, B1 => n200, B2 => n20, ZN 
                           => B_ADD_7_port);
   U292 : OAI22_X1 port map( A1 => OP2(11), A2 => n10, B1 => n173, B2 => n22, 
                           ZN => B_ADD_11_port);
   U293 : OAI22_X1 port map( A1 => OP2(15), A2 => n10, B1 => n177, B2 => n22, 
                           ZN => B_ADD_15_port);
   U294 : OAI22_X1 port map( A1 => OP2(19), A2 => n9, B1 => n181, B2 => n21, ZN
                           => B_ADD_19_port);
   U295 : OAI22_X1 port map( A1 => OP2(23), A2 => n9, B1 => n186, B2 => n21, ZN
                           => B_ADD_23_port);
   U296 : OAI22_X1 port map( A1 => OP2(27), A2 => n9, B1 => n190, B2 => n21, ZN
                           => B_ADD_27_port);
   U297 : OAI22_X1 port map( A1 => OP2(31), A2 => n8, B1 => n195, B2 => n20, ZN
                           => B_ADD_31_port);
   U298 : INV_X1 port map( A => n1, ZN => n30);
   U299 : INV_X1 port map( A => n1, ZN => n29);
   U300 : INV_X1 port map( A => n7, ZN => n31);
   U301 : INV_X1 port map( A => n7, ZN => n32);
   U302 : AOI221_X1 port map( B1 => OP1(10), B2 => n31, C1 => n11, C2 => n49, A
                           => n23, ZN => n151);
   U303 : AOI221_X1 port map( B1 => OP1(11), B2 => n32, C1 => n11, C2 => n50, A
                           => n23, ZN => n149);
   U304 : AOI221_X1 port map( B1 => OP1(12), B2 => n31, C1 => n11, C2 => n51, A
                           => n23, ZN => n147);
   U305 : AOI221_X1 port map( B1 => OP1(13), B2 => n32, C1 => n11, C2 => n52, A
                           => n23, ZN => n145);
   U306 : AOI221_X1 port map( B1 => OP1(14), B2 => n31, C1 => n11, C2 => n53, A
                           => n23, ZN => n143);
   U307 : AOI221_X1 port map( B1 => OP1(15), B2 => n32, C1 => n11, C2 => n54, A
                           => n23, ZN => n141);
   U308 : AOI221_X1 port map( B1 => OP1(16), B2 => n31, C1 => n11, C2 => n55, A
                           => n23, ZN => n139);
   U309 : AOI221_X1 port map( B1 => OP1(1), B2 => n32, C1 => n12, C2 => n59, A 
                           => n24, ZN => n131);
   U310 : AOI221_X1 port map( B1 => OP1(2), B2 => n31, C1 => n13, C2 => n70, A 
                           => n25, ZN => n109);
   U311 : AOI221_X1 port map( B1 => OP1(3), B2 => n31, C1 => n12, C2 => n73, A 
                           => n24, ZN => n103);
   U312 : AOI221_X1 port map( B1 => OP1(4), B2 => n31, C1 => n12, C2 => n74, A 
                           => n24, ZN => n101);
   U313 : AOI221_X1 port map( B1 => OP1(5), B2 => n31, C1 => n12, C2 => n75, A 
                           => n24, ZN => n99);
   U314 : AOI221_X1 port map( B1 => OP1(6), B2 => n31, C1 => n11, C2 => n76, A 
                           => n23, ZN => n97);
   U315 : AOI221_X1 port map( B1 => OP1(7), B2 => n31, C1 => n11, C2 => n77, A 
                           => n23, ZN => n95);
   U316 : AOI221_X1 port map( B1 => OP1(8), B2 => n31, C1 => n11, C2 => n85, A 
                           => n23, ZN => n93);
   U317 : AOI221_X1 port map( B1 => OP1(17), B2 => n32, C1 => n12, C2 => n56, A
                           => n24, ZN => n137);
   U318 : AOI221_X1 port map( B1 => OP1(18), B2 => n32, C1 => n12, C2 => n57, A
                           => n24, ZN => n135);
   U319 : AOI221_X1 port map( B1 => OP1(19), B2 => n32, C1 => n12, C2 => n58, A
                           => n24, ZN => n133);
   U320 : AOI221_X1 port map( B1 => OP1(20), B2 => n32, C1 => n12, C2 => n60, A
                           => n24, ZN => n129);
   U321 : AOI221_X1 port map( B1 => OP1(21), B2 => n32, C1 => n12, C2 => n61, A
                           => n24, ZN => n127);
   U322 : AOI221_X1 port map( B1 => OP1(22), B2 => n32, C1 => n12, C2 => n62, A
                           => n24, ZN => n125);
   U323 : AOI221_X1 port map( B1 => OP1(23), B2 => n32, C1 => n12, C2 => n63, A
                           => n24, ZN => n123);
   U324 : AOI221_X1 port map( B1 => OP1(24), B2 => n32, C1 => n13, C2 => n64, A
                           => n25, ZN => n121);
   U325 : AOI221_X1 port map( B1 => OP1(25), B2 => n32, C1 => n13, C2 => n65, A
                           => n25, ZN => n119);
   U326 : AOI221_X1 port map( B1 => OP1(26), B2 => n32, C1 => n12, C2 => n66, A
                           => n24, ZN => n117);
   U327 : AOI221_X1 port map( B1 => OP1(27), B2 => n32, C1 => n13, C2 => n67, A
                           => n25, ZN => n115);
   U328 : AOI221_X1 port map( B1 => OP1(28), B2 => n31, C1 => n13, C2 => n68, A
                           => n25, ZN => n113);
   U329 : AOI221_X1 port map( B1 => OP1(29), B2 => n31, C1 => n13, C2 => n69, A
                           => n25, ZN => n111);
   U330 : AOI221_X1 port map( B1 => OP1(30), B2 => n31, C1 => n13, C2 => n71, A
                           => n25, ZN => n107);
   U331 : AOI221_X1 port map( B1 => OP1(31), B2 => n31, C1 => n13, C2 => n72, A
                           => n25, ZN => n105);
   U332 : AOI221_X1 port map( B1 => n31, B2 => OP1(9), C1 => n11, C2 => n86, A 
                           => n23, ZN => n90);
   U333 : BUF_X1 port map( A => n81, Z => n43);
   U334 : BUF_X1 port map( A => n81, Z => n44);
   U335 : BUF_X1 port map( A => n81, Z => n45);
   U336 : BUF_X1 port map( A => n81, Z => n46);
   U337 : INV_X1 port map( A => OP2(0), ZN => n171);
   U338 : INV_X1 port map( A => OP2(1), ZN => n182);
   U339 : INV_X1 port map( A => OP2(2), ZN => n193);
   U340 : INV_X1 port map( A => OP2(3), ZN => n196);
   U341 : INV_X1 port map( A => OP2(5), ZN => n198);
   U342 : INV_X1 port map( A => OP2(6), ZN => n199);
   U343 : INV_X1 port map( A => OP2(7), ZN => n200);
   U344 : INV_X1 port map( A => OP2(8), ZN => n201);
   U345 : INV_X1 port map( A => OP2(9), ZN => n202);
   U346 : INV_X1 port map( A => OP2(10), ZN => n172);
   U347 : INV_X1 port map( A => OP2(11), ZN => n173);
   U348 : INV_X1 port map( A => OP2(12), ZN => n174);
   U349 : INV_X1 port map( A => OP2(13), ZN => n175);
   U350 : INV_X1 port map( A => OP2(14), ZN => n176);
   U351 : INV_X1 port map( A => OP2(15), ZN => n177);
   U352 : INV_X1 port map( A => OP2(4), ZN => n197);
   U353 : BUF_X1 port map( A => n92, Z => n23);
   U354 : BUF_X1 port map( A => n92, Z => n24);
   U355 : OAI22_X1 port map( A1 => n153, A2 => n171, B1 => n154, B2 => n48, ZN 
                           => LOGIC_RES_0_port);
   U356 : AOI21_X1 port map( B1 => n13, B2 => n171, A => n25, ZN => n154);
   U357 : AOI221_X1 port map( B1 => OP1(0), B2 => n32, C1 => n11, C2 => n48, A 
                           => n23, ZN => n153);
   U358 : BUF_X1 port map( A => n92, Z => n27);
   U359 : BUF_X1 port map( A => n92, Z => n26);
   U360 : BUF_X1 port map( A => n82, Z => n39);
   U361 : BUF_X1 port map( A => n82, Z => n40);
   U362 : BUF_X1 port map( A => n92, Z => n25);
   U363 : BUF_X1 port map( A => n159, Z => n21);
   U364 : BUF_X1 port map( A => n159, Z => n20);
   U365 : BUF_X1 port map( A => n83, Z => n37);
   U366 : BUF_X1 port map( A => n83, Z => n35);
   U367 : BUF_X1 port map( A => n83, Z => n33);
   U368 : BUF_X1 port map( A => n83, Z => n36);
   U369 : BUF_X1 port map( A => n83, Z => n34);
   U370 : BUF_X1 port map( A => n81, Z => n42);
   U371 : INV_X1 port map( A => OP1(0), ZN => n48);
   U372 : INV_X1 port map( A => OP1(1), ZN => n59);
   U373 : INV_X1 port map( A => OP1(2), ZN => n70);
   U374 : INV_X1 port map( A => OP1(3), ZN => n73);
   U375 : INV_X1 port map( A => OP1(4), ZN => n74);
   U376 : INV_X1 port map( A => OP1(5), ZN => n75);
   U377 : INV_X1 port map( A => OP1(6), ZN => n76);
   U378 : INV_X1 port map( A => OP1(7), ZN => n77);
   U379 : INV_X1 port map( A => OP1(8), ZN => n85);
   U380 : INV_X1 port map( A => OP1(9), ZN => n86);
   U381 : INV_X1 port map( A => OP1(10), ZN => n49);
   U382 : INV_X1 port map( A => OP1(11), ZN => n50);
   U383 : INV_X1 port map( A => OP1(12), ZN => n51);
   U384 : INV_X1 port map( A => OP1(13), ZN => n52);
   U385 : INV_X1 port map( A => OP1(14), ZN => n53);
   U386 : INV_X1 port map( A => OP1(15), ZN => n54);
   U387 : BUF_X1 port map( A => n159, Z => n22);
   U388 : INV_X1 port map( A => OP2(16), ZN => n178);
   U389 : INV_X1 port map( A => OP2(17), ZN => n179);
   U390 : INV_X1 port map( A => OP2(18), ZN => n180);
   U391 : INV_X1 port map( A => OP2(19), ZN => n181);
   U392 : INV_X1 port map( A => OP2(20), ZN => n183);
   U393 : INV_X1 port map( A => OP2(21), ZN => n184);
   U394 : INV_X1 port map( A => OP2(22), ZN => n185);
   U395 : INV_X1 port map( A => OP2(23), ZN => n186);
   U396 : INV_X1 port map( A => OP2(24), ZN => n187);
   U397 : INV_X1 port map( A => OP2(25), ZN => n188);
   U398 : INV_X1 port map( A => OP2(26), ZN => n189);
   U399 : INV_X1 port map( A => OP2(27), ZN => n190);
   U400 : INV_X1 port map( A => OP2(28), ZN => n191);
   U401 : INV_X1 port map( A => OP2(29), ZN => n192);
   U402 : INV_X1 port map( A => OP2(30), ZN => n194);
   U403 : INV_X1 port map( A => OP2(31), ZN => n195);
   U404 : BUF_X1 port map( A => n82, Z => n41);
   U405 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => OPSel_0_port);
   U406 : OAI22_X1 port map( A1 => n103, A2 => n196, B1 => n104, B2 => n73, ZN 
                           => LOGIC_RES_3_port);
   U407 : OAI22_X1 port map( A1 => n101, A2 => n197, B1 => n102, B2 => n74, ZN 
                           => LOGIC_RES_4_port);
   U408 : OAI22_X1 port map( A1 => n93, A2 => n201, B1 => n94, B2 => n85, ZN =>
                           LOGIC_RES_8_port);
   U409 : OAI22_X1 port map( A1 => n131, A2 => n182, B1 => n132, B2 => n59, ZN 
                           => LOGIC_RES_1_port);
   U410 : OAI22_X1 port map( A1 => n109, A2 => n193, B1 => n110, B2 => n70, ZN 
                           => LOGIC_RES_2_port);
   U411 : OAI22_X1 port map( A1 => n147, A2 => n174, B1 => n148, B2 => n51, ZN 
                           => LOGIC_RES_12_port);
   U412 : OAI22_X1 port map( A1 => n139, A2 => n178, B1 => n140, B2 => n55, ZN 
                           => LOGIC_RES_16_port);
   U413 : OAI22_X1 port map( A1 => n129, A2 => n183, B1 => n130, B2 => n60, ZN 
                           => LOGIC_RES_20_port);
   U414 : OAI22_X1 port map( A1 => n121, A2 => n187, B1 => n122, B2 => n64, ZN 
                           => LOGIC_RES_24_port);
   U415 : OAI22_X1 port map( A1 => n113, A2 => n191, B1 => n114, B2 => n68, ZN 
                           => LOGIC_RES_28_port);
   U416 : INV_X1 port map( A => OP1(16), ZN => n55);
   U417 : INV_X1 port map( A => OP1(17), ZN => n56);
   U418 : INV_X1 port map( A => OP1(18), ZN => n57);
   U419 : INV_X1 port map( A => OP1(19), ZN => n58);
   U420 : INV_X1 port map( A => OP1(20), ZN => n60);
   U421 : INV_X1 port map( A => OP1(21), ZN => n61);
   U422 : INV_X1 port map( A => OP1(22), ZN => n62);
   U423 : INV_X1 port map( A => OP1(23), ZN => n63);
   U424 : INV_X1 port map( A => OP1(24), ZN => n64);
   U425 : INV_X1 port map( A => OP1(25), ZN => n65);
   U426 : INV_X1 port map( A => OP1(26), ZN => n66);
   U433 : INV_X1 port map( A => OP1(27), ZN => n67);
   U435 : INV_X1 port map( A => OP1(28), ZN => n68);
   U437 : INV_X1 port map( A => OP1(29), ZN => n69);
   U438 : INV_X1 port map( A => OP1(30), ZN => n71);
   U439 : INV_X1 port map( A => OP1(31), ZN => n72);
   U440 : NAND2_X1 port map( A1 => n157, A2 => n207, ZN => LOGIC_ARITH);
   U441 : INV_X1 port map( A => LEFT_RIGHT, ZN => n207);
   U442 : INV_X1 port map( A => n84, ZN => n208);
   U443 : INV_X1 port map( A => n87, ZN => n206);
   U444 : INV_X1 port map( A => n80, ZN => n205);
   U445 : NOR3_X1 port map( A1 => n212, A2 => ALU_OPC(1), A3 => n210, ZN => 
                           n162);
   U446 : NOR3_X1 port map( A1 => ALU_OPC(1), A2 => ALU_OPC(0), A3 => 
                           ALU_OPC(2), ZN => n80);
   U447 : NAND4_X1 port map( A1 => ALU_OPC(0), A2 => ALU_OPC(3), A3 => n212, A4
                           => n209, ZN => n88);
   U448 : NAND4_X1 port map( A1 => ALU_OPC(3), A2 => ALU_OPC(1), A3 => 
                           ALU_OPC(2), A4 => n204, ZN => n89);
   U449 : INV_X1 port map( A => ALU_OPC(3), ZN => n211);
   U450 : NAND2_X1 port map( A1 => n158, A2 => n39, ZN => LEFT_RIGHT);
   U451 : NOR3_X1 port map( A1 => ALU_OPC(3), A2 => ALU_OPC(0), A3 => 
                           ALU_OPC(2), ZN => n156);
   U452 : NAND4_X1 port map( A1 => ALU_OPC(3), A2 => ALU_OPC(1), A3 => n161, A4
                           => n212, ZN => n157);
   U453 : NOR2_X1 port map( A1 => ALU_OPC(0), A2 => ALU_OPC(2), ZN => n161);
   U454 : INV_X1 port map( A => ALU_OPC(2), ZN => n210);
   U455 : INV_X1 port map( A => ALU_OPC(1), ZN => n209);
   U456 : OAI211_X1 port map( C1 => n166, C2 => n167, A => n209, B => 
                           ALU_OPC(0), ZN => n87);
   U457 : NOR2_X1 port map( A1 => ALU_OPC(2), A2 => n211, ZN => n167);
   U458 : NOR3_X1 port map( A1 => n210, A2 => ALU_OPC(3), A3 => ALU_OPC(4), ZN 
                           => n166);
   U459 : AND3_X1 port map( A1 => ALU_OPC(3), A2 => ALU_OPC(4), A3 => n155, ZN 
                           => n92);
   U460 : NOR3_X1 port map( A1 => n210, A2 => ALU_OPC(0), A3 => ALU_OPC(1), ZN 
                           => n155);
   U461 : INV_X1 port map( A => ALU_OPC(0), ZN => n204);
   U462 : INV_X1 port map( A => ALU_OPC(4), ZN => n212);
   U463 : OAI21_X1 port map( B1 => n78, B2 => n209, A => n79, ZN => 
                           select_zero_sig);
   U464 : AOI21_X1 port map( B1 => ALU_OPC(2), B2 => n211, A => ALU_OPC(0), ZN 
                           => n78);
   U465 : NAND2_X1 port map( A1 => n165, A2 => n89, ZN => OPSel_1_port);
   U466 : NAND4_X1 port map( A1 => ALU_OPC(0), A2 => n211, A3 => n210, A4 => 
                           n209, ZN => n165);
   U467 : NAND2_X1 port map( A1 => n80, A2 => n169, ZN => n159);
   U468 : XNOR2_X1 port map( A => n211, B => ALU_OPC(4), ZN => n169);
   U469 : AND4_X1 port map( A1 => n164, A2 => n88, A3 => n87, A4 => n203, ZN =>
                           n83);
   U470 : INV_X1 port map( A => OPSel_1_port, ZN => n203);
   U471 : OR4_X1 port map( A1 => n211, A2 => n210, A3 => ALU_OPC(1), A4 => 
                           ALU_OPC(0), ZN => n7);
   U472 : AND2_X1 port map( A1 => n160, A2 => n157, ZN => n81);
   U473 : NAND4_X1 port map( A1 => ALU_OPC(4), A2 => ALU_OPC(1), A3 => n210, A4
                           => n204, ZN => n160);
   U474 : NOR3_X1 port map( A1 => ALU_OPC(3), A2 => ALU_OPC(0), A3 => 
                           ALU_OPC(1), ZN => n163);
   U475 : CLKBUF_X1 port map( A => n208, Z => n16);
   U476 : CLKBUF_X1 port map( A => n92, Z => n28);
   U477 : CLKBUF_X1 port map( A => n83, Z => n38);
   U478 : CLKBUF_X1 port map( A => n81, Z => n47);
   COMP_RES_1_port <= '0';
   COMP_RES_2_port <= '0';
   COMP_RES_3_port <= '0';
   COMP_RES_4_port <= '0';
   COMP_RES_5_port <= '0';
   COMP_RES_6_port <= '0';
   COMP_RES_7_port <= '0';
   COMP_RES_8_port <= '0';
   COMP_RES_9_port <= '0';
   COMP_RES_10_port <= '0';
   COMP_RES_11_port <= '0';
   COMP_RES_12_port <= '0';
   COMP_RES_13_port <= '0';
   COMP_RES_14_port <= '0';
   COMP_RES_15_port <= '0';
   COMP_RES_16_port <= '0';
   COMP_RES_17_port <= '0';
   COMP_RES_18_port <= '0';
   COMP_RES_19_port <= '0';
   COMP_RES_20_port <= '0';
   COMP_RES_21_port <= '0';
   COMP_RES_22_port <= '0';
   COMP_RES_23_port <= '0';
   COMP_RES_24_port <= '0';
   COMP_RES_25_port <= '0';
   COMP_RES_26_port <= '0';
   COMP_RES_27_port <= '0';
   COMP_RES_28_port <= '0';
   COMP_RES_29_port <= '0';
   COMP_RES_30_port <= '0';
   COMP_RES_31_port <= '0';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_0 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_0;

architecture SYN_bhv of mux41_NBIT32_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n1, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n6, Z => n72);
   U2 : BUF_X1 port map( A => n6, Z => n73);
   U3 : BUF_X1 port map( A => n4, Z => n78);
   U4 : BUF_X1 port map( A => n4, Z => n79);
   U5 : BUF_X1 port map( A => n7, Z => n1);
   U6 : BUF_X1 port map( A => n7, Z => n70);
   U7 : BUF_X1 port map( A => n5, Z => n75);
   U8 : BUF_X1 port map( A => n5, Z => n76);
   U9 : BUF_X1 port map( A => n6, Z => n74);
   U10 : BUF_X1 port map( A => n4, Z => n80);
   U11 : BUF_X1 port map( A => n7, Z => n71);
   U12 : BUF_X1 port map( A => n5, Z => n77);
   U13 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n6);
   U14 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n7);
   U15 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n4);
   U16 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n5);
   U17 : INV_X1 port map( A => S(0), ZN => n81);
   U18 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => Z(0));
   U19 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n68);
   U20 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n69);
   U21 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => Z(20));
   U22 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => Z(24));
   U23 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => Z(17));
   U24 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n52);
   U25 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n53);
   U26 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => Z(13));
   U27 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n60);
   U28 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN 
                           => n61);
   U29 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => Z(6));
   U30 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n12);
   U31 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n13);
   U32 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => Z(31));
   U33 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN 
                           => n20);
   U34 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN 
                           => n21);
   U35 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => Z(28));
   U36 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n28);
   U37 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n29);
   U38 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => Z(10));
   U39 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => Z(21));
   U40 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n42);
   U41 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n43);
   U42 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => Z(18));
   U43 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n50);
   U44 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n51);
   U45 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => Z(14));
   U46 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n58);
   U47 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN 
                           => n59);
   U48 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => Z(7));
   U49 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n10);
   U50 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n11);
   U51 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => Z(3));
   U52 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN =>
                           n18);
   U53 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN =>
                           n19);
   U54 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => Z(29));
   U55 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n26);
   U56 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n27);
   U57 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => Z(25));
   U58 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n34);
   U59 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n35);
   U60 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Z(9));
   U61 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => Z(11));
   U62 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => Z(22));
   U63 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n40);
   U64 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n41);
   U65 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => Z(19));
   U66 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n48);
   U67 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN 
                           => n49);
   U68 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => Z(15));
   U69 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n56);
   U70 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN 
                           => n57);
   U71 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => Z(8));
   U72 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n8);
   U73 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n9);
   U74 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => Z(4));
   U75 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN =>
                           n16);
   U76 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN =>
                           n17);
   U77 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => Z(2));
   U78 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN =>
                           n24);
   U79 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN =>
                           n25);
   U80 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => Z(26));
   U81 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n32);
   U82 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n33);
   U83 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => Z(23));
   U84 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN 
                           => n38);
   U85 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN 
                           => n39);
   U86 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => Z(1));
   U87 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN => 
                           n46);
   U88 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN =>
                           n47);
   U89 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => Z(16));
   U90 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n54);
   U91 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n55);
   U92 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => Z(12));
   U93 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n62);
   U94 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN 
                           => n63);
   U95 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => Z(5));
   U96 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN =>
                           n14);
   U97 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN =>
                           n15);
   U98 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => Z(30));
   U99 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN 
                           => n22);
   U100 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN
                           => n23);
   U101 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => Z(27));
   U102 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN
                           => n30);
   U103 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN
                           => n31);
   U104 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n64);
   U105 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN
                           => n65);
   U106 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n66);
   U107 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN
                           => n67);
   U108 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN
                           => n44);
   U109 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN
                           => n45);
   U110 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN
                           => n36);
   U111 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN
                           => n37);
   U112 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN 
                           => n2);
   U113 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN 
                           => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FWD_Unit is

   port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB : in 
         std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;  
         FWDA, FWDB : out std_logic_vector (1 downto 0));

end FWD_Unit;

architecture SYN_bhv of FWD_Unit is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42 : std_logic;

begin
   
   U3 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => FWDB(1));
   U4 : AOI21_X1 port map( B1 => n3, B2 => n4, A => n5, ZN => n1);
   U5 : INV_X1 port map( A => n6, ZN => n3);
   U6 : NOR2_X1 port map( A1 => n2, A2 => n7, ZN => FWDB(0));
   U7 : MUX2_X1 port map( A => n6, B => n8, S => n5, Z => n7);
   U8 : AND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => n5);
   U9 : NOR2_X1 port map( A1 => n13, A2 => n14, ZN => n12);
   U10 : XOR2_X1 port map( A => ADD_WR_MEM(4), B => ADD_RS2(4), Z => n14);
   U11 : XOR2_X1 port map( A => ADD_WR_MEM(3), B => ADD_RS2(3), Z => n13);
   U12 : XNOR2_X1 port map( A => ADD_RS2(1), B => ADD_WR_MEM(1), ZN => n11);
   U13 : XNOR2_X1 port map( A => ADD_RS2(2), B => ADD_WR_MEM(2), ZN => n10);
   U14 : XNOR2_X1 port map( A => ADD_RS2(0), B => ADD_WR_MEM(0), ZN => n9);
   U15 : NAND4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           n6);
   U16 : NOR2_X1 port map( A1 => n19, A2 => n20, ZN => n18);
   U17 : XOR2_X1 port map( A => ADD_WR_WB(3), B => ADD_RS2(3), Z => n20);
   U18 : XOR2_X1 port map( A => ADD_WR_WB(2), B => ADD_RS2(2), Z => n19);
   U19 : XNOR2_X1 port map( A => ADD_RS2(4), B => ADD_WR_WB(4), ZN => n17);
   U20 : XNOR2_X1 port map( A => ADD_RS2(1), B => ADD_WR_WB(1), ZN => n16);
   U21 : XNOR2_X1 port map( A => ADD_RS2(0), B => ADD_WR_WB(0), ZN => n15);
   U22 : NOR2_X1 port map( A1 => n21, A2 => n2, ZN => FWDA(1));
   U23 : AOI21_X1 port map( B1 => n22, B2 => n4, A => n23, ZN => n21);
   U24 : OAI21_X1 port map( B1 => n24, B2 => n25, A => RF_WE_WB, ZN => n4);
   U25 : OR2_X1 port map( A1 => ADD_WR_WB(0), A2 => ADD_WR_WB(1), ZN => n25);
   U26 : OR3_X1 port map( A1 => ADD_WR_WB(3), A2 => ADD_WR_WB(4), A3 => 
                           ADD_WR_WB(2), ZN => n24);
   U27 : INV_X1 port map( A => n26, ZN => n22);
   U28 : NOR2_X1 port map( A1 => n2, A2 => n27, ZN => FWDA(0));
   U29 : MUX2_X1 port map( A => n26, B => n8, S => n23, Z => n27);
   U30 : AND4_X1 port map( A1 => n28, A2 => n29, A3 => n30, A4 => n31, ZN => 
                           n23);
   U31 : NOR2_X1 port map( A1 => n32, A2 => n33, ZN => n31);
   U32 : XOR2_X1 port map( A => ADD_WR_MEM(4), B => ADD_RS1(4), Z => n33);
   U33 : XOR2_X1 port map( A => ADD_WR_MEM(3), B => ADD_RS1(3), Z => n32);
   U34 : XNOR2_X1 port map( A => ADD_RS1(1), B => ADD_WR_MEM(1), ZN => n30);
   U35 : XNOR2_X1 port map( A => ADD_RS1(2), B => ADD_WR_MEM(2), ZN => n29);
   U36 : XNOR2_X1 port map( A => ADD_RS1(0), B => ADD_WR_MEM(0), ZN => n28);
   U37 : INV_X1 port map( A => n34, ZN => n8);
   U38 : OAI21_X1 port map( B1 => n35, B2 => n36, A => RF_WE_MEM, ZN => n34);
   U39 : OR2_X1 port map( A1 => ADD_WR_MEM(0), A2 => ADD_WR_MEM(1), ZN => n36);
   U40 : OR3_X1 port map( A1 => ADD_WR_MEM(3), A2 => ADD_WR_MEM(4), A3 => 
                           ADD_WR_MEM(2), ZN => n35);
   U41 : NAND4_X1 port map( A1 => n37, A2 => n38, A3 => n39, A4 => n40, ZN => 
                           n26);
   U42 : NOR2_X1 port map( A1 => n41, A2 => n42, ZN => n40);
   U43 : XOR2_X1 port map( A => ADD_WR_WB(3), B => ADD_RS1(3), Z => n42);
   U44 : XOR2_X1 port map( A => ADD_WR_WB(2), B => ADD_RS1(2), Z => n41);
   U45 : XNOR2_X1 port map( A => ADD_RS1(4), B => ADD_WR_WB(4), ZN => n39);
   U46 : XNOR2_X1 port map( A => ADD_RS1(1), B => ADD_WR_WB(1), ZN => n38);
   U47 : XNOR2_X1 port map( A => ADD_RS1(0), B => ADD_WR_WB(0), ZN => n37);
   U48 : INV_X1 port map( A => RST, ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N2 is

   port( DIN : in std_logic_vector (1 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (1 downto 0));

end regn_N2;

architecture SYN_bhv of regn_N2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   DOUT_reg_1_inst : DFFR_X1 port map( D => n6, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n4);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n5, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n3);
   U2 : OAI21_X1 port map( B1 => n3, B2 => EN, A => n1, ZN => n5);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n1);
   U4 : OAI21_X1 port map( B1 => n4, B2 => EN, A => n2, ZN => n6);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Branch_Cond_Unit_NBIT32 is

   port( RST : in std_logic;  A : in std_logic_vector (31 downto 0);  ALU_OPC :
         in std_logic_vector (0 to 4);  JUMP_TYPE : in std_logic_vector (1 
         downto 0);  PC_SEL : out std_logic_vector (1 downto 0);  ZERO : out 
         std_logic);

end Branch_Cond_Unit_NBIT32;

architecture SYN_bhv of Branch_Cond_Unit_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n1, n2 : std_logic;

begin
   
   U24 : NAND3_X1 port map( A1 => ALU_OPC(2), A2 => n7, A3 => ALU_OPC(1), ZN =>
                           n9);
   U25 : NAND3_X1 port map( A1 => ALU_OPC(1), A2 => ALU_OPC(2), A3 => n20, ZN 
                           => n7);
   U3 : NOR4_X1 port map( A1 => A(23), A2 => A(22), A3 => A(21), A4 => A(20), 
                           ZN => n15);
   U4 : NOR4_X1 port map( A1 => A(9), A2 => A(8), A3 => A(7), A4 => A(6), ZN =>
                           n19);
   U5 : NOR4_X1 port map( A1 => A(1), A2 => A(19), A3 => A(18), A4 => A(17), ZN
                           => n14);
   U6 : NOR4_X1 port map( A1 => A(5), A2 => A(4), A3 => A(3), A4 => A(31), ZN 
                           => n18);
   U7 : NOR4_X1 port map( A1 => A(16), A2 => A(15), A3 => A(14), A4 => A(13), 
                           ZN => n13);
   U8 : NOR4_X1 port map( A1 => A(30), A2 => A(2), A3 => A(29), A4 => A(28), ZN
                           => n17);
   U9 : NOR4_X1 port map( A1 => A(12), A2 => A(11), A3 => A(10), A4 => A(0), ZN
                           => n12);
   U10 : NOR2_X1 port map( A1 => n10, A2 => n11, ZN => n8);
   U11 : NAND4_X1 port map( A1 => n16, A2 => n17, A3 => n18, A4 => n19, ZN => 
                           n10);
   U12 : NAND4_X1 port map( A1 => n12, A2 => n13, A3 => n14, A4 => n15, ZN => 
                           n11);
   U13 : NOR4_X1 port map( A1 => A(27), A2 => A(26), A3 => A(25), A4 => A(24), 
                           ZN => n16);
   U14 : NOR3_X1 port map( A1 => ALU_OPC(4), A2 => ALU_OPC(0), A3 => ALU_OPC(3)
                           , ZN => n20);
   U15 : OAI211_X1 port map( C1 => n5, C2 => n6, A => JUMP_TYPE(0), B => RST, 
                           ZN => n4);
   U16 : NOR2_X1 port map( A1 => n7, A2 => n1, ZN => n6);
   U17 : NOR4_X1 port map( A1 => n9, A2 => n8, A3 => ALU_OPC(0), A4 => 
                           ALU_OPC(3), ZN => n5);
   U18 : INV_X1 port map( A => n8, ZN => n1);
   U19 : NAND2_X1 port map( A1 => JUMP_TYPE(1), A2 => RST, ZN => n3);
   U20 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => ZERO);
   U21 : OAI22_X1 port map( A1 => JUMP_TYPE(0), A2 => n3, B1 => JUMP_TYPE(1), 
                           B2 => n4, ZN => PC_SEL(0));
   U22 : NOR2_X1 port map( A1 => n2, A2 => n3, ZN => PC_SEL(1));
   U23 : INV_X1 port map( A => JUMP_TYPE(0), ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity register_file_NBIT_ADD5_NBIT_DATA32 is

   port( CLK, RST, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RS1, 
         ADD_RS2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_NBIT_ADD5_NBIT_DATA32;

architecture SYN_bhv of register_file_NBIT_ADD5_NBIT_DATA32 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n357, n358, n359, 
      n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, 
      n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, 
      n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, 
      n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, 
      n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, 
      n420, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, 
      n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, 
      n540, n541, n542, n543, n544, n545, n546, n547, n548, n613, n614, n615, 
      n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, 
      n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
      n640, n641, n642, n643, n644, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
      n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, 
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n864, n865, n866, n867, n868, n933, n934, n935, 
      n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, 
      n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, 
      n960, n961, n962, n963, n964, n2506, n2507, n2508, n2509, n2510, n2511, 
      n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, 
      n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, 
      n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, 
      n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, 
      n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, 
      n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, 
      n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, 
      n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, 
      n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, 
      n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, 
      n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, 
      n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, 
      n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, 
      n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, 
      n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, 
      n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, 
      n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, 
      n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, 
      n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, 
      n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, 
      n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, 
      n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, 
      n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, 
      n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, 
      n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, 
      n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, 
      n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, 
      n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, 
      n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, 
      n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, 
      n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, 
      n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, 
      n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, 
      n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, 
      n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, 
      n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, 
      n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, 
      n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, 
      n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, 
      n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, 
      n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, 
      n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, 
      n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, 
      n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, 
      n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, 
      n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, 
      n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, 
      n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, 
      n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, 
      n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, 
      n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, 
      n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, 
      n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, 
      n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, 
      n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, 
      n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, 
      n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, 
      n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, 
      n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, 
      n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, 
      n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, 
      n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, 
      n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, 
      n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, 
      n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, 
      n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, 
      n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, 
      n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, 
      n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, 
      n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, 
      n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, 
      n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, 
      n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, 
      n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, 
      n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, 
      n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, 
      n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, 
      n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, 
      n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, 
      n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, 
      n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, 
      n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, 
      n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, 
      n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, 
      n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, 
      n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, 
      n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, 
      n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, 
      n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, 
      n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, 
      n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, 
      n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, 
      n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, 
      n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, 
      n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, 
      n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, 
      n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, 
      n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, 
      n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, 
      n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, 
      n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, 
      n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, 
      n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, 
      n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, 
      n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n421, n422, n423, n424, n425, n426, n427, 
      n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
      n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, 
      n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n612, n645, n646, n647, 
      n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, 
      n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, 
      n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
      n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, 
      n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, 
      n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, 
      n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, 
      n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, 
      n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, 
      n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, 
      n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, 
      n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, 
      n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, 
      n804, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n965, n966, n967, n968, n969, n970, n971, 
      n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, 
      n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, 
      n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, 
      n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, 
      n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, 
      n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, 
      n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
      n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, 
      n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, 
      n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
      n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, 
      n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, 
      n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, 
      n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, 
      n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, 
      n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, 
      n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, 
      n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, 
      n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
      n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, 
      n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
      n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, 
      n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, 
      n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, 
      n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, 
      n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, 
      n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, 
      n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, 
      n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, 
      n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, 
      n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
      n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, 
      n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, 
      n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, 
      n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, 
      n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, 
      n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, 
      n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
      n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, 
      n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, 
      n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
      n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, 
      n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, 
      n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
      n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, 
      n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, 
      n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
      n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, 
      n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n3562, 
      n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, 
      n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, 
      n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, 
      n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, 
      n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, 
      n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, 
      n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, 
      n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, 
      n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, 
      n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, 
      n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, 
      n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, 
      n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, 
      n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, 
      n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, 
      n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, 
      n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, 
      n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, 
      n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, 
      n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, 
      n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, 
      n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, 
      n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, 
      n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, 
      n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, 
      n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, 
      n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, 
      n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, 
      n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, 
      n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, 
      n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, 
      n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, 
      n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, 
      n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, 
      n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, 
      n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, 
      n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, 
      n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, 
      n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, 
      n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, 
      n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, 
      n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, 
      n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, 
      n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, 
      n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, 
      n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, 
      n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, 
      n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, 
      n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, 
      n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, 
      n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, 
      n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, 
      n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, 
      n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, 
      n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, 
      n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, 
      n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, 
      n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, 
      n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, 
      n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, 
      n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, 
      n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, 
      n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, 
      n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, 
      n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, 
      n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, 
      n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, 
      n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, 
      n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, 
      n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, 
      n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, 
      n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, 
      n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, 
      n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, 
      n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, 
      n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, 
      n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, 
      n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, 
      n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, 
      n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, 
      n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, 
      n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, 
      n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, 
      n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, 
      n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, 
      n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, 
      n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, 
      n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, 
      n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, 
      n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, 
      n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, 
      n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, 
      n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, 
      n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, 
      n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, 
      n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, 
      n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, 
      n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, 
      n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, 
      n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, 
      n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, 
      n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, 
      n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, 
      n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, 
      n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, 
      n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, 
      n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, 
      n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, 
      n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, 
      n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, 
      n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, 
      n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, 
      n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, 
      n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, 
      n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, 
      n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, 
      n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, 
      n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, 
      n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, 
      n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, 
      n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, 
      n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, 
      n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, 
      n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, 
      n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, 
      n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, 
      n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, 
      n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, 
      n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, 
      n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, 
      n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, 
      n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, 
      n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, 
      n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, 
      n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, 
      n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, 
      n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, 
      n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, 
      n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, 
      n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, 
      n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, 
      n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, 
      n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, 
      n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, 
      n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, 
      n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, 
      n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, 
      n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, 
      n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, 
      n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, 
      n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, 
      n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, 
      n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, 
      n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, 
      n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, 
      n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, 
      n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, 
      n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, 
      n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, 
      n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, 
      n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, 
      n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, 
      n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, 
      n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, 
      n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, 
      n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, 
      n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, 
      n5233, n5234, n5235, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, 
      n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, 
      n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, 
      n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, 
      n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, 
      n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, 
      n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, 
      n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, 
      n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, 
      n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, 
      n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, 
      n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, 
      n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, 
      n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, 
      n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, 
      n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, 
      n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, 
      n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, 
      n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, 
      n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, 
      n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, 
      n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, 
      n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, 
      n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, 
      n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, 
      n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, 
      n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, 
      n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, 
      n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, 
      n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, 
      n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, 
      n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, 
      n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, 
      n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, 
      n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, 
      n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, 
      n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, 
      n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, 
      n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, 
      n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, 
      n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, 
      n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, 
      n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580 : 
      std_logic;

begin
   
   REGISTERS_reg_2_31_inst : DFFR_X1 port map( D => n3529, CK => CLK, RN => 
                           n1458, Q => n5235, QN => n_1197);
   REGISTERS_reg_2_30_inst : DFFR_X1 port map( D => n3528, CK => CLK, RN => 
                           n1458, Q => n5234, QN => n_1198);
   REGISTERS_reg_2_29_inst : DFFR_X1 port map( D => n3527, CK => CLK, RN => 
                           n1458, Q => n5233, QN => n_1199);
   REGISTERS_reg_2_28_inst : DFFR_X1 port map( D => n3526, CK => CLK, RN => 
                           n1458, Q => n5232, QN => n_1200);
   REGISTERS_reg_2_27_inst : DFFR_X1 port map( D => n3525, CK => CLK, RN => 
                           n1459, Q => n5231, QN => n_1201);
   REGISTERS_reg_2_26_inst : DFFR_X1 port map( D => n3524, CK => CLK, RN => 
                           n1459, Q => n5230, QN => n_1202);
   REGISTERS_reg_2_25_inst : DFFR_X1 port map( D => n3523, CK => CLK, RN => 
                           n1459, Q => n5229, QN => n_1203);
   REGISTERS_reg_2_24_inst : DFFR_X1 port map( D => n3522, CK => CLK, RN => 
                           n1459, Q => n5228, QN => n_1204);
   REGISTERS_reg_2_23_inst : DFFR_X1 port map( D => n3521, CK => CLK, RN => 
                           n1459, Q => n5227, QN => n_1205);
   REGISTERS_reg_2_22_inst : DFFR_X1 port map( D => n3520, CK => CLK, RN => 
                           n1459, Q => n5226, QN => n_1206);
   REGISTERS_reg_2_21_inst : DFFR_X1 port map( D => n3519, CK => CLK, RN => 
                           n1459, Q => n5225, QN => n_1207);
   REGISTERS_reg_2_20_inst : DFFR_X1 port map( D => n3518, CK => CLK, RN => 
                           n1459, Q => n5224, QN => n_1208);
   REGISTERS_reg_2_19_inst : DFFR_X1 port map( D => n3517, CK => CLK, RN => 
                           n1459, Q => n5223, QN => n_1209);
   REGISTERS_reg_2_18_inst : DFFR_X1 port map( D => n3516, CK => CLK, RN => 
                           n1459, Q => n5222, QN => n_1210);
   REGISTERS_reg_2_17_inst : DFFR_X1 port map( D => n3515, CK => CLK, RN => 
                           n1459, Q => n5221, QN => n_1211);
   REGISTERS_reg_2_16_inst : DFFR_X1 port map( D => n3514, CK => CLK, RN => 
                           n1459, Q => n5220, QN => n_1212);
   REGISTERS_reg_2_15_inst : DFFR_X1 port map( D => n3513, CK => CLK, RN => 
                           n1460, Q => n5219, QN => n_1213);
   REGISTERS_reg_2_14_inst : DFFR_X1 port map( D => n3512, CK => CLK, RN => 
                           n1460, Q => n5218, QN => n_1214);
   REGISTERS_reg_2_13_inst : DFFR_X1 port map( D => n3511, CK => CLK, RN => 
                           n1460, Q => n5217, QN => n_1215);
   REGISTERS_reg_2_12_inst : DFFR_X1 port map( D => n3510, CK => CLK, RN => 
                           n1460, Q => n5216, QN => n_1216);
   REGISTERS_reg_2_11_inst : DFFR_X1 port map( D => n3509, CK => CLK, RN => 
                           n1460, Q => n5215, QN => n_1217);
   REGISTERS_reg_2_10_inst : DFFR_X1 port map( D => n3508, CK => CLK, RN => 
                           n1460, Q => n5214, QN => n_1218);
   REGISTERS_reg_2_9_inst : DFFR_X1 port map( D => n3507, CK => CLK, RN => 
                           n1460, Q => n5213, QN => n_1219);
   REGISTERS_reg_2_8_inst : DFFR_X1 port map( D => n3506, CK => CLK, RN => 
                           n1460, Q => n5212, QN => n_1220);
   REGISTERS_reg_2_7_inst : DFFR_X1 port map( D => n3505, CK => CLK, RN => 
                           n1460, Q => n5211, QN => n_1221);
   REGISTERS_reg_2_6_inst : DFFR_X1 port map( D => n3504, CK => CLK, RN => 
                           n1460, Q => n5210, QN => n_1222);
   REGISTERS_reg_2_5_inst : DFFR_X1 port map( D => n3503, CK => CLK, RN => 
                           n1460, Q => n5209, QN => n_1223);
   REGISTERS_reg_2_4_inst : DFFR_X1 port map( D => n3502, CK => CLK, RN => 
                           n1460, Q => n5208, QN => n_1224);
   REGISTERS_reg_2_3_inst : DFFR_X1 port map( D => n3501, CK => CLK, RN => 
                           n1461, Q => n5207, QN => n_1225);
   REGISTERS_reg_2_2_inst : DFFR_X1 port map( D => n3500, CK => CLK, RN => 
                           n1461, Q => n5206, QN => n_1226);
   REGISTERS_reg_2_1_inst : DFFR_X1 port map( D => n3499, CK => CLK, RN => 
                           n1461, Q => n5205, QN => n_1227);
   REGISTERS_reg_2_0_inst : DFFR_X1 port map( D => n3498, CK => CLK, RN => 
                           n1461, Q => n5204, QN => n_1228);
   REGISTERS_reg_3_31_inst : DFFR_X1 port map( D => n3497, CK => CLK, RN => 
                           n1461, Q => n5203, QN => n2201);
   REGISTERS_reg_3_30_inst : DFFR_X1 port map( D => n3496, CK => CLK, RN => 
                           n1461, Q => n5202, QN => n2179);
   REGISTERS_reg_3_29_inst : DFFR_X1 port map( D => n3495, CK => CLK, RN => 
                           n1461, Q => n5201, QN => n2158);
   REGISTERS_reg_3_28_inst : DFFR_X1 port map( D => n3494, CK => CLK, RN => 
                           n1461, Q => n5200, QN => n2137);
   REGISTERS_reg_3_27_inst : DFFR_X1 port map( D => n3493, CK => CLK, RN => 
                           n1461, Q => n5199, QN => n2116);
   REGISTERS_reg_3_26_inst : DFFR_X1 port map( D => n3492, CK => CLK, RN => 
                           n1461, Q => n5198, QN => n2095);
   REGISTERS_reg_3_25_inst : DFFR_X1 port map( D => n3491, CK => CLK, RN => 
                           n1461, Q => n5197, QN => n2074);
   REGISTERS_reg_3_24_inst : DFFR_X1 port map( D => n3490, CK => CLK, RN => 
                           n1461, Q => n5196, QN => n2053);
   REGISTERS_reg_3_23_inst : DFFR_X1 port map( D => n3489, CK => CLK, RN => 
                           n1462, Q => n5195, QN => n2032);
   REGISTERS_reg_3_22_inst : DFFR_X1 port map( D => n3488, CK => CLK, RN => 
                           n1462, Q => n5194, QN => n2011);
   REGISTERS_reg_3_21_inst : DFFR_X1 port map( D => n3487, CK => CLK, RN => 
                           n1462, Q => n5193, QN => n1991);
   REGISTERS_reg_3_20_inst : DFFR_X1 port map( D => n3486, CK => CLK, RN => 
                           n1462, Q => n5192, QN => n1970);
   REGISTERS_reg_3_19_inst : DFFR_X1 port map( D => n3485, CK => CLK, RN => 
                           n1462, Q => n5191, QN => n1950);
   REGISTERS_reg_3_18_inst : DFFR_X1 port map( D => n3484, CK => CLK, RN => 
                           n1462, Q => n5190, QN => n1930);
   REGISTERS_reg_3_17_inst : DFFR_X1 port map( D => n3483, CK => CLK, RN => 
                           n1462, Q => n5189, QN => n1910);
   REGISTERS_reg_3_16_inst : DFFR_X1 port map( D => n3482, CK => CLK, RN => 
                           n1462, Q => n5188, QN => n1889);
   REGISTERS_reg_3_15_inst : DFFR_X1 port map( D => n3481, CK => CLK, RN => 
                           n1462, Q => n5187, QN => n1870);
   REGISTERS_reg_3_14_inst : DFFR_X1 port map( D => n3480, CK => CLK, RN => 
                           n1462, Q => n5186, QN => n1849);
   REGISTERS_reg_3_13_inst : DFFR_X1 port map( D => n3479, CK => CLK, RN => 
                           n1462, Q => n5185, QN => n1828);
   REGISTERS_reg_3_12_inst : DFFR_X1 port map( D => n3478, CK => CLK, RN => 
                           n1462, Q => n5184, QN => n1808);
   REGISTERS_reg_3_11_inst : DFFR_X1 port map( D => n3477, CK => CLK, RN => 
                           n1463, Q => n5183, QN => n1787);
   REGISTERS_reg_3_10_inst : DFFR_X1 port map( D => n3476, CK => CLK, RN => 
                           n1463, Q => n5182, QN => n1766);
   REGISTERS_reg_3_9_inst : DFFR_X1 port map( D => n3475, CK => CLK, RN => 
                           n1463, Q => n5181, QN => n1745);
   REGISTERS_reg_3_8_inst : DFFR_X1 port map( D => n3474, CK => CLK, RN => 
                           n1463, Q => n5180, QN => n1724);
   REGISTERS_reg_3_7_inst : DFFR_X1 port map( D => n3473, CK => CLK, RN => 
                           n1463, Q => n5179, QN => n1703);
   REGISTERS_reg_3_6_inst : DFFR_X1 port map( D => n3472, CK => CLK, RN => 
                           n1463, Q => n5178, QN => n1682);
   REGISTERS_reg_3_5_inst : DFFR_X1 port map( D => n3471, CK => CLK, RN => 
                           n1463, Q => n5177, QN => n1661);
   REGISTERS_reg_3_4_inst : DFFR_X1 port map( D => n3470, CK => CLK, RN => 
                           n1463, Q => n5176, QN => n1640);
   REGISTERS_reg_3_3_inst : DFFR_X1 port map( D => n3469, CK => CLK, RN => 
                           n1463, Q => n5175, QN => n1620);
   REGISTERS_reg_3_2_inst : DFFR_X1 port map( D => n3468, CK => CLK, RN => 
                           n1463, Q => n5174, QN => n1601);
   REGISTERS_reg_3_1_inst : DFFR_X1 port map( D => n3467, CK => CLK, RN => 
                           n1463, Q => n5173, QN => n1581);
   REGISTERS_reg_3_0_inst : DFFR_X1 port map( D => n3466, CK => CLK, RN => 
                           n1463, Q => n5172, QN => n1556);
   REGISTERS_reg_6_31_inst : DFFR_X1 port map( D => n3401, CK => CLK, RN => 
                           n1469, Q => n5171, QN => n2215);
   REGISTERS_reg_6_30_inst : DFFR_X1 port map( D => n3400, CK => CLK, RN => 
                           n1469, Q => n5170, QN => n2185);
   REGISTERS_reg_6_29_inst : DFFR_X1 port map( D => n3399, CK => CLK, RN => 
                           n1469, Q => n5169, QN => n2164);
   REGISTERS_reg_6_28_inst : DFFR_X1 port map( D => n3398, CK => CLK, RN => 
                           n1469, Q => n5168, QN => n2143);
   REGISTERS_reg_6_27_inst : DFFR_X1 port map( D => n3397, CK => CLK, RN => 
                           n1469, Q => n5167, QN => n2122);
   REGISTERS_reg_6_26_inst : DFFR_X1 port map( D => n3396, CK => CLK, RN => 
                           n1469, Q => n5166, QN => n2101);
   REGISTERS_reg_6_25_inst : DFFR_X1 port map( D => n3395, CK => CLK, RN => 
                           n1469, Q => n5165, QN => n2080);
   REGISTERS_reg_6_24_inst : DFFR_X1 port map( D => n3394, CK => CLK, RN => 
                           n1469, Q => n5164, QN => n2059);
   REGISTERS_reg_6_23_inst : DFFR_X1 port map( D => n3393, CK => CLK, RN => 
                           n1470, Q => n5163, QN => n2038);
   REGISTERS_reg_6_22_inst : DFFR_X1 port map( D => n3392, CK => CLK, RN => 
                           n1470, Q => n5162, QN => n2017);
   REGISTERS_reg_6_21_inst : DFFR_X1 port map( D => n3391, CK => CLK, RN => 
                           n1470, Q => n5161, QN => n1997);
   REGISTERS_reg_6_20_inst : DFFR_X1 port map( D => n3390, CK => CLK, RN => 
                           n1470, Q => n5160, QN => n1976);
   REGISTERS_reg_6_19_inst : DFFR_X1 port map( D => n3389, CK => CLK, RN => 
                           n1470, Q => n5159, QN => n1956);
   REGISTERS_reg_6_18_inst : DFFR_X1 port map( D => n3388, CK => CLK, RN => 
                           n1470, Q => n5158, QN => n1936);
   REGISTERS_reg_6_17_inst : DFFR_X1 port map( D => n3387, CK => CLK, RN => 
                           n1470, Q => n5157, QN => n1916);
   REGISTERS_reg_6_16_inst : DFFR_X1 port map( D => n3386, CK => CLK, RN => 
                           n1470, Q => n5156, QN => n1895);
   REGISTERS_reg_6_15_inst : DFFR_X1 port map( D => n3385, CK => CLK, RN => 
                           n1470, Q => n5155, QN => n1874);
   REGISTERS_reg_6_14_inst : DFFR_X1 port map( D => n3384, CK => CLK, RN => 
                           n1470, Q => n5154, QN => n1855);
   REGISTERS_reg_6_13_inst : DFFR_X1 port map( D => n3383, CK => CLK, RN => 
                           n1470, Q => n5153, QN => n1834);
   REGISTERS_reg_6_12_inst : DFFR_X1 port map( D => n3382, CK => CLK, RN => 
                           n1470, Q => n5152, QN => n1814);
   REGISTERS_reg_6_11_inst : DFFR_X1 port map( D => n3381, CK => CLK, RN => 
                           n1471, Q => n5151, QN => n1793);
   REGISTERS_reg_6_10_inst : DFFR_X1 port map( D => n3380, CK => CLK, RN => 
                           n1471, Q => n5150, QN => n1772);
   REGISTERS_reg_6_9_inst : DFFR_X1 port map( D => n3379, CK => CLK, RN => 
                           n1471, Q => n5149, QN => n1751);
   REGISTERS_reg_6_8_inst : DFFR_X1 port map( D => n3378, CK => CLK, RN => 
                           n1471, Q => n5148, QN => n1730);
   REGISTERS_reg_6_7_inst : DFFR_X1 port map( D => n3377, CK => CLK, RN => 
                           n1471, Q => n5147, QN => n1709);
   REGISTERS_reg_6_6_inst : DFFR_X1 port map( D => n3376, CK => CLK, RN => 
                           n1471, Q => n5146, QN => n1688);
   REGISTERS_reg_6_5_inst : DFFR_X1 port map( D => n3375, CK => CLK, RN => 
                           n1471, Q => n5145, QN => n1667);
   REGISTERS_reg_6_4_inst : DFFR_X1 port map( D => n3374, CK => CLK, RN => 
                           n1471, Q => n5144, QN => n1646);
   REGISTERS_reg_6_3_inst : DFFR_X1 port map( D => n3373, CK => CLK, RN => 
                           n1471, Q => n5143, QN => n1626);
   REGISTERS_reg_6_2_inst : DFFR_X1 port map( D => n3372, CK => CLK, RN => 
                           n1471, Q => n5142, QN => n1605);
   REGISTERS_reg_6_1_inst : DFFR_X1 port map( D => n3371, CK => CLK, RN => 
                           n1471, Q => n5141, QN => n1587);
   REGISTERS_reg_6_0_inst : DFFR_X1 port map( D => n3370, CK => CLK, RN => 
                           n1471, Q => n5140, QN => n1564);
   REGISTERS_reg_7_31_inst : DFFR_X1 port map( D => n3369, CK => CLK, RN => 
                           n1472, Q => n5139, QN => n_1229);
   REGISTERS_reg_7_30_inst : DFFR_X1 port map( D => n3368, CK => CLK, RN => 
                           n1472, Q => n5138, QN => n_1230);
   REGISTERS_reg_7_29_inst : DFFR_X1 port map( D => n3367, CK => CLK, RN => 
                           n1472, Q => n5137, QN => n_1231);
   REGISTERS_reg_7_28_inst : DFFR_X1 port map( D => n3366, CK => CLK, RN => 
                           n1472, Q => n5136, QN => n_1232);
   REGISTERS_reg_7_27_inst : DFFR_X1 port map( D => n3365, CK => CLK, RN => 
                           n1472, Q => n5135, QN => n_1233);
   REGISTERS_reg_7_26_inst : DFFR_X1 port map( D => n3364, CK => CLK, RN => 
                           n1472, Q => n5134, QN => n_1234);
   REGISTERS_reg_7_25_inst : DFFR_X1 port map( D => n3363, CK => CLK, RN => 
                           n1472, Q => n5133, QN => n_1235);
   REGISTERS_reg_7_24_inst : DFFR_X1 port map( D => n3362, CK => CLK, RN => 
                           n1472, Q => n5132, QN => n_1236);
   REGISTERS_reg_7_23_inst : DFFR_X1 port map( D => n3361, CK => CLK, RN => 
                           n1472, Q => n5131, QN => n_1237);
   REGISTERS_reg_7_22_inst : DFFR_X1 port map( D => n3360, CK => CLK, RN => 
                           n1472, Q => n5130, QN => n_1238);
   REGISTERS_reg_7_21_inst : DFFR_X1 port map( D => n3359, CK => CLK, RN => 
                           n1472, Q => n5129, QN => n_1239);
   REGISTERS_reg_7_20_inst : DFFR_X1 port map( D => n3358, CK => CLK, RN => 
                           n1472, Q => n5128, QN => n_1240);
   REGISTERS_reg_7_19_inst : DFFR_X1 port map( D => n3357, CK => CLK, RN => 
                           n1473, Q => n5127, QN => n_1241);
   REGISTERS_reg_7_18_inst : DFFR_X1 port map( D => n3356, CK => CLK, RN => 
                           n1473, Q => n5126, QN => n_1242);
   REGISTERS_reg_7_17_inst : DFFR_X1 port map( D => n3355, CK => CLK, RN => 
                           n1473, Q => n5125, QN => n_1243);
   REGISTERS_reg_7_16_inst : DFFR_X1 port map( D => n3354, CK => CLK, RN => 
                           n1473, Q => n5124, QN => n_1244);
   REGISTERS_reg_7_15_inst : DFFR_X1 port map( D => n3353, CK => CLK, RN => 
                           n1473, Q => n5123, QN => n_1245);
   REGISTERS_reg_7_14_inst : DFFR_X1 port map( D => n3352, CK => CLK, RN => 
                           n1473, Q => n5122, QN => n_1246);
   REGISTERS_reg_7_13_inst : DFFR_X1 port map( D => n3351, CK => CLK, RN => 
                           n1473, Q => n5121, QN => n_1247);
   REGISTERS_reg_7_12_inst : DFFR_X1 port map( D => n3350, CK => CLK, RN => 
                           n1473, Q => n5120, QN => n_1248);
   REGISTERS_reg_7_11_inst : DFFR_X1 port map( D => n3349, CK => CLK, RN => 
                           n1473, Q => n5119, QN => n_1249);
   REGISTERS_reg_7_10_inst : DFFR_X1 port map( D => n3348, CK => CLK, RN => 
                           n1473, Q => n5118, QN => n_1250);
   REGISTERS_reg_7_9_inst : DFFR_X1 port map( D => n3347, CK => CLK, RN => 
                           n1473, Q => n5117, QN => n_1251);
   REGISTERS_reg_7_8_inst : DFFR_X1 port map( D => n3346, CK => CLK, RN => 
                           n1473, Q => n5116, QN => n_1252);
   REGISTERS_reg_7_7_inst : DFFR_X1 port map( D => n3345, CK => CLK, RN => 
                           n1474, Q => n5115, QN => n_1253);
   REGISTERS_reg_7_6_inst : DFFR_X1 port map( D => n3344, CK => CLK, RN => 
                           n1474, Q => n5114, QN => n_1254);
   REGISTERS_reg_7_5_inst : DFFR_X1 port map( D => n3343, CK => CLK, RN => 
                           n1474, Q => n5113, QN => n_1255);
   REGISTERS_reg_7_4_inst : DFFR_X1 port map( D => n3342, CK => CLK, RN => 
                           n1474, Q => n5112, QN => n_1256);
   REGISTERS_reg_7_3_inst : DFFR_X1 port map( D => n3341, CK => CLK, RN => 
                           n1474, Q => n5111, QN => n_1257);
   REGISTERS_reg_7_2_inst : DFFR_X1 port map( D => n3340, CK => CLK, RN => 
                           n1474, Q => n5110, QN => n_1258);
   REGISTERS_reg_7_1_inst : DFFR_X1 port map( D => n3339, CK => CLK, RN => 
                           n1474, Q => n5109, QN => n_1259);
   REGISTERS_reg_7_0_inst : DFFR_X1 port map( D => n3338, CK => CLK, RN => 
                           n1474, Q => n5108, QN => n_1260);
   REGISTERS_reg_8_23_inst : DFFR_X1 port map( D => n3329, CK => CLK, RN => 
                           n1475, Q => n_1261, QN => n237);
   REGISTERS_reg_8_22_inst : DFFR_X1 port map( D => n3328, CK => CLK, RN => 
                           n1475, Q => n_1262, QN => n238);
   REGISTERS_reg_8_20_inst : DFFR_X1 port map( D => n3326, CK => CLK, RN => 
                           n1475, Q => n_1263, QN => n240);
   REGISTERS_reg_8_19_inst : DFFR_X1 port map( D => n3325, CK => CLK, RN => 
                           n1475, Q => n_1264, QN => n241);
   REGISTERS_reg_8_18_inst : DFFR_X1 port map( D => n3324, CK => CLK, RN => 
                           n1475, Q => n_1265, QN => n242);
   REGISTERS_reg_8_17_inst : DFFR_X1 port map( D => n3323, CK => CLK, RN => 
                           n1475, Q => n_1266, QN => n243);
   REGISTERS_reg_8_16_inst : DFFR_X1 port map( D => n3322, CK => CLK, RN => 
                           n1475, Q => n_1267, QN => n244);
   REGISTERS_reg_8_15_inst : DFFR_X1 port map( D => n3321, CK => CLK, RN => 
                           n1476, Q => n_1268, QN => n245);
   REGISTERS_reg_8_14_inst : DFFR_X1 port map( D => n3320, CK => CLK, RN => 
                           n1476, Q => n_1269, QN => n246);
   REGISTERS_reg_8_13_inst : DFFR_X1 port map( D => n3319, CK => CLK, RN => 
                           n1476, Q => n_1270, QN => n247);
   REGISTERS_reg_8_12_inst : DFFR_X1 port map( D => n3318, CK => CLK, RN => 
                           n1476, Q => n_1271, QN => n248);
   REGISTERS_reg_8_11_inst : DFFR_X1 port map( D => n3317, CK => CLK, RN => 
                           n1476, Q => n_1272, QN => n249);
   REGISTERS_reg_8_10_inst : DFFR_X1 port map( D => n3316, CK => CLK, RN => 
                           n1476, Q => n_1273, QN => n250);
   REGISTERS_reg_8_9_inst : DFFR_X1 port map( D => n3315, CK => CLK, RN => 
                           n1476, Q => n_1274, QN => n251);
   REGISTERS_reg_8_8_inst : DFFR_X1 port map( D => n3314, CK => CLK, RN => 
                           n1476, Q => n_1275, QN => n252);
   REGISTERS_reg_8_7_inst : DFFR_X1 port map( D => n3313, CK => CLK, RN => 
                           n1476, Q => n_1276, QN => n253);
   REGISTERS_reg_8_5_inst : DFFR_X1 port map( D => n3311, CK => CLK, RN => 
                           n1476, Q => n_1277, QN => n255);
   REGISTERS_reg_8_4_inst : DFFR_X1 port map( D => n3310, CK => CLK, RN => 
                           n1476, Q => n_1278, QN => n256);
   REGISTERS_reg_8_3_inst : DFFR_X1 port map( D => n3309, CK => CLK, RN => 
                           n1477, Q => n_1279, QN => n257);
   REGISTERS_reg_8_2_inst : DFFR_X1 port map( D => n3308, CK => CLK, RN => 
                           n1477, Q => n_1280, QN => n258);
   REGISTERS_reg_8_1_inst : DFFR_X1 port map( D => n3307, CK => CLK, RN => 
                           n1477, Q => n_1281, QN => n259);
   REGISTERS_reg_8_0_inst : DFFR_X1 port map( D => n3306, CK => CLK, RN => 
                           n1477, Q => n_1282, QN => n260);
   REGISTERS_reg_9_23_inst : DFFR_X1 port map( D => n3297, CK => CLK, RN => 
                           n1478, Q => n212, QN => n269);
   REGISTERS_reg_9_22_inst : DFFR_X1 port map( D => n3296, CK => CLK, RN => 
                           n1478, Q => n211, QN => n270);
   REGISTERS_reg_9_21_inst : DFFR_X1 port map( D => n3295, CK => CLK, RN => 
                           n1478, Q => n210, QN => n271);
   REGISTERS_reg_9_20_inst : DFFR_X1 port map( D => n3294, CK => CLK, RN => 
                           n1478, Q => n209, QN => n272);
   REGISTERS_reg_9_19_inst : DFFR_X1 port map( D => n3293, CK => CLK, RN => 
                           n1478, Q => n208, QN => n273);
   REGISTERS_reg_9_18_inst : DFFR_X1 port map( D => n3292, CK => CLK, RN => 
                           n1478, Q => n207, QN => n274);
   REGISTERS_reg_9_17_inst : DFFR_X1 port map( D => n3291, CK => CLK, RN => 
                           n1478, Q => n206, QN => n275);
   REGISTERS_reg_9_16_inst : DFFR_X1 port map( D => n3290, CK => CLK, RN => 
                           n1478, Q => n205, QN => n276);
   REGISTERS_reg_9_15_inst : DFFR_X1 port map( D => n3289, CK => CLK, RN => 
                           n1478, Q => n204, QN => n277);
   REGISTERS_reg_9_14_inst : DFFR_X1 port map( D => n3288, CK => CLK, RN => 
                           n1478, Q => n217, QN => n278);
   REGISTERS_reg_9_13_inst : DFFR_X1 port map( D => n3287, CK => CLK, RN => 
                           n1478, Q => n216, QN => n279);
   REGISTERS_reg_9_12_inst : DFFR_X1 port map( D => n3286, CK => CLK, RN => 
                           n1478, Q => n215, QN => n280);
   REGISTERS_reg_9_11_inst : DFFR_X1 port map( D => n3285, CK => CLK, RN => 
                           n1479, Q => n214, QN => n281);
   REGISTERS_reg_9_10_inst : DFFR_X1 port map( D => n3284, CK => CLK, RN => 
                           n1479, Q => n203, QN => n282);
   REGISTERS_reg_9_9_inst : DFFR_X1 port map( D => n3283, CK => CLK, RN => 
                           n1479, Q => n213, QN => n283);
   REGISTERS_reg_9_8_inst : DFFR_X1 port map( D => n3282, CK => CLK, RN => 
                           n1479, Q => n202, QN => n284);
   REGISTERS_reg_9_7_inst : DFFR_X1 port map( D => n3281, CK => CLK, RN => 
                           n1479, Q => n201, QN => n285);
   REGISTERS_reg_9_6_inst : DFFR_X1 port map( D => n3280, CK => CLK, RN => 
                           n1479, Q => n200, QN => n286);
   REGISTERS_reg_9_5_inst : DFFR_X1 port map( D => n3279, CK => CLK, RN => 
                           n1479, Q => n199, QN => n287);
   REGISTERS_reg_9_4_inst : DFFR_X1 port map( D => n3278, CK => CLK, RN => 
                           n1479, Q => n198, QN => n288);
   REGISTERS_reg_9_3_inst : DFFR_X1 port map( D => n3277, CK => CLK, RN => 
                           n1479, Q => n197, QN => n289);
   REGISTERS_reg_9_2_inst : DFFR_X1 port map( D => n3276, CK => CLK, RN => 
                           n1479, Q => n196, QN => n290);
   REGISTERS_reg_9_1_inst : DFFR_X1 port map( D => n3275, CK => CLK, RN => 
                           n1479, Q => n195, QN => n291);
   REGISTERS_reg_9_0_inst : DFFR_X1 port map( D => n3274, CK => CLK, RN => 
                           n1479, Q => n194, QN => n292);
   REGISTERS_reg_10_31_inst : DFFR_X1 port map( D => n3273, CK => CLK, RN => 
                           n1480, Q => n5107, QN => n193);
   REGISTERS_reg_10_30_inst : DFFR_X1 port map( D => n3272, CK => CLK, RN => 
                           n1480, Q => n5106, QN => n192);
   REGISTERS_reg_10_29_inst : DFFR_X1 port map( D => n3271, CK => CLK, RN => 
                           n1480, Q => n5105, QN => n191);
   REGISTERS_reg_10_28_inst : DFFR_X1 port map( D => n3270, CK => CLK, RN => 
                           n1480, Q => n5104, QN => n190);
   REGISTERS_reg_10_27_inst : DFFR_X1 port map( D => n3269, CK => CLK, RN => 
                           n1480, Q => n5103, QN => n189);
   REGISTERS_reg_10_26_inst : DFFR_X1 port map( D => n3268, CK => CLK, RN => 
                           n1480, Q => n5102, QN => n188);
   REGISTERS_reg_10_25_inst : DFFR_X1 port map( D => n3267, CK => CLK, RN => 
                           n1480, Q => n5101, QN => n187);
   REGISTERS_reg_10_24_inst : DFFR_X1 port map( D => n3266, CK => CLK, RN => 
                           n1480, Q => n5100, QN => n186);
   REGISTERS_reg_10_23_inst : DFFR_X1 port map( D => n3265, CK => CLK, RN => 
                           n1480, Q => n5099, QN => n185);
   REGISTERS_reg_10_22_inst : DFFR_X1 port map( D => n3264, CK => CLK, RN => 
                           n1480, Q => n5098, QN => n441);
   REGISTERS_reg_10_21_inst : DFFR_X1 port map( D => n3263, CK => CLK, RN => 
                           n1480, Q => n5097, QN => n443);
   REGISTERS_reg_10_20_inst : DFFR_X1 port map( D => n3262, CK => CLK, RN => 
                           n1480, Q => n5096, QN => n453);
   REGISTERS_reg_10_19_inst : DFFR_X1 port map( D => n3261, CK => CLK, RN => 
                           n1481, Q => n5095, QN => n455);
   REGISTERS_reg_10_18_inst : DFFR_X1 port map( D => n3260, CK => CLK, RN => 
                           n1481, Q => n5094, QN => n184);
   REGISTERS_reg_10_17_inst : DFFR_X1 port map( D => n3259, CK => CLK, RN => 
                           n1481, Q => n5093, QN => n445);
   REGISTERS_reg_10_16_inst : DFFR_X1 port map( D => n3258, CK => CLK, RN => 
                           n1481, Q => n5092, QN => n447);
   REGISTERS_reg_10_15_inst : DFFR_X1 port map( D => n3257, CK => CLK, RN => 
                           n1481, Q => n5091, QN => n183);
   REGISTERS_reg_10_14_inst : DFFR_X1 port map( D => n3256, CK => CLK, RN => 
                           n1481, Q => n5090, QN => n182);
   REGISTERS_reg_10_13_inst : DFFR_X1 port map( D => n3255, CK => CLK, RN => 
                           n1481, Q => n5089, QN => n457);
   REGISTERS_reg_10_12_inst : DFFR_X1 port map( D => n3254, CK => CLK, RN => 
                           n1481, Q => n5088, QN => n181);
   REGISTERS_reg_10_11_inst : DFFR_X1 port map( D => n3253, CK => CLK, RN => 
                           n1481, Q => n5087, QN => n459);
   REGISTERS_reg_10_10_inst : DFFR_X1 port map( D => n3252, CK => CLK, RN => 
                           n1481, Q => n5086, QN => n180);
   REGISTERS_reg_10_9_inst : DFFR_X1 port map( D => n3251, CK => CLK, RN => 
                           n1481, Q => n5085, QN => n179);
   REGISTERS_reg_10_8_inst : DFFR_X1 port map( D => n3250, CK => CLK, RN => 
                           n1481, Q => n5084, QN => n178);
   REGISTERS_reg_10_7_inst : DFFR_X1 port map( D => n3249, CK => CLK, RN => 
                           n1482, Q => n5083, QN => n177);
   REGISTERS_reg_10_6_inst : DFFR_X1 port map( D => n3248, CK => CLK, RN => 
                           n1482, Q => n5082, QN => n176);
   REGISTERS_reg_10_5_inst : DFFR_X1 port map( D => n3247, CK => CLK, RN => 
                           n1482, Q => n5081, QN => n175);
   REGISTERS_reg_10_4_inst : DFFR_X1 port map( D => n3246, CK => CLK, RN => 
                           n1482, Q => n5080, QN => n449);
   REGISTERS_reg_10_3_inst : DFFR_X1 port map( D => n3245, CK => CLK, RN => 
                           n1482, Q => n5079, QN => n174);
   REGISTERS_reg_10_2_inst : DFFR_X1 port map( D => n3244, CK => CLK, RN => 
                           n1482, Q => n5078, QN => n173);
   REGISTERS_reg_10_1_inst : DFFR_X1 port map( D => n3243, CK => CLK, RN => 
                           n1482, Q => n5077, QN => n439);
   REGISTERS_reg_10_0_inst : DFFR_X1 port map( D => n3242, CK => CLK, RN => 
                           n1482, Q => n5076, QN => n451);
   REGISTERS_reg_11_31_inst : DFFR_X1 port map( D => n3241, CK => CLK, RN => 
                           n1482, Q => n5075, QN => n342);
   REGISTERS_reg_11_30_inst : DFFR_X1 port map( D => n3240, CK => CLK, RN => 
                           n1482, Q => n5074, QN => n341);
   REGISTERS_reg_11_29_inst : DFFR_X1 port map( D => n3239, CK => CLK, RN => 
                           n1482, Q => n5073, QN => n340);
   REGISTERS_reg_11_28_inst : DFFR_X1 port map( D => n3238, CK => CLK, RN => 
                           n1482, Q => n5072, QN => n339);
   REGISTERS_reg_11_27_inst : DFFR_X1 port map( D => n3237, CK => CLK, RN => 
                           n1483, Q => n5071, QN => n338);
   REGISTERS_reg_11_26_inst : DFFR_X1 port map( D => n3236, CK => CLK, RN => 
                           n1483, Q => n5070, QN => n337);
   REGISTERS_reg_11_25_inst : DFFR_X1 port map( D => n3235, CK => CLK, RN => 
                           n1483, Q => n5069, QN => n336);
   REGISTERS_reg_11_24_inst : DFFR_X1 port map( D => n3234, CK => CLK, RN => 
                           n1483, Q => n5068, QN => n335);
   REGISTERS_reg_11_23_inst : DFFR_X1 port map( D => n3233, CK => CLK, RN => 
                           n1483, Q => n5067, QN => n334);
   REGISTERS_reg_11_22_inst : DFFR_X1 port map( D => n3232, CK => CLK, RN => 
                           n1483, Q => n5066, QN => n442);
   REGISTERS_reg_11_21_inst : DFFR_X1 port map( D => n3231, CK => CLK, RN => 
                           n1483, Q => n5065, QN => n444);
   REGISTERS_reg_11_20_inst : DFFR_X1 port map( D => n3230, CK => CLK, RN => 
                           n1483, Q => n5064, QN => n454);
   REGISTERS_reg_11_19_inst : DFFR_X1 port map( D => n3229, CK => CLK, RN => 
                           n1483, Q => n5063, QN => n456);
   REGISTERS_reg_11_18_inst : DFFR_X1 port map( D => n3228, CK => CLK, RN => 
                           n1483, Q => n5062, QN => n333);
   REGISTERS_reg_11_17_inst : DFFR_X1 port map( D => n3227, CK => CLK, RN => 
                           n1483, Q => n5061, QN => n446);
   REGISTERS_reg_11_16_inst : DFFR_X1 port map( D => n3226, CK => CLK, RN => 
                           n1483, Q => n5060, QN => n448);
   REGISTERS_reg_11_15_inst : DFFR_X1 port map( D => n3225, CK => CLK, RN => 
                           n1484, Q => n5059, QN => n332);
   REGISTERS_reg_11_14_inst : DFFR_X1 port map( D => n3224, CK => CLK, RN => 
                           n1484, Q => n5058, QN => n331);
   REGISTERS_reg_11_13_inst : DFFR_X1 port map( D => n3223, CK => CLK, RN => 
                           n1484, Q => n5057, QN => n458);
   REGISTERS_reg_11_12_inst : DFFR_X1 port map( D => n3222, CK => CLK, RN => 
                           n1484, Q => n5056, QN => n330);
   REGISTERS_reg_11_11_inst : DFFR_X1 port map( D => n3221, CK => CLK, RN => 
                           n1484, Q => n5055, QN => n460);
   REGISTERS_reg_11_10_inst : DFFR_X1 port map( D => n3220, CK => CLK, RN => 
                           n1484, Q => n5054, QN => n329);
   REGISTERS_reg_11_9_inst : DFFR_X1 port map( D => n3219, CK => CLK, RN => 
                           n1484, Q => n5053, QN => n328);
   REGISTERS_reg_11_8_inst : DFFR_X1 port map( D => n3218, CK => CLK, RN => 
                           n1484, Q => n5052, QN => n327);
   REGISTERS_reg_11_7_inst : DFFR_X1 port map( D => n3217, CK => CLK, RN => 
                           n1484, Q => n5051, QN => n326);
   REGISTERS_reg_11_6_inst : DFFR_X1 port map( D => n3216, CK => CLK, RN => 
                           n1484, Q => n5050, QN => n325);
   REGISTERS_reg_11_5_inst : DFFR_X1 port map( D => n3215, CK => CLK, RN => 
                           n1484, Q => n5049, QN => n324);
   REGISTERS_reg_11_4_inst : DFFR_X1 port map( D => n3214, CK => CLK, RN => 
                           n1484, Q => n5048, QN => n450);
   REGISTERS_reg_11_3_inst : DFFR_X1 port map( D => n3213, CK => CLK, RN => 
                           n1485, Q => n5047, QN => n323);
   REGISTERS_reg_11_2_inst : DFFR_X1 port map( D => n3212, CK => CLK, RN => 
                           n1485, Q => n5046, QN => n322);
   REGISTERS_reg_11_1_inst : DFFR_X1 port map( D => n3211, CK => CLK, RN => 
                           n1485, Q => n5045, QN => n440);
   REGISTERS_reg_11_0_inst : DFFR_X1 port map( D => n3210, CK => CLK, RN => 
                           n1485, Q => n5044, QN => n452);
   REGISTERS_reg_12_23_inst : DFFR_X1 port map( D => n3201, CK => CLK, RN => 
                           n1486, Q => n2036, QN => n365);
   REGISTERS_reg_12_22_inst : DFFR_X1 port map( D => n3200, CK => CLK, RN => 
                           n1486, Q => n2015, QN => n366);
   REGISTERS_reg_12_21_inst : DFFR_X1 port map( D => n3199, CK => CLK, RN => 
                           n1486, Q => n1995, QN => n367);
   REGISTERS_reg_12_20_inst : DFFR_X1 port map( D => n3198, CK => CLK, RN => 
                           n1486, Q => n1974, QN => n368);
   REGISTERS_reg_12_19_inst : DFFR_X1 port map( D => n3197, CK => CLK, RN => 
                           n1486, Q => n1954, QN => n369);
   REGISTERS_reg_12_18_inst : DFFR_X1 port map( D => n3196, CK => CLK, RN => 
                           n1486, Q => n1934, QN => n370);
   REGISTERS_reg_12_17_inst : DFFR_X1 port map( D => n3195, CK => CLK, RN => 
                           n1486, Q => n1914, QN => n371);
   REGISTERS_reg_12_16_inst : DFFR_X1 port map( D => n3194, CK => CLK, RN => 
                           n1486, Q => n1893, QN => n372);
   REGISTERS_reg_12_15_inst : DFFR_X1 port map( D => n3193, CK => CLK, RN => 
                           n1486, Q => n221, QN => n373);
   REGISTERS_reg_12_14_inst : DFFR_X1 port map( D => n3192, CK => CLK, RN => 
                           n1486, Q => n1853, QN => n374);
   REGISTERS_reg_12_13_inst : DFFR_X1 port map( D => n3191, CK => CLK, RN => 
                           n1486, Q => n1832, QN => n375);
   REGISTERS_reg_12_12_inst : DFFR_X1 port map( D => n3190, CK => CLK, RN => 
                           n1486, Q => n1812, QN => n376);
   REGISTERS_reg_12_11_inst : DFFR_X1 port map( D => n3189, CK => CLK, RN => 
                           n1487, Q => n1791, QN => n377);
   REGISTERS_reg_12_10_inst : DFFR_X1 port map( D => n3188, CK => CLK, RN => 
                           n1487, Q => n1770, QN => n378);
   REGISTERS_reg_12_9_inst : DFFR_X1 port map( D => n3187, CK => CLK, RN => 
                           n1487, Q => n1749, QN => n379);
   REGISTERS_reg_12_8_inst : DFFR_X1 port map( D => n3186, CK => CLK, RN => 
                           n1487, Q => n1728, QN => n380);
   REGISTERS_reg_12_7_inst : DFFR_X1 port map( D => n3185, CK => CLK, RN => 
                           n1487, Q => n1707, QN => n381);
   REGISTERS_reg_12_6_inst : DFFR_X1 port map( D => n3184, CK => CLK, RN => 
                           n1487, Q => n1686, QN => n382);
   REGISTERS_reg_12_5_inst : DFFR_X1 port map( D => n3183, CK => CLK, RN => 
                           n1487, Q => n1665, QN => n383);
   REGISTERS_reg_12_4_inst : DFFR_X1 port map( D => n3182, CK => CLK, RN => 
                           n1487, Q => n1644, QN => n384);
   REGISTERS_reg_12_3_inst : DFFR_X1 port map( D => n3181, CK => CLK, RN => 
                           n1487, Q => n1624, QN => n385);
   REGISTERS_reg_12_2_inst : DFFR_X1 port map( D => n3180, CK => CLK, RN => 
                           n1487, Q => n219, QN => n386);
   REGISTERS_reg_12_1_inst : DFFR_X1 port map( D => n3179, CK => CLK, RN => 
                           n1487, Q => n1585, QN => n387);
   REGISTERS_reg_12_0_inst : DFFR_X1 port map( D => n3178, CK => CLK, RN => 
                           n1487, Q => n1562, QN => n388);
   REGISTERS_reg_13_23_inst : DFFR_X1 port map( D => n3169, CK => CLK, RN => 
                           n1488, Q => n2034, QN => n397);
   REGISTERS_reg_13_22_inst : DFFR_X1 port map( D => n3168, CK => CLK, RN => 
                           n1488, Q => n2013, QN => n398);
   REGISTERS_reg_13_21_inst : DFFR_X1 port map( D => n3167, CK => CLK, RN => 
                           n1488, Q => n1993, QN => n399);
   REGISTERS_reg_13_20_inst : DFFR_X1 port map( D => n3166, CK => CLK, RN => 
                           n1488, Q => n1972, QN => n400);
   REGISTERS_reg_13_19_inst : DFFR_X1 port map( D => n3165, CK => CLK, RN => 
                           n1489, Q => n1952, QN => n401);
   REGISTERS_reg_13_18_inst : DFFR_X1 port map( D => n3164, CK => CLK, RN => 
                           n1489, Q => n1932, QN => n402);
   REGISTERS_reg_13_17_inst : DFFR_X1 port map( D => n3163, CK => CLK, RN => 
                           n1489, Q => n1912, QN => n403);
   REGISTERS_reg_13_16_inst : DFFR_X1 port map( D => n3162, CK => CLK, RN => 
                           n1489, Q => n1891, QN => n404);
   REGISTERS_reg_13_15_inst : DFFR_X1 port map( D => n3161, CK => CLK, RN => 
                           n1489, Q => n220, QN => n405);
   REGISTERS_reg_13_14_inst : DFFR_X1 port map( D => n3160, CK => CLK, RN => 
                           n1489, Q => n1851, QN => n406);
   REGISTERS_reg_13_13_inst : DFFR_X1 port map( D => n3159, CK => CLK, RN => 
                           n1489, Q => n1830, QN => n407);
   REGISTERS_reg_13_12_inst : DFFR_X1 port map( D => n3158, CK => CLK, RN => 
                           n1489, Q => n1810, QN => n408);
   REGISTERS_reg_13_11_inst : DFFR_X1 port map( D => n3157, CK => CLK, RN => 
                           n1489, Q => n1789, QN => n409);
   REGISTERS_reg_13_10_inst : DFFR_X1 port map( D => n3156, CK => CLK, RN => 
                           n1489, Q => n1768, QN => n410);
   REGISTERS_reg_13_9_inst : DFFR_X1 port map( D => n3155, CK => CLK, RN => 
                           n1489, Q => n1747, QN => n411);
   REGISTERS_reg_13_8_inst : DFFR_X1 port map( D => n3154, CK => CLK, RN => 
                           n1489, Q => n1726, QN => n412);
   REGISTERS_reg_13_7_inst : DFFR_X1 port map( D => n3153, CK => CLK, RN => 
                           n1490, Q => n1705, QN => n413);
   REGISTERS_reg_13_6_inst : DFFR_X1 port map( D => n3152, CK => CLK, RN => 
                           n1490, Q => n1684, QN => n414);
   REGISTERS_reg_13_5_inst : DFFR_X1 port map( D => n3151, CK => CLK, RN => 
                           n1490, Q => n1663, QN => n415);
   REGISTERS_reg_13_4_inst : DFFR_X1 port map( D => n3150, CK => CLK, RN => 
                           n1490, Q => n1642, QN => n416);
   REGISTERS_reg_13_3_inst : DFFR_X1 port map( D => n3149, CK => CLK, RN => 
                           n1490, Q => n1622, QN => n417);
   REGISTERS_reg_13_2_inst : DFFR_X1 port map( D => n3148, CK => CLK, RN => 
                           n1490, Q => n218, QN => n418);
   REGISTERS_reg_13_1_inst : DFFR_X1 port map( D => n3147, CK => CLK, RN => 
                           n1490, Q => n1583, QN => n419);
   REGISTERS_reg_13_0_inst : DFFR_X1 port map( D => n3146, CK => CLK, RN => 
                           n1490, Q => n1558, QN => n420);
   REGISTERS_reg_14_31_inst : DFFR_X1 port map( D => n3145, CK => CLK, RN => 
                           n1490, Q => n5043, QN => n4095);
   REGISTERS_reg_14_30_inst : DFFR_X1 port map( D => n3144, CK => CLK, RN => 
                           n1490, Q => n5042, QN => n4064);
   REGISTERS_reg_14_29_inst : DFFR_X1 port map( D => n3143, CK => CLK, RN => 
                           n1490, Q => n5041, QN => n4038);
   REGISTERS_reg_14_28_inst : DFFR_X1 port map( D => n3142, CK => CLK, RN => 
                           n1490, Q => n5040, QN => n4012);
   REGISTERS_reg_14_27_inst : DFFR_X1 port map( D => n3141, CK => CLK, RN => 
                           n1491, Q => n5039, QN => n3986);
   REGISTERS_reg_14_26_inst : DFFR_X1 port map( D => n3140, CK => CLK, RN => 
                           n1491, Q => n5038, QN => n3960);
   REGISTERS_reg_14_25_inst : DFFR_X1 port map( D => n3139, CK => CLK, RN => 
                           n1491, Q => n5037, QN => n3934);
   REGISTERS_reg_14_24_inst : DFFR_X1 port map( D => n3138, CK => CLK, RN => 
                           n1491, Q => n5036, QN => n3908);
   REGISTERS_reg_14_23_inst : DFFR_X1 port map( D => n3137, CK => CLK, RN => 
                           n1491, Q => n5035, QN => n3882);
   REGISTERS_reg_14_22_inst : DFFR_X1 port map( D => n3136, CK => CLK, RN => 
                           n1491, Q => n5034, QN => n3857);
   REGISTERS_reg_14_21_inst : DFFR_X1 port map( D => n3135, CK => CLK, RN => 
                           n1491, Q => n5033, QN => n3832);
   REGISTERS_reg_14_20_inst : DFFR_X1 port map( D => n3134, CK => CLK, RN => 
                           n1491, Q => n5032, QN => n3807);
   REGISTERS_reg_14_19_inst : DFFR_X1 port map( D => n3133, CK => CLK, RN => 
                           n1491, Q => n5031, QN => n3782);
   REGISTERS_reg_14_18_inst : DFFR_X1 port map( D => n3132, CK => CLK, RN => 
                           n1491, Q => n5030, QN => n3757);
   REGISTERS_reg_14_17_inst : DFFR_X1 port map( D => n3131, CK => CLK, RN => 
                           n1491, Q => n5029, QN => n3732);
   REGISTERS_reg_14_16_inst : DFFR_X1 port map( D => n3130, CK => CLK, RN => 
                           n1491, Q => n5028, QN => n3707);
   REGISTERS_reg_14_15_inst : DFFR_X1 port map( D => n3129, CK => CLK, RN => 
                           n1492, Q => n5027, QN => n3682);
   REGISTERS_reg_14_14_inst : DFFR_X1 port map( D => n3128, CK => CLK, RN => 
                           n1492, Q => n5026, QN => n3657);
   REGISTERS_reg_14_13_inst : DFFR_X1 port map( D => n3127, CK => CLK, RN => 
                           n1492, Q => n5025, QN => n3632);
   REGISTERS_reg_14_12_inst : DFFR_X1 port map( D => n3126, CK => CLK, RN => 
                           n1492, Q => n5024, QN => n3607);
   REGISTERS_reg_14_11_inst : DFFR_X1 port map( D => n3125, CK => CLK, RN => 
                           n1492, Q => n5023, QN => n3582);
   REGISTERS_reg_14_10_inst : DFFR_X1 port map( D => n3124, CK => CLK, RN => 
                           n1492, Q => n5022, QN => n2501);
   REGISTERS_reg_14_9_inst : DFFR_X1 port map( D => n3123, CK => CLK, RN => 
                           n1492, Q => n5021, QN => n2476);
   REGISTERS_reg_14_8_inst : DFFR_X1 port map( D => n3122, CK => CLK, RN => 
                           n1492, Q => n5020, QN => n2451);
   REGISTERS_reg_14_7_inst : DFFR_X1 port map( D => n3121, CK => CLK, RN => 
                           n1492, Q => n5019, QN => n2426);
   REGISTERS_reg_14_6_inst : DFFR_X1 port map( D => n3120, CK => CLK, RN => 
                           n1492, Q => n5018, QN => n2401);
   REGISTERS_reg_14_5_inst : DFFR_X1 port map( D => n3119, CK => CLK, RN => 
                           n1492, Q => n5017, QN => n2376);
   REGISTERS_reg_14_4_inst : DFFR_X1 port map( D => n3118, CK => CLK, RN => 
                           n1492, Q => n5016, QN => n2351);
   REGISTERS_reg_14_3_inst : DFFR_X1 port map( D => n3117, CK => CLK, RN => 
                           n1493, Q => n5015, QN => n2326);
   REGISTERS_reg_14_2_inst : DFFR_X1 port map( D => n3116, CK => CLK, RN => 
                           n1493, Q => n5014, QN => n2301);
   REGISTERS_reg_14_1_inst : DFFR_X1 port map( D => n3115, CK => CLK, RN => 
                           n1493, Q => n5013, QN => n2276);
   REGISTERS_reg_14_0_inst : DFFR_X1 port map( D => n3114, CK => CLK, RN => 
                           n1493, Q => n5012, QN => n2247);
   REGISTERS_reg_15_31_inst : DFFR_X1 port map( D => n3113, CK => CLK, RN => 
                           n1493, Q => n5011, QN => n4093);
   REGISTERS_reg_15_30_inst : DFFR_X1 port map( D => n3112, CK => CLK, RN => 
                           n1493, Q => n5010, QN => n4063);
   REGISTERS_reg_15_29_inst : DFFR_X1 port map( D => n3111, CK => CLK, RN => 
                           n1493, Q => n5009, QN => n4037);
   REGISTERS_reg_15_28_inst : DFFR_X1 port map( D => n3110, CK => CLK, RN => 
                           n1493, Q => n5008, QN => n4011);
   REGISTERS_reg_15_27_inst : DFFR_X1 port map( D => n3109, CK => CLK, RN => 
                           n1493, Q => n5007, QN => n3985);
   REGISTERS_reg_15_26_inst : DFFR_X1 port map( D => n3108, CK => CLK, RN => 
                           n1493, Q => n5006, QN => n3959);
   REGISTERS_reg_15_25_inst : DFFR_X1 port map( D => n3107, CK => CLK, RN => 
                           n1493, Q => n5005, QN => n3933);
   REGISTERS_reg_15_24_inst : DFFR_X1 port map( D => n3106, CK => CLK, RN => 
                           n1493, Q => n5004, QN => n3907);
   REGISTERS_reg_15_23_inst : DFFR_X1 port map( D => n3105, CK => CLK, RN => 
                           n1494, Q => n5003, QN => n3881);
   REGISTERS_reg_15_22_inst : DFFR_X1 port map( D => n3104, CK => CLK, RN => 
                           n1494, Q => n5002, QN => n3856);
   REGISTERS_reg_15_21_inst : DFFR_X1 port map( D => n3103, CK => CLK, RN => 
                           n1494, Q => n5001, QN => n3831);
   REGISTERS_reg_15_20_inst : DFFR_X1 port map( D => n3102, CK => CLK, RN => 
                           n1494, Q => n5000, QN => n3806);
   REGISTERS_reg_15_19_inst : DFFR_X1 port map( D => n3101, CK => CLK, RN => 
                           n1494, Q => n4999, QN => n3781);
   REGISTERS_reg_15_18_inst : DFFR_X1 port map( D => n3100, CK => CLK, RN => 
                           n1494, Q => n4998, QN => n3756);
   REGISTERS_reg_15_17_inst : DFFR_X1 port map( D => n3099, CK => CLK, RN => 
                           n1494, Q => n4997, QN => n3731);
   REGISTERS_reg_15_16_inst : DFFR_X1 port map( D => n3098, CK => CLK, RN => 
                           n1494, Q => n4996, QN => n3706);
   REGISTERS_reg_15_15_inst : DFFR_X1 port map( D => n3097, CK => CLK, RN => 
                           n1494, Q => n4995, QN => n3681);
   REGISTERS_reg_15_14_inst : DFFR_X1 port map( D => n3096, CK => CLK, RN => 
                           n1494, Q => n4994, QN => n3656);
   REGISTERS_reg_15_13_inst : DFFR_X1 port map( D => n3095, CK => CLK, RN => 
                           n1494, Q => n4993, QN => n3631);
   REGISTERS_reg_15_12_inst : DFFR_X1 port map( D => n3094, CK => CLK, RN => 
                           n1494, Q => n4992, QN => n3606);
   REGISTERS_reg_15_11_inst : DFFR_X1 port map( D => n3093, CK => CLK, RN => 
                           n1495, Q => n4991, QN => n3581);
   REGISTERS_reg_15_10_inst : DFFR_X1 port map( D => n3092, CK => CLK, RN => 
                           n1495, Q => n4990, QN => n2500);
   REGISTERS_reg_15_9_inst : DFFR_X1 port map( D => n3091, CK => CLK, RN => 
                           n1495, Q => n4989, QN => n2475);
   REGISTERS_reg_15_8_inst : DFFR_X1 port map( D => n3090, CK => CLK, RN => 
                           n1495, Q => n4988, QN => n2450);
   REGISTERS_reg_15_7_inst : DFFR_X1 port map( D => n3089, CK => CLK, RN => 
                           n1495, Q => n4987, QN => n2425);
   REGISTERS_reg_15_6_inst : DFFR_X1 port map( D => n3088, CK => CLK, RN => 
                           n1495, Q => n4986, QN => n2400);
   REGISTERS_reg_15_5_inst : DFFR_X1 port map( D => n3087, CK => CLK, RN => 
                           n1495, Q => n4985, QN => n2375);
   REGISTERS_reg_15_4_inst : DFFR_X1 port map( D => n3086, CK => CLK, RN => 
                           n1495, Q => n4984, QN => n2350);
   REGISTERS_reg_15_3_inst : DFFR_X1 port map( D => n3085, CK => CLK, RN => 
                           n1495, Q => n4983, QN => n2325);
   REGISTERS_reg_15_2_inst : DFFR_X1 port map( D => n3084, CK => CLK, RN => 
                           n1495, Q => n4982, QN => n2300);
   REGISTERS_reg_15_1_inst : DFFR_X1 port map( D => n3083, CK => CLK, RN => 
                           n1495, Q => n4981, QN => n2275);
   REGISTERS_reg_15_0_inst : DFFR_X1 port map( D => n3082, CK => CLK, RN => 
                           n1495, Q => n4980, QN => n2246);
   REGISTERS_reg_16_23_inst : DFFR_X1 port map( D => n3073, CK => CLK, RN => 
                           n1496, Q => n4232, QN => n_1283);
   REGISTERS_reg_16_22_inst : DFFR_X1 port map( D => n3072, CK => CLK, RN => 
                           n1496, Q => n4233, QN => n_1284);
   REGISTERS_reg_16_21_inst : DFFR_X1 port map( D => n3071, CK => CLK, RN => 
                           n1496, Q => n4234, QN => n_1285);
   REGISTERS_reg_16_20_inst : DFFR_X1 port map( D => n3070, CK => CLK, RN => 
                           n1496, Q => n4235, QN => n_1286);
   REGISTERS_reg_16_19_inst : DFFR_X1 port map( D => n3069, CK => CLK, RN => 
                           n1497, Q => n4236, QN => n_1287);
   REGISTERS_reg_16_18_inst : DFFR_X1 port map( D => n3068, CK => CLK, RN => 
                           n1497, Q => n4237, QN => n_1288);
   REGISTERS_reg_16_17_inst : DFFR_X1 port map( D => n3067, CK => CLK, RN => 
                           n1497, Q => n4238, QN => n_1289);
   REGISTERS_reg_16_16_inst : DFFR_X1 port map( D => n3066, CK => CLK, RN => 
                           n1497, Q => n4239, QN => n_1290);
   REGISTERS_reg_16_15_inst : DFFR_X1 port map( D => n3065, CK => CLK, RN => 
                           n1497, Q => n4240, QN => n_1291);
   REGISTERS_reg_16_14_inst : DFFR_X1 port map( D => n3064, CK => CLK, RN => 
                           n1497, Q => n4241, QN => n_1292);
   REGISTERS_reg_16_13_inst : DFFR_X1 port map( D => n3063, CK => CLK, RN => 
                           n1497, Q => n4242, QN => n_1293);
   REGISTERS_reg_16_12_inst : DFFR_X1 port map( D => n3062, CK => CLK, RN => 
                           n1497, Q => n4243, QN => n_1294);
   REGISTERS_reg_16_11_inst : DFFR_X1 port map( D => n3061, CK => CLK, RN => 
                           n1497, Q => n4244, QN => n_1295);
   REGISTERS_reg_16_10_inst : DFFR_X1 port map( D => n3060, CK => CLK, RN => 
                           n1497, Q => n4245, QN => n_1296);
   REGISTERS_reg_16_9_inst : DFFR_X1 port map( D => n3059, CK => CLK, RN => 
                           n1497, Q => n4246, QN => n_1297);
   REGISTERS_reg_16_8_inst : DFFR_X1 port map( D => n3058, CK => CLK, RN => 
                           n1497, Q => n4247, QN => n_1298);
   REGISTERS_reg_16_7_inst : DFFR_X1 port map( D => n3057, CK => CLK, RN => 
                           n1498, Q => n4248, QN => n_1299);
   REGISTERS_reg_16_6_inst : DFFR_X1 port map( D => n3056, CK => CLK, RN => 
                           n1498, Q => n4249, QN => n_1300);
   REGISTERS_reg_16_5_inst : DFFR_X1 port map( D => n3055, CK => CLK, RN => 
                           n1498, Q => n4250, QN => n_1301);
   REGISTERS_reg_16_4_inst : DFFR_X1 port map( D => n3054, CK => CLK, RN => 
                           n1498, Q => n4251, QN => n_1302);
   REGISTERS_reg_16_3_inst : DFFR_X1 port map( D => n3053, CK => CLK, RN => 
                           n1498, Q => n4252, QN => n_1303);
   REGISTERS_reg_16_2_inst : DFFR_X1 port map( D => n3052, CK => CLK, RN => 
                           n1498, Q => n4253, QN => n_1304);
   REGISTERS_reg_16_1_inst : DFFR_X1 port map( D => n3051, CK => CLK, RN => 
                           n1498, Q => n4254, QN => n_1305);
   REGISTERS_reg_16_0_inst : DFFR_X1 port map( D => n3050, CK => CLK, RN => 
                           n1498, Q => n4255, QN => n_1306);
   REGISTERS_reg_17_23_inst : DFFR_X1 port map( D => n3041, CK => CLK, RN => 
                           n1499, Q => n3898, QN => n525);
   REGISTERS_reg_17_22_inst : DFFR_X1 port map( D => n3040, CK => CLK, RN => 
                           n1499, Q => n3873, QN => n526);
   REGISTERS_reg_17_21_inst : DFFR_X1 port map( D => n3039, CK => CLK, RN => 
                           n1499, Q => n3848, QN => n527);
   REGISTERS_reg_17_20_inst : DFFR_X1 port map( D => n3038, CK => CLK, RN => 
                           n1499, Q => n3823, QN => n528);
   REGISTERS_reg_17_19_inst : DFFR_X1 port map( D => n3037, CK => CLK, RN => 
                           n1499, Q => n3798, QN => n529);
   REGISTERS_reg_17_18_inst : DFFR_X1 port map( D => n3036, CK => CLK, RN => 
                           n1499, Q => n3773, QN => n530);
   REGISTERS_reg_17_17_inst : DFFR_X1 port map( D => n3035, CK => CLK, RN => 
                           n1499, Q => n3748, QN => n531);
   REGISTERS_reg_17_16_inst : DFFR_X1 port map( D => n3034, CK => CLK, RN => 
                           n1499, Q => n3723, QN => n532);
   REGISTERS_reg_17_15_inst : DFFR_X1 port map( D => n3033, CK => CLK, RN => 
                           n1500, Q => n3698, QN => n533);
   REGISTERS_reg_17_14_inst : DFFR_X1 port map( D => n3032, CK => CLK, RN => 
                           n1500, Q => n3673, QN => n534);
   REGISTERS_reg_17_13_inst : DFFR_X1 port map( D => n3031, CK => CLK, RN => 
                           n1500, Q => n3648, QN => n535);
   REGISTERS_reg_17_12_inst : DFFR_X1 port map( D => n3030, CK => CLK, RN => 
                           n1500, Q => n3623, QN => n536);
   REGISTERS_reg_17_11_inst : DFFR_X1 port map( D => n3029, CK => CLK, RN => 
                           n1500, Q => n3598, QN => n537);
   REGISTERS_reg_17_10_inst : DFFR_X1 port map( D => n3028, CK => CLK, RN => 
                           n1500, Q => n3573, QN => n538);
   REGISTERS_reg_17_9_inst : DFFR_X1 port map( D => n3027, CK => CLK, RN => 
                           n1500, Q => n2492, QN => n539);
   REGISTERS_reg_17_8_inst : DFFR_X1 port map( D => n3026, CK => CLK, RN => 
                           n1500, Q => n2467, QN => n540);
   REGISTERS_reg_17_7_inst : DFFR_X1 port map( D => n3025, CK => CLK, RN => 
                           n1500, Q => n2442, QN => n541);
   REGISTERS_reg_17_6_inst : DFFR_X1 port map( D => n3024, CK => CLK, RN => 
                           n1500, Q => n2417, QN => n542);
   REGISTERS_reg_17_5_inst : DFFR_X1 port map( D => n3023, CK => CLK, RN => 
                           n1500, Q => n2392, QN => n543);
   REGISTERS_reg_17_4_inst : DFFR_X1 port map( D => n3022, CK => CLK, RN => 
                           n1500, Q => n2367, QN => n544);
   REGISTERS_reg_17_3_inst : DFFR_X1 port map( D => n3021, CK => CLK, RN => 
                           n1501, Q => n2342, QN => n545);
   REGISTERS_reg_17_2_inst : DFFR_X1 port map( D => n3020, CK => CLK, RN => 
                           n1501, Q => n2317, QN => n546);
   REGISTERS_reg_17_1_inst : DFFR_X1 port map( D => n3019, CK => CLK, RN => 
                           n1501, Q => n2292, QN => n547);
   REGISTERS_reg_17_0_inst : DFFR_X1 port map( D => n3018, CK => CLK, RN => 
                           n1501, Q => n2267, QN => n548);
   REGISTERS_reg_18_31_inst : DFFR_X1 port map( D => n3017, CK => CLK, RN => 
                           n1501, Q => n4979, QN => n_1307);
   REGISTERS_reg_18_30_inst : DFFR_X1 port map( D => n3016, CK => CLK, RN => 
                           n1501, Q => n4978, QN => n_1308);
   REGISTERS_reg_18_29_inst : DFFR_X1 port map( D => n3015, CK => CLK, RN => 
                           n1501, Q => n4977, QN => n_1309);
   REGISTERS_reg_18_28_inst : DFFR_X1 port map( D => n3014, CK => CLK, RN => 
                           n1501, Q => n4976, QN => n_1310);
   REGISTERS_reg_18_27_inst : DFFR_X1 port map( D => n3013, CK => CLK, RN => 
                           n1501, Q => n4975, QN => n_1311);
   REGISTERS_reg_18_26_inst : DFFR_X1 port map( D => n3012, CK => CLK, RN => 
                           n1501, Q => n4974, QN => n_1312);
   REGISTERS_reg_18_25_inst : DFFR_X1 port map( D => n3011, CK => CLK, RN => 
                           n1501, Q => n4973, QN => n_1313);
   REGISTERS_reg_18_24_inst : DFFR_X1 port map( D => n3010, CK => CLK, RN => 
                           n1501, Q => n4972, QN => n_1314);
   REGISTERS_reg_18_23_inst : DFFR_X1 port map( D => n3009, CK => CLK, RN => 
                           n1502, Q => n4971, QN => n_1315);
   REGISTERS_reg_18_22_inst : DFFR_X1 port map( D => n3008, CK => CLK, RN => 
                           n1502, Q => n4970, QN => n_1316);
   REGISTERS_reg_18_21_inst : DFFR_X1 port map( D => n3007, CK => CLK, RN => 
                           n1502, Q => n4969, QN => n_1317);
   REGISTERS_reg_18_20_inst : DFFR_X1 port map( D => n3006, CK => CLK, RN => 
                           n1502, Q => n4968, QN => n_1318);
   REGISTERS_reg_18_19_inst : DFFR_X1 port map( D => n3005, CK => CLK, RN => 
                           n1502, Q => n4967, QN => n_1319);
   REGISTERS_reg_18_18_inst : DFFR_X1 port map( D => n3004, CK => CLK, RN => 
                           n1502, Q => n4966, QN => n_1320);
   REGISTERS_reg_18_17_inst : DFFR_X1 port map( D => n3003, CK => CLK, RN => 
                           n1502, Q => n4965, QN => n_1321);
   REGISTERS_reg_18_16_inst : DFFR_X1 port map( D => n3002, CK => CLK, RN => 
                           n1502, Q => n4964, QN => n_1322);
   REGISTERS_reg_18_15_inst : DFFR_X1 port map( D => n3001, CK => CLK, RN => 
                           n1502, Q => n4963, QN => n_1323);
   REGISTERS_reg_18_14_inst : DFFR_X1 port map( D => n3000, CK => CLK, RN => 
                           n1502, Q => n4962, QN => n_1324);
   REGISTERS_reg_18_13_inst : DFFR_X1 port map( D => n2999, CK => CLK, RN => 
                           n1502, Q => n4961, QN => n_1325);
   REGISTERS_reg_18_12_inst : DFFR_X1 port map( D => n2998, CK => CLK, RN => 
                           n1502, Q => n4960, QN => n_1326);
   REGISTERS_reg_18_11_inst : DFFR_X1 port map( D => n2997, CK => CLK, RN => 
                           n1503, Q => n4959, QN => n_1327);
   REGISTERS_reg_18_10_inst : DFFR_X1 port map( D => n2996, CK => CLK, RN => 
                           n1503, Q => n4958, QN => n_1328);
   REGISTERS_reg_18_9_inst : DFFR_X1 port map( D => n2995, CK => CLK, RN => 
                           n1503, Q => n4957, QN => n_1329);
   REGISTERS_reg_18_8_inst : DFFR_X1 port map( D => n2994, CK => CLK, RN => 
                           n1503, Q => n4956, QN => n_1330);
   REGISTERS_reg_18_7_inst : DFFR_X1 port map( D => n2993, CK => CLK, RN => 
                           n1503, Q => n4955, QN => n_1331);
   REGISTERS_reg_18_6_inst : DFFR_X1 port map( D => n2992, CK => CLK, RN => 
                           n1503, Q => n4954, QN => n_1332);
   REGISTERS_reg_18_5_inst : DFFR_X1 port map( D => n2991, CK => CLK, RN => 
                           n1503, Q => n4953, QN => n_1333);
   REGISTERS_reg_18_4_inst : DFFR_X1 port map( D => n2990, CK => CLK, RN => 
                           n1503, Q => n4952, QN => n_1334);
   REGISTERS_reg_18_3_inst : DFFR_X1 port map( D => n2989, CK => CLK, RN => 
                           n1503, Q => n4951, QN => n_1335);
   REGISTERS_reg_18_2_inst : DFFR_X1 port map( D => n2988, CK => CLK, RN => 
                           n1503, Q => n4950, QN => n_1336);
   REGISTERS_reg_18_1_inst : DFFR_X1 port map( D => n2987, CK => CLK, RN => 
                           n1503, Q => n4949, QN => n_1337);
   REGISTERS_reg_18_0_inst : DFFR_X1 port map( D => n2986, CK => CLK, RN => 
                           n1503, Q => n4948, QN => n_1338);
   REGISTERS_reg_19_31_inst : DFFR_X1 port map( D => n2985, CK => CLK, RN => 
                           n1504, Q => n4947, QN => n4115);
   REGISTERS_reg_19_30_inst : DFFR_X1 port map( D => n2984, CK => CLK, RN => 
                           n1504, Q => n4946, QN => n4076);
   REGISTERS_reg_19_29_inst : DFFR_X1 port map( D => n2983, CK => CLK, RN => 
                           n1504, Q => n4945, QN => n4050);
   REGISTERS_reg_19_28_inst : DFFR_X1 port map( D => n2982, CK => CLK, RN => 
                           n1504, Q => n4944, QN => n4024);
   REGISTERS_reg_19_27_inst : DFFR_X1 port map( D => n2981, CK => CLK, RN => 
                           n1504, Q => n4943, QN => n3998);
   REGISTERS_reg_19_26_inst : DFFR_X1 port map( D => n2980, CK => CLK, RN => 
                           n1504, Q => n4942, QN => n3972);
   REGISTERS_reg_19_25_inst : DFFR_X1 port map( D => n2979, CK => CLK, RN => 
                           n1504, Q => n4941, QN => n3946);
   REGISTERS_reg_19_24_inst : DFFR_X1 port map( D => n2978, CK => CLK, RN => 
                           n1504, Q => n4940, QN => n3920);
   REGISTERS_reg_19_23_inst : DFFR_X1 port map( D => n2977, CK => CLK, RN => 
                           n1504, Q => n4939, QN => n3894);
   REGISTERS_reg_19_22_inst : DFFR_X1 port map( D => n2976, CK => CLK, RN => 
                           n1504, Q => n4938, QN => n3869);
   REGISTERS_reg_19_21_inst : DFFR_X1 port map( D => n2975, CK => CLK, RN => 
                           n1504, Q => n4937, QN => n3844);
   REGISTERS_reg_19_20_inst : DFFR_X1 port map( D => n2974, CK => CLK, RN => 
                           n1504, Q => n4936, QN => n3819);
   REGISTERS_reg_19_19_inst : DFFR_X1 port map( D => n2973, CK => CLK, RN => 
                           n1505, Q => n4935, QN => n3794);
   REGISTERS_reg_19_18_inst : DFFR_X1 port map( D => n2972, CK => CLK, RN => 
                           n1505, Q => n4934, QN => n3769);
   REGISTERS_reg_19_17_inst : DFFR_X1 port map( D => n2971, CK => CLK, RN => 
                           n1505, Q => n4933, QN => n3744);
   REGISTERS_reg_19_16_inst : DFFR_X1 port map( D => n2970, CK => CLK, RN => 
                           n1505, Q => n4932, QN => n3719);
   REGISTERS_reg_19_15_inst : DFFR_X1 port map( D => n2969, CK => CLK, RN => 
                           n1505, Q => n4931, QN => n3694);
   REGISTERS_reg_19_14_inst : DFFR_X1 port map( D => n2968, CK => CLK, RN => 
                           n1505, Q => n4930, QN => n3669);
   REGISTERS_reg_19_13_inst : DFFR_X1 port map( D => n2967, CK => CLK, RN => 
                           n1505, Q => n4929, QN => n3644);
   REGISTERS_reg_19_12_inst : DFFR_X1 port map( D => n2966, CK => CLK, RN => 
                           n1505, Q => n4928, QN => n3619);
   REGISTERS_reg_19_11_inst : DFFR_X1 port map( D => n2965, CK => CLK, RN => 
                           n1505, Q => n4927, QN => n3594);
   REGISTERS_reg_19_10_inst : DFFR_X1 port map( D => n2964, CK => CLK, RN => 
                           n1505, Q => n4926, QN => n3569);
   REGISTERS_reg_19_9_inst : DFFR_X1 port map( D => n2963, CK => CLK, RN => 
                           n1505, Q => n4925, QN => n2488);
   REGISTERS_reg_19_8_inst : DFFR_X1 port map( D => n2962, CK => CLK, RN => 
                           n1505, Q => n4924, QN => n2463);
   REGISTERS_reg_19_7_inst : DFFR_X1 port map( D => n2961, CK => CLK, RN => 
                           n1506, Q => n4923, QN => n2438);
   REGISTERS_reg_19_6_inst : DFFR_X1 port map( D => n2960, CK => CLK, RN => 
                           n1506, Q => n4922, QN => n2413);
   REGISTERS_reg_19_5_inst : DFFR_X1 port map( D => n2959, CK => CLK, RN => 
                           n1506, Q => n4921, QN => n2388);
   REGISTERS_reg_19_4_inst : DFFR_X1 port map( D => n2958, CK => CLK, RN => 
                           n1506, Q => n4920, QN => n2363);
   REGISTERS_reg_19_3_inst : DFFR_X1 port map( D => n2957, CK => CLK, RN => 
                           n1506, Q => n4919, QN => n2338);
   REGISTERS_reg_19_2_inst : DFFR_X1 port map( D => n2956, CK => CLK, RN => 
                           n1506, Q => n4918, QN => n2313);
   REGISTERS_reg_19_1_inst : DFFR_X1 port map( D => n2955, CK => CLK, RN => 
                           n1506, Q => n4917, QN => n2288);
   REGISTERS_reg_19_0_inst : DFFR_X1 port map( D => n2954, CK => CLK, RN => 
                           n1506, Q => n4916, QN => n2261);
   REGISTERS_reg_20_23_inst : DFFR_X1 port map( D => n2945, CK => CLK, RN => 
                           n1507, Q => n_1339, QN => n621);
   REGISTERS_reg_20_22_inst : DFFR_X1 port map( D => n2944, CK => CLK, RN => 
                           n1507, Q => n_1340, QN => n622);
   REGISTERS_reg_20_21_inst : DFFR_X1 port map( D => n2943, CK => CLK, RN => 
                           n1507, Q => n_1341, QN => n623);
   REGISTERS_reg_20_20_inst : DFFR_X1 port map( D => n2942, CK => CLK, RN => 
                           n1507, Q => n_1342, QN => n624);
   REGISTERS_reg_20_19_inst : DFFR_X1 port map( D => n2941, CK => CLK, RN => 
                           n1507, Q => n_1343, QN => n625);
   REGISTERS_reg_20_18_inst : DFFR_X1 port map( D => n2940, CK => CLK, RN => 
                           n1507, Q => n_1344, QN => n626);
   REGISTERS_reg_20_17_inst : DFFR_X1 port map( D => n2939, CK => CLK, RN => 
                           n1507, Q => n_1345, QN => n627);
   REGISTERS_reg_20_16_inst : DFFR_X1 port map( D => n2938, CK => CLK, RN => 
                           n1507, Q => n_1346, QN => n628);
   REGISTERS_reg_20_15_inst : DFFR_X1 port map( D => n2937, CK => CLK, RN => 
                           n1508, Q => n_1347, QN => n629);
   REGISTERS_reg_20_14_inst : DFFR_X1 port map( D => n2936, CK => CLK, RN => 
                           n1508, Q => n_1348, QN => n630);
   REGISTERS_reg_20_13_inst : DFFR_X1 port map( D => n2935, CK => CLK, RN => 
                           n1508, Q => n_1349, QN => n631);
   REGISTERS_reg_20_12_inst : DFFR_X1 port map( D => n2934, CK => CLK, RN => 
                           n1508, Q => n_1350, QN => n632);
   REGISTERS_reg_20_11_inst : DFFR_X1 port map( D => n2933, CK => CLK, RN => 
                           n1508, Q => n_1351, QN => n633);
   REGISTERS_reg_20_10_inst : DFFR_X1 port map( D => n2932, CK => CLK, RN => 
                           n1508, Q => n_1352, QN => n634);
   REGISTERS_reg_20_9_inst : DFFR_X1 port map( D => n2931, CK => CLK, RN => 
                           n1508, Q => n_1353, QN => n635);
   REGISTERS_reg_20_8_inst : DFFR_X1 port map( D => n2930, CK => CLK, RN => 
                           n1508, Q => n_1354, QN => n636);
   REGISTERS_reg_20_7_inst : DFFR_X1 port map( D => n2929, CK => CLK, RN => 
                           n1508, Q => n_1355, QN => n637);
   REGISTERS_reg_20_6_inst : DFFR_X1 port map( D => n2928, CK => CLK, RN => 
                           n1508, Q => n_1356, QN => n638);
   REGISTERS_reg_20_5_inst : DFFR_X1 port map( D => n2927, CK => CLK, RN => 
                           n1508, Q => n_1357, QN => n639);
   REGISTERS_reg_20_4_inst : DFFR_X1 port map( D => n2926, CK => CLK, RN => 
                           n1508, Q => n_1358, QN => n640);
   REGISTERS_reg_20_3_inst : DFFR_X1 port map( D => n2925, CK => CLK, RN => 
                           n1509, Q => n_1359, QN => n641);
   REGISTERS_reg_20_2_inst : DFFR_X1 port map( D => n2924, CK => CLK, RN => 
                           n1509, Q => n_1360, QN => n642);
   REGISTERS_reg_20_1_inst : DFFR_X1 port map( D => n2923, CK => CLK, RN => 
                           n1509, Q => n_1361, QN => n643);
   REGISTERS_reg_20_0_inst : DFFR_X1 port map( D => n2922, CK => CLK, RN => 
                           n1509, Q => n_1362, QN => n644);
   REGISTERS_reg_21_23_inst : DFFR_X1 port map( D => n2913, CK => CLK, RN => 
                           n1510, Q => n4264, QN => n_1363);
   REGISTERS_reg_21_22_inst : DFFR_X1 port map( D => n2912, CK => CLK, RN => 
                           n1510, Q => n4265, QN => n_1364);
   REGISTERS_reg_21_21_inst : DFFR_X1 port map( D => n2911, CK => CLK, RN => 
                           n1510, Q => n4266, QN => n_1365);
   REGISTERS_reg_21_20_inst : DFFR_X1 port map( D => n2910, CK => CLK, RN => 
                           n1510, Q => n4267, QN => n_1366);
   REGISTERS_reg_21_19_inst : DFFR_X1 port map( D => n2909, CK => CLK, RN => 
                           n1510, Q => n4268, QN => n_1367);
   REGISTERS_reg_21_18_inst : DFFR_X1 port map( D => n2908, CK => CLK, RN => 
                           n1510, Q => n4269, QN => n_1368);
   REGISTERS_reg_21_17_inst : DFFR_X1 port map( D => n2907, CK => CLK, RN => 
                           n1510, Q => n4270, QN => n_1369);
   REGISTERS_reg_21_16_inst : DFFR_X1 port map( D => n2906, CK => CLK, RN => 
                           n1510, Q => n4271, QN => n_1370);
   REGISTERS_reg_21_15_inst : DFFR_X1 port map( D => n2905, CK => CLK, RN => 
                           n1510, Q => n4272, QN => n_1371);
   REGISTERS_reg_21_14_inst : DFFR_X1 port map( D => n2904, CK => CLK, RN => 
                           n1510, Q => n4273, QN => n_1372);
   REGISTERS_reg_21_13_inst : DFFR_X1 port map( D => n2903, CK => CLK, RN => 
                           n1510, Q => n4274, QN => n_1373);
   REGISTERS_reg_21_12_inst : DFFR_X1 port map( D => n2902, CK => CLK, RN => 
                           n1510, Q => n4275, QN => n_1374);
   REGISTERS_reg_21_11_inst : DFFR_X1 port map( D => n2901, CK => CLK, RN => 
                           n1511, Q => n4276, QN => n_1375);
   REGISTERS_reg_21_10_inst : DFFR_X1 port map( D => n2900, CK => CLK, RN => 
                           n1511, Q => n4277, QN => n_1376);
   REGISTERS_reg_21_9_inst : DFFR_X1 port map( D => n2899, CK => CLK, RN => 
                           n1511, Q => n4278, QN => n_1377);
   REGISTERS_reg_21_8_inst : DFFR_X1 port map( D => n2898, CK => CLK, RN => 
                           n1511, Q => n4279, QN => n_1378);
   REGISTERS_reg_21_7_inst : DFFR_X1 port map( D => n2897, CK => CLK, RN => 
                           n1511, Q => n4280, QN => n_1379);
   REGISTERS_reg_21_6_inst : DFFR_X1 port map( D => n2896, CK => CLK, RN => 
                           n1511, Q => n4281, QN => n_1380);
   REGISTERS_reg_21_5_inst : DFFR_X1 port map( D => n2895, CK => CLK, RN => 
                           n1511, Q => n4282, QN => n_1381);
   REGISTERS_reg_21_4_inst : DFFR_X1 port map( D => n2894, CK => CLK, RN => 
                           n1511, Q => n4283, QN => n_1382);
   REGISTERS_reg_21_3_inst : DFFR_X1 port map( D => n2893, CK => CLK, RN => 
                           n1511, Q => n4284, QN => n_1383);
   REGISTERS_reg_21_2_inst : DFFR_X1 port map( D => n2892, CK => CLK, RN => 
                           n1511, Q => n4285, QN => n_1384);
   REGISTERS_reg_21_1_inst : DFFR_X1 port map( D => n2891, CK => CLK, RN => 
                           n1511, Q => n4286, QN => n_1385);
   REGISTERS_reg_21_0_inst : DFFR_X1 port map( D => n2890, CK => CLK, RN => 
                           n1511, Q => n4287, QN => n_1386);
   REGISTERS_reg_22_31_inst : DFFR_X1 port map( D => n2889, CK => CLK, RN => 
                           n1512, Q => n4915, QN => n4117);
   REGISTERS_reg_22_30_inst : DFFR_X1 port map( D => n2888, CK => CLK, RN => 
                           n1512, Q => n4914, QN => n4077);
   REGISTERS_reg_22_29_inst : DFFR_X1 port map( D => n2887, CK => CLK, RN => 
                           n1512, Q => n4913, QN => n4051);
   REGISTERS_reg_22_28_inst : DFFR_X1 port map( D => n2886, CK => CLK, RN => 
                           n1512, Q => n4912, QN => n4025);
   REGISTERS_reg_22_27_inst : DFFR_X1 port map( D => n2885, CK => CLK, RN => 
                           n1512, Q => n4911, QN => n3999);
   REGISTERS_reg_22_26_inst : DFFR_X1 port map( D => n2884, CK => CLK, RN => 
                           n1512, Q => n4910, QN => n3973);
   REGISTERS_reg_22_25_inst : DFFR_X1 port map( D => n2883, CK => CLK, RN => 
                           n1512, Q => n4909, QN => n3947);
   REGISTERS_reg_22_24_inst : DFFR_X1 port map( D => n2882, CK => CLK, RN => 
                           n1512, Q => n4908, QN => n3921);
   REGISTERS_reg_22_23_inst : DFFR_X1 port map( D => n2881, CK => CLK, RN => 
                           n1512, Q => n4907, QN => n3895);
   REGISTERS_reg_22_22_inst : DFFR_X1 port map( D => n2880, CK => CLK, RN => 
                           n1512, Q => n4906, QN => n3870);
   REGISTERS_reg_22_21_inst : DFFR_X1 port map( D => n2879, CK => CLK, RN => 
                           n1512, Q => n4905, QN => n3845);
   REGISTERS_reg_22_20_inst : DFFR_X1 port map( D => n2878, CK => CLK, RN => 
                           n1512, Q => n4904, QN => n3820);
   REGISTERS_reg_22_19_inst : DFFR_X1 port map( D => n2877, CK => CLK, RN => 
                           n1513, Q => n4903, QN => n3795);
   REGISTERS_reg_22_18_inst : DFFR_X1 port map( D => n2876, CK => CLK, RN => 
                           n1513, Q => n4902, QN => n3770);
   REGISTERS_reg_22_17_inst : DFFR_X1 port map( D => n2875, CK => CLK, RN => 
                           n1513, Q => n4901, QN => n3745);
   REGISTERS_reg_22_16_inst : DFFR_X1 port map( D => n2874, CK => CLK, RN => 
                           n1513, Q => n4900, QN => n3720);
   REGISTERS_reg_22_15_inst : DFFR_X1 port map( D => n2873, CK => CLK, RN => 
                           n1513, Q => n4899, QN => n3695);
   REGISTERS_reg_22_14_inst : DFFR_X1 port map( D => n2872, CK => CLK, RN => 
                           n1513, Q => n4898, QN => n3670);
   REGISTERS_reg_22_13_inst : DFFR_X1 port map( D => n2871, CK => CLK, RN => 
                           n1513, Q => n4897, QN => n3645);
   REGISTERS_reg_22_12_inst : DFFR_X1 port map( D => n2870, CK => CLK, RN => 
                           n1513, Q => n4896, QN => n3620);
   REGISTERS_reg_22_11_inst : DFFR_X1 port map( D => n2869, CK => CLK, RN => 
                           n1513, Q => n4895, QN => n3595);
   REGISTERS_reg_22_10_inst : DFFR_X1 port map( D => n2868, CK => CLK, RN => 
                           n1513, Q => n4894, QN => n3570);
   REGISTERS_reg_22_9_inst : DFFR_X1 port map( D => n2867, CK => CLK, RN => 
                           n1513, Q => n4893, QN => n2489);
   REGISTERS_reg_22_8_inst : DFFR_X1 port map( D => n2866, CK => CLK, RN => 
                           n1513, Q => n4892, QN => n2464);
   REGISTERS_reg_22_7_inst : DFFR_X1 port map( D => n2865, CK => CLK, RN => 
                           n1514, Q => n4891, QN => n2439);
   REGISTERS_reg_22_6_inst : DFFR_X1 port map( D => n2864, CK => CLK, RN => 
                           n1514, Q => n4890, QN => n2414);
   REGISTERS_reg_22_5_inst : DFFR_X1 port map( D => n2863, CK => CLK, RN => 
                           n1514, Q => n4889, QN => n2389);
   REGISTERS_reg_22_4_inst : DFFR_X1 port map( D => n2862, CK => CLK, RN => 
                           n1514, Q => n4888, QN => n2364);
   REGISTERS_reg_22_3_inst : DFFR_X1 port map( D => n2861, CK => CLK, RN => 
                           n1514, Q => n4887, QN => n2339);
   REGISTERS_reg_22_2_inst : DFFR_X1 port map( D => n2860, CK => CLK, RN => 
                           n1514, Q => n4886, QN => n2314);
   REGISTERS_reg_22_1_inst : DFFR_X1 port map( D => n2859, CK => CLK, RN => 
                           n1514, Q => n4885, QN => n2289);
   REGISTERS_reg_22_0_inst : DFFR_X1 port map( D => n2858, CK => CLK, RN => 
                           n1514, Q => n4884, QN => n2262);
   REGISTERS_reg_23_31_inst : DFFR_X1 port map( D => n2857, CK => CLK, RN => 
                           n1514, Q => n4883, QN => n_1387);
   REGISTERS_reg_23_30_inst : DFFR_X1 port map( D => n2856, CK => CLK, RN => 
                           n1514, Q => n4882, QN => n_1388);
   REGISTERS_reg_23_29_inst : DFFR_X1 port map( D => n2855, CK => CLK, RN => 
                           n1514, Q => n4881, QN => n_1389);
   REGISTERS_reg_23_28_inst : DFFR_X1 port map( D => n2854, CK => CLK, RN => 
                           n1514, Q => n4880, QN => n_1390);
   REGISTERS_reg_23_27_inst : DFFR_X1 port map( D => n2853, CK => CLK, RN => 
                           n1515, Q => n4879, QN => n_1391);
   REGISTERS_reg_23_26_inst : DFFR_X1 port map( D => n2852, CK => CLK, RN => 
                           n1515, Q => n4878, QN => n_1392);
   REGISTERS_reg_23_25_inst : DFFR_X1 port map( D => n2851, CK => CLK, RN => 
                           n1515, Q => n4877, QN => n_1393);
   REGISTERS_reg_23_24_inst : DFFR_X1 port map( D => n2850, CK => CLK, RN => 
                           n1515, Q => n4876, QN => n_1394);
   REGISTERS_reg_23_23_inst : DFFR_X1 port map( D => n2849, CK => CLK, RN => 
                           n1515, Q => n4875, QN => n_1395);
   REGISTERS_reg_23_22_inst : DFFR_X1 port map( D => n2848, CK => CLK, RN => 
                           n1515, Q => n4874, QN => n_1396);
   REGISTERS_reg_23_21_inst : DFFR_X1 port map( D => n2847, CK => CLK, RN => 
                           n1515, Q => n4873, QN => n_1397);
   REGISTERS_reg_23_20_inst : DFFR_X1 port map( D => n2846, CK => CLK, RN => 
                           n1515, Q => n4872, QN => n_1398);
   REGISTERS_reg_23_19_inst : DFFR_X1 port map( D => n2845, CK => CLK, RN => 
                           n1515, Q => n4871, QN => n_1399);
   REGISTERS_reg_23_18_inst : DFFR_X1 port map( D => n2844, CK => CLK, RN => 
                           n1515, Q => n4870, QN => n_1400);
   REGISTERS_reg_23_17_inst : DFFR_X1 port map( D => n2843, CK => CLK, RN => 
                           n1515, Q => n4869, QN => n_1401);
   REGISTERS_reg_23_16_inst : DFFR_X1 port map( D => n2842, CK => CLK, RN => 
                           n1515, Q => n4868, QN => n_1402);
   REGISTERS_reg_23_15_inst : DFFR_X1 port map( D => n2841, CK => CLK, RN => 
                           n1516, Q => n4867, QN => n_1403);
   REGISTERS_reg_23_14_inst : DFFR_X1 port map( D => n2840, CK => CLK, RN => 
                           n1516, Q => n4866, QN => n_1404);
   REGISTERS_reg_23_13_inst : DFFR_X1 port map( D => n2839, CK => CLK, RN => 
                           n1516, Q => n4865, QN => n_1405);
   REGISTERS_reg_23_12_inst : DFFR_X1 port map( D => n2838, CK => CLK, RN => 
                           n1516, Q => n4864, QN => n_1406);
   REGISTERS_reg_23_11_inst : DFFR_X1 port map( D => n2837, CK => CLK, RN => 
                           n1516, Q => n4863, QN => n_1407);
   REGISTERS_reg_23_10_inst : DFFR_X1 port map( D => n2836, CK => CLK, RN => 
                           n1516, Q => n4862, QN => n_1408);
   REGISTERS_reg_23_9_inst : DFFR_X1 port map( D => n2835, CK => CLK, RN => 
                           n1516, Q => n4861, QN => n_1409);
   REGISTERS_reg_23_8_inst : DFFR_X1 port map( D => n2834, CK => CLK, RN => 
                           n1516, Q => n4860, QN => n_1410);
   REGISTERS_reg_23_7_inst : DFFR_X1 port map( D => n2833, CK => CLK, RN => 
                           n1516, Q => n4859, QN => n_1411);
   REGISTERS_reg_23_6_inst : DFFR_X1 port map( D => n2832, CK => CLK, RN => 
                           n1516, Q => n4858, QN => n_1412);
   REGISTERS_reg_23_5_inst : DFFR_X1 port map( D => n2831, CK => CLK, RN => 
                           n1516, Q => n4857, QN => n_1413);
   REGISTERS_reg_23_4_inst : DFFR_X1 port map( D => n2830, CK => CLK, RN => 
                           n1516, Q => n4856, QN => n_1414);
   REGISTERS_reg_23_3_inst : DFFR_X1 port map( D => n2829, CK => CLK, RN => 
                           n1517, Q => n4855, QN => n_1415);
   REGISTERS_reg_23_2_inst : DFFR_X1 port map( D => n2828, CK => CLK, RN => 
                           n1517, Q => n4854, QN => n_1416);
   REGISTERS_reg_23_1_inst : DFFR_X1 port map( D => n2827, CK => CLK, RN => 
                           n1517, Q => n4853, QN => n_1417);
   REGISTERS_reg_23_0_inst : DFFR_X1 port map( D => n2826, CK => CLK, RN => 
                           n1517, Q => n4852, QN => n_1418);
   REGISTERS_reg_24_31_inst : DFFR_X1 port map( D => n2825, CK => CLK, RN => 
                           n1517, Q => n4851, QN => n4104);
   REGISTERS_reg_24_30_inst : DFFR_X1 port map( D => n2824, CK => CLK, RN => 
                           n1517, Q => n4850, QN => n4070);
   REGISTERS_reg_24_29_inst : DFFR_X1 port map( D => n2823, CK => CLK, RN => 
                           n1517, Q => n4849, QN => n4044);
   REGISTERS_reg_24_28_inst : DFFR_X1 port map( D => n2822, CK => CLK, RN => 
                           n1517, Q => n4848, QN => n4018);
   REGISTERS_reg_24_27_inst : DFFR_X1 port map( D => n2821, CK => CLK, RN => 
                           n1517, Q => n4847, QN => n3992);
   REGISTERS_reg_24_26_inst : DFFR_X1 port map( D => n2820, CK => CLK, RN => 
                           n1517, Q => n4846, QN => n3966);
   REGISTERS_reg_24_25_inst : DFFR_X1 port map( D => n2819, CK => CLK, RN => 
                           n1517, Q => n4845, QN => n3940);
   REGISTERS_reg_24_24_inst : DFFR_X1 port map( D => n2818, CK => CLK, RN => 
                           n1517, Q => n4844, QN => n3914);
   REGISTERS_reg_24_23_inst : DFFR_X1 port map( D => n2817, CK => CLK, RN => 
                           n1518, Q => n4843, QN => n3888);
   REGISTERS_reg_24_22_inst : DFFR_X1 port map( D => n2816, CK => CLK, RN => 
                           n1518, Q => n4842, QN => n3863);
   REGISTERS_reg_24_21_inst : DFFR_X1 port map( D => n2815, CK => CLK, RN => 
                           n1518, Q => n4841, QN => n3838);
   REGISTERS_reg_24_20_inst : DFFR_X1 port map( D => n2814, CK => CLK, RN => 
                           n1518, Q => n4840, QN => n3813);
   REGISTERS_reg_24_19_inst : DFFR_X1 port map( D => n2813, CK => CLK, RN => 
                           n1518, Q => n4839, QN => n3788);
   REGISTERS_reg_24_18_inst : DFFR_X1 port map( D => n2812, CK => CLK, RN => 
                           n1518, Q => n4838, QN => n3763);
   REGISTERS_reg_24_17_inst : DFFR_X1 port map( D => n2811, CK => CLK, RN => 
                           n1518, Q => n4837, QN => n3738);
   REGISTERS_reg_24_16_inst : DFFR_X1 port map( D => n2810, CK => CLK, RN => 
                           n1518, Q => n4836, QN => n3713);
   REGISTERS_reg_24_15_inst : DFFR_X1 port map( D => n2809, CK => CLK, RN => 
                           n1518, Q => n4835, QN => n3688);
   REGISTERS_reg_24_14_inst : DFFR_X1 port map( D => n2808, CK => CLK, RN => 
                           n1518, Q => n4834, QN => n3663);
   REGISTERS_reg_24_13_inst : DFFR_X1 port map( D => n2807, CK => CLK, RN => 
                           n1518, Q => n4833, QN => n3638);
   REGISTERS_reg_24_12_inst : DFFR_X1 port map( D => n2806, CK => CLK, RN => 
                           n1518, Q => n4832, QN => n3613);
   REGISTERS_reg_24_11_inst : DFFR_X1 port map( D => n2805, CK => CLK, RN => 
                           n1519, Q => n4831, QN => n3588);
   REGISTERS_reg_24_10_inst : DFFR_X1 port map( D => n2804, CK => CLK, RN => 
                           n1519, Q => n4830, QN => n3563);
   REGISTERS_reg_24_9_inst : DFFR_X1 port map( D => n2803, CK => CLK, RN => 
                           n1519, Q => n4829, QN => n2482);
   REGISTERS_reg_24_8_inst : DFFR_X1 port map( D => n2802, CK => CLK, RN => 
                           n1519, Q => n4828, QN => n2457);
   REGISTERS_reg_24_7_inst : DFFR_X1 port map( D => n2801, CK => CLK, RN => 
                           n1519, Q => n4827, QN => n2432);
   REGISTERS_reg_24_6_inst : DFFR_X1 port map( D => n2800, CK => CLK, RN => 
                           n1519, Q => n4826, QN => n2407);
   REGISTERS_reg_24_5_inst : DFFR_X1 port map( D => n2799, CK => CLK, RN => 
                           n1519, Q => n4825, QN => n2382);
   REGISTERS_reg_24_4_inst : DFFR_X1 port map( D => n2798, CK => CLK, RN => 
                           n1519, Q => n4824, QN => n2357);
   REGISTERS_reg_24_3_inst : DFFR_X1 port map( D => n2797, CK => CLK, RN => 
                           n1519, Q => n4823, QN => n2332);
   REGISTERS_reg_24_2_inst : DFFR_X1 port map( D => n2796, CK => CLK, RN => 
                           n1519, Q => n4822, QN => n2307);
   REGISTERS_reg_24_1_inst : DFFR_X1 port map( D => n2795, CK => CLK, RN => 
                           n1519, Q => n4821, QN => n2282);
   REGISTERS_reg_24_0_inst : DFFR_X1 port map( D => n2794, CK => CLK, RN => 
                           n1519, Q => n4820, QN => n2253);
   REGISTERS_reg_25_31_inst : DFFR_X1 port map( D => n2793, CK => CLK, RN => 
                           n1520, Q => n4819, QN => n_1419);
   REGISTERS_reg_25_30_inst : DFFR_X1 port map( D => n2792, CK => CLK, RN => 
                           n1520, Q => n4818, QN => n_1420);
   REGISTERS_reg_25_29_inst : DFFR_X1 port map( D => n2791, CK => CLK, RN => 
                           n1520, Q => n4817, QN => n_1421);
   REGISTERS_reg_25_28_inst : DFFR_X1 port map( D => n2790, CK => CLK, RN => 
                           n1520, Q => n4816, QN => n_1422);
   REGISTERS_reg_25_27_inst : DFFR_X1 port map( D => n2789, CK => CLK, RN => 
                           n1520, Q => n4815, QN => n_1423);
   REGISTERS_reg_25_26_inst : DFFR_X1 port map( D => n2788, CK => CLK, RN => 
                           n1520, Q => n4814, QN => n_1424);
   REGISTERS_reg_25_25_inst : DFFR_X1 port map( D => n2787, CK => CLK, RN => 
                           n1520, Q => n4813, QN => n_1425);
   REGISTERS_reg_25_24_inst : DFFR_X1 port map( D => n2786, CK => CLK, RN => 
                           n1520, Q => n4812, QN => n_1426);
   REGISTERS_reg_25_23_inst : DFFR_X1 port map( D => n2785, CK => CLK, RN => 
                           n1520, Q => n4811, QN => n_1427);
   REGISTERS_reg_25_22_inst : DFFR_X1 port map( D => n2784, CK => CLK, RN => 
                           n1520, Q => n4810, QN => n_1428);
   REGISTERS_reg_25_21_inst : DFFR_X1 port map( D => n2783, CK => CLK, RN => 
                           n1520, Q => n4809, QN => n_1429);
   REGISTERS_reg_25_20_inst : DFFR_X1 port map( D => n2782, CK => CLK, RN => 
                           n1520, Q => n4808, QN => n_1430);
   REGISTERS_reg_25_19_inst : DFFR_X1 port map( D => n2781, CK => CLK, RN => 
                           n1521, Q => n4807, QN => n_1431);
   REGISTERS_reg_25_18_inst : DFFR_X1 port map( D => n2780, CK => CLK, RN => 
                           n1521, Q => n4806, QN => n_1432);
   REGISTERS_reg_25_17_inst : DFFR_X1 port map( D => n2779, CK => CLK, RN => 
                           n1521, Q => n4805, QN => n_1433);
   REGISTERS_reg_25_16_inst : DFFR_X1 port map( D => n2778, CK => CLK, RN => 
                           n1521, Q => n4804, QN => n_1434);
   REGISTERS_reg_25_15_inst : DFFR_X1 port map( D => n2777, CK => CLK, RN => 
                           n1521, Q => n4803, QN => n_1435);
   REGISTERS_reg_25_14_inst : DFFR_X1 port map( D => n2776, CK => CLK, RN => 
                           n1521, Q => n4802, QN => n_1436);
   REGISTERS_reg_25_13_inst : DFFR_X1 port map( D => n2775, CK => CLK, RN => 
                           n1521, Q => n4801, QN => n_1437);
   REGISTERS_reg_25_12_inst : DFFR_X1 port map( D => n2774, CK => CLK, RN => 
                           n1521, Q => n4800, QN => n_1438);
   REGISTERS_reg_25_11_inst : DFFR_X1 port map( D => n2773, CK => CLK, RN => 
                           n1521, Q => n4799, QN => n_1439);
   REGISTERS_reg_25_10_inst : DFFR_X1 port map( D => n2772, CK => CLK, RN => 
                           n1521, Q => n4798, QN => n_1440);
   REGISTERS_reg_25_9_inst : DFFR_X1 port map( D => n2771, CK => CLK, RN => 
                           n1521, Q => n4797, QN => n_1441);
   REGISTERS_reg_25_8_inst : DFFR_X1 port map( D => n2770, CK => CLK, RN => 
                           n1521, Q => n4796, QN => n_1442);
   REGISTERS_reg_25_7_inst : DFFR_X1 port map( D => n2769, CK => CLK, RN => 
                           n1522, Q => n4795, QN => n_1443);
   REGISTERS_reg_25_6_inst : DFFR_X1 port map( D => n2768, CK => CLK, RN => 
                           n1522, Q => n4794, QN => n_1444);
   REGISTERS_reg_25_5_inst : DFFR_X1 port map( D => n2767, CK => CLK, RN => 
                           n1522, Q => n4793, QN => n_1445);
   REGISTERS_reg_25_4_inst : DFFR_X1 port map( D => n2766, CK => CLK, RN => 
                           n1522, Q => n4792, QN => n_1446);
   REGISTERS_reg_25_3_inst : DFFR_X1 port map( D => n2765, CK => CLK, RN => 
                           n1522, Q => n4791, QN => n_1447);
   REGISTERS_reg_25_2_inst : DFFR_X1 port map( D => n2764, CK => CLK, RN => 
                           n1522, Q => n4790, QN => n_1448);
   REGISTERS_reg_25_1_inst : DFFR_X1 port map( D => n2763, CK => CLK, RN => 
                           n1522, Q => n4789, QN => n_1449);
   REGISTERS_reg_25_0_inst : DFFR_X1 port map( D => n2762, CK => CLK, RN => 
                           n1522, Q => n4788, QN => n_1450);
   REGISTERS_reg_26_23_inst : DFFR_X1 port map( D => n2753, CK => CLK, RN => 
                           n1523, Q => n4296, QN => n813);
   REGISTERS_reg_26_22_inst : DFFR_X1 port map( D => n2752, CK => CLK, RN => 
                           n1523, Q => n4297, QN => n814);
   REGISTERS_reg_26_21_inst : DFFR_X1 port map( D => n2751, CK => CLK, RN => 
                           n1523, Q => n224, QN => n815);
   REGISTERS_reg_26_20_inst : DFFR_X1 port map( D => n2750, CK => CLK, RN => 
                           n1523, Q => n4298, QN => n816);
   REGISTERS_reg_26_19_inst : DFFR_X1 port map( D => n2749, CK => CLK, RN => 
                           n1523, Q => n343, QN => n817);
   REGISTERS_reg_26_18_inst : DFFR_X1 port map( D => n2748, CK => CLK, RN => 
                           n1523, Q => n344, QN => n818);
   REGISTERS_reg_26_17_inst : DFFR_X1 port map( D => n2747, CK => CLK, RN => 
                           n1523, Q => n225, QN => n819);
   REGISTERS_reg_26_16_inst : DFFR_X1 port map( D => n2746, CK => CLK, RN => 
                           n1523, Q => n4299, QN => n820);
   REGISTERS_reg_26_15_inst : DFFR_X1 port map( D => n2745, CK => CLK, RN => 
                           n1524, Q => n345, QN => n821);
   REGISTERS_reg_26_14_inst : DFFR_X1 port map( D => n2744, CK => CLK, RN => 
                           n1524, Q => n4300, QN => n822);
   REGISTERS_reg_26_13_inst : DFFR_X1 port map( D => n2743, CK => CLK, RN => 
                           n1524, Q => n4301, QN => n823);
   REGISTERS_reg_26_12_inst : DFFR_X1 port map( D => n2742, CK => CLK, RN => 
                           n1524, Q => n346, QN => n824);
   REGISTERS_reg_26_11_inst : DFFR_X1 port map( D => n2741, CK => CLK, RN => 
                           n1524, Q => n4302, QN => n825);
   REGISTERS_reg_26_10_inst : DFFR_X1 port map( D => n2740, CK => CLK, RN => 
                           n1524, Q => n226, QN => n826);
   REGISTERS_reg_26_9_inst : DFFR_X1 port map( D => n2739, CK => CLK, RN => 
                           n1524, Q => n4303, QN => n827);
   REGISTERS_reg_26_8_inst : DFFR_X1 port map( D => n2738, CK => CLK, RN => 
                           n1524, Q => n347, QN => n828);
   REGISTERS_reg_26_7_inst : DFFR_X1 port map( D => n2737, CK => CLK, RN => 
                           n1524, Q => n4304, QN => n829);
   REGISTERS_reg_26_6_inst : DFFR_X1 port map( D => n2736, CK => CLK, RN => 
                           n1524, Q => n4305, QN => n830);
   REGISTERS_reg_26_5_inst : DFFR_X1 port map( D => n2735, CK => CLK, RN => 
                           n1524, Q => n351, QN => n831);
   REGISTERS_reg_26_4_inst : DFFR_X1 port map( D => n2734, CK => CLK, RN => 
                           n1524, Q => n348, QN => n832);
   REGISTERS_reg_26_3_inst : DFFR_X1 port map( D => n2733, CK => CLK, RN => 
                           n1525, Q => n349, QN => n833);
   REGISTERS_reg_26_2_inst : DFFR_X1 port map( D => n2732, CK => CLK, RN => 
                           n1525, Q => n4306, QN => n834);
   REGISTERS_reg_26_1_inst : DFFR_X1 port map( D => n2731, CK => CLK, RN => 
                           n1525, Q => n350, QN => n835);
   REGISTERS_reg_26_0_inst : DFFR_X1 port map( D => n2730, CK => CLK, RN => 
                           n1525, Q => n4307, QN => n836);
   REGISTERS_reg_27_23_inst : DFFR_X1 port map( D => n2721, CK => CLK, RN => 
                           n1526, Q => n3891, QN => n845);
   REGISTERS_reg_27_22_inst : DFFR_X1 port map( D => n2720, CK => CLK, RN => 
                           n1526, Q => n3866, QN => n846);
   REGISTERS_reg_27_21_inst : DFFR_X1 port map( D => n2719, CK => CLK, RN => 
                           n1526, Q => n3841, QN => n847);
   REGISTERS_reg_27_20_inst : DFFR_X1 port map( D => n2718, CK => CLK, RN => 
                           n1526, Q => n3816, QN => n848);
   REGISTERS_reg_27_19_inst : DFFR_X1 port map( D => n2717, CK => CLK, RN => 
                           n1526, Q => n3791, QN => n849);
   REGISTERS_reg_27_18_inst : DFFR_X1 port map( D => n2716, CK => CLK, RN => 
                           n1526, Q => n3766, QN => n850);
   REGISTERS_reg_27_17_inst : DFFR_X1 port map( D => n2715, CK => CLK, RN => 
                           n1526, Q => n3741, QN => n851);
   REGISTERS_reg_27_16_inst : DFFR_X1 port map( D => n2714, CK => CLK, RN => 
                           n1526, Q => n3716, QN => n852);
   REGISTERS_reg_27_15_inst : DFFR_X1 port map( D => n2713, CK => CLK, RN => 
                           n1526, Q => n3691, QN => n853);
   REGISTERS_reg_27_14_inst : DFFR_X1 port map( D => n2712, CK => CLK, RN => 
                           n1526, Q => n3666, QN => n854);
   REGISTERS_reg_27_13_inst : DFFR_X1 port map( D => n2711, CK => CLK, RN => 
                           n1526, Q => n3641, QN => n855);
   REGISTERS_reg_27_12_inst : DFFR_X1 port map( D => n2710, CK => CLK, RN => 
                           n1526, Q => n3616, QN => n856);
   REGISTERS_reg_27_11_inst : DFFR_X1 port map( D => n2709, CK => CLK, RN => 
                           n1527, Q => n3591, QN => n857);
   REGISTERS_reg_27_10_inst : DFFR_X1 port map( D => n2708, CK => CLK, RN => 
                           n1527, Q => n3566, QN => n858);
   REGISTERS_reg_27_9_inst : DFFR_X1 port map( D => n2707, CK => CLK, RN => 
                           n1527, Q => n2485, QN => n859);
   REGISTERS_reg_27_8_inst : DFFR_X1 port map( D => n2706, CK => CLK, RN => 
                           n1527, Q => n2460, QN => n860);
   REGISTERS_reg_27_7_inst : DFFR_X1 port map( D => n2705, CK => CLK, RN => 
                           n1527, Q => n2435, QN => n861);
   REGISTERS_reg_27_6_inst : DFFR_X1 port map( D => n2704, CK => CLK, RN => 
                           n1527, Q => n2410, QN => n862);
   REGISTERS_reg_27_5_inst : DFFR_X1 port map( D => n2703, CK => CLK, RN => 
                           n1527, Q => n2385, QN => n863);
   REGISTERS_reg_27_4_inst : DFFR_X1 port map( D => n2702, CK => CLK, RN => 
                           n1527, Q => n2360, QN => n864);
   REGISTERS_reg_27_3_inst : DFFR_X1 port map( D => n2701, CK => CLK, RN => 
                           n1527, Q => n2335, QN => n865);
   REGISTERS_reg_27_2_inst : DFFR_X1 port map( D => n2700, CK => CLK, RN => 
                           n1527, Q => n2310, QN => n866);
   REGISTERS_reg_27_1_inst : DFFR_X1 port map( D => n2699, CK => CLK, RN => 
                           n1527, Q => n2285, QN => n867);
   REGISTERS_reg_27_0_inst : DFFR_X1 port map( D => n2698, CK => CLK, RN => 
                           n1527, Q => n2256, QN => n868);
   REGISTERS_reg_28_31_inst : DFFR_X1 port map( D => n2697, CK => CLK, RN => 
                           n1528, Q => n4787, QN => n4112);
   REGISTERS_reg_28_30_inst : DFFR_X1 port map( D => n2696, CK => CLK, RN => 
                           n1528, Q => n4786, QN => n4074);
   REGISTERS_reg_28_29_inst : DFFR_X1 port map( D => n2695, CK => CLK, RN => 
                           n1528, Q => n4785, QN => n4048);
   REGISTERS_reg_28_28_inst : DFFR_X1 port map( D => n2694, CK => CLK, RN => 
                           n1528, Q => n4784, QN => n4022);
   REGISTERS_reg_28_27_inst : DFFR_X1 port map( D => n2693, CK => CLK, RN => 
                           n1528, Q => n4783, QN => n3996);
   REGISTERS_reg_28_26_inst : DFFR_X1 port map( D => n2692, CK => CLK, RN => 
                           n1528, Q => n4782, QN => n3970);
   REGISTERS_reg_28_25_inst : DFFR_X1 port map( D => n2691, CK => CLK, RN => 
                           n1528, Q => n4781, QN => n3944);
   REGISTERS_reg_28_24_inst : DFFR_X1 port map( D => n2690, CK => CLK, RN => 
                           n1528, Q => n4780, QN => n3918);
   REGISTERS_reg_28_23_inst : DFFR_X1 port map( D => n2689, CK => CLK, RN => 
                           n1528, Q => n4779, QN => n3892);
   REGISTERS_reg_28_22_inst : DFFR_X1 port map( D => n2688, CK => CLK, RN => 
                           n1528, Q => n4778, QN => n3867);
   REGISTERS_reg_28_21_inst : DFFR_X1 port map( D => n2687, CK => CLK, RN => 
                           n1528, Q => n4777, QN => n3842);
   REGISTERS_reg_28_20_inst : DFFR_X1 port map( D => n2686, CK => CLK, RN => 
                           n1528, Q => n4776, QN => n3817);
   REGISTERS_reg_28_19_inst : DFFR_X1 port map( D => n2685, CK => CLK, RN => 
                           n1529, Q => n4775, QN => n3792);
   REGISTERS_reg_28_18_inst : DFFR_X1 port map( D => n2684, CK => CLK, RN => 
                           n1529, Q => n4774, QN => n3767);
   REGISTERS_reg_28_17_inst : DFFR_X1 port map( D => n2683, CK => CLK, RN => 
                           n1529, Q => n4773, QN => n3742);
   REGISTERS_reg_28_16_inst : DFFR_X1 port map( D => n2682, CK => CLK, RN => 
                           n1529, Q => n4772, QN => n3717);
   REGISTERS_reg_28_15_inst : DFFR_X1 port map( D => n2681, CK => CLK, RN => 
                           n1529, Q => n4771, QN => n3692);
   REGISTERS_reg_28_14_inst : DFFR_X1 port map( D => n2680, CK => CLK, RN => 
                           n1529, Q => n4770, QN => n3667);
   REGISTERS_reg_28_13_inst : DFFR_X1 port map( D => n2679, CK => CLK, RN => 
                           n1529, Q => n4769, QN => n3642);
   REGISTERS_reg_28_12_inst : DFFR_X1 port map( D => n2678, CK => CLK, RN => 
                           n1529, Q => n4768, QN => n3617);
   REGISTERS_reg_28_11_inst : DFFR_X1 port map( D => n2677, CK => CLK, RN => 
                           n1529, Q => n4767, QN => n3592);
   REGISTERS_reg_28_10_inst : DFFR_X1 port map( D => n2676, CK => CLK, RN => 
                           n1529, Q => n4766, QN => n3567);
   REGISTERS_reg_28_9_inst : DFFR_X1 port map( D => n2675, CK => CLK, RN => 
                           n1529, Q => n4765, QN => n2486);
   REGISTERS_reg_28_8_inst : DFFR_X1 port map( D => n2674, CK => CLK, RN => 
                           n1529, Q => n4764, QN => n2461);
   REGISTERS_reg_28_7_inst : DFFR_X1 port map( D => n2673, CK => CLK, RN => 
                           n1530, Q => n4763, QN => n2436);
   REGISTERS_reg_28_6_inst : DFFR_X1 port map( D => n2672, CK => CLK, RN => 
                           n1530, Q => n4762, QN => n2411);
   REGISTERS_reg_28_5_inst : DFFR_X1 port map( D => n2671, CK => CLK, RN => 
                           n1530, Q => n4761, QN => n2386);
   REGISTERS_reg_28_4_inst : DFFR_X1 port map( D => n2670, CK => CLK, RN => 
                           n1530, Q => n4760, QN => n2361);
   REGISTERS_reg_28_3_inst : DFFR_X1 port map( D => n2669, CK => CLK, RN => 
                           n1530, Q => n4759, QN => n2336);
   REGISTERS_reg_28_2_inst : DFFR_X1 port map( D => n2668, CK => CLK, RN => 
                           n1530, Q => n4758, QN => n2311);
   REGISTERS_reg_28_1_inst : DFFR_X1 port map( D => n2667, CK => CLK, RN => 
                           n1530, Q => n4757, QN => n2286);
   REGISTERS_reg_28_0_inst : DFFR_X1 port map( D => n2666, CK => CLK, RN => 
                           n1530, Q => n4756, QN => n2257);
   REGISTERS_reg_29_31_inst : DFFR_X1 port map( D => n2665, CK => CLK, RN => 
                           n1530, Q => n4755, QN => n321);
   REGISTERS_reg_29_30_inst : DFFR_X1 port map( D => n2664, CK => CLK, RN => 
                           n1530, Q => n4754, QN => n320);
   REGISTERS_reg_29_29_inst : DFFR_X1 port map( D => n2663, CK => CLK, RN => 
                           n1530, Q => n4753, QN => n319);
   REGISTERS_reg_29_28_inst : DFFR_X1 port map( D => n2662, CK => CLK, RN => 
                           n1530, Q => n4752, QN => n318);
   REGISTERS_reg_29_27_inst : DFFR_X1 port map( D => n2661, CK => CLK, RN => 
                           n1531, Q => n4751, QN => n317);
   REGISTERS_reg_29_26_inst : DFFR_X1 port map( D => n2660, CK => CLK, RN => 
                           n1531, Q => n4750, QN => n316);
   REGISTERS_reg_29_25_inst : DFFR_X1 port map( D => n2659, CK => CLK, RN => 
                           n1531, Q => n4749, QN => n315);
   REGISTERS_reg_29_24_inst : DFFR_X1 port map( D => n2658, CK => CLK, RN => 
                           n1531, Q => n4748, QN => n314);
   REGISTERS_reg_29_23_inst : DFFR_X1 port map( D => n2657, CK => CLK, RN => 
                           n1531, Q => n4747, QN => n313);
   REGISTERS_reg_29_22_inst : DFFR_X1 port map( D => n2656, CK => CLK, RN => 
                           n1531, Q => n4746, QN => n312);
   REGISTERS_reg_29_21_inst : DFFR_X1 port map( D => n2655, CK => CLK, RN => 
                           n1531, Q => n4745, QN => n311);
   REGISTERS_reg_29_20_inst : DFFR_X1 port map( D => n2654, CK => CLK, RN => 
                           n1531, Q => n4744, QN => n310);
   REGISTERS_reg_29_19_inst : DFFR_X1 port map( D => n2653, CK => CLK, RN => 
                           n1531, Q => n4743, QN => n309);
   REGISTERS_reg_29_18_inst : DFFR_X1 port map( D => n2652, CK => CLK, RN => 
                           n1531, Q => n4742, QN => n308);
   REGISTERS_reg_29_17_inst : DFFR_X1 port map( D => n2651, CK => CLK, RN => 
                           n1531, Q => n4741, QN => n307);
   REGISTERS_reg_29_16_inst : DFFR_X1 port map( D => n2650, CK => CLK, RN => 
                           n1531, Q => n4740, QN => n306);
   REGISTERS_reg_29_15_inst : DFFR_X1 port map( D => n2649, CK => CLK, RN => 
                           n1532, Q => n4739, QN => n305);
   REGISTERS_reg_29_14_inst : DFFR_X1 port map( D => n2648, CK => CLK, RN => 
                           n1532, Q => n4738, QN => n304);
   REGISTERS_reg_29_13_inst : DFFR_X1 port map( D => n2647, CK => CLK, RN => 
                           n1532, Q => n4737, QN => n303);
   REGISTERS_reg_29_12_inst : DFFR_X1 port map( D => n2646, CK => CLK, RN => 
                           n1532, Q => n4736, QN => n461);
   REGISTERS_reg_29_11_inst : DFFR_X1 port map( D => n2645, CK => CLK, RN => 
                           n1532, Q => n4735, QN => n302);
   REGISTERS_reg_29_10_inst : DFFR_X1 port map( D => n2644, CK => CLK, RN => 
                           n1532, Q => n4734, QN => n301);
   REGISTERS_reg_29_9_inst : DFFR_X1 port map( D => n2643, CK => CLK, RN => 
                           n1532, Q => n4733, QN => n300);
   REGISTERS_reg_29_8_inst : DFFR_X1 port map( D => n2642, CK => CLK, RN => 
                           n1532, Q => n4732, QN => n299);
   REGISTERS_reg_29_7_inst : DFFR_X1 port map( D => n2641, CK => CLK, RN => 
                           n1532, Q => n4731, QN => n298);
   REGISTERS_reg_29_6_inst : DFFR_X1 port map( D => n2640, CK => CLK, RN => 
                           n1532, Q => n4730, QN => n297);
   REGISTERS_reg_29_5_inst : DFFR_X1 port map( D => n2639, CK => CLK, RN => 
                           n1532, Q => n4729, QN => n296);
   REGISTERS_reg_29_4_inst : DFFR_X1 port map( D => n2638, CK => CLK, RN => 
                           n1532, Q => n4728, QN => n295);
   REGISTERS_reg_29_3_inst : DFFR_X1 port map( D => n2637, CK => CLK, RN => 
                           n1533, Q => n4727, QN => n294);
   REGISTERS_reg_29_2_inst : DFFR_X1 port map( D => n2636, CK => CLK, RN => 
                           n1533, Q => n4726, QN => n293);
   REGISTERS_reg_29_1_inst : DFFR_X1 port map( D => n2635, CK => CLK, RN => 
                           n1533, Q => n4725, QN => n228);
   REGISTERS_reg_29_0_inst : DFFR_X1 port map( D => n2634, CK => CLK, RN => 
                           n1533, Q => n4724, QN => n227);
   REGISTERS_reg_30_23_inst : DFFR_X1 port map( D => n2625, CK => CLK, RN => 
                           n1534, Q => n_1451, QN => n941);
   REGISTERS_reg_30_22_inst : DFFR_X1 port map( D => n2624, CK => CLK, RN => 
                           n1534, Q => n_1452, QN => n942);
   REGISTERS_reg_30_21_inst : DFFR_X1 port map( D => n2623, CK => CLK, RN => 
                           n1534, Q => n_1453, QN => n943);
   REGISTERS_reg_30_20_inst : DFFR_X1 port map( D => n2622, CK => CLK, RN => 
                           n1534, Q => n_1454, QN => n944);
   REGISTERS_reg_30_19_inst : DFFR_X1 port map( D => n2621, CK => CLK, RN => 
                           n1534, Q => n_1455, QN => n945);
   REGISTERS_reg_30_18_inst : DFFR_X1 port map( D => n2620, CK => CLK, RN => 
                           n1534, Q => n_1456, QN => n946);
   REGISTERS_reg_30_17_inst : DFFR_X1 port map( D => n2619, CK => CLK, RN => 
                           n1534, Q => n_1457, QN => n947);
   REGISTERS_reg_30_16_inst : DFFR_X1 port map( D => n2618, CK => CLK, RN => 
                           n1534, Q => n_1458, QN => n948);
   REGISTERS_reg_30_15_inst : DFFR_X1 port map( D => n2617, CK => CLK, RN => 
                           n1534, Q => n_1459, QN => n949);
   REGISTERS_reg_30_14_inst : DFFR_X1 port map( D => n2616, CK => CLK, RN => 
                           n1534, Q => n_1460, QN => n950);
   REGISTERS_reg_30_13_inst : DFFR_X1 port map( D => n2615, CK => CLK, RN => 
                           n1534, Q => n_1461, QN => n951);
   REGISTERS_reg_30_12_inst : DFFR_X1 port map( D => n2614, CK => CLK, RN => 
                           n1534, Q => n_1462, QN => n952);
   REGISTERS_reg_30_11_inst : DFFR_X1 port map( D => n2613, CK => CLK, RN => 
                           n1535, Q => n_1463, QN => n953);
   REGISTERS_reg_30_10_inst : DFFR_X1 port map( D => n2612, CK => CLK, RN => 
                           n1535, Q => n_1464, QN => n954);
   REGISTERS_reg_30_9_inst : DFFR_X1 port map( D => n2611, CK => CLK, RN => 
                           n1535, Q => n_1465, QN => n955);
   REGISTERS_reg_30_8_inst : DFFR_X1 port map( D => n2610, CK => CLK, RN => 
                           n1535, Q => n_1466, QN => n956);
   REGISTERS_reg_30_7_inst : DFFR_X1 port map( D => n2609, CK => CLK, RN => 
                           n1535, Q => n_1467, QN => n957);
   REGISTERS_reg_30_6_inst : DFFR_X1 port map( D => n2608, CK => CLK, RN => 
                           n1535, Q => n_1468, QN => n958);
   REGISTERS_reg_30_5_inst : DFFR_X1 port map( D => n2607, CK => CLK, RN => 
                           n1535, Q => n_1469, QN => n959);
   REGISTERS_reg_30_4_inst : DFFR_X1 port map( D => n2606, CK => CLK, RN => 
                           n1535, Q => n_1470, QN => n960);
   REGISTERS_reg_30_3_inst : DFFR_X1 port map( D => n2605, CK => CLK, RN => 
                           n1535, Q => n_1471, QN => n961);
   REGISTERS_reg_30_2_inst : DFFR_X1 port map( D => n2604, CK => CLK, RN => 
                           n1535, Q => n_1472, QN => n962);
   REGISTERS_reg_30_1_inst : DFFR_X1 port map( D => n2603, CK => CLK, RN => 
                           n1535, Q => n_1473, QN => n963);
   REGISTERS_reg_30_0_inst : DFFR_X1 port map( D => n2602, CK => CLK, RN => 
                           n1535, Q => n_1474, QN => n964);
   REGISTERS_reg_31_23_inst : DFFR_X1 port map( D => n2593, CK => CLK, RN => 
                           n1536, Q => n4316, QN => n_1475);
   REGISTERS_reg_31_22_inst : DFFR_X1 port map( D => n2592, CK => CLK, RN => 
                           n1536, Q => n4317, QN => n_1476);
   REGISTERS_reg_31_21_inst : DFFR_X1 port map( D => n2591, CK => CLK, RN => 
                           n1536, Q => n4318, QN => n_1477);
   REGISTERS_reg_31_20_inst : DFFR_X1 port map( D => n2590, CK => CLK, RN => 
                           n1536, Q => n4319, QN => n_1478);
   REGISTERS_reg_31_19_inst : DFFR_X1 port map( D => n2589, CK => CLK, RN => 
                           n1537, Q => n4320, QN => n_1479);
   REGISTERS_reg_31_18_inst : DFFR_X1 port map( D => n2588, CK => CLK, RN => 
                           n1537, Q => n4321, QN => n_1480);
   REGISTERS_reg_31_17_inst : DFFR_X1 port map( D => n2587, CK => CLK, RN => 
                           n1537, Q => n4322, QN => n_1481);
   REGISTERS_reg_31_16_inst : DFFR_X1 port map( D => n2586, CK => CLK, RN => 
                           n1537, Q => n4323, QN => n_1482);
   REGISTERS_reg_31_15_inst : DFFR_X1 port map( D => n2585, CK => CLK, RN => 
                           n1537, Q => n4324, QN => n_1483);
   REGISTERS_reg_31_14_inst : DFFR_X1 port map( D => n2584, CK => CLK, RN => 
                           n1537, Q => n4325, QN => n_1484);
   REGISTERS_reg_31_13_inst : DFFR_X1 port map( D => n2583, CK => CLK, RN => 
                           n1537, Q => n4326, QN => n_1485);
   REGISTERS_reg_31_12_inst : DFFR_X1 port map( D => n2582, CK => CLK, RN => 
                           n1537, Q => n4327, QN => n_1486);
   REGISTERS_reg_31_11_inst : DFFR_X1 port map( D => n2581, CK => CLK, RN => 
                           n1537, Q => n4328, QN => n_1487);
   REGISTERS_reg_31_10_inst : DFFR_X1 port map( D => n2580, CK => CLK, RN => 
                           n1537, Q => n4329, QN => n_1488);
   REGISTERS_reg_31_9_inst : DFFR_X1 port map( D => n2579, CK => CLK, RN => 
                           n1537, Q => n4330, QN => n_1489);
   REGISTERS_reg_31_8_inst : DFFR_X1 port map( D => n2578, CK => CLK, RN => 
                           n1537, Q => n4331, QN => n_1490);
   REGISTERS_reg_31_7_inst : DFFR_X1 port map( D => n2577, CK => CLK, RN => 
                           n1538, Q => n4332, QN => n_1491);
   REGISTERS_reg_31_6_inst : DFFR_X1 port map( D => n2576, CK => CLK, RN => 
                           n1538, Q => n4333, QN => n_1492);
   REGISTERS_reg_31_5_inst : DFFR_X1 port map( D => n2575, CK => CLK, RN => 
                           n1538, Q => n4334, QN => n_1493);
   REGISTERS_reg_31_4_inst : DFFR_X1 port map( D => n2574, CK => CLK, RN => 
                           n1538, Q => n4335, QN => n_1494);
   REGISTERS_reg_31_3_inst : DFFR_X1 port map( D => n2573, CK => CLK, RN => 
                           n1538, Q => n4336, QN => n_1495);
   REGISTERS_reg_31_2_inst : DFFR_X1 port map( D => n2572, CK => CLK, RN => 
                           n1538, Q => n4337, QN => n_1496);
   REGISTERS_reg_31_1_inst : DFFR_X1 port map( D => n2571, CK => CLK, RN => 
                           n1538, Q => n4338, QN => n_1497);
   REGISTERS_reg_31_0_inst : DFFR_X1 port map( D => n2570, CK => CLK, RN => 
                           n1538, Q => n4339, QN => n_1498);
   OUT2_reg_31_inst : DFF_X1 port map( D => n2569, CK => CLK, Q => OUT2(31), QN
                           => n4723);
   OUT2_reg_30_inst : DFF_X1 port map( D => n2568, CK => CLK, Q => OUT2(30), QN
                           => n4722);
   OUT2_reg_29_inst : DFF_X1 port map( D => n2567, CK => CLK, Q => OUT2(29), QN
                           => n4721);
   OUT2_reg_28_inst : DFF_X1 port map( D => n2566, CK => CLK, Q => OUT2(28), QN
                           => n4720);
   OUT2_reg_27_inst : DFF_X1 port map( D => n2565, CK => CLK, Q => OUT2(27), QN
                           => n4719);
   OUT2_reg_26_inst : DFF_X1 port map( D => n2564, CK => CLK, Q => OUT2(26), QN
                           => n4718);
   OUT2_reg_25_inst : DFF_X1 port map( D => n2563, CK => CLK, Q => OUT2(25), QN
                           => n4717);
   OUT2_reg_24_inst : DFF_X1 port map( D => n2562, CK => CLK, Q => OUT2(24), QN
                           => n4716);
   OUT2_reg_23_inst : DFF_X1 port map( D => n2561, CK => CLK, Q => OUT2(23), QN
                           => n4715);
   OUT2_reg_22_inst : DFF_X1 port map( D => n2560, CK => CLK, Q => OUT2(22), QN
                           => n4714);
   OUT2_reg_21_inst : DFF_X1 port map( D => n2559, CK => CLK, Q => OUT2(21), QN
                           => n4713);
   OUT2_reg_20_inst : DFF_X1 port map( D => n2558, CK => CLK, Q => OUT2(20), QN
                           => n4712);
   OUT2_reg_19_inst : DFF_X1 port map( D => n2557, CK => CLK, Q => OUT2(19), QN
                           => n4711);
   OUT2_reg_18_inst : DFF_X1 port map( D => n2556, CK => CLK, Q => OUT2(18), QN
                           => n4710);
   OUT2_reg_17_inst : DFF_X1 port map( D => n2555, CK => CLK, Q => OUT2(17), QN
                           => n4709);
   OUT2_reg_16_inst : DFF_X1 port map( D => n2554, CK => CLK, Q => OUT2(16), QN
                           => n4708);
   OUT2_reg_15_inst : DFF_X1 port map( D => n2553, CK => CLK, Q => OUT2(15), QN
                           => n4707);
   OUT2_reg_14_inst : DFF_X1 port map( D => n2552, CK => CLK, Q => OUT2(14), QN
                           => n4706);
   OUT2_reg_13_inst : DFF_X1 port map( D => n2551, CK => CLK, Q => OUT2(13), QN
                           => n4705);
   OUT2_reg_12_inst : DFF_X1 port map( D => n2550, CK => CLK, Q => OUT2(12), QN
                           => n4704);
   OUT2_reg_11_inst : DFF_X1 port map( D => n2549, CK => CLK, Q => OUT2(11), QN
                           => n4703);
   OUT2_reg_10_inst : DFF_X1 port map( D => n2548, CK => CLK, Q => OUT2(10), QN
                           => n4702);
   OUT2_reg_9_inst : DFF_X1 port map( D => n2547, CK => CLK, Q => OUT2(9), QN 
                           => n4701);
   OUT2_reg_8_inst : DFF_X1 port map( D => n2546, CK => CLK, Q => OUT2(8), QN 
                           => n4700);
   OUT2_reg_7_inst : DFF_X1 port map( D => n2545, CK => CLK, Q => OUT2(7), QN 
                           => n4699);
   OUT2_reg_6_inst : DFF_X1 port map( D => n2544, CK => CLK, Q => OUT2(6), QN 
                           => n4698);
   OUT2_reg_5_inst : DFF_X1 port map( D => n2543, CK => CLK, Q => OUT2(5), QN 
                           => n4697);
   OUT2_reg_4_inst : DFF_X1 port map( D => n2542, CK => CLK, Q => OUT2(4), QN 
                           => n4696);
   OUT2_reg_3_inst : DFF_X1 port map( D => n2541, CK => CLK, Q => OUT2(3), QN 
                           => n4695);
   OUT2_reg_2_inst : DFF_X1 port map( D => n2540, CK => CLK, Q => OUT2(2), QN 
                           => n4694);
   OUT2_reg_1_inst : DFF_X1 port map( D => n2539, CK => CLK, Q => OUT2(1), QN 
                           => n4693);
   OUT2_reg_0_inst : DFF_X1 port map( D => n2538, CK => CLK, Q => OUT2(0), QN 
                           => n4692);
   OUT1_reg_31_inst : DFF_X1 port map( D => n2537, CK => CLK, Q => OUT1(31), QN
                           => n4691);
   OUT1_reg_30_inst : DFF_X1 port map( D => n2536, CK => CLK, Q => OUT1(30), QN
                           => n4690);
   OUT1_reg_29_inst : DFF_X1 port map( D => n2535, CK => CLK, Q => OUT1(29), QN
                           => n4689);
   OUT1_reg_28_inst : DFF_X1 port map( D => n2534, CK => CLK, Q => OUT1(28), QN
                           => n4688);
   OUT1_reg_27_inst : DFF_X1 port map( D => n2533, CK => CLK, Q => OUT1(27), QN
                           => n4687);
   OUT1_reg_26_inst : DFF_X1 port map( D => n2532, CK => CLK, Q => OUT1(26), QN
                           => n4686);
   OUT1_reg_25_inst : DFF_X1 port map( D => n2531, CK => CLK, Q => OUT1(25), QN
                           => n4685);
   OUT1_reg_24_inst : DFF_X1 port map( D => n2530, CK => CLK, Q => OUT1(24), QN
                           => n4684);
   OUT1_reg_23_inst : DFF_X1 port map( D => n2529, CK => CLK, Q => OUT1(23), QN
                           => n4683);
   OUT1_reg_22_inst : DFF_X1 port map( D => n2528, CK => CLK, Q => OUT1(22), QN
                           => n4682);
   OUT1_reg_21_inst : DFF_X1 port map( D => n2527, CK => CLK, Q => OUT1(21), QN
                           => n4681);
   OUT1_reg_20_inst : DFF_X1 port map( D => n2526, CK => CLK, Q => OUT1(20), QN
                           => n4680);
   OUT1_reg_19_inst : DFF_X1 port map( D => n2525, CK => CLK, Q => OUT1(19), QN
                           => n4679);
   OUT1_reg_18_inst : DFF_X1 port map( D => n2524, CK => CLK, Q => OUT1(18), QN
                           => n4678);
   OUT1_reg_17_inst : DFF_X1 port map( D => n2523, CK => CLK, Q => OUT1(17), QN
                           => n4677);
   OUT1_reg_16_inst : DFF_X1 port map( D => n2522, CK => CLK, Q => OUT1(16), QN
                           => n4676);
   OUT1_reg_15_inst : DFF_X1 port map( D => n2521, CK => CLK, Q => OUT1(15), QN
                           => n4675);
   OUT1_reg_14_inst : DFF_X1 port map( D => n2520, CK => CLK, Q => OUT1(14), QN
                           => n4674);
   OUT1_reg_13_inst : DFF_X1 port map( D => n2519, CK => CLK, Q => OUT1(13), QN
                           => n4673);
   OUT1_reg_12_inst : DFF_X1 port map( D => n2518, CK => CLK, Q => OUT1(12), QN
                           => n4672);
   OUT1_reg_11_inst : DFF_X1 port map( D => n2517, CK => CLK, Q => OUT1(11), QN
                           => n4671);
   OUT1_reg_10_inst : DFF_X1 port map( D => n2516, CK => CLK, Q => OUT1(10), QN
                           => n4670);
   OUT1_reg_9_inst : DFF_X1 port map( D => n2515, CK => CLK, Q => OUT1(9), QN 
                           => n4669);
   OUT1_reg_8_inst : DFF_X1 port map( D => n2514, CK => CLK, Q => OUT1(8), QN 
                           => n4668);
   OUT1_reg_7_inst : DFF_X1 port map( D => n2513, CK => CLK, Q => OUT1(7), QN 
                           => n4667);
   OUT1_reg_6_inst : DFF_X1 port map( D => n2512, CK => CLK, Q => OUT1(6), QN 
                           => n4666);
   OUT1_reg_5_inst : DFF_X1 port map( D => n2511, CK => CLK, Q => OUT1(5), QN 
                           => n4665);
   OUT1_reg_4_inst : DFF_X1 port map( D => n2510, CK => CLK, Q => OUT1(4), QN 
                           => n4664);
   OUT1_reg_3_inst : DFF_X1 port map( D => n2509, CK => CLK, Q => OUT1(3), QN 
                           => n4663);
   OUT1_reg_2_inst : DFF_X1 port map( D => n2508, CK => CLK, Q => OUT1(2), QN 
                           => n4662);
   OUT1_reg_0_inst : DFF_X1 port map( D => n2506, CK => CLK, Q => OUT1(0), QN 
                           => n4660);
   REGISTERS_reg_8_21_inst : DFFR_X1 port map( D => n3327, CK => CLK, RN => 
                           n1475, Q => n_1499, QN => n239);
   REGISTERS_reg_5_31_inst : DFFR_X1 port map( D => n3433, CK => CLK, RN => 
                           n1466, Q => n4192, QN => n133);
   REGISTERS_reg_5_30_inst : DFFR_X1 port map( D => n3432, CK => CLK, RN => 
                           n1466, Q => n4193, QN => n134);
   REGISTERS_reg_5_29_inst : DFFR_X1 port map( D => n3431, CK => CLK, RN => 
                           n1466, Q => n4194, QN => n135);
   REGISTERS_reg_5_28_inst : DFFR_X1 port map( D => n3430, CK => CLK, RN => 
                           n1466, Q => n4195, QN => n136);
   REGISTERS_reg_5_27_inst : DFFR_X1 port map( D => n3429, CK => CLK, RN => 
                           n1467, Q => n4196, QN => n137);
   REGISTERS_reg_5_26_inst : DFFR_X1 port map( D => n3428, CK => CLK, RN => 
                           n1467, Q => n4197, QN => n138);
   REGISTERS_reg_5_25_inst : DFFR_X1 port map( D => n3427, CK => CLK, RN => 
                           n1467, Q => n4198, QN => n139);
   REGISTERS_reg_5_24_inst : DFFR_X1 port map( D => n3426, CK => CLK, RN => 
                           n1467, Q => n4199, QN => n140);
   REGISTERS_reg_4_31_inst : DFFR_X1 port map( D => n3465, CK => CLK, RN => 
                           n1464, Q => n4160, QN => n101);
   REGISTERS_reg_4_30_inst : DFFR_X1 port map( D => n3464, CK => CLK, RN => 
                           n1464, Q => n4161, QN => n102);
   REGISTERS_reg_4_29_inst : DFFR_X1 port map( D => n3463, CK => CLK, RN => 
                           n1464, Q => n4162, QN => n103);
   REGISTERS_reg_4_28_inst : DFFR_X1 port map( D => n3462, CK => CLK, RN => 
                           n1464, Q => n4163, QN => n104);
   REGISTERS_reg_4_27_inst : DFFR_X1 port map( D => n3461, CK => CLK, RN => 
                           n1464, Q => n4164, QN => n105);
   REGISTERS_reg_4_26_inst : DFFR_X1 port map( D => n3460, CK => CLK, RN => 
                           n1464, Q => n4165, QN => n106);
   REGISTERS_reg_4_25_inst : DFFR_X1 port map( D => n3459, CK => CLK, RN => 
                           n1464, Q => n4166, QN => n107);
   REGISTERS_reg_4_24_inst : DFFR_X1 port map( D => n3458, CK => CLK, RN => 
                           n1464, Q => n4167, QN => n108);
   REGISTERS_reg_1_31_inst : DFFR_X1 port map( D => n3561, CK => CLK, RN => 
                           n1456, Q => n4128, QN => n_1500);
   REGISTERS_reg_1_30_inst : DFFR_X1 port map( D => n3560, CK => CLK, RN => 
                           n1456, Q => n4129, QN => n_1501);
   REGISTERS_reg_1_29_inst : DFFR_X1 port map( D => n3559, CK => CLK, RN => 
                           n1456, Q => n4130, QN => n_1502);
   REGISTERS_reg_1_28_inst : DFFR_X1 port map( D => n3558, CK => CLK, RN => 
                           n1456, Q => n4131, QN => n_1503);
   REGISTERS_reg_1_27_inst : DFFR_X1 port map( D => n3557, CK => CLK, RN => 
                           n1456, Q => n4132, QN => n_1504);
   REGISTERS_reg_1_26_inst : DFFR_X1 port map( D => n3556, CK => CLK, RN => 
                           n1456, Q => n4133, QN => n_1505);
   REGISTERS_reg_1_25_inst : DFFR_X1 port map( D => n3555, CK => CLK, RN => 
                           n1456, Q => n4134, QN => n_1506);
   REGISTERS_reg_1_24_inst : DFFR_X1 port map( D => n3554, CK => CLK, RN => 
                           n1456, Q => n4135, QN => n_1507);
   REGISTERS_reg_21_31_inst : DFFR_X1 port map( D => n2921, CK => CLK, RN => 
                           n1509, Q => n4256, QN => n_1508);
   REGISTERS_reg_21_30_inst : DFFR_X1 port map( D => n2920, CK => CLK, RN => 
                           n1509, Q => n4257, QN => n_1509);
   REGISTERS_reg_21_29_inst : DFFR_X1 port map( D => n2919, CK => CLK, RN => 
                           n1509, Q => n4258, QN => n_1510);
   REGISTERS_reg_21_28_inst : DFFR_X1 port map( D => n2918, CK => CLK, RN => 
                           n1509, Q => n4259, QN => n_1511);
   REGISTERS_reg_21_27_inst : DFFR_X1 port map( D => n2917, CK => CLK, RN => 
                           n1509, Q => n4260, QN => n_1512);
   REGISTERS_reg_21_26_inst : DFFR_X1 port map( D => n2916, CK => CLK, RN => 
                           n1509, Q => n4261, QN => n_1513);
   REGISTERS_reg_21_25_inst : DFFR_X1 port map( D => n2915, CK => CLK, RN => 
                           n1509, Q => n4262, QN => n_1514);
   REGISTERS_reg_21_24_inst : DFFR_X1 port map( D => n2914, CK => CLK, RN => 
                           n1509, Q => n4263, QN => n_1515);
   REGISTERS_reg_16_31_inst : DFFR_X1 port map( D => n3081, CK => CLK, RN => 
                           n1496, Q => n4224, QN => n_1516);
   REGISTERS_reg_16_30_inst : DFFR_X1 port map( D => n3080, CK => CLK, RN => 
                           n1496, Q => n4225, QN => n_1517);
   REGISTERS_reg_16_29_inst : DFFR_X1 port map( D => n3079, CK => CLK, RN => 
                           n1496, Q => n4226, QN => n_1518);
   REGISTERS_reg_16_28_inst : DFFR_X1 port map( D => n3078, CK => CLK, RN => 
                           n1496, Q => n4227, QN => n_1519);
   REGISTERS_reg_16_27_inst : DFFR_X1 port map( D => n3077, CK => CLK, RN => 
                           n1496, Q => n4228, QN => n_1520);
   REGISTERS_reg_16_26_inst : DFFR_X1 port map( D => n3076, CK => CLK, RN => 
                           n1496, Q => n4229, QN => n_1521);
   REGISTERS_reg_16_25_inst : DFFR_X1 port map( D => n3075, CK => CLK, RN => 
                           n1496, Q => n4230, QN => n_1522);
   REGISTERS_reg_16_24_inst : DFFR_X1 port map( D => n3074, CK => CLK, RN => 
                           n1496, Q => n4231, QN => n_1523);
   REGISTERS_reg_31_31_inst : DFFR_X1 port map( D => n2601, CK => CLK, RN => 
                           n1536, Q => n4308, QN => n_1524);
   REGISTERS_reg_31_30_inst : DFFR_X1 port map( D => n2600, CK => CLK, RN => 
                           n1536, Q => n4309, QN => n_1525);
   REGISTERS_reg_31_29_inst : DFFR_X1 port map( D => n2599, CK => CLK, RN => 
                           n1536, Q => n4310, QN => n_1526);
   REGISTERS_reg_31_28_inst : DFFR_X1 port map( D => n2598, CK => CLK, RN => 
                           n1536, Q => n4311, QN => n_1527);
   REGISTERS_reg_31_27_inst : DFFR_X1 port map( D => n2597, CK => CLK, RN => 
                           n1536, Q => n4312, QN => n_1528);
   REGISTERS_reg_31_26_inst : DFFR_X1 port map( D => n2596, CK => CLK, RN => 
                           n1536, Q => n4313, QN => n_1529);
   REGISTERS_reg_31_25_inst : DFFR_X1 port map( D => n2595, CK => CLK, RN => 
                           n1536, Q => n4314, QN => n_1530);
   REGISTERS_reg_31_24_inst : DFFR_X1 port map( D => n2594, CK => CLK, RN => 
                           n1536, Q => n4315, QN => n_1531);
   REGISTERS_reg_26_31_inst : DFFR_X1 port map( D => n2761, CK => CLK, RN => 
                           n1522, Q => n4288, QN => n805);
   REGISTERS_reg_26_30_inst : DFFR_X1 port map( D => n2760, CK => CLK, RN => 
                           n1522, Q => n4289, QN => n806);
   REGISTERS_reg_26_29_inst : DFFR_X1 port map( D => n2759, CK => CLK, RN => 
                           n1522, Q => n4290, QN => n807);
   REGISTERS_reg_26_28_inst : DFFR_X1 port map( D => n2758, CK => CLK, RN => 
                           n1522, Q => n4291, QN => n808);
   REGISTERS_reg_26_27_inst : DFFR_X1 port map( D => n2757, CK => CLK, RN => 
                           n1523, Q => n4292, QN => n809);
   REGISTERS_reg_26_26_inst : DFFR_X1 port map( D => n2756, CK => CLK, RN => 
                           n1523, Q => n4293, QN => n810);
   REGISTERS_reg_26_25_inst : DFFR_X1 port map( D => n2755, CK => CLK, RN => 
                           n1523, Q => n4294, QN => n811);
   REGISTERS_reg_26_24_inst : DFFR_X1 port map( D => n2754, CK => CLK, RN => 
                           n1523, Q => n4295, QN => n812);
   REGISTERS_reg_5_23_inst : DFFR_X1 port map( D => n3425, CK => CLK, RN => 
                           n1467, Q => n4200, QN => n141);
   REGISTERS_reg_5_22_inst : DFFR_X1 port map( D => n3424, CK => CLK, RN => 
                           n1467, Q => n4201, QN => n142);
   REGISTERS_reg_5_21_inst : DFFR_X1 port map( D => n3423, CK => CLK, RN => 
                           n1467, Q => n4202, QN => n143);
   REGISTERS_reg_5_20_inst : DFFR_X1 port map( D => n3422, CK => CLK, RN => 
                           n1467, Q => n4203, QN => n144);
   REGISTERS_reg_5_19_inst : DFFR_X1 port map( D => n3421, CK => CLK, RN => 
                           n1467, Q => n4204, QN => n145);
   REGISTERS_reg_5_18_inst : DFFR_X1 port map( D => n3420, CK => CLK, RN => 
                           n1467, Q => n4205, QN => n146);
   REGISTERS_reg_5_17_inst : DFFR_X1 port map( D => n3419, CK => CLK, RN => 
                           n1467, Q => n4206, QN => n147);
   REGISTERS_reg_5_16_inst : DFFR_X1 port map( D => n3418, CK => CLK, RN => 
                           n1467, Q => n4207, QN => n148);
   REGISTERS_reg_5_15_inst : DFFR_X1 port map( D => n3417, CK => CLK, RN => 
                           n1468, Q => n4208, QN => n149);
   REGISTERS_reg_5_14_inst : DFFR_X1 port map( D => n3416, CK => CLK, RN => 
                           n1468, Q => n4209, QN => n150);
   REGISTERS_reg_5_13_inst : DFFR_X1 port map( D => n3415, CK => CLK, RN => 
                           n1468, Q => n4210, QN => n151);
   REGISTERS_reg_5_12_inst : DFFR_X1 port map( D => n3414, CK => CLK, RN => 
                           n1468, Q => n4211, QN => n152);
   REGISTERS_reg_5_11_inst : DFFR_X1 port map( D => n3413, CK => CLK, RN => 
                           n1468, Q => n4212, QN => n153);
   REGISTERS_reg_5_10_inst : DFFR_X1 port map( D => n3412, CK => CLK, RN => 
                           n1468, Q => n4213, QN => n154);
   REGISTERS_reg_5_9_inst : DFFR_X1 port map( D => n3411, CK => CLK, RN => 
                           n1468, Q => n4214, QN => n155);
   REGISTERS_reg_5_8_inst : DFFR_X1 port map( D => n3410, CK => CLK, RN => 
                           n1468, Q => n4215, QN => n156);
   REGISTERS_reg_5_7_inst : DFFR_X1 port map( D => n3409, CK => CLK, RN => 
                           n1468, Q => n4216, QN => n157);
   REGISTERS_reg_5_6_inst : DFFR_X1 port map( D => n3408, CK => CLK, RN => 
                           n1468, Q => n4217, QN => n158);
   REGISTERS_reg_5_5_inst : DFFR_X1 port map( D => n3407, CK => CLK, RN => 
                           n1468, Q => n4218, QN => n159);
   REGISTERS_reg_5_4_inst : DFFR_X1 port map( D => n3406, CK => CLK, RN => 
                           n1468, Q => n4219, QN => n160);
   REGISTERS_reg_5_3_inst : DFFR_X1 port map( D => n3405, CK => CLK, RN => 
                           n1469, Q => n4220, QN => n161);
   REGISTERS_reg_5_2_inst : DFFR_X1 port map( D => n3404, CK => CLK, RN => 
                           n1469, Q => n4221, QN => n162);
   REGISTERS_reg_5_1_inst : DFFR_X1 port map( D => n3403, CK => CLK, RN => 
                           n1469, Q => n4222, QN => n163);
   REGISTERS_reg_5_0_inst : DFFR_X1 port map( D => n3402, CK => CLK, RN => 
                           n1469, Q => n4223, QN => n164);
   REGISTERS_reg_4_23_inst : DFFR_X1 port map( D => n3457, CK => CLK, RN => 
                           n1464, Q => n4168, QN => n109);
   REGISTERS_reg_4_22_inst : DFFR_X1 port map( D => n3456, CK => CLK, RN => 
                           n1464, Q => n4169, QN => n110);
   REGISTERS_reg_4_21_inst : DFFR_X1 port map( D => n3455, CK => CLK, RN => 
                           n1464, Q => n4170, QN => n111);
   REGISTERS_reg_4_20_inst : DFFR_X1 port map( D => n3454, CK => CLK, RN => 
                           n1464, Q => n4171, QN => n112);
   REGISTERS_reg_4_19_inst : DFFR_X1 port map( D => n3453, CK => CLK, RN => 
                           n1465, Q => n4172, QN => n113);
   REGISTERS_reg_4_18_inst : DFFR_X1 port map( D => n3452, CK => CLK, RN => 
                           n1465, Q => n4173, QN => n114);
   REGISTERS_reg_4_17_inst : DFFR_X1 port map( D => n3451, CK => CLK, RN => 
                           n1465, Q => n4174, QN => n115);
   REGISTERS_reg_4_16_inst : DFFR_X1 port map( D => n3450, CK => CLK, RN => 
                           n1465, Q => n4175, QN => n116);
   REGISTERS_reg_4_15_inst : DFFR_X1 port map( D => n3449, CK => CLK, RN => 
                           n1465, Q => n4176, QN => n117);
   REGISTERS_reg_4_14_inst : DFFR_X1 port map( D => n3448, CK => CLK, RN => 
                           n1465, Q => n4177, QN => n118);
   REGISTERS_reg_4_13_inst : DFFR_X1 port map( D => n3447, CK => CLK, RN => 
                           n1465, Q => n4178, QN => n119);
   REGISTERS_reg_4_12_inst : DFFR_X1 port map( D => n3446, CK => CLK, RN => 
                           n1465, Q => n4179, QN => n120);
   REGISTERS_reg_4_11_inst : DFFR_X1 port map( D => n3445, CK => CLK, RN => 
                           n1465, Q => n4180, QN => n121);
   REGISTERS_reg_4_10_inst : DFFR_X1 port map( D => n3444, CK => CLK, RN => 
                           n1465, Q => n4181, QN => n122);
   REGISTERS_reg_4_9_inst : DFFR_X1 port map( D => n3443, CK => CLK, RN => 
                           n1465, Q => n4182, QN => n123);
   REGISTERS_reg_4_8_inst : DFFR_X1 port map( D => n3442, CK => CLK, RN => 
                           n1465, Q => n4183, QN => n124);
   REGISTERS_reg_4_7_inst : DFFR_X1 port map( D => n3441, CK => CLK, RN => 
                           n1466, Q => n4184, QN => n125);
   REGISTERS_reg_4_6_inst : DFFR_X1 port map( D => n3440, CK => CLK, RN => 
                           n1466, Q => n4185, QN => n126);
   REGISTERS_reg_4_5_inst : DFFR_X1 port map( D => n3439, CK => CLK, RN => 
                           n1466, Q => n4186, QN => n127);
   REGISTERS_reg_4_4_inst : DFFR_X1 port map( D => n3438, CK => CLK, RN => 
                           n1466, Q => n4187, QN => n128);
   REGISTERS_reg_4_3_inst : DFFR_X1 port map( D => n3437, CK => CLK, RN => 
                           n1466, Q => n4188, QN => n129);
   REGISTERS_reg_4_2_inst : DFFR_X1 port map( D => n3436, CK => CLK, RN => 
                           n1466, Q => n4189, QN => n130);
   REGISTERS_reg_4_1_inst : DFFR_X1 port map( D => n3435, CK => CLK, RN => 
                           n1466, Q => n4190, QN => n131);
   REGISTERS_reg_4_0_inst : DFFR_X1 port map( D => n3434, CK => CLK, RN => 
                           n1466, Q => n4191, QN => n132);
   REGISTERS_reg_1_23_inst : DFFR_X1 port map( D => n3553, CK => CLK, RN => 
                           n1456, Q => n4136, QN => n_1532);
   REGISTERS_reg_1_22_inst : DFFR_X1 port map( D => n3552, CK => CLK, RN => 
                           n1456, Q => n4137, QN => n_1533);
   REGISTERS_reg_1_21_inst : DFFR_X1 port map( D => n3551, CK => CLK, RN => 
                           n1456, Q => n4138, QN => n_1534);
   REGISTERS_reg_1_20_inst : DFFR_X1 port map( D => n3550, CK => CLK, RN => 
                           n1456, Q => n4139, QN => n_1535);
   REGISTERS_reg_1_19_inst : DFFR_X1 port map( D => n3549, CK => CLK, RN => 
                           n1457, Q => n4140, QN => n_1536);
   REGISTERS_reg_1_18_inst : DFFR_X1 port map( D => n3548, CK => CLK, RN => 
                           n1457, Q => n4141, QN => n_1537);
   REGISTERS_reg_1_17_inst : DFFR_X1 port map( D => n3547, CK => CLK, RN => 
                           n1457, Q => n4142, QN => n_1538);
   REGISTERS_reg_1_16_inst : DFFR_X1 port map( D => n3546, CK => CLK, RN => 
                           n1457, Q => n4143, QN => n_1539);
   REGISTERS_reg_1_15_inst : DFFR_X1 port map( D => n3545, CK => CLK, RN => 
                           n1457, Q => n4144, QN => n_1540);
   REGISTERS_reg_1_14_inst : DFFR_X1 port map( D => n3544, CK => CLK, RN => 
                           n1457, Q => n4145, QN => n_1541);
   REGISTERS_reg_1_13_inst : DFFR_X1 port map( D => n3543, CK => CLK, RN => 
                           n1457, Q => n4146, QN => n_1542);
   REGISTERS_reg_1_12_inst : DFFR_X1 port map( D => n3542, CK => CLK, RN => 
                           n1457, Q => n4147, QN => n_1543);
   REGISTERS_reg_1_11_inst : DFFR_X1 port map( D => n3541, CK => CLK, RN => 
                           n1457, Q => n4148, QN => n_1544);
   REGISTERS_reg_1_10_inst : DFFR_X1 port map( D => n3540, CK => CLK, RN => 
                           n1457, Q => n4149, QN => n_1545);
   REGISTERS_reg_1_9_inst : DFFR_X1 port map( D => n3539, CK => CLK, RN => 
                           n1457, Q => n4150, QN => n_1546);
   REGISTERS_reg_1_8_inst : DFFR_X1 port map( D => n3538, CK => CLK, RN => 
                           n1457, Q => n4151, QN => n_1547);
   REGISTERS_reg_1_7_inst : DFFR_X1 port map( D => n3537, CK => CLK, RN => 
                           n1458, Q => n4152, QN => n_1548);
   REGISTERS_reg_1_6_inst : DFFR_X1 port map( D => n3536, CK => CLK, RN => 
                           n1458, Q => n4153, QN => n_1549);
   REGISTERS_reg_1_5_inst : DFFR_X1 port map( D => n3535, CK => CLK, RN => 
                           n1458, Q => n4154, QN => n_1550);
   REGISTERS_reg_1_4_inst : DFFR_X1 port map( D => n3534, CK => CLK, RN => 
                           n1458, Q => n4155, QN => n_1551);
   REGISTERS_reg_1_3_inst : DFFR_X1 port map( D => n3533, CK => CLK, RN => 
                           n1458, Q => n4156, QN => n_1552);
   REGISTERS_reg_1_2_inst : DFFR_X1 port map( D => n3532, CK => CLK, RN => 
                           n1458, Q => n4157, QN => n_1553);
   REGISTERS_reg_1_1_inst : DFFR_X1 port map( D => n3531, CK => CLK, RN => 
                           n1458, Q => n4158, QN => n_1554);
   REGISTERS_reg_1_0_inst : DFFR_X1 port map( D => n3530, CK => CLK, RN => 
                           n1458, Q => n4159, QN => n_1555);
   REGISTERS_reg_13_31_inst : DFFR_X1 port map( D => n3177, CK => CLK, RN => 
                           n1488, Q => n2206, QN => n389);
   REGISTERS_reg_13_30_inst : DFFR_X1 port map( D => n3176, CK => CLK, RN => 
                           n1488, Q => n2181, QN => n390);
   REGISTERS_reg_13_29_inst : DFFR_X1 port map( D => n3175, CK => CLK, RN => 
                           n1488, Q => n2160, QN => n391);
   REGISTERS_reg_13_28_inst : DFFR_X1 port map( D => n3174, CK => CLK, RN => 
                           n1488, Q => n2139, QN => n392);
   REGISTERS_reg_13_27_inst : DFFR_X1 port map( D => n3173, CK => CLK, RN => 
                           n1488, Q => n2118, QN => n393);
   REGISTERS_reg_13_26_inst : DFFR_X1 port map( D => n3172, CK => CLK, RN => 
                           n1488, Q => n2097, QN => n394);
   REGISTERS_reg_13_25_inst : DFFR_X1 port map( D => n3171, CK => CLK, RN => 
                           n1488, Q => n2076, QN => n395);
   REGISTERS_reg_13_24_inst : DFFR_X1 port map( D => n3170, CK => CLK, RN => 
                           n1488, Q => n2055, QN => n396);
   REGISTERS_reg_12_31_inst : DFFR_X1 port map( D => n3209, CK => CLK, RN => 
                           n1485, Q => n2210, QN => n357);
   REGISTERS_reg_12_30_inst : DFFR_X1 port map( D => n3208, CK => CLK, RN => 
                           n1485, Q => n2183, QN => n358);
   REGISTERS_reg_12_29_inst : DFFR_X1 port map( D => n3207, CK => CLK, RN => 
                           n1485, Q => n2162, QN => n359);
   REGISTERS_reg_12_28_inst : DFFR_X1 port map( D => n3206, CK => CLK, RN => 
                           n1485, Q => n2141, QN => n360);
   REGISTERS_reg_12_27_inst : DFFR_X1 port map( D => n3205, CK => CLK, RN => 
                           n1485, Q => n2120, QN => n361);
   REGISTERS_reg_12_26_inst : DFFR_X1 port map( D => n3204, CK => CLK, RN => 
                           n1485, Q => n2099, QN => n362);
   REGISTERS_reg_12_25_inst : DFFR_X1 port map( D => n3203, CK => CLK, RN => 
                           n1485, Q => n2078, QN => n363);
   REGISTERS_reg_12_24_inst : DFFR_X1 port map( D => n3202, CK => CLK, RN => 
                           n1485, Q => n2057, QN => n364);
   REGISTERS_reg_20_31_inst : DFFR_X1 port map( D => n2953, CK => CLK, RN => 
                           n1506, Q => n_1556, QN => n613);
   REGISTERS_reg_20_30_inst : DFFR_X1 port map( D => n2952, CK => CLK, RN => 
                           n1506, Q => n_1557, QN => n614);
   REGISTERS_reg_20_29_inst : DFFR_X1 port map( D => n2951, CK => CLK, RN => 
                           n1506, Q => n_1558, QN => n615);
   REGISTERS_reg_20_28_inst : DFFR_X1 port map( D => n2950, CK => CLK, RN => 
                           n1506, Q => n_1559, QN => n616);
   REGISTERS_reg_20_27_inst : DFFR_X1 port map( D => n2949, CK => CLK, RN => 
                           n1507, Q => n_1560, QN => n617);
   REGISTERS_reg_20_26_inst : DFFR_X1 port map( D => n2948, CK => CLK, RN => 
                           n1507, Q => n_1561, QN => n618);
   REGISTERS_reg_20_25_inst : DFFR_X1 port map( D => n2947, CK => CLK, RN => 
                           n1507, Q => n_1562, QN => n619);
   REGISTERS_reg_20_24_inst : DFFR_X1 port map( D => n2946, CK => CLK, RN => 
                           n1507, Q => n_1563, QN => n620);
   REGISTERS_reg_9_31_inst : DFFR_X1 port map( D => n3305, CK => CLK, RN => 
                           n1477, Q => n4085, QN => n261);
   REGISTERS_reg_9_30_inst : DFFR_X1 port map( D => n3304, CK => CLK, RN => 
                           n1477, Q => n4059, QN => n262);
   REGISTERS_reg_9_29_inst : DFFR_X1 port map( D => n3303, CK => CLK, RN => 
                           n1477, Q => n4033, QN => n263);
   REGISTERS_reg_9_28_inst : DFFR_X1 port map( D => n3302, CK => CLK, RN => 
                           n1477, Q => n4007, QN => n264);
   REGISTERS_reg_9_27_inst : DFFR_X1 port map( D => n3301, CK => CLK, RN => 
                           n1477, Q => n3981, QN => n265);
   REGISTERS_reg_9_26_inst : DFFR_X1 port map( D => n3300, CK => CLK, RN => 
                           n1477, Q => n3955, QN => n266);
   REGISTERS_reg_9_25_inst : DFFR_X1 port map( D => n3299, CK => CLK, RN => 
                           n1477, Q => n3929, QN => n267);
   REGISTERS_reg_9_24_inst : DFFR_X1 port map( D => n3298, CK => CLK, RN => 
                           n1477, Q => n3903, QN => n268);
   REGISTERS_reg_17_31_inst : DFFR_X1 port map( D => n3049, CK => CLK, RN => 
                           n1498, Q => n4123, QN => n517);
   REGISTERS_reg_17_30_inst : DFFR_X1 port map( D => n3048, CK => CLK, RN => 
                           n1498, Q => n4080, QN => n518);
   REGISTERS_reg_17_29_inst : DFFR_X1 port map( D => n3047, CK => CLK, RN => 
                           n1498, Q => n4054, QN => n519);
   REGISTERS_reg_17_28_inst : DFFR_X1 port map( D => n3046, CK => CLK, RN => 
                           n1498, Q => n4028, QN => n520);
   REGISTERS_reg_17_27_inst : DFFR_X1 port map( D => n3045, CK => CLK, RN => 
                           n1499, Q => n4002, QN => n521);
   REGISTERS_reg_17_26_inst : DFFR_X1 port map( D => n3044, CK => CLK, RN => 
                           n1499, Q => n3976, QN => n522);
   REGISTERS_reg_17_25_inst : DFFR_X1 port map( D => n3043, CK => CLK, RN => 
                           n1499, Q => n3950, QN => n523);
   REGISTERS_reg_17_24_inst : DFFR_X1 port map( D => n3042, CK => CLK, RN => 
                           n1499, Q => n3924, QN => n524);
   REGISTERS_reg_8_31_inst : DFFR_X1 port map( D => n3337, CK => CLK, RN => 
                           n1474, Q => n_1564, QN => n229);
   REGISTERS_reg_8_30_inst : DFFR_X1 port map( D => n3336, CK => CLK, RN => 
                           n1474, Q => n_1565, QN => n230);
   REGISTERS_reg_8_29_inst : DFFR_X1 port map( D => n3335, CK => CLK, RN => 
                           n1474, Q => n_1566, QN => n231);
   REGISTERS_reg_8_28_inst : DFFR_X1 port map( D => n3334, CK => CLK, RN => 
                           n1474, Q => n_1567, QN => n232);
   REGISTERS_reg_8_27_inst : DFFR_X1 port map( D => n3333, CK => CLK, RN => 
                           n1475, Q => n_1568, QN => n233);
   REGISTERS_reg_8_26_inst : DFFR_X1 port map( D => n3332, CK => CLK, RN => 
                           n1475, Q => n_1569, QN => n234);
   REGISTERS_reg_8_25_inst : DFFR_X1 port map( D => n3331, CK => CLK, RN => 
                           n1475, Q => n_1570, QN => n235);
   REGISTERS_reg_8_24_inst : DFFR_X1 port map( D => n3330, CK => CLK, RN => 
                           n1475, Q => n_1571, QN => n236);
   REGISTERS_reg_30_31_inst : DFFR_X1 port map( D => n2633, CK => CLK, RN => 
                           n1533, Q => n_1572, QN => n933);
   REGISTERS_reg_30_30_inst : DFFR_X1 port map( D => n2632, CK => CLK, RN => 
                           n1533, Q => n_1573, QN => n934);
   REGISTERS_reg_30_29_inst : DFFR_X1 port map( D => n2631, CK => CLK, RN => 
                           n1533, Q => n_1574, QN => n935);
   REGISTERS_reg_30_28_inst : DFFR_X1 port map( D => n2630, CK => CLK, RN => 
                           n1533, Q => n_1575, QN => n936);
   REGISTERS_reg_30_27_inst : DFFR_X1 port map( D => n2629, CK => CLK, RN => 
                           n1533, Q => n_1576, QN => n937);
   REGISTERS_reg_30_26_inst : DFFR_X1 port map( D => n2628, CK => CLK, RN => 
                           n1533, Q => n_1577, QN => n938);
   REGISTERS_reg_30_25_inst : DFFR_X1 port map( D => n2627, CK => CLK, RN => 
                           n1533, Q => n_1578, QN => n939);
   REGISTERS_reg_30_24_inst : DFFR_X1 port map( D => n2626, CK => CLK, RN => 
                           n1533, Q => n_1579, QN => n940);
   REGISTERS_reg_27_31_inst : DFFR_X1 port map( D => n2729, CK => CLK, RN => 
                           n1525, Q => n4110, QN => n837);
   REGISTERS_reg_27_30_inst : DFFR_X1 port map( D => n2728, CK => CLK, RN => 
                           n1525, Q => n4073, QN => n838);
   REGISTERS_reg_27_29_inst : DFFR_X1 port map( D => n2727, CK => CLK, RN => 
                           n1525, Q => n4047, QN => n839);
   REGISTERS_reg_27_28_inst : DFFR_X1 port map( D => n2726, CK => CLK, RN => 
                           n1525, Q => n4021, QN => n840);
   REGISTERS_reg_27_27_inst : DFFR_X1 port map( D => n2725, CK => CLK, RN => 
                           n1525, Q => n3995, QN => n841);
   REGISTERS_reg_27_26_inst : DFFR_X1 port map( D => n2724, CK => CLK, RN => 
                           n1525, Q => n3969, QN => n842);
   REGISTERS_reg_27_25_inst : DFFR_X1 port map( D => n2723, CK => CLK, RN => 
                           n1525, Q => n3943, QN => n843);
   REGISTERS_reg_27_24_inst : DFFR_X1 port map( D => n2722, CK => CLK, RN => 
                           n1525, Q => n3917, QN => n844);
   REGISTERS_reg_8_6_inst : DFFR_X2 port map( D => n3312, CK => CLK, RN => 
                           n1476, Q => n_1580, QN => n254);
   OUT1_reg_1_inst : DFF_X2 port map( D => n2507, CK => CLK, Q => OUT1(1), QN 
                           => n4661);
   U2 : AND2_X1 port map( A1 => n1030, A2 => n973, ZN => n1);
   U3 : AND2_X1 port map( A1 => n1030, A2 => n973, ZN => n2);
   U4 : AND2_X2 port map( A1 => n1030, A2 => n973, ZN => n932);
   U5 : AND3_X1 port map( A1 => ADD_RS1(0), A2 => n706, A3 => n1560, ZN => 
                           n1028);
   U6 : AND2_X1 port map( A1 => n1182, A2 => n4256, ZN => n3);
   U7 : AND2_X1 port map( A1 => n1179, A2 => n4224, ZN => n4);
   U8 : NOR3_X1 port map( A1 => n3, A2 => n4, A3 => n2231, ZN => n2235);
   U9 : CLKBUF_X1 port map( A => n4656, Z => n5);
   U10 : BUF_X2 port map( A => n990, Z => n1182);
   U11 : BUF_X2 port map( A => n992, Z => n1179);
   U12 : BUF_X2 port map( A => n4088, Z => n1205);
   U13 : CLKBUF_X3 port map( A => n2225, Z => n1159);
   U14 : CLKBUF_X3 port map( A => n4091, Z => n6);
   U15 : BUF_X1 port map( A => n4091, Z => n1214);
   U16 : CLKBUF_X1 port map( A => n1036, Z => n7);
   U17 : CLKBUF_X3 port map( A => n4090, Z => n8);
   U18 : BUF_X1 port map( A => n4090, Z => n1211);
   U19 : CLKBUF_X3 port map( A => n4099, Z => n1230);
   U20 : BUF_X1 port map( A => n166, Z => n55);
   U21 : BUF_X1 port map( A => n968, Z => n9);
   U22 : BUF_X1 port map( A => n968, Z => n1198);
   U23 : AND2_X2 port map( A1 => n1554, A2 => n784, ZN => n705);
   U24 : OR2_X1 port map( A1 => n1071, A2 => n1072, ZN => n10);
   U25 : OR2_X1 port map( A1 => n1069, A2 => n1070, ZN => n11);
   U26 : OR2_X1 port map( A1 => n686, A2 => n687, ZN => n12);
   U27 : OR2_X1 port map( A1 => n602, A2 => n603, ZN => n13);
   U28 : OR2_X1 port map( A1 => n907, A2 => n906, ZN => n14);
   U29 : OR2_X1 port map( A1 => n919, A2 => n918, ZN => n15);
   U30 : OR2_X1 port map( A1 => n1042, A2 => n1041, ZN => n16);
   U31 : OR2_X1 port map( A1 => n1038, A2 => n1037, ZN => n17);
   U32 : OR2_X1 port map( A1 => n910, A2 => n911, ZN => n18);
   U33 : OR2_X1 port map( A1 => n1065, A2 => n1066, ZN => n19);
   U34 : OR2_X1 port map( A1 => n1057, A2 => n1058, ZN => n20);
   U35 : OR2_X1 port map( A1 => n765, A2 => n766, ZN => n21);
   U36 : OR2_X1 port map( A1 => n779, A2 => n780, ZN => n22);
   U37 : OR2_X1 port map( A1 => n1051, A2 => n1052, ZN => n23);
   U38 : OR2_X1 port map( A1 => n900, A2 => n901, ZN => n24);
   U39 : OR2_X1 port map( A1 => n904, A2 => n905, ZN => n25);
   U40 : OR2_X1 port map( A1 => n898, A2 => n899, ZN => n26);
   U41 : OR2_X1 port map( A1 => n777, A2 => n778, ZN => n27);
   U42 : OR2_X1 port map( A1 => n767, A2 => n768, ZN => n28);
   U43 : OR2_X1 port map( A1 => n1059, A2 => n1060, ZN => n29);
   U44 : OR2_X1 port map( A1 => n902, A2 => n903, ZN => n30);
   U45 : OR2_X1 port map( A1 => n1049, A2 => n1050, ZN => n31);
   U46 : OR2_X1 port map( A1 => n894, A2 => n895, ZN => n32);
   U47 : BUF_X1 port map( A => n2209, Z => n507);
   U48 : NOR2_X1 port map( A1 => n2149, A2 => n21, ZN => n2156);
   U49 : NOR2_X1 port map( A1 => n2128, A2 => n31, ZN => n2135);
   U50 : NOR2_X1 port map( A1 => n2107, A2 => n28, ZN => n2114);
   U51 : NOR2_X1 port map( A1 => n1778, A2 => n26, ZN => n1785);
   U52 : NOR2_X1 port map( A1 => n1757, A2 => n30, ZN => n1764);
   U53 : BUF_X2 port map( A => n977, Z => n33);
   U54 : CLKBUF_X3 port map( A => n4118, Z => n1261);
   U55 : OR2_X1 port map( A1 => n385, A2 => n1214, ZN => n34);
   U56 : OR2_X1 port map( A1 => n417, A2 => n1211, ZN => n35);
   U57 : NAND3_X1 port map( A1 => n34, A2 => n35, A3 => n2323, ZN => n2330);
   U58 : AND2_X1 port map( A1 => n1181, A2 => n4274, ZN => n36);
   U59 : AND2_X1 port map( A1 => n1178, A2 => n4242, ZN => n37);
   U60 : NOR3_X1 port map( A1 => n36, A2 => n37, A3 => n1842, ZN => n1845);
   U61 : BUF_X2 port map( A => n967, Z => n1201);
   U62 : AND2_X1 port map( A1 => n4797, A2 => n1253, ZN => n38);
   U63 : AND2_X1 port map( A1 => n1250, A2 => n4330, ZN => n39);
   U64 : NOR3_X1 port map( A1 => n38, A2 => n39, A3 => n2487, ZN => n2495);
   U65 : AND2_X1 port map( A1 => ADD_RS1(2), A2 => n1553, ZN => n887);
   U66 : CLKBUF_X3 port map( A => n1003, Z => n1186);
   U67 : CLKBUF_X3 port map( A => n1003, Z => n1187);
   U68 : NOR2_X1 port map( A1 => n1694, A2 => n19, ZN => n1701);
   U69 : AND2_X2 port map( A1 => n973, A2 => n695, ZN => n40);
   U70 : CLKBUF_X3 port map( A => n4088, Z => n1207);
   U71 : OR2_X1 port map( A1 => n1230, A2 => n186, ZN => n41);
   U72 : OR2_X1 port map( A1 => n1227, A2 => n335, ZN => n42);
   U73 : NAND3_X1 port map( A1 => n41, A2 => n42, A3 => n3909, ZN => n3910);
   U74 : OR2_X1 port map( A1 => n1228, A2 => n178, ZN => n43);
   U75 : OR2_X1 port map( A1 => n1225, A2 => n327, ZN => n44);
   U76 : NAND3_X1 port map( A1 => n43, A2 => n44, A3 => n2452, ZN => n2453);
   U77 : OR2_X1 port map( A1 => n1229, A2 => n175, ZN => n45);
   U78 : OR2_X1 port map( A1 => n1225, A2 => n324, ZN => n46);
   U79 : NAND3_X1 port map( A1 => n45, A2 => n46, A3 => n2377, ZN => n2378);
   U80 : OR2_X1 port map( A1 => n1228, A2 => n185, ZN => n47);
   U81 : OR2_X1 port map( A1 => n1226, A2 => n334, ZN => n48);
   U82 : NAND3_X1 port map( A1 => n47, A2 => n48, A3 => n3883, ZN => n3884);
   U83 : BUF_X1 port map( A => ADD_RS1(3), Z => n1054);
   U84 : NOR2_X1 port map( A1 => n4020, A2 => n12, ZN => n4032);
   U85 : BUF_X1 port map( A => ADD_RS2(4), Z => n889);
   U86 : NOR2_X1 port map( A1 => n3765, A2 => n15, ZN => n3777);
   U87 : OR2_X1 port map( A1 => n1936, A2 => n1140, ZN => n49);
   U88 : OR2_X1 port map( A1 => n114, A2 => n1137, ZN => n50);
   U89 : NAND3_X1 port map( A1 => n49, A2 => n50, A3 => n1935, ZN => n1937);
   U90 : BUF_X1 port map( A => n494, Z => n51);
   U91 : BUF_X1 port map( A => n494, Z => n1121);
   U92 : BUF_X1 port map( A => n970, Z => n52);
   U93 : BUF_X1 port map( A => n970, Z => n1120);
   U94 : BUF_X2 port map( A => n970, Z => n508);
   U95 : BUF_X2 port map( A => n482, Z => n1016);
   U96 : NOR2_X1 port map( A1 => n53, A2 => n2238, ZN => n1000);
   U97 : OR3_X1 port map( A1 => ADD_RS2(4), A2 => ADD_RS2(3), A3 => ADD_RS2(0),
                           ZN => n53);
   U98 : CLKBUF_X1 port map( A => n1028, Z => n1015);
   U99 : BUF_X2 port map( A => n166, Z => n54);
   U100 : BUF_X2 port map( A => n965, Z => n56);
   U101 : BUF_X2 port map( A => n965, Z => n57);
   U102 : AND2_X1 port map( A1 => n1077, A2 => n705, ZN => n166);
   U103 : NOR2_X1 port map( A1 => n3640, A2 => n16, ZN => n3652);
   U104 : OR2_X1 port map( A1 => n1874, A2 => n1140, ZN => n58);
   U105 : OR2_X1 port map( A1 => n117, A2 => n1137, ZN => n59);
   U106 : NAND3_X1 port map( A1 => n58, A2 => n59, A3 => n1873, ZN => n1875);
   U107 : OR2_X1 port map( A1 => n3959, A2 => n1127, ZN => n60);
   U108 : OR2_X1 port map( A1 => n266, A2 => n678, ZN => n61);
   U109 : NAND3_X1 port map( A1 => n60, A2 => n61, A3 => n2096, ZN => n2104);
   U110 : BUF_X2 port map( A => n494, Z => n512);
   U111 : OR2_X1 port map( A1 => n3681, A2 => n1128, ZN => n62);
   U112 : OR2_X1 port map( A1 => n277, A2 => n1126, ZN => n63);
   U113 : NAND3_X1 port map( A1 => n1871, A2 => n63, A3 => n62, ZN => n1877);
   U114 : OR2_X1 port map( A1 => n1997, A2 => n1140, ZN => n64);
   U115 : OR2_X1 port map( A1 => n111, A2 => n1137, ZN => n65);
   U116 : NAND3_X1 port map( A1 => n64, A2 => n65, A3 => n1996, ZN => n1998);
   U117 : NOR2_X1 port map( A1 => n2086, A2 => n23, ZN => n2093);
   U118 : BUF_X2 port map( A => n967, Z => n66);
   U119 : AND2_X2 port map( A1 => n974, A2 => n2265, ZN => n967);
   U120 : NOR2_X1 port map( A1 => n2434, A2 => n11, ZN => n2446);
   U121 : NOR2_X1 port map( A1 => n1736, A2 => n20, ZN => n1743);
   U122 : OR2_X1 port map( A1 => n1730, A2 => n1139, ZN => n67);
   U123 : OR2_X1 port map( A1 => n124, A2 => n1136, ZN => n68);
   U124 : NAND3_X1 port map( A1 => n67, A2 => n68, A3 => n1729, ZN => n1731);
   U125 : NOR2_X1 port map( A1 => n1715, A2 => n29, ZN => n1722);
   U126 : OR2_X1 port map( A1 => n1709, A2 => n1139, ZN => n69);
   U127 : OR2_X1 port map( A1 => n125, A2 => n1136, ZN => n70);
   U128 : NAND3_X1 port map( A1 => n69, A2 => n70, A3 => n1708, ZN => n1710);
   U129 : NOR2_X1 port map( A1 => n1611, A2 => n27, ZN => n1618);
   U130 : OR2_X1 port map( A1 => n1605, A2 => n1139, ZN => n71);
   U131 : OR2_X1 port map( A1 => n130, A2 => n1136, ZN => n72);
   U132 : NAND3_X1 port map( A1 => n71, A2 => n72, A3 => n1604, ZN => n1606);
   U133 : NOR2_X1 port map( A1 => n2044, A2 => n24, ZN => n2051);
   U134 : OR2_X1 port map( A1 => n2038, A2 => n1140, ZN => n73);
   U135 : OR2_X1 port map( A1 => n109, A2 => n1137, ZN => n74);
   U136 : NAND3_X1 port map( A1 => n73, A2 => n74, A3 => n2037, ZN => n2039);
   U137 : NOR2_X1 port map( A1 => n2023, A2 => n25, ZN => n2030);
   U138 : OR2_X1 port map( A1 => n2017, A2 => n1140, ZN => n75);
   U139 : OR2_X1 port map( A1 => n110, A2 => n1137, ZN => n76);
   U140 : NAND3_X1 port map( A1 => n75, A2 => n76, A3 => n2016, ZN => n2018);
   U141 : NOR2_X1 port map( A1 => n1982, A2 => n18, ZN => n1989);
   U142 : NOR3_X1 port map( A1 => n4656, A2 => n4645, A3 => n4657, ZN => n77);
   U143 : NOR3_X1 port map( A1 => n4657, A2 => n4645, A3 => n5, ZN => n78);
   U144 : AND2_X1 port map( A1 => n1268, A2 => n4278, ZN => n79);
   U145 : AND2_X1 port map( A1 => n1265, A2 => n4246, ZN => n80);
   U146 : NOR3_X1 port map( A1 => n79, A2 => n80, A3 => n2490, ZN => n2494);
   U147 : OR2_X1 port map( A1 => n635, A2 => n1262, ZN => n81);
   U148 : OR2_X1 port map( A1 => n1259, A2 => n2489, ZN => n82);
   U149 : OR2_X1 port map( A1 => n590, A2 => n2488, ZN => n83);
   U150 : NAND3_X1 port map( A1 => n81, A2 => n82, A3 => n83, ZN => n2490);
   U151 : BUF_X2 port map( A => n986, Z => n1268);
   U152 : BUF_X2 port map( A => n985, Z => n1265);
   U153 : BUF_X1 port map( A => ADD_RS1(3), Z => n84);
   U154 : OR2_X1 port map( A1 => n376, A2 => n1213, ZN => n85);
   U155 : OR2_X1 port map( A1 => n408, A2 => n8, ZN => n86);
   U156 : NAND3_X1 port map( A1 => n85, A2 => n86, A3 => n3604, ZN => n3611);
   U157 : CLKBUF_X1 port map( A => n998, Z => n87);
   U158 : NOR2_X1 port map( A1 => n1861, A2 => n22, ZN => n1868);
   U159 : NOR2_X1 port map( A1 => n1799, A2 => n32, ZN => n1806);
   U160 : OR2_X1 port map( A1 => n1230, A2 => n187, ZN => n88);
   U161 : OR2_X1 port map( A1 => n1227, A2 => n336, ZN => n89);
   U162 : NAND3_X1 port map( A1 => n88, A2 => n89, A3 => n3935, ZN => n3936);
   U163 : BUF_X2 port map( A => n4098, Z => n1227);
   U164 : NOR2_X1 port map( A1 => n4046, A2 => n13, ZN => n4058);
   U165 : OR2_X1 port map( A1 => n1205, A2 => n319, ZN => n90);
   U166 : OR2_X1 port map( A1 => n231, A2 => n1204, ZN => n91);
   U167 : NAND3_X1 port map( A1 => n90, A2 => n91, A3 => n4034, ZN => n4043);
   U168 : BUF_X2 port map( A => n4087, Z => n1204);
   U169 : OR2_X1 port map( A1 => n1205, A2 => n308, ZN => n92);
   U170 : OR2_X1 port map( A1 => n242, A2 => n1203, ZN => n93);
   U171 : NAND3_X1 port map( A1 => n92, A2 => n93, A3 => n3753, ZN => n3762);
   U172 : OR2_X1 port map( A1 => n1205, A2 => n303, ZN => n94);
   U173 : OR2_X1 port map( A1 => n247, A2 => n1203, ZN => n95);
   U174 : NAND3_X1 port map( A1 => n94, A2 => n95, A3 => n3628, ZN => n3637);
   U175 : NOR2_X1 port map( A1 => n2409, A2 => n10, ZN => n2421);
   U176 : OR2_X1 port map( A1 => n1228, A2 => n176, ZN => n96);
   U177 : OR2_X1 port map( A1 => n1225, A2 => n325, ZN => n97);
   U178 : NAND3_X1 port map( A1 => n96, A2 => n97, A3 => n2402, ZN => n2403);
   U179 : NOR2_X1 port map( A1 => n3665, A2 => n17, ZN => n3677);
   U180 : OR2_X1 port map( A1 => n1230, A2 => n182, ZN => n98);
   U181 : OR2_X1 port map( A1 => n1226, A2 => n331, ZN => n99);
   U182 : NAND3_X1 port map( A1 => n98, A2 => n99, A3 => n3658, ZN => n3659);
   U183 : OR2_X1 port map( A1 => n1229, A2 => n184, ZN => n100);
   U184 : OR2_X1 port map( A1 => n1226, A2 => n333, ZN => n165);
   U185 : NAND3_X1 port map( A1 => n100, A2 => n165, A3 => n3758, ZN => n3759);
   U186 : AND2_X1 port map( A1 => n1077, A2 => n705, ZN => n965);
   U187 : NOR2_X1 port map( A1 => n3890, A2 => n14, ZN => n3902);
   U188 : OR2_X1 port map( A1 => n1205, A2 => n313, ZN => n167);
   U189 : OR2_X1 port map( A1 => n237, A2 => n1203, ZN => n168);
   U190 : NAND3_X1 port map( A1 => n167, A2 => n168, A3 => n3878, ZN => n3887);
   U191 : OR2_X1 port map( A1 => n1205, A2 => n297, ZN => n169);
   U192 : OR2_X1 port map( A1 => n254, A2 => n1202, ZN => n170);
   U193 : NAND3_X1 port map( A1 => n169, A2 => n170, A3 => n2397, ZN => n2406);
   U194 : CLKBUF_X3 port map( A => n4087, Z => n1202);
   U195 : BUF_X2 port map( A => n4111, Z => n1245);
   U196 : AND2_X1 port map( A1 => ADD_RS1(2), A2 => n784, ZN => n171);
   U197 : AND2_X1 port map( A1 => ADD_RS1(0), A2 => n1002, ZN => n172);
   U198 : AND2_X1 port map( A1 => n4004, A2 => n4003, ZN => n222);
   U199 : AND2_X1 port map( A1 => n3952, A2 => n3951, ZN => n223);
   U200 : NAND2_X1 port map( A1 => n693, A2 => n694, ZN => n352);
   U201 : OR2_X1 port map( A1 => n709, A2 => n708, ZN => n353);
   U202 : OR2_X1 port map( A1 => n1107, A2 => n1108, ZN => n354);
   U203 : OR2_X1 port map( A1 => n908, A2 => n909, ZN => n355);
   U204 : OR2_X1 port map( A1 => n1103, A2 => n1104, ZN => n356);
   U205 : OR2_X1 port map( A1 => n912, A2 => n913, ZN => n421);
   U206 : OR2_X1 port map( A1 => n920, A2 => n921, ZN => n422);
   U207 : OR2_X1 port map( A1 => n923, A2 => n924, ZN => n423);
   U208 : OR2_X1 port map( A1 => n1095, A2 => n1096, ZN => n424);
   U209 : OR2_X1 port map( A1 => n1109, A2 => n1110, ZN => n425);
   U210 : OR2_X1 port map( A1 => n914, A2 => n915, ZN => n426);
   U211 : OR2_X1 port map( A1 => n916, A2 => n917, ZN => n427);
   U212 : OR2_X1 port map( A1 => n1043, A2 => n1044, ZN => n428);
   U213 : OR2_X1 port map( A1 => n772, A2 => n771, ZN => n429);
   U214 : OR2_X1 port map( A1 => n1105, A2 => n1106, ZN => n430);
   U215 : OR2_X1 port map( A1 => n1064, A2 => n1063, ZN => n431);
   U216 : OR2_X1 port map( A1 => n897, A2 => n896, ZN => n432);
   U217 : OR2_X1 port map( A1 => n758, A2 => n757, ZN => n433);
   U218 : OR2_X1 port map( A1 => n683, A2 => n682, ZN => n434);
   U219 : OR2_X1 port map( A1 => n761, A2 => n762, ZN => n435);
   U220 : OR2_X1 port map( A1 => n774, A2 => n773, ZN => n436);
   U221 : OR2_X1 port map( A1 => n770, A2 => n769, ZN => n437);
   U222 : OR2_X1 port map( A1 => n782, A2 => n781, ZN => n438);
   U223 : AND2_X1 port map( A1 => ENABLE, A2 => n1538, ZN => n462);
   U224 : CLKBUF_X3 port map( A => n4113, Z => n1248);
   U225 : AND4_X1 port map( A1 => n979, A2 => n2260, A3 => n1274, A4 => n926, 
                           ZN => n463);
   U226 : OR2_X1 port map( A1 => n1048, A2 => n1047, ZN => n464);
   U227 : BUF_X2 port map( A => n988, Z => n1281);
   U228 : AND2_X1 port map( A1 => n3978, A2 => n3977, ZN => n465);
   U229 : AND2_X1 port map( A1 => n3926, A2 => n3925, ZN => n466);
   U230 : BUF_X2 port map( A => n988, Z => n1283);
   U231 : BUF_X1 port map( A => n972, Z => n739);
   U232 : BUF_X1 port map( A => n1208, Z => n892);
   U233 : OR2_X1 port map( A1 => n785, A2 => n786, ZN => n467);
   U234 : AND2_X2 port map( A1 => n1554, A2 => n1553, ZN => n468);
   U235 : AND2_X1 port map( A1 => n4030, A2 => n4029, ZN => n469);
   U236 : AND2_X2 port map( A1 => n1031, A2 => n705, ZN => n888);
   U237 : AND3_X1 port map( A1 => n4648, A2 => n4646, A3 => n4647, ZN => n470);
   U238 : AND2_X1 port map( A1 => n4081, A2 => n4082, ZN => n471);
   U239 : AND3_X1 port map( A1 => n4648, A2 => n4646, A3 => n4647, ZN => n1006)
                           ;
   U240 : AND2_X1 port map( A1 => n4056, A2 => n4055, ZN => n472);
   U241 : CLKBUF_X1 port map( A => n976, Z => n473);
   U242 : BUF_X1 port map( A => ADD_RS2(0), Z => n882);
   U243 : NOR2_X1 port map( A1 => n474, A2 => n475, ZN => n1968);
   U244 : NAND3_X1 port map( A1 => n515, A2 => n516, A3 => n549, ZN => n474);
   U245 : OR2_X1 port map( A1 => n1067, A2 => n1068, ZN => n475);
   U246 : NOR2_X1 port map( A1 => n476, A2 => n477, ZN => n1948);
   U247 : NAND3_X1 port map( A1 => n499, A2 => n500, A3 => n501, ZN => n476);
   U248 : OR2_X1 port map( A1 => n1075, A2 => n1076, ZN => n477);
   U249 : NOR2_X1 port map( A1 => n478, A2 => n479, ZN => n1826);
   U250 : NAND3_X1 port map( A1 => n793, A2 => n794, A3 => n795, ZN => n478);
   U251 : OR2_X1 port map( A1 => n1100, A2 => n1099, ZN => n479);
   U252 : CLKBUF_X3 port map( A => n4111, Z => n480);
   U253 : BUF_X1 port map( A => n2208, Z => n1132);
   U254 : BUF_X1 port map( A => n968, Z => n1196);
   U255 : AND2_X1 port map( A1 => n705, A2 => n692, ZN => n481);
   U256 : AND2_X1 port map( A1 => n705, A2 => n880, ZN => n482);
   U257 : AND2_X1 port map( A1 => n705, A2 => n880, ZN => n877);
   U258 : AND2_X1 port map( A1 => n172, A2 => n887, ZN => n483);
   U259 : AND2_X1 port map( A1 => n172, A2 => n887, ZN => n484);
   U260 : AND2_X1 port map( A1 => n172, A2 => n887, ZN => n972);
   U261 : BUF_X1 port map( A => n2209, Z => n1134);
   U262 : AND2_X2 port map( A1 => n2260, A2 => n883, ZN => n987);
   U263 : AND2_X2 port map( A1 => n2260, A2 => n883, ZN => n704);
   U264 : AND2_X2 port map( A1 => n2260, A2 => n883, ZN => n589);
   U265 : NAND2_X1 port map( A1 => n886, A2 => n468, ZN => n485);
   U266 : CLKBUF_X1 port map( A => n972, Z => n486);
   U267 : CLKBUF_X1 port map( A => n972, Z => n487);
   U268 : INV_X1 port map( A => ADD_RS2(3), ZN => n488);
   U269 : BUF_X1 port map( A => n702, Z => n489);
   U270 : BUF_X1 port map( A => n702, Z => n490);
   U271 : BUF_X1 port map( A => n702, Z => n577);
   U272 : NOR2_X1 port map( A1 => n2284, A2 => n354, ZN => n2296);
   U273 : OR2_X1 port map( A1 => n1229, A2 => n439, ZN => n491);
   U274 : OR2_X1 port map( A1 => n1225, A2 => n440, ZN => n492);
   U275 : NAND3_X1 port map( A1 => n491, A2 => n492, A3 => n2277, ZN => n2278);
   U276 : AND2_X1 port map( A1 => n1028, A2 => n171, ZN => n493);
   U277 : AND2_X1 port map( A1 => n1028, A2 => n171, ZN => n494);
   U278 : AND2_X1 port map( A1 => n1028, A2 => n171, ZN => n970);
   U279 : BUF_X1 port map( A => n968, Z => n495);
   U280 : BUF_X1 port map( A => n968, Z => n496);
   U281 : CLKBUF_X3 port map( A => n4088, Z => n1206);
   U282 : BUF_X1 port map( A => n484, Z => n497);
   U283 : CLKBUF_X3 port map( A => n4119, Z => n1262);
   U284 : CLKBUF_X3 port map( A => n4119, Z => n1263);
   U285 : CLKBUF_X3 port map( A => n4119, Z => n1264);
   U286 : BUF_X1 port map( A => n4116, Z => n1257);
   U287 : NAND4_X1 port map( A1 => n926, A2 => n878, A3 => n1274, A4 => n980, 
                           ZN => n498);
   U288 : BUF_X1 port map( A => n1036, Z => n878);
   U289 : OR2_X1 port map( A1 => n1941, A2 => n1146, ZN => n499);
   U290 : OR2_X1 port map( A1 => n818, A2 => n1149, ZN => n500);
   U291 : OR2_X1 port map( A1 => n3763, A2 => n1143, ZN => n501);
   U292 : NOR2_X1 port map( A1 => n502, A2 => n503, ZN => n1638);
   U293 : NAND3_X1 port map( A1 => n796, A2 => n797, A3 => n798, ZN => n502);
   U294 : OR2_X1 port map( A1 => n1087, A2 => n1086, ZN => n503);
   U295 : BUF_X1 port map( A => n702, Z => n578);
   U296 : NOR2_X1 port map( A1 => n3865, A2 => n355, ZN => n3877);
   U297 : OR2_X1 port map( A1 => n1229, A2 => n441, ZN => n504);
   U298 : OR2_X1 port map( A1 => n1226, A2 => n442, ZN => n505);
   U299 : NAND3_X1 port map( A1 => n504, A2 => n505, A3 => n3858, ZN => n3859);
   U300 : INV_X1 port map( A => n1561, ZN => n1014);
   U301 : CLKBUF_X3 port map( A => n2208, Z => n506);
   U302 : CLKBUF_X3 port map( A => n4113, Z => n509);
   U303 : NOR2_X1 port map( A1 => n2309, A2 => n356, ZN => n2321);
   U304 : OR2_X1 port map( A1 => n386, A2 => n1214, ZN => n510);
   U305 : OR2_X1 port map( A1 => n418, A2 => n1211, ZN => n511);
   U306 : NAND3_X1 port map( A1 => n510, A2 => n511, A3 => n2298, ZN => n2305);
   U307 : CLKBUF_X3 port map( A => n4091, Z => n1213);
   U308 : CLKBUF_X3 port map( A => n4090, Z => n1210);
   U309 : NOR2_X1 port map( A1 => n4109, A2 => n435, ZN => n4127);
   U310 : AND2_X1 port map( A1 => n4791, A2 => n1253, ZN => n513);
   U311 : AND2_X1 port map( A1 => n1250, A2 => n4336, ZN => n514);
   U312 : NOR3_X1 port map( A1 => n513, A2 => n2337, A3 => n514, ZN => n2345);
   U313 : BUF_X2 port map( A => n977, Z => n1253);
   U314 : BUF_X2 port map( A => n989, Z => n1250);
   U315 : OR2_X1 port map( A1 => n1961, A2 => n1146, ZN => n515);
   U316 : OR2_X1 port map( A1 => n817, A2 => n1149, ZN => n516);
   U317 : OR2_X1 port map( A1 => n3788, A2 => n1143, ZN => n549);
   U318 : AND3_X1 port map( A1 => n1560, A2 => n706, A3 => n881, ZN => n1031);
   U319 : BUF_X1 port map( A => n702, Z => n579);
   U320 : OR2_X1 port map( A1 => n161, A2 => n1117, ZN => n550);
   U321 : OR2_X1 port map( A1 => n1620, A2 => n2200, ZN => n551);
   U322 : NAND3_X1 port map( A1 => n550, A2 => n551, A3 => n1619, ZN => n1630);
   U323 : NOR2_X1 port map( A1 => n3840, A2 => n421, ZN => n3852);
   U324 : OR2_X1 port map( A1 => n1230, A2 => n443, ZN => n552);
   U325 : OR2_X1 port map( A1 => n1226, A2 => n444, ZN => n553);
   U326 : NAND3_X1 port map( A1 => n552, A2 => n553, A3 => n3833, ZN => n3834);
   U327 : NOR2_X1 port map( A1 => n3740, A2 => n422, ZN => n3752);
   U328 : OR2_X1 port map( A1 => n1228, A2 => n445, ZN => n554);
   U329 : OR2_X1 port map( A1 => n1226, A2 => n446, ZN => n555);
   U330 : NAND3_X1 port map( A1 => n554, A2 => n555, A3 => n3733, ZN => n3734);
   U331 : NOR2_X1 port map( A1 => n3715, A2 => n423, ZN => n3727);
   U332 : OR2_X1 port map( A1 => n1229, A2 => n447, ZN => n556);
   U333 : OR2_X1 port map( A1 => n1226, A2 => n448, ZN => n557);
   U334 : NAND3_X1 port map( A1 => n556, A2 => n557, A3 => n3708, ZN => n3709);
   U335 : NOR2_X1 port map( A1 => n2359, A2 => n424, ZN => n2371);
   U336 : OR2_X1 port map( A1 => n1228, A2 => n449, ZN => n558);
   U337 : OR2_X1 port map( A1 => n1225, A2 => n450, ZN => n559);
   U338 : NAND3_X1 port map( A1 => n558, A2 => n559, A3 => n2352, ZN => n2353);
   U339 : NOR2_X1 port map( A1 => n2255, A2 => n425, ZN => n2271);
   U340 : OR2_X1 port map( A1 => n1230, A2 => n451, ZN => n560);
   U341 : OR2_X1 port map( A1 => n1225, A2 => n452, ZN => n561);
   U342 : NAND3_X1 port map( A1 => n560, A2 => n561, A3 => n2248, ZN => n2249);
   U343 : CLKBUF_X3 port map( A => n4099, Z => n1228);
   U344 : CLKBUF_X3 port map( A => n4098, Z => n1225);
   U345 : NOR2_X1 port map( A1 => n3815, A2 => n426, ZN => n3827);
   U346 : OR2_X1 port map( A1 => n1230, A2 => n453, ZN => n562);
   U347 : OR2_X1 port map( A1 => n1226, A2 => n454, ZN => n563);
   U348 : NAND3_X1 port map( A1 => n562, A2 => n563, A3 => n3808, ZN => n3809);
   U349 : NOR2_X1 port map( A1 => n3790, A2 => n427, ZN => n3802);
   U350 : OR2_X1 port map( A1 => n1228, A2 => n455, ZN => n564);
   U351 : OR2_X1 port map( A1 => n1226, A2 => n456, ZN => n565);
   U352 : NAND3_X1 port map( A1 => n564, A2 => n565, A3 => n3783, ZN => n3784);
   U353 : CLKBUF_X3 port map( A => n4098, Z => n1226);
   U354 : OR2_X1 port map( A1 => n3581, A2 => n1129, ZN => n566);
   U355 : OR2_X1 port map( A1 => n281, A2 => n1125, ZN => n567);
   U356 : NAND3_X1 port map( A1 => n566, A2 => n567, A3 => n1788, ZN => n1796);
   U357 : OR2_X1 port map( A1 => n2475, A2 => n1128, ZN => n568);
   U358 : OR2_X1 port map( A1 => n283, A2 => n1125, ZN => n569);
   U359 : NAND3_X1 port map( A1 => n568, A2 => n569, A3 => n1746, ZN => n1754);
   U360 : OR2_X1 port map( A1 => n3656, A2 => n1127, ZN => n570);
   U361 : OR2_X1 port map( A1 => n278, A2 => n1126, ZN => n571);
   U362 : NAND3_X1 port map( A1 => n570, A2 => n571, A3 => n1850, ZN => n1858);
   U363 : OR2_X1 port map( A1 => n3631, A2 => n1128, ZN => n572);
   U364 : OR2_X1 port map( A1 => n279, A2 => n1126, ZN => n573);
   U365 : NAND3_X1 port map( A1 => n1829, A2 => n573, A3 => n572, ZN => n1837);
   U366 : NOR2_X1 port map( A1 => n1673, A2 => n467, ZN => n1680);
   U367 : OR2_X1 port map( A1 => n831, A2 => n1148, ZN => n574);
   U368 : OR2_X1 port map( A1 => n1672, A2 => n1145, ZN => n575);
   U369 : OR2_X1 port map( A1 => n2382, A2 => n1142, ZN => n576);
   U370 : NAND3_X1 port map( A1 => n575, A2 => n574, A3 => n576, ZN => n1673);
   U371 : CLKBUF_X3 port map( A => n2220, Z => n1142);
   U372 : BUF_X2 port map( A => n783, Z => n668);
   U373 : BUF_X2 port map( A => n482, Z => n1123);
   U374 : NOR2_X1 port map( A1 => n2224, A2 => n434, ZN => n2237);
   U375 : OR2_X1 port map( A1 => n805, A2 => n1150, ZN => n580);
   U376 : OR2_X1 port map( A1 => n2222, A2 => n1147, ZN => n581);
   U377 : OR2_X1 port map( A1 => n4104, A2 => n1144, ZN => n582);
   U378 : NAND3_X1 port map( A1 => n580, A2 => n581, A3 => n582, ZN => n2224);
   U379 : OR2_X1 port map( A1 => n1646, A2 => n1139, ZN => n583);
   U380 : OR2_X1 port map( A1 => n128, A2 => n1136, ZN => n584);
   U381 : NAND3_X1 port map( A1 => n583, A2 => n584, A3 => n1645, ZN => n1647);
   U382 : CLKBUF_X3 port map( A => n4118, Z => n1260);
   U383 : OR2_X1 port map( A1 => n3606, A2 => n1129, ZN => n585);
   U384 : OR2_X1 port map( A1 => n280, A2 => n1126, ZN => n586);
   U385 : NAND3_X1 port map( A1 => n1809, A2 => n586, A3 => n585, ZN => n1817);
   U386 : CLKBUF_X3 port map( A => n4111, Z => n1246);
   U387 : OR2_X1 port map( A1 => n1587, A2 => n1139, ZN => n587);
   U388 : OR2_X1 port map( A1 => n131, A2 => n1136, ZN => n588);
   U389 : NAND3_X1 port map( A1 => n587, A2 => n588, A3 => n1586, ZN => n1588);
   U390 : CLKBUF_X3 port map( A => n4116, Z => n590);
   U391 : CLKBUF_X1 port map( A => n1092, Z => n763);
   U392 : NOR2_X1 port map( A1 => n3690, A2 => n353, ZN => n3702);
   U393 : OR2_X1 port map( A1 => n821, A2 => n1238, ZN => n591);
   U394 : OR2_X1 port map( A1 => n3689, A2 => n1235, ZN => n592);
   U395 : OR2_X1 port map( A1 => n1232, A2 => n3688, ZN => n593);
   U396 : NAND3_X1 port map( A1 => n592, A2 => n591, A3 => n593, ZN => n3690);
   U397 : CLKBUF_X3 port map( A => n4108, Z => n1238);
   U398 : CLKBUF_X3 port map( A => n4106, Z => n1235);
   U399 : CLKBUF_X3 port map( A => n4105, Z => n1232);
   U400 : AND2_X1 port map( A1 => n4882, A2 => n1244, ZN => n594);
   U401 : AND2_X1 port map( A1 => n1242, A2 => n4073, ZN => n595);
   U402 : NOR3_X1 port map( A1 => n4072, A2 => n595, A3 => n594, ZN => n4084);
   U403 : NOR2_X1 port map( A1 => n2065, A2 => n429, ZN => n2072);
   U404 : OR2_X1 port map( A1 => n812, A2 => n1150, ZN => n596);
   U405 : OR2_X1 port map( A1 => n2064, A2 => n1147, ZN => n597);
   U406 : OR2_X1 port map( A1 => n3914, A2 => n1144, ZN => n598);
   U407 : NAND3_X1 port map( A1 => n597, A2 => n596, A3 => n598, ZN => n2065);
   U408 : CLKBUF_X3 port map( A => n2226, Z => n1161);
   U409 : CLKBUF_X3 port map( A => n2226, Z => n1160);
   U410 : NOR2_X1 port map( A1 => n2170, A2 => n433, ZN => n2177);
   U411 : OR2_X1 port map( A1 => n807, A2 => n1150, ZN => n599);
   U412 : OR2_X1 port map( A1 => n2169, A2 => n1147, ZN => n600);
   U413 : OR2_X1 port map( A1 => n4044, A2 => n1144, ZN => n601);
   U414 : NAND3_X1 port map( A1 => n600, A2 => n599, A3 => n601, ZN => n2170);
   U415 : BUF_X2 port map( A => n2223, Z => n1150);
   U416 : BUF_X2 port map( A => n2221, Z => n1147);
   U417 : AND2_X1 port map( A1 => n4881, A2 => n1244, ZN => n602);
   U418 : AND2_X1 port map( A1 => n1242, A2 => n4047, ZN => n603);
   U419 : AND2_X1 port map( A1 => n1077, A2 => n887, ZN => n966);
   U420 : NOR2_X1 port map( A1 => n3615, A2 => n428, ZN => n3627);
   U421 : OR2_X1 port map( A1 => n1205, A2 => n461, ZN => n604);
   U422 : OR2_X1 port map( A1 => n248, A2 => n1203, ZN => n605);
   U423 : NAND3_X1 port map( A1 => n604, A2 => n605, A3 => n3603, ZN => n3612);
   U424 : CLKBUF_X3 port map( A => n4087, Z => n1203);
   U425 : NOR2_X1 port map( A1 => n1570, A2 => n430, ZN => n1579);
   U426 : AND2_X1 port map( A1 => n1270, A2 => n4259, ZN => n606);
   U427 : AND2_X1 port map( A1 => n1267, A2 => n4227, ZN => n607);
   U428 : NOR3_X1 port map( A1 => n4026, A2 => n607, A3 => n606, ZN => n4030);
   U429 : OR2_X1 port map( A1 => n616, A2 => n1264, ZN => n608);
   U430 : OR2_X1 port map( A1 => n1261, A2 => n4025, ZN => n609);
   U431 : OR2_X1 port map( A1 => n1256, A2 => n4024, ZN => n610);
   U432 : NAND3_X1 port map( A1 => n608, A2 => n609, A3 => n610, ZN => n4026);
   U433 : AND2_X1 port map( A1 => n1270, A2 => n4260, ZN => n611);
   U434 : AND2_X1 port map( A1 => n1267, A2 => n4228, ZN => n612);
   U435 : NOR3_X1 port map( A1 => n4000, A2 => n612, A3 => n611, ZN => n4004);
   U436 : OR2_X1 port map( A1 => n617, A2 => n1264, ZN => n645);
   U437 : OR2_X1 port map( A1 => n1261, A2 => n3999, ZN => n646);
   U438 : OR2_X1 port map( A1 => n3998, A2 => n1258, ZN => n647);
   U439 : NAND3_X1 port map( A1 => n645, A2 => n646, A3 => n647, ZN => n4000);
   U440 : AND2_X1 port map( A1 => n1270, A2 => n4261, ZN => n648);
   U441 : AND2_X1 port map( A1 => n1267, A2 => n4229, ZN => n649);
   U442 : NOR3_X1 port map( A1 => n648, A2 => n649, A3 => n3974, ZN => n3978);
   U443 : OR2_X1 port map( A1 => n618, A2 => n1264, ZN => n650);
   U444 : OR2_X1 port map( A1 => n1261, A2 => n3973, ZN => n651);
   U445 : OR2_X1 port map( A1 => n3972, A2 => n1257, ZN => n652);
   U446 : NAND3_X1 port map( A1 => n650, A2 => n651, A3 => n652, ZN => n3974);
   U447 : AND2_X1 port map( A1 => n1270, A2 => n4262, ZN => n653);
   U448 : AND2_X1 port map( A1 => n1267, A2 => n4230, ZN => n654);
   U449 : NOR3_X1 port map( A1 => n653, A2 => n654, A3 => n3948, ZN => n3952);
   U450 : OR2_X1 port map( A1 => n619, A2 => n1264, ZN => n655);
   U451 : OR2_X1 port map( A1 => n1261, A2 => n3947, ZN => n656);
   U452 : OR2_X1 port map( A1 => n3946, A2 => n1257, ZN => n657);
   U453 : NAND3_X1 port map( A1 => n655, A2 => n656, A3 => n657, ZN => n3948);
   U454 : AND2_X1 port map( A1 => n1270, A2 => n4263, ZN => n658);
   U455 : AND2_X1 port map( A1 => n1267, A2 => n4231, ZN => n659);
   U456 : NOR3_X1 port map( A1 => n658, A2 => n659, A3 => n3922, ZN => n3926);
   U457 : OR2_X1 port map( A1 => n620, A2 => n1264, ZN => n660);
   U458 : OR2_X1 port map( A1 => n1261, A2 => n3921, ZN => n661);
   U459 : OR2_X1 port map( A1 => n3920, A2 => n1257, ZN => n662);
   U460 : NAND3_X1 port map( A1 => n660, A2 => n661, A3 => n662, ZN => n3922);
   U461 : BUF_X2 port map( A => n986, Z => n1270);
   U462 : BUF_X2 port map( A => n985, Z => n1267);
   U463 : AND2_X1 port map( A1 => n1156, A2 => n4882, ZN => n663);
   U464 : AND2_X1 port map( A1 => n1151, A2 => n4073, ZN => n664);
   U465 : NOR3_X1 port map( A1 => n2191, A2 => n664, A3 => n663, ZN => n2198);
   U466 : NOR2_X1 port map( A1 => n3968, A2 => n436, ZN => n3980);
   U467 : OR2_X1 port map( A1 => n810, A2 => n1239, ZN => n665);
   U468 : OR2_X1 port map( A1 => n3967, A2 => n1236, ZN => n666);
   U469 : OR2_X1 port map( A1 => n1233, A2 => n3966, ZN => n667);
   U470 : NAND3_X1 port map( A1 => n666, A2 => n665, A3 => n667, ZN => n3968);
   U471 : AND2_X1 port map( A1 => n1077, A2 => n887, ZN => n702);
   U472 : BUF_X2 port map( A => n783, Z => n669);
   U473 : NOR2_X1 port map( A1 => n2459, A2 => n431, ZN => n2471);
   U474 : OR2_X1 port map( A1 => n828, A2 => n1237, ZN => n670);
   U475 : OR2_X1 port map( A1 => n2458, A2 => n1234, ZN => n671);
   U476 : OR2_X1 port map( A1 => n1231, A2 => n2457, ZN => n672);
   U477 : NAND3_X1 port map( A1 => n671, A2 => n670, A3 => n672, ZN => n2459);
   U478 : NOR2_X1 port map( A1 => n2384, A2 => n432, ZN => n2396);
   U479 : OR2_X1 port map( A1 => n831, A2 => n1237, ZN => n673);
   U480 : OR2_X1 port map( A1 => n2383, A2 => n1234, ZN => n674);
   U481 : OR2_X1 port map( A1 => n1231, A2 => n2382, ZN => n675);
   U482 : NAND3_X1 port map( A1 => n674, A2 => n673, A3 => n675, ZN => n2384);
   U483 : CLKBUF_X3 port map( A => n4108, Z => n1237);
   U484 : CLKBUF_X3 port map( A => n4106, Z => n1234);
   U485 : CLKBUF_X3 port map( A => n4105, Z => n1231);
   U486 : NOR2_X1 port map( A1 => n3994, A2 => n437, ZN => n4006);
   U487 : OR2_X1 port map( A1 => n1222, A2 => n3986, ZN => n676);
   U488 : OR2_X1 port map( A1 => n1221, A2 => n3985, ZN => n677);
   U489 : NAND3_X1 port map( A1 => n676, A2 => n677, A3 => n3984, ZN => n3989);
   U490 : BUF_X2 port map( A => n4096, Z => n1224);
   U491 : BUF_X2 port map( A => n4094, Z => n1221);
   U492 : BUF_X2 port map( A => n485, Z => n678);
   U493 : NOR2_X1 port map( A1 => n3916, A2 => n438, ZN => n3928);
   U494 : OR2_X1 port map( A1 => n812, A2 => n1239, ZN => n679);
   U495 : OR2_X1 port map( A1 => n3915, A2 => n1236, ZN => n680);
   U496 : OR2_X1 port map( A1 => n1233, A2 => n3914, ZN => n681);
   U497 : NAND3_X1 port map( A1 => n680, A2 => n679, A3 => n681, ZN => n3916);
   U498 : BUF_X2 port map( A => n4108, Z => n1239);
   U499 : BUF_X2 port map( A => n4106, Z => n1236);
   U500 : BUF_X2 port map( A => n4105, Z => n1233);
   U501 : AND2_X1 port map( A1 => n1028, A2 => n468, ZN => n783);
   U502 : NOR2_X1 port map( A1 => n3590, A2 => n464, ZN => n3602);
   U503 : AND2_X1 port map( A1 => n1155, A2 => n4883, ZN => n682);
   U504 : AND2_X1 port map( A1 => n1151, A2 => n4110, ZN => n683);
   U505 : OR2_X1 port map( A1 => n2185, A2 => n1141, ZN => n684);
   U506 : OR2_X1 port map( A1 => n102, A2 => n1138, ZN => n685);
   U507 : NAND3_X1 port map( A1 => n684, A2 => n685, A3 => n2184, ZN => n2186);
   U508 : BUF_X2 port map( A => n2214, Z => n1141);
   U509 : BUF_X2 port map( A => n2213, Z => n1138);
   U510 : NAND3_X1 port map( A1 => n472, A2 => n4057, A3 => n4058, ZN => n2567)
                           ;
   U511 : NAND3_X1 port map( A1 => n4032, A2 => n4031, A3 => n469, ZN => n2566)
                           ;
   U512 : AND2_X1 port map( A1 => n4880, A2 => n1244, ZN => n686);
   U513 : AND2_X1 port map( A1 => n1242, A2 => n4021, ZN => n687);
   U514 : AND4_X1 port map( A1 => n978, A2 => n171, A3 => n1186, A4 => n875, ZN
                           => n982);
   U515 : CLKBUF_X3 port map( A => n4099, Z => n1229);
   U516 : BUF_X1 port map( A => n968, Z => n688);
   U517 : AND2_X2 port map( A1 => n2265, A2 => n884, ZN => n968);
   U518 : AND2_X1 port map( A1 => n884, A2 => n1036, ZN => n689);
   U519 : AND3_X1 port map( A1 => n4652, A2 => n4653, A3 => n4654, ZN => n690);
   U520 : AND3_X1 port map( A1 => n4652, A2 => n4653, A3 => n4654, ZN => n1005)
                           ;
   U521 : BUF_X1 port map( A => n483, Z => n691);
   U522 : AND3_X1 port map( A1 => n1054, A2 => ADD_RS1(0), A3 => n1560, ZN => 
                           n692);
   U523 : NAND2_X1 port map( A1 => n1151, A2 => n2360, ZN => n693);
   U524 : NAND2_X1 port map( A1 => n1156, A2 => n4856, ZN => n694);
   U525 : NOR3_X1 port map( A1 => ADD_RS2(0), A2 => ADD_RS2(4), A3 => 
                           ADD_RS2(3), ZN => n695);
   U526 : INV_X1 port map( A => ADD_RS2(2), ZN => n696);
   U527 : BUF_X2 port map( A => n967, Z => n697);
   U528 : NOR2_X1 port map( A1 => n2240, A2 => ADD_RS2(1), ZN => n1036);
   U529 : CLKBUF_X3 port map( A => n2225, Z => n1157);
   U530 : CLKBUF_X3 port map( A => n2225, Z => n1158);
   U531 : AND2_X1 port map( A1 => n1166, A2 => n4791, ZN => n698);
   U532 : AND2_X1 port map( A1 => n1163, A2 => n4336, ZN => n699);
   U533 : NOR3_X1 port map( A1 => n698, A2 => n699, A3 => n1632, ZN => n1637);
   U534 : BUF_X2 port map( A => n991, Z => n1166);
   U535 : BUF_X2 port map( A => n996, Z => n1163);
   U536 : BUF_X1 port map( A => n968, Z => n1197);
   U537 : BUF_X2 port map( A => n481, Z => n1124);
   U538 : AND2_X1 port map( A1 => n4862, A2 => n1243, ZN => n700);
   U539 : AND2_X1 port map( A1 => n1240, A2 => n3566, ZN => n701);
   U540 : NOR3_X1 port map( A1 => n3565, A2 => n701, A3 => n700, ZN => n3577);
   U541 : CLKBUF_X2 port map( A => n2220, Z => n1143);
   U542 : CLKBUF_X3 port map( A => n2230, Z => n1176);
   U543 : AND2_X1 port map( A1 => n1036, A2 => n695, ZN => n879);
   U544 : BUF_X2 port map( A => n2220, Z => n1144);
   U545 : INV_X1 port map( A => n2241, ZN => n703);
   U546 : NAND3_X1 port map( A1 => n4084, A2 => n4083, A3 => n471, ZN => n2568)
                           ;
   U547 : INV_X1 port map( A => ADD_RS1(3), ZN => n706);
   U548 : BUF_X1 port map( A => n2226, Z => n707);
   U549 : AND2_X1 port map( A1 => n4867, A2 => n463, ZN => n708);
   U550 : AND2_X1 port map( A1 => n1241, A2 => n3691, ZN => n709);
   U551 : AND2_X1 port map( A1 => n883, A2 => n973, ZN => n710);
   U552 : AND2_X1 port map( A1 => n1181, A2 => n4266, ZN => n711);
   U553 : AND2_X1 port map( A1 => n1178, A2 => n4234, ZN => n712);
   U554 : NOR3_X1 port map( A1 => n711, A2 => n712, A3 => n2004, ZN => n2007);
   U555 : OR2_X1 port map( A1 => n623, A2 => n1176, ZN => n713);
   U556 : OR2_X1 port map( A1 => n3845, A2 => n1172, ZN => n714);
   U557 : OR2_X1 port map( A1 => n3844, A2 => n1169, ZN => n715);
   U558 : NAND3_X1 port map( A1 => n713, A2 => n714, A3 => n715, ZN => n2004);
   U559 : AND2_X1 port map( A1 => n1180, A2 => n4286, ZN => n716);
   U560 : AND2_X1 port map( A1 => n1177, A2 => n4254, ZN => n717);
   U561 : NOR3_X1 port map( A1 => n716, A2 => n717, A3 => n1594, ZN => n1597);
   U562 : OR2_X1 port map( A1 => n643, A2 => n1176, ZN => n718);
   U563 : OR2_X1 port map( A1 => n2289, A2 => n1172, ZN => n719);
   U564 : OR2_X1 port map( A1 => n2288, A2 => n1169, ZN => n720);
   U565 : NAND3_X1 port map( A1 => n718, A2 => n719, A3 => n720, ZN => n1594);
   U566 : AND2_X1 port map( A1 => n1181, A2 => n4268, ZN => n721);
   U567 : AND2_X1 port map( A1 => n1178, A2 => n4236, ZN => n722);
   U568 : NOR3_X1 port map( A1 => n721, A2 => n722, A3 => n1963, ZN => n1966);
   U569 : OR2_X1 port map( A1 => n625, A2 => n1174, ZN => n723);
   U570 : OR2_X1 port map( A1 => n3795, A2 => n1171, ZN => n724);
   U571 : OR2_X1 port map( A1 => n3794, A2 => n1170, ZN => n725);
   U572 : NAND3_X1 port map( A1 => n723, A2 => n724, A3 => n725, ZN => n1963);
   U573 : AND2_X1 port map( A1 => n1168, A2 => n4813, ZN => n726);
   U574 : AND2_X1 port map( A1 => n1165, A2 => n4314, ZN => n727);
   U575 : NOR3_X1 port map( A1 => n726, A2 => n727, A3 => n2087, ZN => n2092);
   U576 : BUF_X2 port map( A => n991, Z => n1168);
   U577 : BUF_X2 port map( A => n996, Z => n1165);
   U578 : AND2_X1 port map( A1 => n1181, A2 => n4269, ZN => n728);
   U579 : AND2_X1 port map( A1 => n1178, A2 => n4237, ZN => n729);
   U580 : NOR3_X1 port map( A1 => n728, A2 => n729, A3 => n1943, ZN => n1946);
   U581 : OR2_X1 port map( A1 => n626, A2 => n1174, ZN => n730);
   U582 : OR2_X1 port map( A1 => n3770, A2 => n1172, ZN => n731);
   U583 : OR2_X1 port map( A1 => n3769, A2 => n1170, ZN => n732);
   U584 : NAND3_X1 port map( A1 => n730, A2 => n731, A3 => n732, ZN => n1943);
   U585 : AND2_X1 port map( A1 => n1181, A2 => n4270, ZN => n733);
   U586 : AND2_X1 port map( A1 => n1178, A2 => n4238, ZN => n734);
   U587 : NOR3_X1 port map( A1 => n733, A2 => n734, A3 => n1923, ZN => n1926);
   U588 : OR2_X1 port map( A1 => n627, A2 => n1174, ZN => n735);
   U589 : OR2_X1 port map( A1 => n3745, A2 => n1173, ZN => n736);
   U590 : OR2_X1 port map( A1 => n3744, A2 => n1170, ZN => n737);
   U591 : NAND3_X1 port map( A1 => n735, A2 => n736, A3 => n737, ZN => n1923);
   U592 : BUF_X1 port map( A => n483, Z => n738);
   U593 : AND2_X1 port map( A1 => n1181, A2 => n4271, ZN => n740);
   U594 : AND2_X1 port map( A1 => n1178, A2 => n4239, ZN => n741);
   U595 : NOR3_X1 port map( A1 => n740, A2 => n741, A3 => n1903, ZN => n1906);
   U596 : OR2_X1 port map( A1 => n628, A2 => n1174, ZN => n742);
   U597 : OR2_X1 port map( A1 => n3720, A2 => n1173, ZN => n743);
   U598 : OR2_X1 port map( A1 => n3719, A2 => n1169, ZN => n744);
   U599 : NAND3_X1 port map( A1 => n742, A2 => n743, A3 => n744, ZN => n1903);
   U600 : BUF_X2 port map( A => n990, Z => n1181);
   U601 : BUF_X2 port map( A => n992, Z => n1178);
   U602 : AND2_X1 port map( A1 => n1180, A2 => n4287, ZN => n745);
   U603 : AND2_X1 port map( A1 => n1177, A2 => n4255, ZN => n746);
   U604 : NOR3_X1 port map( A1 => n745, A2 => n746, A3 => n1573, ZN => n1577);
   U605 : OR2_X1 port map( A1 => n644, A2 => n1175, ZN => n747);
   U606 : OR2_X1 port map( A1 => n2262, A2 => n1171, ZN => n748);
   U607 : OR2_X1 port map( A1 => n2261, A2 => n1169, ZN => n749);
   U608 : NAND3_X1 port map( A1 => n747, A2 => n748, A3 => n749, ZN => n1573);
   U609 : BUF_X2 port map( A => n990, Z => n1180);
   U610 : BUF_X2 port map( A => n992, Z => n1177);
   U611 : AND2_X1 port map( A1 => n695, A2 => n973, ZN => n750);
   U612 : OR2_X1 port map( A1 => n4093, A2 => n1128, ZN => n751);
   U613 : OR2_X1 port map( A1 => n261, A2 => n485, ZN => n752);
   U614 : NAND3_X1 port map( A1 => n2203, A2 => n752, A3 => n751, ZN => n2218);
   U615 : OR2_X1 port map( A1 => n4063, A2 => n1127, ZN => n753);
   U616 : OR2_X1 port map( A1 => n262, A2 => n485, ZN => n754);
   U617 : NAND3_X1 port map( A1 => n2180, A2 => n754, A3 => n753, ZN => n2188);
   U618 : BUF_X2 port map( A => n2205, Z => n1129);
   U619 : INV_X1 port map( A => ADD_RS2(4), ZN => n755);
   U620 : BUF_X2 port map( A => n1000, Z => n1217);
   U621 : INV_X1 port map( A => n84, ZN => n756);
   U622 : AND2_X1 port map( A1 => n1154, A2 => n4881, ZN => n757);
   U623 : AND2_X1 port map( A1 => n1152, A2 => n4047, ZN => n758);
   U624 : AND2_X2 port map( A1 => n880, A2 => n887, ZN => n759);
   U625 : AND2_X2 port map( A1 => n692, A2 => n887, ZN => n760);
   U626 : AND2_X1 port map( A1 => n692, A2 => n887, ZN => n1029);
   U627 : BUF_X2 port map( A => n1000, Z => n1218);
   U628 : AND2_X1 port map( A1 => n4883, A2 => n1244, ZN => n761);
   U629 : AND2_X1 port map( A1 => n1242, A2 => n4110, ZN => n762);
   U630 : INV_X1 port map( A => n1554, ZN => n764);
   U631 : BUF_X1 port map( A => ADD_RS1(4), Z => n1092);
   U632 : AND2_X1 port map( A1 => n1155, A2 => n4880, ZN => n765);
   U633 : AND2_X1 port map( A1 => n1152, A2 => n4021, ZN => n766);
   U634 : AND2_X1 port map( A1 => n1156, A2 => n4878, ZN => n767);
   U635 : AND2_X1 port map( A1 => n1153, A2 => n3969, ZN => n768);
   U636 : NAND3_X1 port map( A1 => n4006, A2 => n4005, A3 => n222, ZN => n2565)
                           ;
   U637 : AND2_X1 port map( A1 => n4879, A2 => n1244, ZN => n769);
   U638 : AND2_X1 port map( A1 => n1242, A2 => n3995, ZN => n770);
   U639 : AND2_X1 port map( A1 => n1156, A2 => n4876, ZN => n771);
   U640 : AND2_X1 port map( A1 => n1153, A2 => n3917, ZN => n772);
   U641 : BUF_X2 port map( A => n982, Z => n1156);
   U642 : BUF_X2 port map( A => n981, Z => n1153);
   U643 : NAND3_X1 port map( A1 => n3980, A2 => n3979, A3 => n465, ZN => n2564)
                           ;
   U644 : AND2_X1 port map( A1 => n4878, A2 => n1244, ZN => n773);
   U645 : AND2_X1 port map( A1 => n1242, A2 => n3969, ZN => n774);
   U646 : NAND3_X1 port map( A1 => n3954, A2 => n3953, A3 => n223, ZN => n2563)
                           ;
   U647 : AND2_X1 port map( A1 => n4877, A2 => n1244, ZN => n775);
   U648 : AND2_X1 port map( A1 => n1242, A2 => n3943, ZN => n776);
   U649 : NOR3_X1 port map( A1 => n3942, A2 => n776, A3 => n775, ZN => n3954);
   U650 : AND2_X1 port map( A1 => n1156, A2 => n4854, ZN => n777);
   U651 : AND2_X1 port map( A1 => n1151, A2 => n2310, ZN => n778);
   U652 : AND2_X1 port map( A1 => n1154, A2 => n4866, ZN => n779);
   U653 : AND2_X1 port map( A1 => n1152, A2 => n3666, ZN => n780);
   U654 : NAND3_X1 port map( A1 => n3928, A2 => n3927, A3 => n466, ZN => n2562)
                           ;
   U655 : AND2_X1 port map( A1 => n4876, A2 => n1244, ZN => n781);
   U656 : AND2_X1 port map( A1 => n1242, A2 => n3917, ZN => n782);
   U657 : BUF_X2 port map( A => n984, Z => n1244);
   U658 : BUF_X2 port map( A => n983, Z => n1242);
   U659 : BUF_X1 port map( A => ADD_RS1(1), Z => n784);
   U660 : AND2_X2 port map( A1 => n1028, A2 => n468, ZN => n969);
   U661 : AND2_X1 port map( A1 => n1155, A2 => n4857, ZN => n785);
   U662 : AND2_X1 port map( A1 => n1153, A2 => n2385, ZN => n786);
   U663 : NAND3_X1 port map( A1 => n787, A2 => n788, A3 => n789, ZN => n2340);
   U664 : OR2_X1 port map( A1 => n641, A2 => n1262, ZN => n787);
   U665 : OR2_X1 port map( A1 => n1260, A2 => n2339, ZN => n788);
   U666 : OR2_X1 port map( A1 => n590, A2 => n2338, ZN => n789);
   U667 : NOR3_X1 port map( A1 => n4656, A2 => n4645, A3 => n4657, ZN => n4655)
                           ;
   U668 : AND2_X1 port map( A1 => n2470, A2 => n2468, ZN => n790);
   U669 : AND2_X1 port map( A1 => n2445, A2 => n2443, ZN => n791);
   U670 : AND2_X1 port map( A1 => n2395, A2 => n2393, ZN => n792);
   U671 : OR2_X1 port map( A1 => n824, A2 => n1149, ZN => n793);
   U672 : OR2_X1 port map( A1 => n1819, A2 => n1146, ZN => n794);
   U673 : OR2_X1 port map( A1 => n3613, A2 => n1143, ZN => n795);
   U674 : OR2_X1 port map( A1 => n833, A2 => n1148, ZN => n796);
   U675 : OR2_X1 port map( A1 => n1631, A2 => n1145, ZN => n797);
   U676 : OR2_X1 port map( A1 => n2332, A2 => n1142, ZN => n798);
   U677 : OR2_X1 port map( A1 => n835, A2 => n1148, ZN => n799);
   U678 : OR2_X1 port map( A1 => n1592, A2 => n1145, ZN => n800);
   U679 : OR2_X1 port map( A1 => n2282, A2 => n1142, ZN => n801);
   U680 : NOR2_X1 port map( A1 => n802, A2 => n803, ZN => n1599);
   U681 : NAND3_X1 port map( A1 => n800, A2 => n799, A3 => n801, ZN => n802);
   U682 : OR2_X1 port map( A1 => n1102, A2 => n1101, ZN => n803);
   U683 : AND2_X1 port map( A1 => n804, A2 => n922, ZN => n2009);
   U684 : NOR3_X1 port map( A1 => n1011, A2 => n1010, A3 => n1012, ZN => n804);
   U685 : AND2_X1 port map( A1 => n869, A2 => n927, ZN => n1928);
   U686 : NOR3_X1 port map( A1 => n1008, A2 => n1007, A3 => n1009, ZN => n869);
   U687 : NAND3_X1 port map( A1 => n870, A2 => n871, A3 => n872, ZN => n1652);
   U688 : OR2_X1 port map( A1 => n1651, A2 => n1145, ZN => n870);
   U689 : OR2_X1 port map( A1 => n832, A2 => n1148, ZN => n871);
   U690 : OR2_X1 port map( A1 => n2357, A2 => n1142, ZN => n872);
   U691 : BUF_X2 port map( A => n1000, Z => n1216);
   U692 : BUF_X2 port map( A => n967, Z => n1199);
   U693 : AND3_X1 port map( A1 => n2344, A2 => n2343, A3 => n2345, ZN => n873);
   U694 : NAND2_X1 port map( A1 => n1005, A2 => n1027, ZN => n874);
   U695 : NAND2_X1 port map( A1 => n690, A2 => n77, ZN => n875);
   U696 : NAND4_X1 port map( A1 => n1574, A2 => n705, A3 => n1187, A4 => n978, 
                           ZN => n876);
   U697 : NAND2_X1 port map( A1 => n4655, A2 => n1005, ZN => n1574);
   U698 : CLKBUF_X3 port map( A => n2230, Z => n1175);
   U699 : CLKBUF_X3 port map( A => n2229, Z => n1173);
   U700 : CLKBUF_X3 port map( A => n2230, Z => n1174);
   U701 : AND2_X2 port map( A1 => n884, A2 => n1036, ZN => n998);
   U702 : CLKBUF_X3 port map( A => n2228, Z => n1170);
   U703 : CLKBUF_X3 port map( A => n2229, Z => n1172);
   U704 : AND2_X1 port map( A1 => n695, A2 => n1036, ZN => n997);
   U705 : CLKBUF_X3 port map( A => n2228, Z => n1169);
   U706 : CLKBUF_X3 port map( A => n2229, Z => n1171);
   U707 : AND3_X1 port map( A1 => n1054, A2 => ADD_RS1(0), A3 => n1560, ZN => 
                           n880);
   U708 : CLKBUF_X1 port map( A => n4116, Z => n1256);
   U709 : CLKBUF_X3 port map( A => n4116, Z => n1258);
   U710 : INV_X1 port map( A => ADD_RS1(0), ZN => n881);
   U711 : AND3_X1 port map( A1 => n882, A2 => n1062, A3 => n2243, ZN => n883);
   U712 : AND3_X1 port map( A1 => n2243, A2 => n882, A3 => n488, ZN => n884);
   U713 : AND3_X1 port map( A1 => n882, A2 => n755, A3 => n1061, ZN => n1030);
   U714 : CLKBUF_X1 port map( A => ADD_RS2(3), Z => n885);
   U715 : AND3_X1 port map( A1 => ADD_RS1(0), A2 => n1054, A3 => n1560, ZN => 
                           n886);
   U716 : BUF_X1 port map( A => n1077, Z => n1053);
   U717 : CLKBUF_X1 port map( A => ADD_RS1(0), Z => n890);
   U718 : CLKBUF_X1 port map( A => n889, Z => n891);
   U719 : NOR3_X1 port map( A1 => n4650, A2 => n4651, A3 => n4645, ZN => n893);
   U720 : NOR3_X1 port map( A1 => n4650, A2 => n4651, A3 => n4645, ZN => n4649)
                           ;
   U721 : BUF_X2 port map( A => n967, Z => n1200);
   U722 : BUF_X2 port map( A => n997, Z => n1209);
   U723 : CLKBUF_X3 port map( A => n4118, Z => n1259);
   U724 : BUF_X2 port map( A => n997, Z => n1208);
   U725 : BUF_X2 port map( A => n481, Z => n1024);
   U726 : AND2_X1 port map( A1 => n1155, A2 => n4863, ZN => n894);
   U727 : AND2_X1 port map( A1 => n1153, A2 => n3591, ZN => n895);
   U728 : AND2_X1 port map( A1 => n4857, A2 => n1243, ZN => n896);
   U729 : AND2_X1 port map( A1 => n1240, A2 => n2385, ZN => n897);
   U730 : BUF_X2 port map( A => n984, Z => n1243);
   U731 : BUF_X2 port map( A => n983, Z => n1240);
   U732 : AND2_X1 port map( A1 => n1154, A2 => n4862, ZN => n898);
   U733 : AND2_X1 port map( A1 => n1151, A2 => n3566, ZN => n899);
   U734 : AND2_X1 port map( A1 => n1154, A2 => n4875, ZN => n900);
   U735 : AND2_X1 port map( A1 => n1151, A2 => n3891, ZN => n901);
   U736 : AND2_X1 port map( A1 => n1155, A2 => n4861, ZN => n902);
   U737 : AND2_X1 port map( A1 => n1153, A2 => n2485, ZN => n903);
   U738 : BUF_X2 port map( A => n981, Z => n1151);
   U739 : AND2_X1 port map( A1 => n1155, A2 => n4874, ZN => n904);
   U740 : AND2_X1 port map( A1 => n1151, A2 => n3866, ZN => n905);
   U741 : AND2_X1 port map( A1 => n4875, A2 => n463, ZN => n906);
   U742 : AND2_X1 port map( A1 => n1241, A2 => n3891, ZN => n907);
   U743 : AND2_X1 port map( A1 => n4874, A2 => n463, ZN => n908);
   U744 : AND2_X1 port map( A1 => n1241, A2 => n3866, ZN => n909);
   U745 : AND2_X1 port map( A1 => n1156, A2 => n4872, ZN => n910);
   U746 : AND2_X1 port map( A1 => n1152, A2 => n3816, ZN => n911);
   U747 : BUF_X2 port map( A => n982, Z => n1155);
   U748 : BUF_X2 port map( A => n981, Z => n1152);
   U749 : AND2_X1 port map( A1 => n4873, A2 => n463, ZN => n912);
   U750 : AND2_X1 port map( A1 => n1241, A2 => n3841, ZN => n913);
   U751 : AND2_X1 port map( A1 => n4872, A2 => n463, ZN => n914);
   U752 : AND2_X1 port map( A1 => n1241, A2 => n3816, ZN => n915);
   U753 : AND2_X1 port map( A1 => n4871, A2 => n463, ZN => n916);
   U754 : AND2_X1 port map( A1 => n1241, A2 => n3791, ZN => n917);
   U755 : BUF_X2 port map( A => n983, Z => n1241);
   U756 : AND2_X1 port map( A1 => n4870, A2 => n463, ZN => n918);
   U757 : AND2_X1 port map( A1 => n1241, A2 => n3766, ZN => n919);
   U758 : AND2_X1 port map( A1 => n4869, A2 => n463, ZN => n920);
   U759 : AND2_X1 port map( A1 => n1241, A2 => n3741, ZN => n921);
   U760 : NOR2_X1 port map( A1 => n1033, A2 => n1032, ZN => n922);
   U761 : AND2_X1 port map( A1 => n4868, A2 => n463, ZN => n923);
   U762 : AND2_X1 port map( A1 => n1241, A2 => n3716, ZN => n924);
   U763 : NAND2_X1 port map( A1 => n1006, A2 => n893, ZN => n925);
   U764 : NAND2_X1 port map( A1 => n4649, A2 => n470, ZN => n926);
   U765 : NAND2_X1 port map( A1 => n1006, A2 => n4649, ZN => n2264);
   U766 : NOR2_X1 port map( A1 => n1079, A2 => n1078, ZN => n927);
   U767 : NOR2_X1 port map( A1 => n1652, A2 => n352, ZN => n1659);
   U768 : OR2_X1 port map( A1 => n1134, A2 => n3832, ZN => n928);
   U769 : OR2_X1 port map( A1 => n239, A2 => n1132, ZN => n929);
   U770 : NAND3_X1 port map( A1 => n928, A2 => n929, A3 => n1994, ZN => n1999);
   U771 : BUF_X2 port map( A => n982, Z => n1154);
   U772 : CLKBUF_X1 port map( A => n1004, Z => n1276);
   U773 : BUF_X2 port map( A => n1004, Z => n1275);
   U774 : BUF_X1 port map( A => n1539, Z => n1538);
   U775 : BUF_X1 port map( A => n483, Z => n1113);
   U776 : BUF_X1 port map( A => n484, Z => n1112);
   U777 : BUF_X1 port map( A => n484, Z => n1111);
   U778 : BUF_X1 port map( A => n1449, Z => n1539);
   U779 : BUF_X1 port map( A => n1449, Z => n1540);
   U780 : BUF_X1 port map( A => n1449, Z => n1541);
   U781 : BUF_X1 port map( A => n1450, Z => n1542);
   U782 : BUF_X1 port map( A => n1450, Z => n1543);
   U783 : BUF_X1 port map( A => n1450, Z => n1544);
   U784 : BUF_X1 port map( A => n1451, Z => n1545);
   U785 : BUF_X1 port map( A => n1451, Z => n1546);
   U786 : BUF_X1 port map( A => n1451, Z => n1547);
   U787 : BUF_X1 port map( A => n1452, Z => n1548);
   U788 : BUF_X1 port map( A => n1452, Z => n1549);
   U789 : BUF_X1 port map( A => n1452, Z => n1550);
   U790 : BUF_X1 port map( A => n1453, Z => n1551);
   U791 : BUF_X1 port map( A => n1453, Z => n1552);
   U792 : BUF_X2 port map( A => n4096, Z => n1223);
   U793 : BUF_X2 port map( A => n4096, Z => n1222);
   U794 : BUF_X1 port map( A => n985, Z => n1266);
   U795 : BUF_X1 port map( A => n994, Z => n1278);
   U796 : BUF_X1 port map( A => n996, Z => n1164);
   U797 : BUF_X1 port map( A => n993, Z => n1190);
   U798 : BUF_X1 port map( A => n993, Z => n1191);
   U799 : BUF_X1 port map( A => n989, Z => n1251);
   U800 : BUF_X1 port map( A => n994, Z => n1279);
   U801 : BUF_X1 port map( A => n977, Z => n1254);
   U802 : BUF_X1 port map( A => n988, Z => n1282);
   U803 : BUF_X1 port map( A => n986, Z => n1269);
   U804 : BUF_X1 port map( A => n991, Z => n1167);
   U805 : BUF_X1 port map( A => n995, Z => n1193);
   U806 : BUF_X1 port map( A => n995, Z => n1194);
   U807 : BUF_X2 port map( A => n4094, Z => n1220);
   U808 : BUF_X2 port map( A => n4094, Z => n1219);
   U809 : AND2_X1 port map( A1 => n1002, A2 => n1572, ZN => n930);
   U810 : BUF_X1 port map( A => n4113, Z => n1249);
   U811 : BUF_X1 port map( A => n4111, Z => n1247);
   U812 : BUF_X1 port map( A => n989, Z => n1252);
   U813 : BUF_X1 port map( A => n993, Z => n1192);
   U814 : BUF_X1 port map( A => n994, Z => n1280);
   U815 : BUF_X1 port map( A => n977, Z => n1255);
   U816 : BUF_X1 port map( A => n2226, Z => n1162);
   U817 : BUF_X1 port map( A => n4091, Z => n1215);
   U818 : BUF_X1 port map( A => n4090, Z => n1212);
   U819 : BUF_X1 port map( A => n995, Z => n1195);
   U820 : AND2_X1 port map( A1 => n973, A2 => n695, ZN => n931);
   U821 : AND3_X1 port map( A1 => n763, A2 => n1572, A3 => n756, ZN => n971);
   U822 : BUF_X1 port map( A => n1454, Z => n1451);
   U823 : BUF_X1 port map( A => n1454, Z => n1452);
   U824 : BUF_X1 port map( A => n1455, Z => n1449);
   U825 : BUF_X1 port map( A => n1455, Z => n1450);
   U826 : BUF_X1 port map( A => n1454, Z => n1453);
   U827 : AND2_X2 port map( A1 => n696, A2 => ADD_RS2(1), ZN => n973);
   U828 : BUF_X1 port map( A => n4576, Z => n1362);
   U829 : BUF_X1 port map( A => n4576, Z => n1363);
   U830 : BUF_X1 port map( A => n4611, Z => n1371);
   U831 : BUF_X1 port map( A => n4611, Z => n1372);
   U832 : BUF_X1 port map( A => n4359, Z => n1305);
   U833 : BUF_X1 port map( A => n4359, Z => n1306);
   U834 : BUF_X1 port map( A => n4499, Z => n1332);
   U835 : BUF_X1 port map( A => n4499, Z => n1333);
   U836 : BUF_X1 port map( A => n4394, Z => n1308);
   U837 : BUF_X1 port map( A => n4394, Z => n1309);
   U838 : BUF_X1 port map( A => n4534, Z => n1341);
   U839 : BUF_X1 port map( A => n4534, Z => n1342);
   U840 : BUF_X1 port map( A => n4462, Z => n1320);
   U841 : BUF_X1 port map( A => n4462, Z => n1321);
   U842 : BUF_X1 port map( A => n4429, Z => n1317);
   U843 : BUF_X1 port map( A => n4429, Z => n1318);
   U844 : BUF_X1 port map( A => n4569, Z => n1353);
   U845 : BUF_X1 port map( A => n4569, Z => n1354);
   U846 : BUF_X1 port map( A => n4573, Z => n1359);
   U847 : BUF_X1 port map( A => n4573, Z => n1360);
   U848 : BUF_X1 port map( A => n4571, Z => n1356);
   U849 : BUF_X1 port map( A => n4571, Z => n1357);
   U850 : BUF_X1 port map( A => n4643, Z => n1374);
   U851 : BUF_X1 port map( A => n4643, Z => n1375);
   U852 : BUF_X1 port map( A => n4609, Z => n1368);
   U853 : BUF_X1 port map( A => n4609, Z => n1369);
   U854 : BUF_X1 port map( A => n4608, Z => n1365);
   U855 : BUF_X1 port map( A => n4608, Z => n1366);
   U856 : BUF_X1 port map( A => n4496, Z => n1329);
   U857 : BUF_X1 port map( A => n4496, Z => n1330);
   U858 : BUF_X1 port map( A => n4532, Z => n1338);
   U859 : BUF_X1 port map( A => n4532, Z => n1339);
   U860 : BUF_X1 port map( A => n4531, Z => n1335);
   U861 : BUF_X1 port map( A => n4531, Z => n1336);
   U862 : BUF_X1 port map( A => n4427, Z => n1314);
   U863 : BUF_X1 port map( A => n4427, Z => n1315);
   U864 : BUF_X1 port map( A => n4426, Z => n1311);
   U865 : BUF_X1 port map( A => n4426, Z => n1312);
   U866 : BUF_X1 port map( A => n4568, Z => n1350);
   U867 : BUF_X1 port map( A => n4568, Z => n1351);
   U868 : BUF_X1 port map( A => n4567, Z => n1347);
   U869 : BUF_X1 port map( A => n4567, Z => n1348);
   U870 : BUF_X1 port map( A => n4566, Z => n1344);
   U871 : BUF_X1 port map( A => n4566, Z => n1345);
   U872 : BUF_X1 port map( A => n4495, Z => n1326);
   U873 : BUF_X1 port map( A => n4495, Z => n1327);
   U874 : BUF_X1 port map( A => n4494, Z => n1323);
   U875 : BUF_X1 port map( A => n4494, Z => n1324);
   U876 : BUF_X1 port map( A => n4345, Z => n1290);
   U877 : BUF_X1 port map( A => n4345, Z => n1291);
   U878 : BUF_X1 port map( A => n4343, Z => n1287);
   U879 : BUF_X1 port map( A => n4343, Z => n1288);
   U880 : BUF_X1 port map( A => n4340, Z => n1284);
   U881 : BUF_X1 port map( A => n4340, Z => n1285);
   U882 : BUF_X1 port map( A => n4353, Z => n1302);
   U883 : BUF_X1 port map( A => n4353, Z => n1303);
   U884 : BUF_X1 port map( A => n4351, Z => n1299);
   U885 : BUF_X1 port map( A => n4351, Z => n1300);
   U886 : BUF_X1 port map( A => n4349, Z => n1296);
   U887 : BUF_X1 port map( A => n4349, Z => n1297);
   U888 : BUF_X1 port map( A => n4347, Z => n1293);
   U889 : BUF_X1 port map( A => n4347, Z => n1294);
   U890 : BUF_X1 port map( A => n1004, Z => n1274);
   U891 : BUF_X2 port map( A => n4121, Z => n1271);
   U892 : BUF_X2 port map( A => n2232, Z => n1183);
   U893 : BUF_X2 port map( A => n2232, Z => n1184);
   U894 : BUF_X2 port map( A => n4121, Z => n1272);
   U895 : BUF_X1 port map( A => n1004, Z => n1277);
   U896 : BUF_X1 port map( A => n1003, Z => n1189);
   U897 : BUF_X1 port map( A => n1003, Z => n1188);
   U898 : AND3_X1 port map( A1 => ADD_RS2(3), A2 => n755, A3 => n882, ZN => 
                           n974);
   U899 : AND3_X1 port map( A1 => ADD_RS2(3), A2 => n2259, A3 => n2243, ZN => 
                           n975);
   U900 : AND2_X1 port map( A1 => ADD_RS2(3), A2 => n999, ZN => n976);
   U901 : AND4_X1 port map( A1 => n703, A2 => n473, A3 => n1274, A4 => n926, ZN
                           => n977);
   U902 : AND3_X1 port map( A1 => n763, A2 => ADD_RS1(0), A3 => n756, ZN => 
                           n978);
   U903 : AND2_X1 port map( A1 => n999, A2 => n1062, ZN => n979);
   U904 : AND3_X1 port map( A1 => n2259, A2 => n885, A3 => n891, ZN => n980);
   U905 : BUF_X1 port map( A => n4576, Z => n1364);
   U906 : BUF_X1 port map( A => n4611, Z => n1373);
   U907 : BUF_X1 port map( A => n4359, Z => n1307);
   U908 : BUF_X1 port map( A => n4499, Z => n1334);
   U909 : BUF_X1 port map( A => n4394, Z => n1310);
   U910 : BUF_X1 port map( A => n4534, Z => n1343);
   U911 : BUF_X1 port map( A => n4462, Z => n1322);
   U912 : BUF_X1 port map( A => n4429, Z => n1319);
   U913 : BUF_X1 port map( A => n4569, Z => n1355);
   U914 : BUF_X1 port map( A => n4573, Z => n1361);
   U915 : BUF_X1 port map( A => n4571, Z => n1358);
   U916 : BUF_X1 port map( A => n4643, Z => n1376);
   U917 : BUF_X1 port map( A => n4609, Z => n1370);
   U918 : BUF_X1 port map( A => n4608, Z => n1367);
   U919 : BUF_X1 port map( A => n4496, Z => n1331);
   U920 : BUF_X1 port map( A => n4532, Z => n1340);
   U921 : BUF_X1 port map( A => n4531, Z => n1337);
   U922 : BUF_X1 port map( A => n4427, Z => n1316);
   U923 : BUF_X1 port map( A => n4426, Z => n1313);
   U924 : BUF_X1 port map( A => n4345, Z => n1292);
   U925 : BUF_X1 port map( A => n4343, Z => n1289);
   U926 : BUF_X1 port map( A => n4340, Z => n1286);
   U927 : BUF_X1 port map( A => n4568, Z => n1352);
   U928 : BUF_X1 port map( A => n4567, Z => n1349);
   U929 : BUF_X1 port map( A => n4566, Z => n1346);
   U930 : BUF_X1 port map( A => n4495, Z => n1328);
   U931 : BUF_X1 port map( A => n4494, Z => n1325);
   U932 : BUF_X1 port map( A => n4353, Z => n1304);
   U933 : BUF_X1 port map( A => n4351, Z => n1301);
   U934 : BUF_X1 port map( A => n4349, Z => n1298);
   U935 : BUF_X1 port map( A => n4347, Z => n1295);
   U936 : AND4_X1 port map( A1 => n874, A2 => n172, A3 => n1186, A4 => n705, ZN
                           => n981);
   U937 : AND4_X1 port map( A1 => n473, A2 => n973, A3 => n1274, A4 => n925, ZN
                           => n983);
   U938 : AND4_X1 port map( A1 => n979, A2 => n2260, A3 => n1274, A4 => n926, 
                           ZN => n984);
   U939 : BUF_X1 port map( A => n2232, Z => n1185);
   U940 : BUF_X1 port map( A => n4121, Z => n1273);
   U941 : AND4_X1 port map( A1 => n1001, A2 => n703, A3 => n1274, A4 => n925, 
                           ZN => n985);
   U942 : AND4_X1 port map( A1 => n979, A2 => n878, A3 => n1274, A4 => n925, ZN
                           => n986);
   U943 : AND4_X1 port map( A1 => n1001, A2 => n973, A3 => n1275, A4 => n925, 
                           ZN => n988);
   U944 : AND4_X1 port map( A1 => n473, A2 => n2260, A3 => n1274, A4 => n925, 
                           ZN => n989);
   U945 : AND4_X1 port map( A1 => n1574, A2 => n887, A3 => n1186, A4 => n978, 
                           ZN => n990);
   U946 : AND4_X1 port map( A1 => n172, A2 => n468, A3 => n1186, A4 => n875, ZN
                           => n991);
   U947 : AND4_X1 port map( A1 => n1574, A2 => n468, A3 => n1186, A4 => n971, 
                           ZN => n992);
   U948 : AND4_X1 port map( A1 => n978, A2 => n468, A3 => n1187, A4 => n875, ZN
                           => n993);
   U949 : AND4_X1 port map( A1 => n979, A2 => n703, A3 => n1275, A4 => n926, ZN
                           => n994);
   U950 : AND4_X1 port map( A1 => n1574, A2 => n705, A3 => n1187, A4 => n971, 
                           ZN => n995);
   U951 : AND4_X1 port map( A1 => n172, A2 => n171, A3 => n1186, A4 => n875, ZN
                           => n996);
   U952 : AND2_X1 port map( A1 => n889, A2 => n882, ZN => n999);
   U953 : AND3_X1 port map( A1 => n891, A2 => n2259, A3 => n1062, ZN => n1001);
   U954 : AND2_X1 port map( A1 => ADD_RS1(4), A2 => ADD_RS1(3), ZN => n1002);
   U955 : BUF_X1 port map( A => RST, Z => n1454);
   U956 : BUF_X1 port map( A => RST, Z => n1455);
   U957 : AND2_X1 port map( A1 => RD1, A2 => n462, ZN => n1003);
   U958 : AND2_X1 port map( A1 => RD2, A2 => n462, ZN => n1004);
   U959 : INV_X1 port map( A => DATAIN(0), ZN => n1378);
   U960 : INV_X1 port map( A => DATAIN(1), ZN => n1380);
   U961 : INV_X1 port map( A => DATAIN(2), ZN => n1382);
   U962 : INV_X1 port map( A => DATAIN(3), ZN => n1384);
   U963 : INV_X1 port map( A => DATAIN(4), ZN => n1386);
   U964 : INV_X1 port map( A => DATAIN(5), ZN => n1388);
   U965 : INV_X1 port map( A => DATAIN(6), ZN => n1390);
   U966 : INV_X1 port map( A => DATAIN(7), ZN => n1392);
   U967 : INV_X1 port map( A => DATAIN(8), ZN => n1394);
   U968 : INV_X1 port map( A => DATAIN(12), ZN => n1402);
   U969 : INV_X1 port map( A => DATAIN(13), ZN => n1404);
   U970 : INV_X1 port map( A => DATAIN(14), ZN => n1406);
   U971 : INV_X1 port map( A => DATAIN(15), ZN => n1408);
   U972 : INV_X1 port map( A => DATAIN(16), ZN => n1410);
   U973 : INV_X1 port map( A => DATAIN(17), ZN => n1412);
   U974 : INV_X1 port map( A => DATAIN(18), ZN => n1414);
   U975 : INV_X1 port map( A => DATAIN(19), ZN => n1416);
   U976 : INV_X1 port map( A => DATAIN(21), ZN => n1420);
   U977 : INV_X1 port map( A => DATAIN(22), ZN => n1422);
   U978 : INV_X1 port map( A => DATAIN(23), ZN => n1424);
   U979 : INV_X1 port map( A => DATAIN(25), ZN => n1430);
   U980 : INV_X1 port map( A => DATAIN(26), ZN => n1433);
   U981 : INV_X1 port map( A => DATAIN(27), ZN => n1436);
   U982 : INV_X1 port map( A => DATAIN(28), ZN => n1439);
   U983 : INV_X1 port map( A => DATAIN(29), ZN => n1442);
   U984 : INV_X1 port map( A => DATAIN(30), ZN => n1445);
   U985 : INV_X1 port map( A => DATAIN(31), ZN => n1448);
   U986 : INV_X1 port map( A => DATAIN(10), ZN => n1398);
   U987 : INV_X1 port map( A => DATAIN(20), ZN => n1418);
   U988 : INV_X1 port map( A => DATAIN(24), ZN => n1427);
   U989 : INV_X1 port map( A => DATAIN(11), ZN => n1400);
   U990 : INV_X1 port map( A => DATAIN(9), ZN => n1396);
   U991 : AOI221_X1 port map( B1 => n1268, B2 => n4280, C1 => n1265, C2 => 
                           n4248, A => n2440, ZN => n2444);
   U992 : AOI221_X1 port map( B1 => n1268, B2 => n4279, C1 => n1265, C2 => 
                           n4247, A => n2465, ZN => n2469);
   U993 : AOI221_X1 port map( B1 => n1268, B2 => n4282, C1 => n1265, C2 => 
                           n4250, A => n2390, ZN => n2394);
   U994 : NOR2_X1 port map( A1 => n819, A2 => n1149, ZN => n1007);
   U995 : NOR2_X1 port map( A1 => n1921, A2 => n1146, ZN => n1008);
   U996 : NOR2_X1 port map( A1 => n3738, A2 => n1143, ZN => n1009);
   U997 : NOR2_X1 port map( A1 => n815, A2 => n1149, ZN => n1010);
   U998 : NOR2_X1 port map( A1 => n2002, A2 => n1146, ZN => n1011);
   U999 : NOR2_X1 port map( A1 => n3838, A2 => n1143, ZN => n1012);
   U1000 : AND3_X1 port map( A1 => n3574, A2 => n3575, A3 => n3576, ZN => n1013
                           );
   U1001 : AND2_X1 port map( A1 => n1268, A2 => n4277, ZN => n1017);
   U1002 : AND2_X1 port map( A1 => n1265, A2 => n4245, ZN => n1018);
   U1003 : NOR3_X1 port map( A1 => n1017, A2 => n1018, A3 => n3571, ZN => n3575
                           );
   U1004 : OR2_X1 port map( A1 => n634, A2 => n1262, ZN => n1019);
   U1005 : OR2_X1 port map( A1 => n1261, A2 => n3570, ZN => n1020);
   U1006 : OR2_X1 port map( A1 => n590, A2 => n3569, ZN => n1021);
   U1007 : NAND3_X1 port map( A1 => n1019, A2 => n1020, A3 => n1021, ZN => 
                           n3571);
   U1008 : NOR3_X1 port map( A1 => n1092, A2 => n706, A3 => ADD_RS1(0), ZN => 
                           n1077);
   U1009 : AND3_X1 port map( A1 => n2494, A2 => n2493, A3 => n2495, ZN => n1022
                           );
   U1010 : BUF_X1 port map( A => n877, Z => n1023);
   U1011 : BUF_X1 port map( A => n877, Z => n1122);
   U1012 : AND2_X1 port map( A1 => n1268, A2 => n4284, ZN => n1025);
   U1013 : AND2_X1 port map( A1 => n1265, A2 => n4252, ZN => n1026);
   U1014 : NOR3_X1 port map( A1 => n1025, A2 => n1026, A3 => n2340, ZN => n2344
                           );
   U1015 : NOR3_X1 port map( A1 => n4656, A2 => n4645, A3 => n4657, ZN => n1027
                           );
   U1016 : AND2_X1 port map( A1 => n1155, A2 => n4873, ZN => n1032);
   U1017 : AND2_X1 port map( A1 => n1153, A2 => n3841, ZN => n1033);
   U1018 : OR2_X1 port map( A1 => n373, A2 => n1214, ZN => n1034);
   U1019 : OR2_X1 port map( A1 => n405, A2 => n1211, ZN => n1035);
   U1020 : NAND3_X1 port map( A1 => n1034, A2 => n1035, A3 => n3679, ZN => 
                           n3686);
   U1021 : AND2_X1 port map( A1 => n4866, A2 => n463, ZN => n1037);
   U1022 : AND2_X1 port map( A1 => n1241, A2 => n3666, ZN => n1038);
   U1023 : OR2_X1 port map( A1 => n1228, A2 => n457, ZN => n1039);
   U1024 : OR2_X1 port map( A1 => n1226, A2 => n458, ZN => n1040);
   U1025 : NAND3_X1 port map( A1 => n1039, A2 => n1040, A3 => n3633, ZN => 
                           n3634);
   U1026 : AND2_X1 port map( A1 => n4865, A2 => n463, ZN => n1041);
   U1027 : AND2_X1 port map( A1 => n1241, A2 => n3641, ZN => n1042);
   U1028 : AND2_X1 port map( A1 => n4864, A2 => n463, ZN => n1043);
   U1029 : AND2_X1 port map( A1 => n1241, A2 => n3616, ZN => n1044);
   U1030 : OR2_X1 port map( A1 => n1229, A2 => n459, ZN => n1045);
   U1031 : OR2_X1 port map( A1 => n1225, A2 => n460, ZN => n1046);
   U1032 : NAND3_X1 port map( A1 => n1045, A2 => n1046, A3 => n3583, ZN => 
                           n3584);
   U1033 : AND2_X1 port map( A1 => n4863, A2 => n1243, ZN => n1047);
   U1034 : AND2_X1 port map( A1 => n1240, A2 => n3591, ZN => n1048);
   U1035 : NAND2_X1 port map( A1 => n1013, A2 => n3577, ZN => n2548);
   U1036 : AND2_X1 port map( A1 => n1156, A2 => n4879, ZN => n1049);
   U1037 : AND2_X1 port map( A1 => n1153, A2 => n3995, ZN => n1050);
   U1038 : AND2_X1 port map( A1 => n1156, A2 => n4877, ZN => n1051);
   U1039 : AND2_X1 port map( A1 => n1151, A2 => n3943, ZN => n1052);
   U1040 : NAND2_X1 port map( A1 => n2496, A2 => n1022, ZN => n2547);
   U1041 : AND2_X1 port map( A1 => n4861, A2 => n1243, ZN => n1055);
   U1042 : AND2_X1 port map( A1 => n1240, A2 => n2485, ZN => n1056);
   U1043 : NOR3_X1 port map( A1 => n2484, A2 => n1056, A3 => n1055, ZN => n2496
                           );
   U1044 : AND2_X1 port map( A1 => n1155, A2 => n4860, ZN => n1057);
   U1045 : AND2_X1 port map( A1 => n1152, A2 => n2460, ZN => n1058);
   U1046 : AND2_X1 port map( A1 => n1154, A2 => n4859, ZN => n1059);
   U1047 : AND2_X1 port map( A1 => n1153, A2 => n2435, ZN => n1060);
   U1048 : INV_X1 port map( A => ADD_RS2(3), ZN => n1061);
   U1049 : INV_X1 port map( A => ADD_RS2(3), ZN => n1062);
   U1050 : NAND3_X1 port map( A1 => n790, A2 => n2471, A3 => n2469, ZN => n2546
                           );
   U1051 : AND2_X1 port map( A1 => n4860, A2 => n1243, ZN => n1063);
   U1052 : AND2_X1 port map( A1 => n1240, A2 => n2460, ZN => n1064);
   U1053 : AND2_X1 port map( A1 => n1154, A2 => n4858, ZN => n1065);
   U1054 : AND2_X1 port map( A1 => n1152, A2 => n2410, ZN => n1066);
   U1055 : AND2_X1 port map( A1 => n1154, A2 => n4871, ZN => n1067);
   U1056 : AND2_X1 port map( A1 => n1151, A2 => n3791, ZN => n1068);
   U1057 : NAND3_X1 port map( A1 => n2446, A2 => n791, A3 => n2444, ZN => n2545
                           );
   U1058 : AND2_X1 port map( A1 => n4859, A2 => n1243, ZN => n1069);
   U1059 : AND2_X1 port map( A1 => n1240, A2 => n2435, ZN => n1070);
   U1060 : AND2_X1 port map( A1 => n4858, A2 => n1243, ZN => n1071);
   U1061 : AND2_X1 port map( A1 => n1240, A2 => n2410, ZN => n1072);
   U1062 : OR2_X1 port map( A1 => n2376, A2 => n1134, ZN => n1073);
   U1063 : OR2_X1 port map( A1 => n255, A2 => n1132, ZN => n1074);
   U1064 : NAND3_X1 port map( A1 => n1073, A2 => n1074, A3 => n1664, ZN => 
                           n1669);
   U1065 : AND2_X1 port map( A1 => n1155, A2 => n4870, ZN => n1075);
   U1066 : AND2_X1 port map( A1 => n1152, A2 => n3766, ZN => n1076);
   U1067 : AND2_X1 port map( A1 => n1154, A2 => n4869, ZN => n1078);
   U1068 : AND2_X1 port map( A1 => n1152, A2 => n3741, ZN => n1079);
   U1069 : OR2_X1 port map( A1 => n1895, A2 => n1140, ZN => n1080);
   U1070 : OR2_X1 port map( A1 => n116, A2 => n1137, ZN => n1081);
   U1071 : NAND3_X1 port map( A1 => n1894, A2 => n1081, A3 => n1080, ZN => 
                           n1896);
   U1072 : AND2_X1 port map( A1 => n1154, A2 => n4868, ZN => n1082);
   U1073 : AND2_X1 port map( A1 => n1152, A2 => n3716, ZN => n1083);
   U1074 : NOR3_X1 port map( A1 => n1901, A2 => n1083, A3 => n1082, ZN => n1908
                           );
   U1075 : AND2_X1 port map( A1 => n1155, A2 => n4867, ZN => n1084);
   U1076 : AND2_X1 port map( A1 => n1153, A2 => n3691, ZN => n1085);
   U1077 : NOR3_X1 port map( A1 => n1880, A2 => n1085, A3 => n1084, ZN => n1887
                           );
   U1078 : AND2_X1 port map( A1 => n1154, A2 => n4855, ZN => n1086);
   U1079 : AND2_X1 port map( A1 => n1152, A2 => n2335, ZN => n1087);
   U1080 : OR2_X1 port map( A1 => n3657, A2 => n1134, ZN => n1088);
   U1081 : OR2_X1 port map( A1 => n1132, A2 => n246, ZN => n1089);
   U1082 : NAND3_X1 port map( A1 => n1088, A2 => n1089, A3 => n1852, ZN => 
                           n1857);
   U1083 : NAND3_X1 port map( A1 => n792, A2 => n2396, A3 => n2394, ZN => n2543
                           );
   U1084 : AND2_X1 port map( A1 => n1156, A2 => n4865, ZN => n1090);
   U1085 : AND2_X1 port map( A1 => n1151, A2 => n3641, ZN => n1091);
   U1086 : NOR3_X1 port map( A1 => n1840, A2 => n1091, A3 => n1090, ZN => n1847
                           );
   U1087 : OR2_X1 port map( A1 => n2301, A2 => n1134, ZN => n1093);
   U1088 : OR2_X1 port map( A1 => n258, A2 => n1132, ZN => n1094);
   U1089 : NAND3_X1 port map( A1 => n1093, A2 => n1094, A3 => n1603, ZN => 
                           n1607);
   U1090 : AND2_X1 port map( A1 => n4856, A2 => n1243, ZN => n1095);
   U1091 : AND2_X1 port map( A1 => n1240, A2 => n2360, ZN => n1096);
   U1092 : NAND2_X1 port map( A1 => n2346, A2 => n873, ZN => n2541);
   U1093 : AND2_X1 port map( A1 => n4855, A2 => n1243, ZN => n1097);
   U1094 : AND2_X1 port map( A1 => n1240, A2 => n2335, ZN => n1098);
   U1095 : NOR3_X1 port map( A1 => n2334, A2 => n1098, A3 => n1097, ZN => n2346
                           );
   U1096 : AND2_X1 port map( A1 => n1156, A2 => n4864, ZN => n1099);
   U1097 : AND2_X1 port map( A1 => n1153, A2 => n3616, ZN => n1100);
   U1098 : AND2_X1 port map( A1 => n1154, A2 => n4853, ZN => n1101);
   U1099 : AND2_X1 port map( A1 => n1153, A2 => n2285, ZN => n1102);
   U1100 : AND2_X1 port map( A1 => n4854, A2 => n1243, ZN => n1103);
   U1101 : AND2_X1 port map( A1 => n1240, A2 => n2310, ZN => n1104);
   U1102 : AND2_X1 port map( A1 => n1156, A2 => n4852, ZN => n1105);
   U1103 : AND2_X1 port map( A1 => n1151, A2 => n2256, ZN => n1106);
   U1104 : AND2_X1 port map( A1 => n4853, A2 => n1243, ZN => n1107);
   U1105 : AND2_X1 port map( A1 => n1240, A2 => n2285, ZN => n1108);
   U1106 : AND2_X1 port map( A1 => n4852, A2 => n1243, ZN => n1109);
   U1107 : AND2_X1 port map( A1 => n1240, A2 => n2256, ZN => n1110);
   U1108 : CLKBUF_X3 port map( A => n2200, Z => n1114);
   U1109 : CLKBUF_X3 port map( A => n2200, Z => n1115);
   U1110 : CLKBUF_X3 port map( A => n2200, Z => n1116);
   U1111 : CLKBUF_X3 port map( A => n2202, Z => n1117);
   U1112 : CLKBUF_X3 port map( A => n2202, Z => n1118);
   U1113 : CLKBUF_X3 port map( A => n2202, Z => n1119);
   U1114 : CLKBUF_X3 port map( A => n2204, Z => n1125);
   U1115 : CLKBUF_X3 port map( A => n2204, Z => n1126);
   U1116 : CLKBUF_X3 port map( A => n2205, Z => n1127);
   U1117 : CLKBUF_X3 port map( A => n2205, Z => n1128);
   U1118 : CLKBUF_X3 port map( A => n2208, Z => n1130);
   U1119 : CLKBUF_X3 port map( A => n2208, Z => n1131);
   U1120 : CLKBUF_X3 port map( A => n2209, Z => n1133);
   U1121 : CLKBUF_X3 port map( A => n2209, Z => n1135);
   U1122 : CLKBUF_X3 port map( A => n2213, Z => n1136);
   U1123 : CLKBUF_X3 port map( A => n2213, Z => n1137);
   U1124 : CLKBUF_X3 port map( A => n2214, Z => n1139);
   U1125 : CLKBUF_X3 port map( A => n2214, Z => n1140);
   U1126 : CLKBUF_X3 port map( A => n2221, Z => n1145);
   U1127 : CLKBUF_X3 port map( A => n2221, Z => n1146);
   U1128 : CLKBUF_X3 port map( A => n2223, Z => n1148);
   U1129 : CLKBUF_X3 port map( A => n2223, Z => n1149);
   U1130 : INV_X1 port map( A => n1378, ZN => n1377);
   U1131 : INV_X1 port map( A => n1380, ZN => n1379);
   U1132 : INV_X1 port map( A => n1382, ZN => n1381);
   U1133 : INV_X1 port map( A => n1384, ZN => n1383);
   U1134 : INV_X1 port map( A => n1386, ZN => n1385);
   U1135 : INV_X1 port map( A => n1388, ZN => n1387);
   U1136 : INV_X1 port map( A => n1390, ZN => n1389);
   U1137 : INV_X1 port map( A => n1392, ZN => n1391);
   U1138 : INV_X1 port map( A => n1394, ZN => n1393);
   U1139 : INV_X1 port map( A => n1396, ZN => n1395);
   U1140 : INV_X1 port map( A => n1398, ZN => n1397);
   U1141 : INV_X1 port map( A => n1400, ZN => n1399);
   U1142 : INV_X1 port map( A => n1402, ZN => n1401);
   U1143 : INV_X1 port map( A => n1404, ZN => n1403);
   U1144 : INV_X1 port map( A => n1406, ZN => n1405);
   U1145 : INV_X1 port map( A => n1408, ZN => n1407);
   U1146 : INV_X1 port map( A => n1410, ZN => n1409);
   U1147 : INV_X1 port map( A => n1412, ZN => n1411);
   U1148 : INV_X1 port map( A => n1414, ZN => n1413);
   U1149 : INV_X1 port map( A => n1416, ZN => n1415);
   U1150 : INV_X1 port map( A => n1418, ZN => n1417);
   U1151 : INV_X1 port map( A => n1420, ZN => n1419);
   U1152 : INV_X1 port map( A => n1422, ZN => n1421);
   U1153 : INV_X1 port map( A => n1424, ZN => n1423);
   U1154 : INV_X1 port map( A => n1427, ZN => n1425);
   U1155 : INV_X1 port map( A => n1427, ZN => n1426);
   U1156 : INV_X1 port map( A => n1430, ZN => n1428);
   U1157 : INV_X1 port map( A => n1430, ZN => n1429);
   U1158 : INV_X1 port map( A => n1433, ZN => n1431);
   U1159 : INV_X1 port map( A => n1433, ZN => n1432);
   U1160 : INV_X1 port map( A => n1436, ZN => n1434);
   U1161 : INV_X1 port map( A => n1436, ZN => n1435);
   U1162 : INV_X1 port map( A => n1439, ZN => n1437);
   U1163 : INV_X1 port map( A => n1439, ZN => n1438);
   U1164 : INV_X1 port map( A => n1442, ZN => n1440);
   U1165 : INV_X1 port map( A => n1442, ZN => n1441);
   U1166 : INV_X1 port map( A => n1445, ZN => n1443);
   U1167 : INV_X1 port map( A => n1445, ZN => n1444);
   U1168 : INV_X1 port map( A => n1448, ZN => n1446);
   U1169 : INV_X1 port map( A => n1448, ZN => n1447);
   U1170 : CLKBUF_X1 port map( A => n1552, Z => n1456);
   U1171 : CLKBUF_X1 port map( A => n1552, Z => n1457);
   U1172 : CLKBUF_X1 port map( A => n1552, Z => n1458);
   U1173 : CLKBUF_X1 port map( A => n1552, Z => n1459);
   U1174 : CLKBUF_X1 port map( A => n1552, Z => n1460);
   U1175 : CLKBUF_X1 port map( A => n1551, Z => n1461);
   U1176 : CLKBUF_X1 port map( A => n1551, Z => n1462);
   U1177 : CLKBUF_X1 port map( A => n1551, Z => n1463);
   U1178 : CLKBUF_X1 port map( A => n1551, Z => n1464);
   U1179 : CLKBUF_X1 port map( A => n1551, Z => n1465);
   U1180 : CLKBUF_X1 port map( A => n1551, Z => n1466);
   U1181 : CLKBUF_X1 port map( A => n1550, Z => n1467);
   U1182 : CLKBUF_X1 port map( A => n1550, Z => n1468);
   U1183 : CLKBUF_X1 port map( A => n1550, Z => n1469);
   U1184 : CLKBUF_X1 port map( A => n1550, Z => n1470);
   U1185 : CLKBUF_X1 port map( A => n1550, Z => n1471);
   U1186 : CLKBUF_X1 port map( A => n1550, Z => n1472);
   U1187 : CLKBUF_X1 port map( A => n1549, Z => n1473);
   U1188 : CLKBUF_X1 port map( A => n1549, Z => n1474);
   U1189 : CLKBUF_X1 port map( A => n1549, Z => n1475);
   U1190 : CLKBUF_X1 port map( A => n1549, Z => n1476);
   U1191 : CLKBUF_X1 port map( A => n1549, Z => n1477);
   U1192 : CLKBUF_X1 port map( A => n1549, Z => n1478);
   U1193 : CLKBUF_X1 port map( A => n1548, Z => n1479);
   U1194 : CLKBUF_X1 port map( A => n1548, Z => n1480);
   U1195 : CLKBUF_X1 port map( A => n1548, Z => n1481);
   U1196 : CLKBUF_X1 port map( A => n1548, Z => n1482);
   U1197 : CLKBUF_X1 port map( A => n1548, Z => n1483);
   U1198 : CLKBUF_X1 port map( A => n1548, Z => n1484);
   U1199 : CLKBUF_X1 port map( A => n1547, Z => n1485);
   U1200 : CLKBUF_X1 port map( A => n1547, Z => n1486);
   U1201 : CLKBUF_X1 port map( A => n1547, Z => n1487);
   U1202 : CLKBUF_X1 port map( A => n1547, Z => n1488);
   U1203 : CLKBUF_X1 port map( A => n1547, Z => n1489);
   U1204 : CLKBUF_X1 port map( A => n1547, Z => n1490);
   U1205 : CLKBUF_X1 port map( A => n1546, Z => n1491);
   U1206 : CLKBUF_X1 port map( A => n1546, Z => n1492);
   U1207 : CLKBUF_X1 port map( A => n1546, Z => n1493);
   U1208 : CLKBUF_X1 port map( A => n1546, Z => n1494);
   U1209 : CLKBUF_X1 port map( A => n1546, Z => n1495);
   U1210 : CLKBUF_X1 port map( A => n1546, Z => n1496);
   U1211 : CLKBUF_X1 port map( A => n1545, Z => n1497);
   U1212 : CLKBUF_X1 port map( A => n1545, Z => n1498);
   U1213 : CLKBUF_X1 port map( A => n1545, Z => n1499);
   U1214 : CLKBUF_X1 port map( A => n1545, Z => n1500);
   U1215 : CLKBUF_X1 port map( A => n1545, Z => n1501);
   U1216 : CLKBUF_X1 port map( A => n1545, Z => n1502);
   U1217 : CLKBUF_X1 port map( A => n1544, Z => n1503);
   U1218 : CLKBUF_X1 port map( A => n1544, Z => n1504);
   U1219 : CLKBUF_X1 port map( A => n1544, Z => n1505);
   U1220 : CLKBUF_X1 port map( A => n1544, Z => n1506);
   U1221 : CLKBUF_X1 port map( A => n1544, Z => n1507);
   U1222 : CLKBUF_X1 port map( A => n1544, Z => n1508);
   U1223 : CLKBUF_X1 port map( A => n1543, Z => n1509);
   U1224 : CLKBUF_X1 port map( A => n1543, Z => n1510);
   U1225 : CLKBUF_X1 port map( A => n1543, Z => n1511);
   U1226 : CLKBUF_X1 port map( A => n1543, Z => n1512);
   U1227 : CLKBUF_X1 port map( A => n1543, Z => n1513);
   U1228 : CLKBUF_X1 port map( A => n1543, Z => n1514);
   U1229 : CLKBUF_X1 port map( A => n1542, Z => n1515);
   U1230 : CLKBUF_X1 port map( A => n1542, Z => n1516);
   U1231 : CLKBUF_X1 port map( A => n1542, Z => n1517);
   U1232 : CLKBUF_X1 port map( A => n1542, Z => n1518);
   U1233 : CLKBUF_X1 port map( A => n1542, Z => n1519);
   U1234 : CLKBUF_X1 port map( A => n1542, Z => n1520);
   U1235 : CLKBUF_X1 port map( A => n1541, Z => n1521);
   U1236 : CLKBUF_X1 port map( A => n1541, Z => n1522);
   U1237 : CLKBUF_X1 port map( A => n1541, Z => n1523);
   U1238 : CLKBUF_X1 port map( A => n1541, Z => n1524);
   U1239 : CLKBUF_X1 port map( A => n1541, Z => n1525);
   U1240 : CLKBUF_X1 port map( A => n1541, Z => n1526);
   U1241 : CLKBUF_X1 port map( A => n1540, Z => n1527);
   U1242 : CLKBUF_X1 port map( A => n1540, Z => n1528);
   U1243 : CLKBUF_X1 port map( A => n1540, Z => n1529);
   U1244 : CLKBUF_X1 port map( A => n1540, Z => n1530);
   U1245 : CLKBUF_X1 port map( A => n1540, Z => n1531);
   U1246 : CLKBUF_X1 port map( A => n1540, Z => n1532);
   U1247 : CLKBUF_X1 port map( A => n1539, Z => n1533);
   U1248 : CLKBUF_X1 port map( A => n1539, Z => n1534);
   U1249 : CLKBUF_X1 port map( A => n1539, Z => n1535);
   U1250 : CLKBUF_X1 port map( A => n1539, Z => n1536);
   U1251 : CLKBUF_X1 port map( A => n1539, Z => n1537);
   U1252 : INV_X1 port map( A => ADD_RS1(2), ZN => n1554);
   U1253 : INV_X1 port map( A => n890, ZN => n1572);
   U1254 : NAND4_X1 port map( A1 => n930, A2 => n705, A3 => n1186, A4 => n875, 
                           ZN => n2223);
   U1255 : INV_X1 port map( A => ADD_RS1(4), ZN => n1560);
   U1256 : INV_X1 port map( A => ADD_RS1(1), ZN => n1553);
   U1257 : NAND2_X1 port map( A1 => n1015, A2 => n887, ZN => n2202);
   U1258 : NAND2_X1 port map( A1 => n1015, A2 => n705, ZN => n2200);
   U1259 : AOI22_X1 port map( A1 => n969, A2 => n4159, B1 => n739, B2 => n4724,
                           ZN => n1555);
   U1260 : OAI221_X1 port map( B1 => n164, B2 => n1117, C1 => n1556, C2 => 
                           n1115, A => n1555, ZN => n1568);
   U1261 : NAND2_X1 port map( A1 => n886, A2 => n171, ZN => n2205);
   U1262 : NAND2_X1 port map( A1 => n886, A2 => n468, ZN => n2204);
   U1263 : AOI22_X1 port map( A1 => n1124, A2 => n5044, B1 => n512, B2 => n5108
                           , ZN => n1557);
   U1264 : OAI221_X1 port map( B1 => n2246, B2 => n1129, C1 => n292, C2 => 
                           n1125, A => n1557, ZN => n1567);
   U1265 : NAND2_X1 port map( A1 => n1053, A2 => n171, ZN => n2209);
   U1266 : NAND2_X1 port map( A1 => n1053, A2 => n468, ZN => n2208);
   U1267 : AOI22_X1 port map( A1 => n56, A2 => n5076, B1 => n760, B2 => n1558, 
                           ZN => n1559);
   U1268 : OAI221_X1 port map( B1 => n2247, B2 => n1135, C1 => n260, C2 => 
                           n1130, A => n1559, ZN => n1566);
   U1269 : NAND2_X1 port map( A1 => n1031, A2 => n171, ZN => n2214);
   U1270 : NAND2_X1 port map( A1 => n1031, A2 => n887, ZN => n2213);
   U1271 : NAND2_X1 port map( A1 => n1031, A2 => n705, ZN => n1561);
   U1272 : INV_X1 port map( A => n1561, ZN => n2211);
   U1273 : AOI22_X1 port map( A1 => n1014, A2 => n5204, B1 => n489, B2 => n1562
                           , ZN => n1563);
   U1274 : OAI221_X1 port map( B1 => n1564, B2 => n1139, C1 => n132, C2 => 
                           n1136, A => n1563, ZN => n1565);
   U1275 : NOR4_X1 port map( A1 => n1568, A2 => n1567, A3 => n1565, A4 => n1566
                           , ZN => n1569);
   U1276 : NAND2_X1 port map( A1 => n1574, A2 => n1187, ZN => n2221);
   U1277 : NAND4_X1 port map( A1 => n874, A2 => n468, A3 => n1186, A4 => n930, 
                           ZN => n2220);
   U1278 : OAI222_X1 port map( A1 => n836, A2 => n1148, B1 => n1569, B2 => 
                           n1145, C1 => n2253, C2 => n1142, ZN => n1570);
   U1279 : NAND4_X1 port map( A1 => n875, A2 => n887, A3 => n1186, A4 => n930, 
                           ZN => n2226);
   U1280 : NAND4_X1 port map( A1 => n874, A2 => n171, A3 => n1186, A4 => n930, 
                           ZN => n2225);
   U1281 : OAI22_X1 port map( A1 => n2257, A2 => n707, B1 => n964, B2 => n1157,
                           ZN => n1571);
   U1282 : AOI221_X1 port map( B1 => n1166, B2 => n4788, C1 => n1163, C2 => 
                           n4339, A => n1571, ZN => n1578);
   U1283 : NAND4_X1 port map( A1 => n1574, A2 => n887, A3 => n1186, A4 => n971,
                           ZN => n2230);
   U1284 : NAND4_X1 port map( A1 => n874, A2 => n171, A3 => n1186, A4 => n971, 
                           ZN => n2229);
   U1285 : NAND4_X1 port map( A1 => n874, A2 => n705, A3 => n1187, A4 => n978, 
                           ZN => n2228);
   U1286 : NAND3_X1 port map( A1 => n1187, A2 => n78, A3 => n690, ZN => n2232);
   U1287 : OAI22_X1 port map( A1 => n4660, A2 => n1187, B1 => n1378, B2 => 
                           n1183, ZN => n1575);
   U1288 : AOI221_X1 port map( B1 => n1193, B2 => n4948, C1 => n1190, C2 => 
                           n2267, A => n1575, ZN => n1576);
   U1289 : NAND4_X1 port map( A1 => n1579, A2 => n1577, A3 => n1576, A4 => 
                           n1578, ZN => n2506);
   U1290 : AOI22_X1 port map( A1 => n969, A2 => n4158, B1 => n486, B2 => n4725,
                           ZN => n1580);
   U1291 : OAI221_X1 port map( B1 => n163, B2 => n1118, C1 => n1581, C2 => 
                           n1115, A => n1580, ZN => n1591);
   U1292 : AOI22_X1 port map( A1 => n1122, A2 => n5045, B1 => n493, B2 => n5109
                           , ZN => n1582);
   U1293 : OAI221_X1 port map( B1 => n2275, B2 => n1127, C1 => n291, C2 => 
                           n1125, A => n1582, ZN => n1590);
   U1294 : AOI22_X1 port map( A1 => n54, A2 => n5077, B1 => n759, B2 => n1583, 
                           ZN => n1584);
   U1295 : OAI221_X1 port map( B1 => n2276, B2 => n1133, C1 => n259, C2 => 
                           n1130, A => n1584, ZN => n1589);
   U1296 : AOI22_X1 port map( A1 => n1014, A2 => n5205, B1 => n966, B2 => n1585
                           , ZN => n1586);
   U1297 : NOR4_X1 port map( A1 => n1591, A2 => n1589, A3 => n1590, A4 => n1588
                           , ZN => n1592);
   U1298 : OAI22_X1 port map( A1 => n2286, A2 => n1161, B1 => n963, B2 => n1157
                           , ZN => n1593);
   U1299 : AOI221_X1 port map( B1 => n1166, B2 => n4789, C1 => n1163, C2 => 
                           n4338, A => n1593, ZN => n1598);
   U1300 : OAI22_X1 port map( A1 => n4661, A2 => n1189, B1 => n1380, B2 => 
                           n1183, ZN => n1595);
   U1301 : AOI221_X1 port map( B1 => n1193, B2 => n4949, C1 => n1190, C2 => 
                           n2292, A => n1595, ZN => n1596);
   U1302 : NAND4_X1 port map( A1 => n1599, A2 => n1597, A3 => n1596, A4 => 
                           n1598, ZN => n2507);
   U1303 : AOI22_X1 port map( A1 => n969, A2 => n4157, B1 => n486, B2 => n4726,
                           ZN => n1600);
   U1304 : OAI221_X1 port map( B1 => n162, B2 => n1118, C1 => n1601, C2 => 
                           n1115, A => n1600, ZN => n1609);
   U1305 : AOI22_X1 port map( A1 => n1123, A2 => n5046, B1 => n493, B2 => n5110
                           , ZN => n1602);
   U1306 : OAI221_X1 port map( B1 => n2300, B2 => n1127, C1 => n290, C2 => 
                           n1125, A => n1602, ZN => n1608);
   U1307 : AOI22_X1 port map( A1 => n56, A2 => n5078, B1 => n1029, B2 => n218, 
                           ZN => n1603);
   U1308 : AOI22_X1 port map( A1 => n888, A2 => n5206, B1 => n579, B2 => n219, 
                           ZN => n1604);
   U1309 : NOR4_X1 port map( A1 => n1609, A2 => n1608, A3 => n1606, A4 => n1607
                           , ZN => n1610);
   U1310 : OAI222_X1 port map( A1 => n834, A2 => n1148, B1 => n1610, B2 => 
                           n1145, C1 => n2307, C2 => n1142, ZN => n1611);
   U1311 : OAI22_X1 port map( A1 => n2311, A2 => n1160, B1 => n962, B2 => n1157
                           , ZN => n1612);
   U1312 : AOI221_X1 port map( B1 => n1166, B2 => n4790, C1 => n1163, C2 => 
                           n4337, A => n1612, ZN => n1617);
   U1313 : OAI222_X1 port map( A1 => n642, A2 => n1175, B1 => n2314, B2 => 
                           n1173, C1 => n2313, C2 => n1169, ZN => n1613);
   U1314 : AOI221_X1 port map( B1 => n1180, B2 => n4285, C1 => n1177, C2 => 
                           n4253, A => n1613, ZN => n1616);
   U1315 : OAI22_X1 port map( A1 => n4662, A2 => n1189, B1 => n1382, B2 => 
                           n1183, ZN => n1614);
   U1316 : AOI221_X1 port map( B1 => n1193, B2 => n4950, C1 => n1190, C2 => 
                           n2317, A => n1614, ZN => n1615);
   U1317 : NAND4_X1 port map( A1 => n1618, A2 => n1615, A3 => n1617, A4 => 
                           n1616, ZN => n2508);
   U1318 : AOI22_X1 port map( A1 => n969, A2 => n4156, B1 => n738, B2 => n4727,
                           ZN => n1619);
   U1319 : AOI22_X1 port map( A1 => n1122, A2 => n5047, B1 => n493, B2 => n5111
                           , ZN => n1621);
   U1320 : OAI221_X1 port map( B1 => n2325, B2 => n1127, C1 => n289, C2 => 
                           n1125, A => n1621, ZN => n1629);
   U1321 : AOI22_X1 port map( A1 => n56, A2 => n5079, B1 => n760, B2 => n1622, 
                           ZN => n1623);
   U1322 : OAI221_X1 port map( B1 => n507, B2 => n2326, C1 => n257, C2 => n1131
                           , A => n1623, ZN => n1628);
   U1323 : AOI22_X1 port map( A1 => n888, A2 => n5207, B1 => n966, B2 => n1624,
                           ZN => n1625);
   U1324 : OAI221_X1 port map( B1 => n1626, B2 => n1139, C1 => n129, C2 => 
                           n1136, A => n1625, ZN => n1627);
   U1325 : NOR4_X1 port map( A1 => n1630, A2 => n1628, A3 => n1629, A4 => n1627
                           , ZN => n1631);
   U1326 : OAI22_X1 port map( A1 => n2336, A2 => n707, B1 => n961, B2 => n1157,
                           ZN => n1632);
   U1327 : OAI222_X1 port map( A1 => n641, A2 => n1175, B1 => n2339, B2 => 
                           n1173, C1 => n2338, C2 => n1169, ZN => n1633);
   U1328 : AOI221_X1 port map( B1 => n1180, B2 => n4284, C1 => n1177, C2 => 
                           n4252, A => n1633, ZN => n1636);
   U1329 : OAI22_X1 port map( A1 => n4663, A2 => n1189, B1 => n1384, B2 => 
                           n1183, ZN => n1634);
   U1330 : AOI221_X1 port map( B1 => n1193, B2 => n4951, C1 => n1190, C2 => 
                           n2342, A => n1634, ZN => n1635);
   U1331 : NAND4_X1 port map( A1 => n1636, A2 => n1637, A3 => n1638, A4 => 
                           n1635, ZN => n2509);
   U1332 : AOI22_X1 port map( A1 => n669, A2 => n4155, B1 => n1111, B2 => n4728
                           , ZN => n1639);
   U1333 : OAI221_X1 port map( B1 => n160, B2 => n1118, C1 => n1640, C2 => 
                           n1114, A => n1639, ZN => n1650);
   U1334 : AOI22_X1 port map( A1 => n1122, A2 => n5048, B1 => n493, B2 => n5112
                           , ZN => n1641);
   U1335 : OAI221_X1 port map( B1 => n2350, B2 => n1129, C1 => n288, C2 => 
                           n1125, A => n1641, ZN => n1649);
   U1336 : AOI22_X1 port map( A1 => n55, A2 => n5080, B1 => n759, B2 => n1642, 
                           ZN => n1643);
   U1337 : OAI221_X1 port map( B1 => n1133, B2 => n2351, C1 => n256, C2 => 
                           n1131, A => n1643, ZN => n1648);
   U1338 : AOI22_X1 port map( A1 => n1014, A2 => n5208, B1 => n966, B2 => n1644
                           , ZN => n1645);
   U1339 : NOR4_X1 port map( A1 => n1650, A2 => n1648, A3 => n1649, A4 => n1647
                           , ZN => n1651);
   U1340 : OAI22_X1 port map( A1 => n2361, A2 => n707, B1 => n960, B2 => n1157,
                           ZN => n1653);
   U1341 : AOI221_X1 port map( B1 => n1166, B2 => n4792, C1 => n1163, C2 => 
                           n4335, A => n1653, ZN => n1658);
   U1342 : OAI222_X1 port map( A1 => n640, A2 => n1176, B1 => n2364, B2 => 
                           n1173, C1 => n2363, C2 => n1169, ZN => n1654);
   U1343 : AOI221_X1 port map( B1 => n1180, B2 => n4283, C1 => n1177, C2 => 
                           n4251, A => n1654, ZN => n1657);
   U1344 : OAI22_X1 port map( A1 => n4664, A2 => n1189, B1 => n1386, B2 => 
                           n1183, ZN => n1655);
   U1345 : AOI221_X1 port map( B1 => n1193, B2 => n4952, C1 => n1190, C2 => 
                           n2367, A => n1655, ZN => n1656);
   U1346 : NAND4_X1 port map( A1 => n1657, A2 => n1659, A3 => n1656, A4 => 
                           n1658, ZN => n2510);
   U1347 : AOI22_X1 port map( A1 => n668, A2 => n4154, B1 => n739, B2 => n4729,
                           ZN => n1660);
   U1348 : OAI221_X1 port map( B1 => n159, B2 => n1119, C1 => n1661, C2 => 
                           n1114, A => n1660, ZN => n1671);
   U1349 : AOI22_X1 port map( A1 => n1023, A2 => n5049, B1 => n52, B2 => n5113,
                           ZN => n1662);
   U1350 : OAI221_X1 port map( B1 => n2375, B2 => n1128, C1 => n287, C2 => 
                           n1125, A => n1662, ZN => n1670);
   U1351 : AOI22_X1 port map( A1 => n56, A2 => n5081, B1 => n1029, B2 => n1663,
                           ZN => n1664);
   U1352 : AOI22_X1 port map( A1 => n2211, A2 => n5209, B1 => n966, B2 => n1665
                           , ZN => n1666);
   U1353 : OAI221_X1 port map( B1 => n1667, B2 => n1139, C1 => n127, C2 => 
                           n1136, A => n1666, ZN => n1668);
   U1354 : NOR4_X1 port map( A1 => n1671, A2 => n1670, A3 => n1668, A4 => n1669
                           , ZN => n1672);
   U1355 : OAI22_X1 port map( A1 => n2386, A2 => n1161, B1 => n959, B2 => n1157
                           , ZN => n1674);
   U1356 : AOI221_X1 port map( B1 => n1166, B2 => n4793, C1 => n1163, C2 => 
                           n4334, A => n1674, ZN => n1679);
   U1357 : OAI222_X1 port map( A1 => n639, A2 => n1175, B1 => n2389, B2 => 
                           n1173, C1 => n2388, C2 => n1169, ZN => n1675);
   U1358 : AOI221_X1 port map( B1 => n1180, B2 => n4282, C1 => n1177, C2 => 
                           n4250, A => n1675, ZN => n1678);
   U1359 : OAI22_X1 port map( A1 => n4665, A2 => n1189, B1 => n1388, B2 => 
                           n1183, ZN => n1676);
   U1360 : AOI221_X1 port map( B1 => n1193, B2 => n4953, C1 => n1190, C2 => 
                           n2392, A => n1676, ZN => n1677);
   U1361 : NAND4_X1 port map( A1 => n1678, A2 => n1680, A3 => n1677, A4 => 
                           n1679, ZN => n2511);
   U1362 : AOI22_X1 port map( A1 => n969, A2 => n4153, B1 => n738, B2 => n4730,
                           ZN => n1681);
   U1363 : OAI221_X1 port map( B1 => n158, B2 => n1117, C1 => n1682, C2 => 
                           n1114, A => n1681, ZN => n1692);
   U1364 : AOI22_X1 port map( A1 => n1024, A2 => n5050, B1 => n1120, B2 => 
                           n5114, ZN => n1683);
   U1365 : OAI221_X1 port map( B1 => n2400, B2 => n1129, C1 => n286, C2 => 
                           n1125, A => n1683, ZN => n1691);
   U1366 : AOI22_X1 port map( A1 => n57, A2 => n5082, B1 => n759, B2 => n1684, 
                           ZN => n1685);
   U1367 : OAI221_X1 port map( B1 => n2401, B2 => n1135, C1 => n254, C2 => 
                           n1130, A => n1685, ZN => n1690);
   U1368 : AOI22_X1 port map( A1 => n888, A2 => n5210, B1 => n966, B2 => n1686,
                           ZN => n1687);
   U1369 : OAI221_X1 port map( B1 => n1688, B2 => n1139, C1 => n126, C2 => 
                           n1136, A => n1687, ZN => n1689);
   U1370 : NOR4_X1 port map( A1 => n1692, A2 => n1691, A3 => n1690, A4 => n1689
                           , ZN => n1693);
   U1371 : OAI222_X1 port map( A1 => n830, A2 => n1148, B1 => n1693, B2 => 
                           n1145, C1 => n2407, C2 => n1142, ZN => n1694);
   U1372 : OAI22_X1 port map( A1 => n2411, A2 => n1161, B1 => n958, B2 => n1157
                           , ZN => n1695);
   U1373 : AOI221_X1 port map( B1 => n1166, B2 => n4794, C1 => n1163, C2 => 
                           n4333, A => n1695, ZN => n1700);
   U1374 : OAI222_X1 port map( A1 => n638, A2 => n1174, B1 => n1171, B2 => 
                           n2414, C1 => n2413, C2 => n1169, ZN => n1696);
   U1375 : AOI221_X1 port map( B1 => n1180, B2 => n4281, C1 => n1177, C2 => 
                           n4249, A => n1696, ZN => n1699);
   U1376 : OAI22_X1 port map( A1 => n4666, A2 => n1189, B1 => n1390, B2 => 
                           n1183, ZN => n1697);
   U1377 : AOI221_X1 port map( B1 => n1193, B2 => n4954, C1 => n1190, C2 => 
                           n2417, A => n1697, ZN => n1698);
   U1378 : NAND4_X1 port map( A1 => n1699, A2 => n1701, A3 => n1700, A4 => 
                           n1698, ZN => n2512);
   U1379 : AOI22_X1 port map( A1 => n669, A2 => n4152, B1 => n738, B2 => n4731,
                           ZN => n1702);
   U1380 : OAI221_X1 port map( B1 => n157, B2 => n1118, C1 => n1703, C2 => 
                           n1114, A => n1702, ZN => n1713);
   U1381 : AOI22_X1 port map( A1 => n1024, A2 => n5051, B1 => n508, B2 => n5115
                           , ZN => n1704);
   U1382 : OAI221_X1 port map( B1 => n2425, B2 => n1129, C1 => n285, C2 => 
                           n1125, A => n1704, ZN => n1712);
   U1383 : AOI22_X1 port map( A1 => n54, A2 => n5083, B1 => n1029, B2 => n1705,
                           ZN => n1706);
   U1384 : OAI221_X1 port map( B1 => n2426, B2 => n1133, C1 => n253, C2 => n506
                           , A => n1706, ZN => n1711);
   U1385 : AOI22_X1 port map( A1 => n888, A2 => n5211, B1 => n578, B2 => n1707,
                           ZN => n1708);
   U1386 : NOR4_X1 port map( A1 => n1713, A2 => n1712, A3 => n1710, A4 => n1711
                           , ZN => n1714);
   U1387 : OAI222_X1 port map( A1 => n829, A2 => n1148, B1 => n1714, B2 => 
                           n1145, C1 => n2432, C2 => n1142, ZN => n1715);
   U1388 : OAI22_X1 port map( A1 => n2436, A2 => n1162, B1 => n957, B2 => n1157
                           , ZN => n1716);
   U1389 : AOI221_X1 port map( B1 => n1166, B2 => n4795, C1 => n1163, C2 => 
                           n4332, A => n1716, ZN => n1721);
   U1390 : OAI222_X1 port map( A1 => n637, A2 => n1174, B1 => n1171, B2 => 
                           n2439, C1 => n2438, C2 => n1169, ZN => n1717);
   U1391 : AOI221_X1 port map( B1 => n1180, B2 => n4280, C1 => n1177, C2 => 
                           n4248, A => n1717, ZN => n1720);
   U1392 : OAI22_X1 port map( A1 => n4667, A2 => n1189, B1 => n1392, B2 => 
                           n1183, ZN => n1718);
   U1393 : AOI221_X1 port map( B1 => n1193, B2 => n4955, C1 => n1190, C2 => 
                           n2442, A => n1718, ZN => n1719);
   U1394 : NAND4_X1 port map( A1 => n1722, A2 => n1721, A3 => n1719, A4 => 
                           n1720, ZN => n2513);
   U1395 : AOI22_X1 port map( A1 => n669, A2 => n4151, B1 => n739, B2 => n4732,
                           ZN => n1723);
   U1396 : OAI221_X1 port map( B1 => n156, B2 => n1118, C1 => n1724, C2 => 
                           n1116, A => n1723, ZN => n1734);
   U1397 : AOI22_X1 port map( A1 => n1123, A2 => n5052, B1 => n52, B2 => n5116,
                           ZN => n1725);
   U1398 : OAI221_X1 port map( B1 => n2450, B2 => n1128, C1 => n284, C2 => 
                           n1125, A => n1725, ZN => n1733);
   U1399 : AOI22_X1 port map( A1 => n54, A2 => n5084, B1 => n760, B2 => n1726, 
                           ZN => n1727);
   U1400 : OAI221_X1 port map( B1 => n2451, B2 => n1135, C1 => n252, C2 => 
                           n1130, A => n1727, ZN => n1732);
   U1401 : AOI22_X1 port map( A1 => n1014, A2 => n5212, B1 => n577, B2 => n1728
                           , ZN => n1729);
   U1402 : NOR4_X1 port map( A1 => n1734, A2 => n1733, A3 => n1731, A4 => n1732
                           , ZN => n1735);
   U1403 : OAI222_X1 port map( A1 => n828, A2 => n1148, B1 => n1735, B2 => 
                           n1145, C1 => n2457, C2 => n1142, ZN => n1736);
   U1404 : OAI22_X1 port map( A1 => n2461, A2 => n707, B1 => n956, B2 => n1157,
                           ZN => n1737);
   U1405 : AOI221_X1 port map( B1 => n1166, B2 => n4796, C1 => n1163, C2 => 
                           n4331, A => n1737, ZN => n1742);
   U1406 : OAI222_X1 port map( A1 => n636, A2 => n1175, B1 => n2464, B2 => 
                           n1172, C1 => n2463, C2 => n1169, ZN => n1738);
   U1407 : AOI221_X1 port map( B1 => n1180, B2 => n4279, C1 => n1177, C2 => 
                           n4247, A => n1738, ZN => n1741);
   U1408 : OAI22_X1 port map( A1 => n4668, A2 => n1189, B1 => n1394, B2 => 
                           n1183, ZN => n1739);
   U1409 : AOI221_X1 port map( B1 => n1193, B2 => n4956, C1 => n1190, C2 => 
                           n2467, A => n1739, ZN => n1740);
   U1410 : NAND4_X1 port map( A1 => n1743, A2 => n1742, A3 => n1740, A4 => 
                           n1741, ZN => n2514);
   U1411 : AOI22_X1 port map( A1 => n969, A2 => n4150, B1 => n739, B2 => n4733,
                           ZN => n1744);
   U1412 : OAI221_X1 port map( B1 => n155, B2 => n1118, C1 => n1745, C2 => 
                           n1116, A => n1744, ZN => n1755);
   U1413 : AOI22_X1 port map( A1 => n1016, A2 => n5053, B1 => n1121, B2 => 
                           n5117, ZN => n1746);
   U1414 : AOI22_X1 port map( A1 => n54, A2 => n5085, B1 => n760, B2 => n1747, 
                           ZN => n1748);
   U1415 : OAI221_X1 port map( B1 => n2476, B2 => n1133, C1 => n251, C2 => 
                           n1131, A => n1748, ZN => n1753);
   U1416 : AOI22_X1 port map( A1 => n888, A2 => n5213, B1 => n578, B2 => n1749,
                           ZN => n1750);
   U1417 : OAI221_X1 port map( B1 => n1751, B2 => n1139, C1 => n123, C2 => 
                           n1136, A => n1750, ZN => n1752);
   U1418 : NOR4_X1 port map( A1 => n1755, A2 => n1752, A3 => n1753, A4 => n1754
                           , ZN => n1756);
   U1419 : OAI222_X1 port map( A1 => n827, A2 => n1148, B1 => n1756, B2 => 
                           n1145, C1 => n2482, C2 => n1142, ZN => n1757);
   U1420 : OAI22_X1 port map( A1 => n2486, A2 => n1161, B1 => n955, B2 => n1157
                           , ZN => n1758);
   U1421 : AOI221_X1 port map( B1 => n1166, B2 => n4797, C1 => n1163, C2 => 
                           n4330, A => n1758, ZN => n1763);
   U1422 : OAI222_X1 port map( A1 => n635, A2 => n1176, B1 => n2489, B2 => 
                           n1173, C1 => n2488, C2 => n1169, ZN => n1759);
   U1423 : AOI221_X1 port map( B1 => n1180, B2 => n4278, C1 => n1177, C2 => 
                           n4246, A => n1759, ZN => n1762);
   U1424 : OAI22_X1 port map( A1 => n4669, A2 => n1189, B1 => n1396, B2 => 
                           n1183, ZN => n1760);
   U1425 : AOI221_X1 port map( B1 => n1193, B2 => n4957, C1 => n1190, C2 => 
                           n2492, A => n1760, ZN => n1761);
   U1426 : NAND4_X1 port map( A1 => n1762, A2 => n1761, A3 => n1763, A4 => 
                           n1764, ZN => n2515);
   U1427 : AOI22_X1 port map( A1 => n669, A2 => n4149, B1 => n487, B2 => n4734,
                           ZN => n1765);
   U1428 : OAI221_X1 port map( B1 => n154, B2 => n1118, C1 => n1766, C2 => 
                           n1115, A => n1765, ZN => n1776);
   U1429 : AOI22_X1 port map( A1 => n1016, A2 => n5054, B1 => n1121, B2 => 
                           n5118, ZN => n1767);
   U1430 : OAI221_X1 port map( B1 => n2500, B2 => n1128, C1 => n282, C2 => 
                           n1125, A => n1767, ZN => n1775);
   U1431 : AOI22_X1 port map( A1 => n54, A2 => n5086, B1 => n759, B2 => n1768, 
                           ZN => n1769);
   U1432 : OAI221_X1 port map( B1 => n2501, B2 => n1135, C1 => n250, C2 => 
                           n1130, A => n1769, ZN => n1774);
   U1433 : AOI22_X1 port map( A1 => n888, A2 => n5214, B1 => n966, B2 => n1770,
                           ZN => n1771);
   U1434 : OAI221_X1 port map( B1 => n1772, B2 => n1139, C1 => n122, C2 => 
                           n1136, A => n1771, ZN => n1773);
   U1435 : NOR4_X1 port map( A1 => n1776, A2 => n1775, A3 => n1774, A4 => n1773
                           , ZN => n1777);
   U1436 : OAI222_X1 port map( A1 => n826, A2 => n1148, B1 => n1777, B2 => 
                           n1145, C1 => n3563, C2 => n1142, ZN => n1778);
   U1437 : OAI22_X1 port map( A1 => n3567, A2 => n1161, B1 => n954, B2 => n1157
                           , ZN => n1779);
   U1438 : AOI221_X1 port map( B1 => n1166, B2 => n4798, C1 => n1163, C2 => 
                           n4329, A => n1779, ZN => n1784);
   U1439 : OAI222_X1 port map( A1 => n634, A2 => n1174, B1 => n3570, B2 => 
                           n1173, C1 => n3569, C2 => n1170, ZN => n1780);
   U1440 : AOI221_X1 port map( B1 => n1180, B2 => n4277, C1 => n1177, C2 => 
                           n4245, A => n1780, ZN => n1783);
   U1441 : OAI22_X1 port map( A1 => n4670, A2 => n1189, B1 => n1398, B2 => 
                           n1183, ZN => n1781);
   U1442 : AOI221_X1 port map( B1 => n1193, B2 => n4958, C1 => n1190, C2 => 
                           n3573, A => n1781, ZN => n1782);
   U1443 : NAND4_X1 port map( A1 => n1783, A2 => n1782, A3 => n1784, A4 => 
                           n1785, ZN => n2516);
   U1444 : AOI22_X1 port map( A1 => n969, A2 => n4148, B1 => n497, B2 => n4735,
                           ZN => n1786);
   U1445 : OAI221_X1 port map( B1 => n153, B2 => n1118, C1 => n1787, C2 => 
                           n1114, A => n1786, ZN => n1797);
   U1446 : AOI22_X1 port map( A1 => n1024, A2 => n5055, B1 => n493, B2 => n5119
                           , ZN => n1788);
   U1447 : AOI22_X1 port map( A1 => n55, A2 => n5087, B1 => n1029, B2 => n1789,
                           ZN => n1790);
   U1448 : OAI221_X1 port map( B1 => n3582, B2 => n1133, C1 => n249, C2 => 
                           n1130, A => n1790, ZN => n1795);
   U1449 : AOI22_X1 port map( A1 => n1014, A2 => n5215, B1 => n579, B2 => n1791
                           , ZN => n1792);
   U1450 : OAI221_X1 port map( B1 => n1793, B2 => n1139, C1 => n121, C2 => 
                           n1136, A => n1792, ZN => n1794);
   U1451 : NOR4_X1 port map( A1 => n1797, A2 => n1794, A3 => n1796, A4 => n1795
                           , ZN => n1798);
   U1452 : OAI222_X1 port map( A1 => n825, A2 => n1148, B1 => n1798, B2 => 
                           n1145, C1 => n3588, C2 => n1142, ZN => n1799);
   U1453 : OAI22_X1 port map( A1 => n3592, A2 => n1162, B1 => n953, B2 => n1157
                           , ZN => n1800);
   U1454 : AOI221_X1 port map( B1 => n1166, B2 => n4799, C1 => n1163, C2 => 
                           n4328, A => n1800, ZN => n1805);
   U1455 : OAI222_X1 port map( A1 => n633, A2 => n1175, B1 => n3595, B2 => 
                           n1172, C1 => n3594, C2 => n1170, ZN => n1801);
   U1456 : AOI221_X1 port map( B1 => n1180, B2 => n4276, C1 => n1177, C2 => 
                           n4244, A => n1801, ZN => n1804);
   U1457 : OAI22_X1 port map( A1 => n4671, A2 => n1189, B1 => n1400, B2 => 
                           n1183, ZN => n1802);
   U1458 : AOI221_X1 port map( B1 => n1193, B2 => n4959, C1 => n1190, C2 => 
                           n3598, A => n1802, ZN => n1803);
   U1459 : NAND4_X1 port map( A1 => n1804, A2 => n1806, A3 => n1803, A4 => 
                           n1805, ZN => n2517);
   U1460 : AOI22_X1 port map( A1 => n668, A2 => n4147, B1 => n691, B2 => n4736,
                           ZN => n1807);
   U1461 : OAI221_X1 port map( B1 => n152, B2 => n1119, C1 => n1808, C2 => 
                           n1114, A => n1807, ZN => n1818);
   U1462 : AOI22_X1 port map( A1 => n1124, A2 => n5056, B1 => n493, B2 => n5120
                           , ZN => n1809);
   U1463 : AOI22_X1 port map( A1 => n54, A2 => n5088, B1 => n759, B2 => n1810, 
                           ZN => n1811);
   U1464 : OAI221_X1 port map( B1 => n507, B2 => n3607, C1 => n248, C2 => n1131
                           , A => n1811, ZN => n1816);
   U1465 : AOI22_X1 port map( A1 => n888, A2 => n5216, B1 => n966, B2 => n1812,
                           ZN => n1813);
   U1466 : OAI221_X1 port map( B1 => n1814, B2 => n1140, C1 => n120, C2 => 
                           n1137, A => n1813, ZN => n1815);
   U1467 : NOR4_X1 port map( A1 => n1818, A2 => n1816, A3 => n1817, A4 => n1815
                           , ZN => n1819);
   U1468 : OAI22_X1 port map( A1 => n3617, A2 => n707, B1 => n952, B2 => n1158,
                           ZN => n1820);
   U1469 : AOI221_X1 port map( B1 => n1167, B2 => n4800, C1 => n1164, C2 => 
                           n4327, A => n1820, ZN => n1825);
   U1470 : OAI222_X1 port map( A1 => n632, A2 => n1176, B1 => n3620, B2 => 
                           n1171, C1 => n3619, C2 => n1170, ZN => n1821);
   U1471 : AOI221_X1 port map( B1 => n1181, B2 => n4275, C1 => n1178, C2 => 
                           n4243, A => n1821, ZN => n1824);
   U1472 : OAI22_X1 port map( A1 => n4672, A2 => n1189, B1 => n1402, B2 => 
                           n1184, ZN => n1822);
   U1473 : AOI221_X1 port map( B1 => n1194, B2 => n4960, C1 => n1191, C2 => 
                           n3623, A => n1822, ZN => n1823);
   U1474 : NAND4_X1 port map( A1 => n1824, A2 => n1825, A3 => n1826, A4 => 
                           n1823, ZN => n2518);
   U1475 : AOI22_X1 port map( A1 => n969, A2 => n4146, B1 => n1111, B2 => n4737
                           , ZN => n1827);
   U1476 : OAI221_X1 port map( B1 => n151, B2 => n1117, C1 => n1828, C2 => 
                           n1115, A => n1827, ZN => n1838);
   U1477 : AOI22_X1 port map( A1 => n1124, A2 => n5057, B1 => n52, B2 => n5121,
                           ZN => n1829);
   U1478 : AOI22_X1 port map( A1 => n56, A2 => n5089, B1 => n1029, B2 => n1830,
                           ZN => n1831);
   U1479 : OAI221_X1 port map( B1 => n3632, B2 => n1135, C1 => n247, C2 => 
                           n1130, A => n1831, ZN => n1836);
   U1480 : AOI22_X1 port map( A1 => n888, A2 => n5217, B1 => n966, B2 => n1832,
                           ZN => n1833);
   U1481 : OAI221_X1 port map( B1 => n1834, B2 => n1140, C1 => n119, C2 => 
                           n1137, A => n1833, ZN => n1835);
   U1482 : NOR4_X1 port map( A1 => n1838, A2 => n1836, A3 => n1837, A4 => n1835
                           , ZN => n1839);
   U1483 : OAI222_X1 port map( A1 => n823, A2 => n1149, B1 => n1839, B2 => 
                           n1146, C1 => n3638, C2 => n1143, ZN => n1840);
   U1484 : OAI22_X1 port map( A1 => n3642, A2 => n1161, B1 => n951, B2 => n1158
                           , ZN => n1841);
   U1485 : AOI221_X1 port map( B1 => n1167, B2 => n4801, C1 => n1164, C2 => 
                           n4326, A => n1841, ZN => n1846);
   U1486 : OAI222_X1 port map( A1 => n631, A2 => n1174, B1 => n3645, B2 => 
                           n1171, C1 => n3644, C2 => n1170, ZN => n1842);
   U1487 : OAI22_X1 port map( A1 => n4673, A2 => n1189, B1 => n1404, B2 => 
                           n1184, ZN => n1843);
   U1488 : AOI221_X1 port map( B1 => n1194, B2 => n4961, C1 => n1191, C2 => 
                           n3648, A => n1843, ZN => n1844);
   U1489 : NAND4_X1 port map( A1 => n1847, A2 => n1845, A3 => n1844, A4 => 
                           n1846, ZN => n2519);
   U1490 : AOI22_X1 port map( A1 => n669, A2 => n4145, B1 => n1113, B2 => n4738
                           , ZN => n1848);
   U1491 : OAI221_X1 port map( B1 => n150, B2 => n1119, C1 => n1849, C2 => 
                           n1116, A => n1848, ZN => n1859);
   U1492 : AOI22_X1 port map( A1 => n1024, A2 => n5058, B1 => n493, B2 => n5122
                           , ZN => n1850);
   U1493 : AOI22_X1 port map( A1 => n54, A2 => n5090, B1 => n759, B2 => n1851, 
                           ZN => n1852);
   U1494 : AOI22_X1 port map( A1 => n1014, A2 => n5218, B1 => n490, B2 => n1853
                           , ZN => n1854);
   U1495 : OAI221_X1 port map( B1 => n1855, B2 => n1140, C1 => n118, C2 => 
                           n1137, A => n1854, ZN => n1856);
   U1496 : NOR4_X1 port map( A1 => n1859, A2 => n1856, A3 => n1858, A4 => n1857
                           , ZN => n1860);
   U1497 : OAI222_X1 port map( A1 => n822, A2 => n1149, B1 => n1860, B2 => 
                           n1146, C1 => n3663, C2 => n1143, ZN => n1861);
   U1498 : OAI22_X1 port map( A1 => n3667, A2 => n1162, B1 => n950, B2 => n1158
                           , ZN => n1862);
   U1499 : AOI221_X1 port map( B1 => n1167, B2 => n4802, C1 => n1164, C2 => 
                           n4325, A => n1862, ZN => n1867);
   U1500 : OAI222_X1 port map( A1 => n630, A2 => n1176, B1 => n3670, B2 => 
                           n1171, C1 => n3669, C2 => n1170, ZN => n1863);
   U1501 : AOI221_X1 port map( B1 => n1181, B2 => n4273, C1 => n1178, C2 => 
                           n4241, A => n1863, ZN => n1866);
   U1502 : OAI22_X1 port map( A1 => n4674, A2 => n1188, B1 => n1406, B2 => 
                           n1184, ZN => n1864);
   U1503 : AOI221_X1 port map( B1 => n1194, B2 => n4962, C1 => n1191, C2 => 
                           n3673, A => n1864, ZN => n1865);
   U1504 : NAND4_X1 port map( A1 => n1866, A2 => n1868, A3 => n1867, A4 => 
                           n1865, ZN => n2520);
   U1505 : AOI22_X1 port map( A1 => n969, A2 => n4144, B1 => n1112, B2 => n4739
                           , ZN => n1869);
   U1506 : OAI221_X1 port map( B1 => n149, B2 => n1119, C1 => n1870, C2 => 
                           n1114, A => n1869, ZN => n1878);
   U1507 : AOI22_X1 port map( A1 => n1024, A2 => n5059, B1 => n508, B2 => n5123
                           , ZN => n1871);
   U1508 : AOI22_X1 port map( A1 => n54, A2 => n5091, B1 => n760, B2 => n220, 
                           ZN => n1872);
   U1509 : OAI221_X1 port map( B1 => n3682, B2 => n1135, C1 => n245, C2 => n506
                           , A => n1872, ZN => n1876);
   U1510 : AOI22_X1 port map( A1 => n2211, A2 => n5219, B1 => n489, B2 => n221,
                           ZN => n1873);
   U1511 : NOR4_X1 port map( A1 => n1878, A2 => n1876, A3 => n1877, A4 => n1875
                           , ZN => n1879);
   U1512 : OAI222_X1 port map( A1 => n821, A2 => n1149, B1 => n1879, B2 => 
                           n1146, C1 => n3688, C2 => n1143, ZN => n1880);
   U1513 : OAI22_X1 port map( A1 => n3692, A2 => n1161, B1 => n949, B2 => n1158
                           , ZN => n1881);
   U1514 : AOI221_X1 port map( B1 => n1167, B2 => n4803, C1 => n1164, C2 => 
                           n4324, A => n1881, ZN => n1886);
   U1515 : OAI222_X1 port map( A1 => n629, A2 => n1176, B1 => n3695, B2 => 
                           n1171, C1 => n3694, C2 => n1170, ZN => n1882);
   U1516 : AOI221_X1 port map( B1 => n1181, B2 => n4272, C1 => n1178, C2 => 
                           n4240, A => n1882, ZN => n1885);
   U1517 : OAI22_X1 port map( A1 => n4675, A2 => n1188, B1 => n1408, B2 => 
                           n1184, ZN => n1883);
   U1518 : AOI221_X1 port map( B1 => n1194, B2 => n4963, C1 => n1191, C2 => 
                           n3698, A => n1883, ZN => n1884);
   U1519 : NAND4_X1 port map( A1 => n1887, A2 => n1884, A3 => n1886, A4 => 
                           n1885, ZN => n2521);
   U1520 : AOI22_X1 port map( A1 => n669, A2 => n4143, B1 => n486, B2 => n4740,
                           ZN => n1888);
   U1521 : OAI221_X1 port map( B1 => n148, B2 => n1117, C1 => n1889, C2 => 
                           n1115, A => n1888, ZN => n1899);
   U1522 : AOI22_X1 port map( A1 => n1123, A2 => n5060, B1 => n493, B2 => n5124
                           , ZN => n1890);
   U1523 : OAI221_X1 port map( B1 => n3706, B2 => n1129, C1 => n276, C2 => 
                           n1126, A => n1890, ZN => n1898);
   U1524 : AOI22_X1 port map( A1 => n55, A2 => n5092, B1 => n1029, B2 => n1891,
                           ZN => n1892);
   U1525 : OAI221_X1 port map( B1 => n3707, B2 => n1134, C1 => n506, C2 => n244
                           , A => n1892, ZN => n1897);
   U1526 : AOI22_X1 port map( A1 => n2211, A2 => n5220, B1 => n489, B2 => n1893
                           , ZN => n1894);
   U1527 : NOR4_X1 port map( A1 => n1899, A2 => n1898, A3 => n1897, A4 => n1896
                           , ZN => n1900);
   U1528 : OAI222_X1 port map( A1 => n820, A2 => n1149, B1 => n1900, B2 => 
                           n1146, C1 => n3713, C2 => n1143, ZN => n1901);
   U1529 : OAI22_X1 port map( A1 => n3717, A2 => n1162, B1 => n948, B2 => n1158
                           , ZN => n1902);
   U1530 : AOI221_X1 port map( B1 => n1167, B2 => n4804, C1 => n1164, C2 => 
                           n4323, A => n1902, ZN => n1907);
   U1531 : OAI22_X1 port map( A1 => n4676, A2 => n1188, B1 => n1410, B2 => 
                           n1184, ZN => n1904);
   U1532 : AOI221_X1 port map( B1 => n1194, B2 => n4964, C1 => n1191, C2 => 
                           n3723, A => n1904, ZN => n1905);
   U1533 : NAND4_X1 port map( A1 => n1908, A2 => n1907, A3 => n1905, A4 => 
                           n1906, ZN => n2522);
   U1534 : AOI22_X1 port map( A1 => n669, A2 => n4142, B1 => n487, B2 => n4741,
                           ZN => n1909);
   U1535 : OAI221_X1 port map( B1 => n147, B2 => n1119, C1 => n1910, C2 => 
                           n1115, A => n1909, ZN => n1920);
   U1536 : AOI22_X1 port map( A1 => n1024, A2 => n5061, B1 => n1120, B2 => 
                           n5125, ZN => n1911);
   U1537 : OAI221_X1 port map( B1 => n3731, B2 => n1128, C1 => n275, C2 => 
                           n1126, A => n1911, ZN => n1919);
   U1538 : AOI22_X1 port map( A1 => n57, A2 => n5093, B1 => n1029, B2 => n1912,
                           ZN => n1913);
   U1539 : OAI221_X1 port map( B1 => n507, B2 => n3732, C1 => n243, C2 => n1131
                           , A => n1913, ZN => n1918);
   U1540 : AOI22_X1 port map( A1 => n888, A2 => n5221, B1 => n966, B2 => n1914,
                           ZN => n1915);
   U1541 : OAI221_X1 port map( B1 => n1916, B2 => n1140, C1 => n115, C2 => 
                           n1137, A => n1915, ZN => n1917);
   U1542 : NOR4_X1 port map( A1 => n1920, A2 => n1919, A3 => n1917, A4 => n1918
                           , ZN => n1921);
   U1543 : OAI22_X1 port map( A1 => n3742, A2 => n707, B1 => n947, B2 => n1158,
                           ZN => n1922);
   U1544 : AOI221_X1 port map( B1 => n1167, B2 => n4805, C1 => n1164, C2 => 
                           n4322, A => n1922, ZN => n1927);
   U1545 : OAI22_X1 port map( A1 => n4677, A2 => n1188, B1 => n1412, B2 => 
                           n1184, ZN => n1924);
   U1546 : AOI221_X1 port map( B1 => n1194, B2 => n4965, C1 => n1191, C2 => 
                           n3748, A => n1924, ZN => n1925);
   U1547 : NAND4_X1 port map( A1 => n1928, A2 => n1927, A3 => n1925, A4 => 
                           n1926, ZN => n2523);
   U1548 : AOI22_X1 port map( A1 => n669, A2 => n4141, B1 => n691, B2 => n4742,
                           ZN => n1929);
   U1549 : OAI221_X1 port map( B1 => n146, B2 => n1119, C1 => n1930, C2 => 
                           n1116, A => n1929, ZN => n1940);
   U1550 : AOI22_X1 port map( A1 => n1122, A2 => n5062, B1 => n508, B2 => n5126
                           , ZN => n1931);
   U1551 : OAI221_X1 port map( B1 => n3756, B2 => n1127, C1 => n274, C2 => 
                           n1126, A => n1931, ZN => n1939);
   U1552 : AOI22_X1 port map( A1 => n54, A2 => n5094, B1 => n1029, B2 => n1932,
                           ZN => n1933);
   U1553 : OAI221_X1 port map( B1 => n3757, B2 => n1135, C1 => n242, C2 => 
                           n1131, A => n1933, ZN => n1938);
   U1554 : AOI22_X1 port map( A1 => n888, A2 => n5222, B1 => n578, B2 => n1934,
                           ZN => n1935);
   U1555 : NOR4_X1 port map( A1 => n1940, A2 => n1939, A3 => n1938, A4 => n1937
                           , ZN => n1941);
   U1556 : OAI22_X1 port map( A1 => n3767, A2 => n1161, B1 => n946, B2 => n1158
                           , ZN => n1942);
   U1557 : AOI221_X1 port map( B1 => n1167, B2 => n4806, C1 => n1164, C2 => 
                           n4321, A => n1942, ZN => n1947);
   U1558 : OAI22_X1 port map( A1 => n4678, A2 => n1188, B1 => n1414, B2 => 
                           n1184, ZN => n1944);
   U1559 : AOI221_X1 port map( B1 => n1194, B2 => n4966, C1 => n1191, C2 => 
                           n3773, A => n1944, ZN => n1945);
   U1560 : NAND4_X1 port map( A1 => n1948, A2 => n1947, A3 => n1945, A4 => 
                           n1946, ZN => n2524);
   U1561 : AOI22_X1 port map( A1 => n969, A2 => n4140, B1 => n691, B2 => n4743,
                           ZN => n1949);
   U1562 : OAI221_X1 port map( B1 => n145, B2 => n1118, C1 => n1950, C2 => 
                           n1115, A => n1949, ZN => n1960);
   U1563 : AOI22_X1 port map( A1 => n1123, A2 => n5063, B1 => n51, B2 => n5127,
                           ZN => n1951);
   U1564 : OAI221_X1 port map( B1 => n3781, B2 => n1129, C1 => n273, C2 => 
                           n1126, A => n1951, ZN => n1959);
   U1565 : AOI22_X1 port map( A1 => n55, A2 => n5095, B1 => n759, B2 => n1952, 
                           ZN => n1953);
   U1566 : OAI221_X1 port map( B1 => n3782, B2 => n507, C1 => n241, C2 => n1131
                           , A => n1953, ZN => n1958);
   U1567 : AOI22_X1 port map( A1 => n2211, A2 => n5223, B1 => n966, B2 => n1954
                           , ZN => n1955);
   U1568 : OAI221_X1 port map( B1 => n1956, B2 => n1140, C1 => n113, C2 => 
                           n1137, A => n1955, ZN => n1957);
   U1569 : NOR4_X1 port map( A1 => n1960, A2 => n1959, A3 => n1957, A4 => n1958
                           , ZN => n1961);
   U1570 : OAI22_X1 port map( A1 => n3792, A2 => n1161, B1 => n945, B2 => n1158
                           , ZN => n1962);
   U1571 : AOI221_X1 port map( B1 => n1167, B2 => n4807, C1 => n1164, C2 => 
                           n4320, A => n1962, ZN => n1967);
   U1572 : OAI22_X1 port map( A1 => n4679, A2 => n1188, B1 => n1416, B2 => 
                           n1184, ZN => n1964);
   U1573 : AOI221_X1 port map( B1 => n1194, B2 => n4967, C1 => n1191, C2 => 
                           n3798, A => n1964, ZN => n1965);
   U1574 : NAND4_X1 port map( A1 => n1968, A2 => n1966, A3 => n1965, A4 => 
                           n1967, ZN => n2525);
   U1575 : AOI22_X1 port map( A1 => n669, A2 => n4139, B1 => n497, B2 => n4744,
                           ZN => n1969);
   U1576 : OAI221_X1 port map( B1 => n144, B2 => n1119, C1 => n1970, C2 => 
                           n1116, A => n1969, ZN => n1980);
   U1577 : AOI22_X1 port map( A1 => n1023, A2 => n5064, B1 => n508, B2 => n5128
                           , ZN => n1971);
   U1578 : OAI221_X1 port map( B1 => n3806, B2 => n1127, C1 => n272, C2 => 
                           n1126, A => n1971, ZN => n1979);
   U1579 : AOI22_X1 port map( A1 => n56, A2 => n5096, B1 => n1029, B2 => n1972,
                           ZN => n1973);
   U1580 : OAI221_X1 port map( B1 => n3807, B2 => n1135, C1 => n240, C2 => n506
                           , A => n1973, ZN => n1978);
   U1581 : AOI22_X1 port map( A1 => n1014, A2 => n5224, B1 => n578, B2 => n1974
                           , ZN => n1975);
   U1582 : OAI221_X1 port map( B1 => n1976, B2 => n1140, C1 => n112, C2 => 
                           n1137, A => n1975, ZN => n1977);
   U1583 : NOR4_X1 port map( A1 => n1980, A2 => n1979, A3 => n1977, A4 => n1978
                           , ZN => n1981);
   U1584 : OAI222_X1 port map( A1 => n816, A2 => n1149, B1 => n1981, B2 => 
                           n1146, C1 => n3813, C2 => n1143, ZN => n1982);
   U1585 : OAI22_X1 port map( A1 => n3817, A2 => n1161, B1 => n944, B2 => n1158
                           , ZN => n1983);
   U1586 : AOI221_X1 port map( B1 => n1167, B2 => n4808, C1 => n1164, C2 => 
                           n4319, A => n1983, ZN => n1988);
   U1587 : OAI222_X1 port map( A1 => n624, A2 => n1175, B1 => n3820, B2 => 
                           n1171, C1 => n3819, C2 => n1170, ZN => n1984);
   U1588 : AOI221_X1 port map( B1 => n1181, B2 => n4267, C1 => n1178, C2 => 
                           n4235, A => n1984, ZN => n1987);
   U1589 : OAI22_X1 port map( A1 => n4680, A2 => n1188, B1 => n1418, B2 => 
                           n1184, ZN => n1985);
   U1590 : AOI221_X1 port map( B1 => n1194, B2 => n4968, C1 => n1191, C2 => 
                           n3823, A => n1985, ZN => n1986);
   U1591 : NAND4_X1 port map( A1 => n1989, A2 => n1986, A3 => n1988, A4 => 
                           n1987, ZN => n2526);
   U1592 : AOI22_X1 port map( A1 => n969, A2 => n4138, B1 => n1113, B2 => n4745
                           , ZN => n1990);
   U1593 : OAI221_X1 port map( B1 => n143, B2 => n1118, C1 => n1991, C2 => 
                           n1116, A => n1990, ZN => n2001);
   U1594 : AOI22_X1 port map( A1 => n1124, A2 => n5065, B1 => n51, B2 => n5129,
                           ZN => n1992);
   U1595 : OAI221_X1 port map( B1 => n3831, B2 => n1129, C1 => n271, C2 => 
                           n1126, A => n1992, ZN => n2000);
   U1596 : AOI22_X1 port map( A1 => n56, A2 => n5097, B1 => n760, B2 => n1993, 
                           ZN => n1994);
   U1597 : AOI22_X1 port map( A1 => n1014, A2 => n5225, B1 => n579, B2 => n1995
                           , ZN => n1996);
   U1598 : NOR4_X1 port map( A1 => n2001, A2 => n2000, A3 => n1999, A4 => n1998
                           , ZN => n2002);
   U1599 : OAI22_X1 port map( A1 => n3842, A2 => n1162, B1 => n943, B2 => n1158
                           , ZN => n2003);
   U1600 : AOI221_X1 port map( B1 => n1167, B2 => n4809, C1 => n1164, C2 => 
                           n4318, A => n2003, ZN => n2008);
   U1601 : OAI22_X1 port map( A1 => n4681, A2 => n1188, B1 => n1420, B2 => 
                           n1184, ZN => n2005);
   U1602 : AOI221_X1 port map( B1 => n1194, B2 => n4969, C1 => n1191, C2 => 
                           n3848, A => n2005, ZN => n2006);
   U1603 : NAND4_X1 port map( A1 => n2009, A2 => n2008, A3 => n2006, A4 => 
                           n2007, ZN => n2527);
   U1604 : AOI22_X1 port map( A1 => n669, A2 => n4137, B1 => n738, B2 => n4746,
                           ZN => n2010);
   U1605 : OAI221_X1 port map( B1 => n142, B2 => n1119, C1 => n2011, C2 => 
                           n1114, A => n2010, ZN => n2021);
   U1606 : AOI22_X1 port map( A1 => n1124, A2 => n5066, B1 => n493, B2 => n5130
                           , ZN => n2012);
   U1607 : OAI221_X1 port map( B1 => n3856, B2 => n1128, C1 => n270, C2 => 
                           n1126, A => n2012, ZN => n2020);
   U1608 : AOI22_X1 port map( A1 => n54, A2 => n5098, B1 => n760, B2 => n2013, 
                           ZN => n2014);
   U1609 : OAI221_X1 port map( B1 => n3857, B2 => n1133, C1 => n238, C2 => 
                           n1130, A => n2014, ZN => n2019);
   U1610 : AOI22_X1 port map( A1 => n1014, A2 => n5226, B1 => n490, B2 => n2015
                           , ZN => n2016);
   U1611 : NOR4_X1 port map( A1 => n2021, A2 => n2020, A3 => n2018, A4 => n2019
                           , ZN => n2022);
   U1612 : OAI222_X1 port map( A1 => n814, A2 => n1149, B1 => n2022, B2 => 
                           n1146, C1 => n3863, C2 => n1143, ZN => n2023);
   U1613 : OAI22_X1 port map( A1 => n3867, A2 => n1160, B1 => n942, B2 => n1158
                           , ZN => n2024);
   U1614 : AOI221_X1 port map( B1 => n1167, B2 => n4810, C1 => n1164, C2 => 
                           n4317, A => n2024, ZN => n2029);
   U1615 : OAI222_X1 port map( A1 => n622, A2 => n1175, B1 => n3870, B2 => 
                           n1172, C1 => n3869, C2 => n1170, ZN => n2025);
   U1616 : AOI221_X1 port map( B1 => n1181, B2 => n4265, C1 => n1178, C2 => 
                           n4233, A => n2025, ZN => n2028);
   U1617 : OAI22_X1 port map( A1 => n4682, A2 => n1188, B1 => n1422, B2 => 
                           n1184, ZN => n2026);
   U1618 : AOI221_X1 port map( B1 => n1194, B2 => n4970, C1 => n1191, C2 => 
                           n3873, A => n2026, ZN => n2027);
   U1619 : NAND4_X1 port map( A1 => n2030, A2 => n2029, A3 => n2027, A4 => 
                           n2028, ZN => n2528);
   U1620 : AOI22_X1 port map( A1 => n969, A2 => n4136, B1 => n487, B2 => n4747,
                           ZN => n2031);
   U1621 : OAI221_X1 port map( B1 => n141, B2 => n1119, C1 => n2032, C2 => 
                           n1116, A => n2031, ZN => n2042);
   U1622 : AOI22_X1 port map( A1 => n1124, A2 => n5067, B1 => n512, B2 => n5131
                           , ZN => n2033);
   U1623 : OAI221_X1 port map( B1 => n3881, B2 => n1127, C1 => n269, C2 => 
                           n1126, A => n2033, ZN => n2041);
   U1624 : AOI22_X1 port map( A1 => n54, A2 => n5099, B1 => n759, B2 => n2034, 
                           ZN => n2035);
   U1625 : OAI221_X1 port map( B1 => n3882, B2 => n1133, C1 => n237, C2 => n506
                           , A => n2035, ZN => n2040);
   U1626 : AOI22_X1 port map( A1 => n1014, A2 => n5227, B1 => n577, B2 => n2036
                           , ZN => n2037);
   U1627 : NOR4_X1 port map( A1 => n2042, A2 => n2041, A3 => n2039, A4 => n2040
                           , ZN => n2043);
   U1628 : OAI222_X1 port map( A1 => n813, A2 => n1149, B1 => n2043, B2 => 
                           n1146, C1 => n3888, C2 => n1143, ZN => n2044);
   U1629 : OAI22_X1 port map( A1 => n3892, A2 => n1160, B1 => n941, B2 => n1158
                           , ZN => n2045);
   U1630 : AOI221_X1 port map( B1 => n1167, B2 => n4811, C1 => n1164, C2 => 
                           n4316, A => n2045, ZN => n2050);
   U1631 : OAI222_X1 port map( A1 => n621, A2 => n1176, B1 => n3895, B2 => 
                           n1172, C1 => n3894, C2 => n1170, ZN => n2046);
   U1632 : AOI221_X1 port map( B1 => n1181, B2 => n4264, C1 => n1178, C2 => 
                           n4232, A => n2046, ZN => n2049);
   U1633 : OAI22_X1 port map( A1 => n4683, A2 => n1188, B1 => n1424, B2 => 
                           n1184, ZN => n2047);
   U1634 : AOI221_X1 port map( B1 => n1194, B2 => n4971, C1 => n1191, C2 => 
                           n3898, A => n2047, ZN => n2048);
   U1635 : NAND4_X1 port map( A1 => n2051, A2 => n2050, A3 => n2048, A4 => 
                           n2049, ZN => n2529);
   U1636 : AOI22_X1 port map( A1 => n969, A2 => n4135, B1 => n1113, B2 => n4748
                           , ZN => n2052);
   U1637 : OAI221_X1 port map( B1 => n140, B2 => n1119, C1 => n2053, C2 => 
                           n1114, A => n2052, ZN => n2063);
   U1638 : AOI22_X1 port map( A1 => n1016, A2 => n5068, B1 => n512, B2 => n5132
                           , ZN => n2054);
   U1639 : OAI221_X1 port map( B1 => n3907, B2 => n1129, C1 => n268, C2 => n678
                           , A => n2054, ZN => n2062);
   U1640 : AOI22_X1 port map( A1 => n56, A2 => n5100, B1 => n760, B2 => n2055, 
                           ZN => n2056);
   U1641 : OAI221_X1 port map( B1 => n3908, B2 => n1133, C1 => n236, C2 => 
                           n1131, A => n2056, ZN => n2061);
   U1642 : AOI22_X1 port map( A1 => n888, A2 => n5228, B1 => n490, B2 => n2057,
                           ZN => n2058);
   U1643 : OAI221_X1 port map( B1 => n2059, B2 => n1141, C1 => n108, C2 => 
                           n1138, A => n2058, ZN => n2060);
   U1644 : NOR4_X1 port map( A1 => n2063, A2 => n2062, A3 => n2060, A4 => n2061
                           , ZN => n2064);
   U1645 : OAI22_X1 port map( A1 => n3918, A2 => n1160, B1 => n940, B2 => n1159
                           , ZN => n2066);
   U1646 : AOI221_X1 port map( B1 => n1168, B2 => n4812, C1 => n1165, C2 => 
                           n4315, A => n2066, ZN => n2071);
   U1647 : OAI222_X1 port map( A1 => n620, A2 => n1175, B1 => n3921, B2 => 
                           n1172, C1 => n3920, C2 => n876, ZN => n2067);
   U1648 : AOI221_X1 port map( B1 => n1182, B2 => n4263, C1 => n1179, C2 => 
                           n4231, A => n2067, ZN => n2070);
   U1649 : OAI22_X1 port map( A1 => n4684, A2 => n1188, B1 => n1427, B2 => 
                           n1185, ZN => n2068);
   U1650 : AOI221_X1 port map( B1 => n1195, B2 => n4972, C1 => n1192, C2 => 
                           n3924, A => n2068, ZN => n2069);
   U1651 : NAND4_X1 port map( A1 => n2072, A2 => n2071, A3 => n2069, A4 => 
                           n2070, ZN => n2530);
   U1652 : AOI22_X1 port map( A1 => n669, A2 => n4134, B1 => n1112, B2 => n4749
                           , ZN => n2073);
   U1653 : OAI221_X1 port map( B1 => n139, B2 => n1119, C1 => n2074, C2 => 
                           n1116, A => n2073, ZN => n2084);
   U1654 : AOI22_X1 port map( A1 => n1123, A2 => n5069, B1 => n52, B2 => n5133,
                           ZN => n2075);
   U1655 : OAI221_X1 port map( B1 => n3933, B2 => n1127, C1 => n267, C2 => n678
                           , A => n2075, ZN => n2083);
   U1656 : AOI22_X1 port map( A1 => n56, A2 => n5101, B1 => n760, B2 => n2076, 
                           ZN => n2077);
   U1657 : OAI221_X1 port map( B1 => n3934, B2 => n1133, C1 => n235, C2 => 
                           n1130, A => n2077, ZN => n2082);
   U1658 : AOI22_X1 port map( A1 => n1014, A2 => n5229, B1 => n490, B2 => n2078
                           , ZN => n2079);
   U1659 : OAI221_X1 port map( B1 => n2080, B2 => n1141, C1 => n107, C2 => 
                           n1138, A => n2079, ZN => n2081);
   U1660 : NOR4_X1 port map( A1 => n2084, A2 => n2083, A3 => n2081, A4 => n2082
                           , ZN => n2085);
   U1661 : OAI222_X1 port map( A1 => n811, A2 => n1150, B1 => n2085, B2 => 
                           n1147, C1 => n3940, C2 => n1144, ZN => n2086);
   U1662 : OAI22_X1 port map( A1 => n3944, A2 => n1162, B1 => n939, B2 => n1159
                           , ZN => n2087);
   U1663 : OAI222_X1 port map( A1 => n619, A2 => n1176, B1 => n3947, B2 => 
                           n1172, C1 => n3946, C2 => n876, ZN => n2088);
   U1664 : AOI221_X1 port map( B1 => n1182, B2 => n4262, C1 => n1179, C2 => 
                           n4230, A => n2088, ZN => n2091);
   U1665 : OAI22_X1 port map( A1 => n4685, A2 => n1187, B1 => n1430, B2 => 
                           n1185, ZN => n2089);
   U1666 : AOI221_X1 port map( B1 => n1195, B2 => n4973, C1 => n1192, C2 => 
                           n3950, A => n2089, ZN => n2090);
   U1667 : NAND4_X1 port map( A1 => n2093, A2 => n2092, A3 => n2090, A4 => 
                           n2091, ZN => n2531);
   U1668 : AOI22_X1 port map( A1 => n668, A2 => n4133, B1 => n1113, B2 => n4750
                           , ZN => n2094);
   U1669 : OAI221_X1 port map( B1 => n138, B2 => n1119, C1 => n2095, C2 => 
                           n1114, A => n2094, ZN => n2105);
   U1670 : AOI22_X1 port map( A1 => n1016, A2 => n5070, B1 => n1120, B2 => 
                           n5134, ZN => n2096);
   U1671 : AOI22_X1 port map( A1 => n57, A2 => n5102, B1 => n1029, B2 => n2097,
                           ZN => n2098);
   U1672 : OAI221_X1 port map( B1 => n3960, B2 => n1135, C1 => n234, C2 => n506
                           , A => n2098, ZN => n2103);
   U1673 : AOI22_X1 port map( A1 => n888, A2 => n5230, B1 => n577, B2 => n2099,
                           ZN => n2100);
   U1674 : OAI221_X1 port map( B1 => n2101, B2 => n1141, C1 => n106, C2 => 
                           n1138, A => n2100, ZN => n2102);
   U1675 : NOR4_X1 port map( A1 => n2105, A2 => n2102, A3 => n2103, A4 => n2104
                           , ZN => n2106);
   U1676 : OAI222_X1 port map( A1 => n810, A2 => n1150, B1 => n2106, B2 => 
                           n1147, C1 => n3966, C2 => n1144, ZN => n2107);
   U1677 : OAI22_X1 port map( A1 => n3970, A2 => n1160, B1 => n938, B2 => n1159
                           , ZN => n2108);
   U1678 : AOI221_X1 port map( B1 => n1168, B2 => n4814, C1 => n1165, C2 => 
                           n4313, A => n2108, ZN => n2113);
   U1679 : OAI222_X1 port map( A1 => n618, A2 => n1176, B1 => n3973, B2 => 
                           n1173, C1 => n3972, C2 => n876, ZN => n2109);
   U1680 : AOI221_X1 port map( B1 => n1182, B2 => n4261, C1 => n1179, C2 => 
                           n4229, A => n2109, ZN => n2112);
   U1681 : OAI22_X1 port map( A1 => n4686, A2 => n1187, B1 => n1433, B2 => 
                           n1185, ZN => n2110);
   U1682 : AOI221_X1 port map( B1 => n1195, B2 => n4974, C1 => n1192, C2 => 
                           n3976, A => n2110, ZN => n2111);
   U1683 : NAND4_X1 port map( A1 => n2112, A2 => n2113, A3 => n2111, A4 => 
                           n2114, ZN => n2532);
   U1684 : AOI22_X1 port map( A1 => n969, A2 => n4132, B1 => n497, B2 => n4751,
                           ZN => n2115);
   U1685 : OAI221_X1 port map( B1 => n137, B2 => n1118, C1 => n2116, C2 => 
                           n1115, A => n2115, ZN => n2126);
   U1686 : AOI22_X1 port map( A1 => n1023, A2 => n5071, B1 => n493, B2 => n5135
                           , ZN => n2117);
   U1687 : OAI221_X1 port map( B1 => n3985, B2 => n1128, C1 => n265, C2 => n678
                           , A => n2117, ZN => n2125);
   U1688 : AOI22_X1 port map( A1 => n57, A2 => n5103, B1 => n759, B2 => n2118, 
                           ZN => n2119);
   U1689 : OAI221_X1 port map( B1 => n3986, B2 => n1133, C1 => n233, C2 => n506
                           , A => n2119, ZN => n2124);
   U1690 : AOI22_X1 port map( A1 => n888, A2 => n5231, B1 => n966, B2 => n2120,
                           ZN => n2121);
   U1691 : OAI221_X1 port map( B1 => n2122, B2 => n1141, C1 => n105, C2 => 
                           n1138, A => n2121, ZN => n2123);
   U1692 : NOR4_X1 port map( A1 => n2126, A2 => n2125, A3 => n2124, A4 => n2123
                           , ZN => n2127);
   U1693 : OAI222_X1 port map( A1 => n809, A2 => n1150, B1 => n2127, B2 => 
                           n1147, C1 => n3992, C2 => n1144, ZN => n2128);
   U1694 : OAI22_X1 port map( A1 => n3996, A2 => n1160, B1 => n937, B2 => n1159
                           , ZN => n2129);
   U1695 : AOI221_X1 port map( B1 => n1168, B2 => n4815, C1 => n1165, C2 => 
                           n4312, A => n2129, ZN => n2134);
   U1696 : OAI222_X1 port map( A1 => n617, A2 => n1174, B1 => n1173, B2 => 
                           n3999, C1 => n3998, C2 => n876, ZN => n2130);
   U1697 : AOI221_X1 port map( B1 => n1182, B2 => n4260, C1 => n1179, C2 => 
                           n4228, A => n2130, ZN => n2133);
   U1698 : OAI22_X1 port map( A1 => n4687, A2 => n1187, B1 => n1436, B2 => 
                           n1185, ZN => n2131);
   U1699 : AOI221_X1 port map( B1 => n1195, B2 => n4975, C1 => n1192, C2 => 
                           n4002, A => n2131, ZN => n2132);
   U1700 : NAND4_X1 port map( A1 => n2133, A2 => n2132, A3 => n2135, A4 => 
                           n2134, ZN => n2533);
   U1701 : AOI22_X1 port map( A1 => n969, A2 => n4131, B1 => n1111, B2 => n4752
                           , ZN => n2136);
   U1702 : OAI221_X1 port map( B1 => n136, B2 => n1118, C1 => n2137, C2 => 
                           n1116, A => n2136, ZN => n2147);
   U1703 : AOI22_X1 port map( A1 => n1023, A2 => n5072, B1 => n1121, B2 => 
                           n5136, ZN => n2138);
   U1704 : OAI221_X1 port map( B1 => n4011, B2 => n1129, C1 => n264, C2 => n678
                           , A => n2138, ZN => n2146);
   U1705 : AOI22_X1 port map( A1 => n57, A2 => n5104, B1 => n759, B2 => n2139, 
                           ZN => n2140);
   U1706 : OAI221_X1 port map( B1 => n4012, B2 => n1133, C1 => n232, C2 => n506
                           , A => n2140, ZN => n2145);
   U1707 : AOI22_X1 port map( A1 => n888, A2 => n5232, B1 => n966, B2 => n2141,
                           ZN => n2142);
   U1708 : OAI221_X1 port map( B1 => n2143, B2 => n1141, C1 => n104, C2 => 
                           n1138, A => n2142, ZN => n2144);
   U1709 : NOR4_X1 port map( A1 => n2147, A2 => n2146, A3 => n2145, A4 => n2144
                           , ZN => n2148);
   U1710 : OAI222_X1 port map( A1 => n808, A2 => n1150, B1 => n2148, B2 => 
                           n1147, C1 => n4018, C2 => n1144, ZN => n2149);
   U1711 : OAI22_X1 port map( A1 => n4022, A2 => n1160, B1 => n936, B2 => n1159
                           , ZN => n2150);
   U1712 : AOI221_X1 port map( B1 => n1168, B2 => n4816, C1 => n1165, C2 => 
                           n4311, A => n2150, ZN => n2155);
   U1713 : OAI222_X1 port map( A1 => n616, A2 => n1175, B1 => n4025, B2 => 
                           n1172, C1 => n4024, C2 => n876, ZN => n2151);
   U1714 : AOI221_X1 port map( B1 => n1182, B2 => n4259, C1 => n1179, C2 => 
                           n4227, A => n2151, ZN => n2154);
   U1715 : OAI22_X1 port map( A1 => n4688, A2 => n1187, B1 => n1439, B2 => 
                           n1185, ZN => n2152);
   U1716 : AOI221_X1 port map( B1 => n1195, B2 => n4976, C1 => n1192, C2 => 
                           n4028, A => n2152, ZN => n2153);
   U1717 : NAND4_X1 port map( A1 => n2154, A2 => n2155, A3 => n2153, A4 => 
                           n2156, ZN => n2534);
   U1718 : AOI22_X1 port map( A1 => n668, A2 => n4130, B1 => n1112, B2 => n4753
                           , ZN => n2157);
   U1719 : OAI221_X1 port map( B1 => n135, B2 => n1118, C1 => n2158, C2 => 
                           n1116, A => n2157, ZN => n2168);
   U1720 : AOI22_X1 port map( A1 => n1123, A2 => n5073, B1 => n51, B2 => n5137,
                           ZN => n2159);
   U1721 : OAI221_X1 port map( B1 => n4037, B2 => n1128, C1 => n263, C2 => n678
                           , A => n2159, ZN => n2167);
   U1722 : AOI22_X1 port map( A1 => n56, A2 => n5105, B1 => n1029, B2 => n2160,
                           ZN => n2161);
   U1723 : OAI221_X1 port map( B1 => n4038, B2 => n507, C1 => n231, C2 => n506,
                           A => n2161, ZN => n2166);
   U1724 : AOI22_X1 port map( A1 => n2211, A2 => n5233, B1 => n577, B2 => n2162
                           , ZN => n2163);
   U1725 : OAI221_X1 port map( B1 => n2164, B2 => n1141, C1 => n103, C2 => 
                           n1138, A => n2163, ZN => n2165);
   U1726 : NOR4_X1 port map( A1 => n2168, A2 => n2167, A3 => n2165, A4 => n2166
                           , ZN => n2169);
   U1727 : OAI22_X1 port map( A1 => n4048, A2 => n1160, B1 => n935, B2 => n1159
                           , ZN => n2171);
   U1728 : AOI221_X1 port map( B1 => n1168, B2 => n4817, C1 => n1165, C2 => 
                           n4310, A => n2171, ZN => n2176);
   U1729 : OAI222_X1 port map( A1 => n615, A2 => n1174, B1 => n1171, B2 => 
                           n4051, C1 => n4050, C2 => n876, ZN => n2172);
   U1730 : AOI221_X1 port map( B1 => n1182, B2 => n4258, C1 => n1179, C2 => 
                           n4226, A => n2172, ZN => n2175);
   U1731 : OAI22_X1 port map( A1 => n4689, A2 => n1187, B1 => n1442, B2 => 
                           n1185, ZN => n2173);
   U1732 : AOI221_X1 port map( B1 => n1195, B2 => n4977, C1 => n1192, C2 => 
                           n4054, A => n2173, ZN => n2174);
   U1733 : NAND4_X1 port map( A1 => n2177, A2 => n2176, A3 => n2174, A4 => 
                           n2175, ZN => n2535);
   U1734 : AOI22_X1 port map( A1 => n969, A2 => n4129, B1 => n1111, B2 => n4754
                           , ZN => n2178);
   U1735 : OAI221_X1 port map( B1 => n134, B2 => n1117, C1 => n2179, C2 => 
                           n1115, A => n2178, ZN => n2189);
   U1736 : AOI22_X1 port map( A1 => n1016, A2 => n5074, B1 => n512, B2 => n5138
                           , ZN => n2180);
   U1737 : AOI22_X1 port map( A1 => n57, A2 => n5106, B1 => n759, B2 => n2181, 
                           ZN => n2182);
   U1738 : OAI221_X1 port map( B1 => n4064, B2 => n1135, C1 => n230, C2 => n506
                           , A => n2182, ZN => n2187);
   U1739 : AOI22_X1 port map( A1 => n2211, A2 => n5234, B1 => n966, B2 => n2183
                           , ZN => n2184);
   U1740 : NOR4_X1 port map( A1 => n2189, A2 => n2187, A3 => n2188, A4 => n2186
                           , ZN => n2190);
   U1741 : OAI222_X1 port map( A1 => n806, A2 => n1150, B1 => n2190, B2 => 
                           n1147, C1 => n4070, C2 => n1144, ZN => n2191);
   U1742 : OAI22_X1 port map( A1 => n4074, A2 => n1160, B1 => n934, B2 => n1159
                           , ZN => n2192);
   U1743 : AOI221_X1 port map( B1 => n1168, B2 => n4818, C1 => n1165, C2 => 
                           n4309, A => n2192, ZN => n2197);
   U1744 : OAI222_X1 port map( A1 => n614, A2 => n1174, B1 => n1171, B2 => 
                           n4077, C1 => n4076, C2 => n876, ZN => n2193);
   U1745 : AOI221_X1 port map( B1 => n1182, B2 => n4257, C1 => n1179, C2 => 
                           n4225, A => n2193, ZN => n2196);
   U1746 : OAI22_X1 port map( A1 => n4690, A2 => n1187, B1 => n1445, B2 => 
                           n1185, ZN => n2194);
   U1747 : AOI221_X1 port map( B1 => n1195, B2 => n4978, C1 => n1192, C2 => 
                           n4080, A => n2194, ZN => n2195);
   U1748 : NAND4_X1 port map( A1 => n2198, A2 => n2197, A3 => n2195, A4 => 
                           n2196, ZN => n2536);
   U1749 : AOI22_X1 port map( A1 => n668, A2 => n4128, B1 => n497, B2 => n4755,
                           ZN => n2199);
   U1750 : OAI221_X1 port map( B1 => n133, B2 => n1119, C1 => n2201, C2 => 
                           n1115, A => n2199, ZN => n2219);
   U1751 : AOI22_X1 port map( A1 => n1023, A2 => n5075, B1 => n508, B2 => n5139
                           , ZN => n2203);
   U1752 : AOI22_X1 port map( A1 => n55, A2 => n5107, B1 => n760, B2 => n2206, 
                           ZN => n2207);
   U1753 : OAI221_X1 port map( B1 => n4095, B2 => n1135, C1 => n229, C2 => 
                           n1130, A => n2207, ZN => n2217);
   U1754 : AOI22_X1 port map( A1 => n2211, A2 => n5235, B1 => n579, B2 => n2210
                           , ZN => n2212);
   U1755 : OAI221_X1 port map( B1 => n2215, B2 => n1141, C1 => n101, C2 => 
                           n1138, A => n2212, ZN => n2216);
   U1756 : NOR4_X1 port map( A1 => n2219, A2 => n2218, A3 => n2216, A4 => n2217
                           , ZN => n2222);
   U1757 : OAI22_X1 port map( A1 => n4112, A2 => n1160, B1 => n933, B2 => n1159
                           , ZN => n2227);
   U1758 : AOI221_X1 port map( B1 => n1168, B2 => n4819, C1 => n1165, C2 => 
                           n4308, A => n2227, ZN => n2236);
   U1759 : OAI222_X1 port map( A1 => n613, A2 => n1176, B1 => n4117, B2 => 
                           n1173, C1 => n4115, C2 => n876, ZN => n2231);
   U1760 : OAI22_X1 port map( A1 => n4691, A2 => n1188, B1 => n1448, B2 => 
                           n1185, ZN => n2233);
   U1761 : AOI221_X1 port map( B1 => n1195, B2 => n4979, C1 => n1192, C2 => 
                           n4123, A => n2233, ZN => n2234);
   U1762 : NAND4_X1 port map( A1 => n2237, A2 => n2236, A3 => n2234, A4 => 
                           n2235, ZN => n2537);
   U1763 : NAND2_X1 port map( A1 => ADD_RS2(1), A2 => ADD_RS2(2), ZN => n2238);
   U1764 : INV_X1 port map( A => n2238, ZN => n2260);
   U1765 : INV_X1 port map( A => ADD_RS2(2), ZN => n2240);
   U1766 : INV_X1 port map( A => ADD_RS2(0), ZN => n2259);
   U1767 : NAND4_X1 port map( A1 => n980, A2 => n973, A3 => n1274, A4 => n926, 
                           ZN => n4108);
   U1768 : INV_X1 port map( A => ADD_RS2(1), ZN => n2239);
   U1769 : NAND2_X1 port map( A1 => n976, A2 => n878, ZN => n4088);
   U1770 : NAND2_X1 port map( A1 => n2239, A2 => n2240, ZN => n2241);
   U1771 : INV_X1 port map( A => n2241, ZN => n2265);
   U1772 : INV_X1 port map( A => ADD_RS2(4), ZN => n2243);
   U1773 : NAND2_X1 port map( A1 => n975, A2 => n2265, ZN => n4087);
   U1774 : AOI22_X1 port map( A1 => n1200, A2 => n194, B1 => n1198, B2 => n4159
                           , ZN => n2242);
   U1775 : OAI221_X1 port map( B1 => n1207, B2 => n227, C1 => n260, C2 => n1202
                           , A => n2242, ZN => n2252);
   U1776 : NAND2_X1 port map( A1 => n975, A2 => n1036, ZN => n4091);
   U1777 : NAND2_X1 port map( A1 => n7, A2 => n974, ZN => n4090);
   U1778 : AOI22_X1 port map( A1 => n689, A2 => n4223, B1 => n879, B2 => n4191,
                           ZN => n2244);
   U1779 : OAI221_X1 port map( B1 => n388, B2 => n6, C1 => n420, C2 => n1210, A
                           => n2244, ZN => n2251);
   U1780 : NAND2_X1 port map( A1 => n975, A2 => n2260, ZN => n4096);
   U1781 : NAND2_X1 port map( A1 => n2260, A2 => n974, ZN => n4094);
   U1782 : AOI22_X1 port map( A1 => n5108, A2 => n704, B1 => n5140, B2 => n1216
                           , ZN => n2245);
   U1783 : OAI221_X1 port map( B1 => n1223, B2 => n2247, C1 => n1219, C2 => 
                           n2246, A => n2245, ZN => n2250);
   U1784 : NAND2_X1 port map( A1 => n975, A2 => n973, ZN => n4099);
   U1785 : NAND2_X1 port map( A1 => n974, A2 => n973, ZN => n4098);
   U1786 : AOI22_X1 port map( A1 => n5172, A2 => n932, B1 => n5204, B2 => n750,
                           ZN => n2248);
   U1787 : NOR4_X1 port map( A1 => n2252, A2 => n2251, A3 => n2250, A4 => n2249
                           , ZN => n2254);
   U1788 : NAND2_X1 port map( A1 => n1275, A2 => n926, ZN => n4106);
   U1789 : NAND4_X1 port map( A1 => n980, A2 => n703, A3 => n1274, A4 => n925, 
                           ZN => n4105);
   U1790 : OAI222_X1 port map( A1 => n836, A2 => n1237, B1 => n2254, B2 => 
                           n1234, C1 => n1231, C2 => n2253, ZN => n2255);
   U1791 : NAND4_X1 port map( A1 => n980, A2 => n878, A3 => n1274, A4 => n926, 
                           ZN => n4113);
   U1792 : NAND4_X1 port map( A1 => n925, A2 => n2260, A3 => n1274, A4 => n980,
                           ZN => n4111);
   U1793 : OAI22_X1 port map( A1 => n509, A2 => n2257, B1 => n964, B2 => n480, 
                           ZN => n2258);
   U1794 : AOI221_X1 port map( B1 => n4788, B2 => n1255, C1 => n1250, C2 => 
                           n4339, A => n2258, ZN => n2270);
   U1795 : NAND4_X1 port map( A1 => n2264, A2 => n878, A3 => n1274, A4 => n1001
                           , ZN => n4119);
   U1796 : NAND4_X1 port map( A1 => n2264, A2 => n2260, A3 => n1274, A4 => 
                           n1001, ZN => n4118);
   U1797 : NAND4_X1 port map( A1 => n2264, A2 => n973, A3 => n1275, A4 => n979,
                           ZN => n4116);
   U1798 : OAI222_X1 port map( A1 => n644, A2 => n1262, B1 => n1259, B2 => 
                           n2262, C1 => n1258, C2 => n2261, ZN => n2263);
   U1799 : AOI221_X1 port map( B1 => n1268, B2 => n4287, C1 => n1265, C2 => 
                           n4255, A => n2263, ZN => n2269);
   U1800 : NAND3_X1 port map( A1 => n1275, A2 => n893, A3 => n470, ZN => n4121)
                           ;
   U1801 : OAI22_X1 port map( A1 => n4692, A2 => n1275, B1 => n1378, B2 => 
                           n1271, ZN => n2266);
   U1802 : AOI221_X1 port map( B1 => n4948, B2 => n1281, C1 => n1278, C2 => 
                           n2267, A => n2266, ZN => n2268);
   U1803 : NAND4_X1 port map( A1 => n2271, A2 => n2270, A3 => n2269, A4 => 
                           n2268, ZN => n2538);
   U1804 : AOI22_X1 port map( A1 => n1201, A2 => n195, B1 => n495, B2 => n4158,
                           ZN => n2272);
   U1805 : OAI221_X1 port map( B1 => n1206, B2 => n228, C1 => n259, C2 => n1202
                           , A => n2272, ZN => n2281);
   U1806 : AOI22_X1 port map( A1 => n689, A2 => n4222, B1 => n879, B2 => n4190,
                           ZN => n2273);
   U1807 : OAI221_X1 port map( B1 => n387, B2 => n1213, C1 => n419, C2 => n1212
                           , A => n2273, ZN => n2280);
   U1808 : AOI22_X1 port map( A1 => n5109, A2 => n589, B1 => n5141, B2 => n1216
                           , ZN => n2274);
   U1809 : OAI221_X1 port map( B1 => n1222, B2 => n2276, C1 => n1219, C2 => 
                           n2275, A => n2274, ZN => n2279);
   U1810 : AOI22_X1 port map( A1 => n5173, A2 => n2, B1 => n5205, B2 => n931, 
                           ZN => n2277);
   U1811 : NOR4_X1 port map( A1 => n2281, A2 => n2280, A3 => n2279, A4 => n2278
                           , ZN => n2283);
   U1812 : OAI222_X1 port map( A1 => n835, A2 => n1237, B1 => n2283, B2 => 
                           n1234, C1 => n1231, C2 => n2282, ZN => n2284);
   U1813 : OAI22_X1 port map( A1 => n1249, A2 => n2286, B1 => n963, B2 => n1246
                           , ZN => n2287);
   U1814 : AOI221_X1 port map( B1 => n4789, B2 => n33, C1 => n1250, C2 => n4338
                           , A => n2287, ZN => n2295);
   U1815 : OAI222_X1 port map( A1 => n643, A2 => n1262, B1 => n1259, B2 => 
                           n2289, C1 => n1256, C2 => n2288, ZN => n2290);
   U1816 : AOI221_X1 port map( B1 => n1268, B2 => n4286, C1 => n1265, C2 => 
                           n4254, A => n2290, ZN => n2294);
   U1817 : OAI22_X1 port map( A1 => n4693, A2 => n1277, B1 => n1380, B2 => 
                           n1271, ZN => n2291);
   U1818 : AOI221_X1 port map( B1 => n4949, B2 => n1281, C1 => n1278, C2 => 
                           n2292, A => n2291, ZN => n2293);
   U1819 : NAND4_X1 port map( A1 => n2296, A2 => n2295, A3 => n2294, A4 => 
                           n2293, ZN => n2539);
   U1820 : AOI22_X1 port map( A1 => n1200, A2 => n196, B1 => n1196, B2 => n4157
                           , ZN => n2297);
   U1821 : OAI221_X1 port map( B1 => n1207, B2 => n293, C1 => n258, C2 => n1202
                           , A => n2297, ZN => n2306);
   U1822 : AOI22_X1 port map( A1 => n998, A2 => n4221, B1 => n879, B2 => n4189,
                           ZN => n2298);
   U1823 : AOI22_X1 port map( A1 => n5110, A2 => n704, B1 => n5142, B2 => n1216
                           , ZN => n2299);
   U1824 : OAI221_X1 port map( B1 => n1224, B2 => n2301, C1 => n1219, C2 => 
                           n2300, A => n2299, ZN => n2304);
   U1825 : AOI22_X1 port map( A1 => n5174, A2 => n932, B1 => n5206, B2 => n931,
                           ZN => n2302);
   U1826 : OAI221_X1 port map( B1 => n1230, B2 => n173, C1 => n1225, C2 => n322
                           , A => n2302, ZN => n2303);
   U1827 : NOR4_X1 port map( A1 => n2306, A2 => n2303, A3 => n2305, A4 => n2304
                           , ZN => n2308);
   U1828 : OAI222_X1 port map( A1 => n834, A2 => n1237, B1 => n2308, B2 => 
                           n1234, C1 => n1231, C2 => n2307, ZN => n2309);
   U1829 : OAI22_X1 port map( A1 => n1248, A2 => n2311, B1 => n962, B2 => n1246
                           , ZN => n2312);
   U1830 : AOI221_X1 port map( B1 => n4790, B2 => n33, C1 => n1250, C2 => n4337
                           , A => n2312, ZN => n2320);
   U1831 : OAI222_X1 port map( A1 => n642, A2 => n1262, B1 => n1260, B2 => 
                           n2314, C1 => n1256, C2 => n2313, ZN => n2315);
   U1832 : AOI221_X1 port map( B1 => n1268, B2 => n4285, C1 => n1265, C2 => 
                           n4253, A => n2315, ZN => n2319);
   U1833 : OAI22_X1 port map( A1 => n4694, A2 => n1277, B1 => n1382, B2 => 
                           n1271, ZN => n2316);
   U1834 : AOI221_X1 port map( B1 => n4950, B2 => n1281, C1 => n1278, C2 => 
                           n2317, A => n2316, ZN => n2318);
   U1835 : NAND4_X1 port map( A1 => n2321, A2 => n2320, A3 => n2319, A4 => 
                           n2318, ZN => n2540);
   U1836 : AOI22_X1 port map( A1 => n66, A2 => n197, B1 => n1196, B2 => n4156, 
                           ZN => n2322);
   U1837 : OAI221_X1 port map( B1 => n1206, B2 => n294, C1 => n257, C2 => n1202
                           , A => n2322, ZN => n2331);
   U1838 : AOI22_X1 port map( A1 => n998, A2 => n4220, B1 => n879, B2 => n4188,
                           ZN => n2323);
   U1839 : AOI22_X1 port map( A1 => n5111, A2 => n987, B1 => n5143, B2 => n1216
                           , ZN => n2324);
   U1840 : OAI221_X1 port map( B1 => n1222, B2 => n2326, C1 => n1219, C2 => 
                           n2325, A => n2324, ZN => n2329);
   U1841 : AOI22_X1 port map( A1 => n5175, A2 => n1, B1 => n5207, B2 => n40, ZN
                           => n2327);
   U1842 : OAI221_X1 port map( B1 => n1230, B2 => n174, C1 => n1225, C2 => n323
                           , A => n2327, ZN => n2328);
   U1843 : NOR4_X1 port map( A1 => n2331, A2 => n2328, A3 => n2330, A4 => n2329
                           , ZN => n2333);
   U1844 : OAI222_X1 port map( A1 => n833, A2 => n1237, B1 => n2333, B2 => 
                           n1234, C1 => n1231, C2 => n2332, ZN => n2334);
   U1845 : OAI22_X1 port map( A1 => n509, A2 => n2336, B1 => n961, B2 => n1247,
                           ZN => n2337);
   U1846 : OAI22_X1 port map( A1 => n4695, A2 => n1277, B1 => n1384, B2 => 
                           n1271, ZN => n2341);
   U1847 : AOI221_X1 port map( B1 => n4951, B2 => n1281, C1 => n1278, C2 => 
                           n2342, A => n2341, ZN => n2343);
   U1848 : AOI22_X1 port map( A1 => n697, A2 => n198, B1 => n9, B2 => n4155, ZN
                           => n2347);
   U1849 : OAI221_X1 port map( B1 => n1207, B2 => n295, C1 => n256, C2 => n1202
                           , A => n2347, ZN => n2356);
   U1850 : AOI22_X1 port map( A1 => n998, A2 => n4219, B1 => n879, B2 => n4187,
                           ZN => n2348);
   U1851 : OAI221_X1 port map( B1 => n384, B2 => n1215, C1 => n416, C2 => n8, A
                           => n2348, ZN => n2355);
   U1852 : AOI22_X1 port map( A1 => n5112, A2 => n987, B1 => n5144, B2 => n1216
                           , ZN => n2349);
   U1853 : OAI221_X1 port map( B1 => n1224, B2 => n2351, C1 => n1219, C2 => 
                           n2350, A => n2349, ZN => n2354);
   U1854 : AOI22_X1 port map( A1 => n5176, A2 => n1, B1 => n5208, B2 => n750, 
                           ZN => n2352);
   U1855 : NOR4_X1 port map( A1 => n2356, A2 => n2355, A3 => n2354, A4 => n2353
                           , ZN => n2358);
   U1856 : OAI222_X1 port map( A1 => n832, A2 => n1237, B1 => n2358, B2 => 
                           n1234, C1 => n1231, C2 => n2357, ZN => n2359);
   U1857 : OAI22_X1 port map( A1 => n509, A2 => n2361, B1 => n960, B2 => n1246,
                           ZN => n2362);
   U1858 : AOI221_X1 port map( B1 => n4792, B2 => n1254, C1 => n1250, C2 => 
                           n4335, A => n2362, ZN => n2370);
   U1859 : OAI222_X1 port map( A1 => n640, A2 => n1262, B1 => n1259, B2 => 
                           n2364, C1 => n590, C2 => n2363, ZN => n2365);
   U1860 : AOI221_X1 port map( B1 => n1268, B2 => n4283, C1 => n1265, C2 => 
                           n4251, A => n2365, ZN => n2369);
   U1861 : OAI22_X1 port map( A1 => n4696, A2 => n1277, B1 => n1386, B2 => 
                           n1271, ZN => n2366);
   U1862 : AOI221_X1 port map( B1 => n4952, B2 => n1281, C1 => n1278, C2 => 
                           n2367, A => n2366, ZN => n2368);
   U1863 : NAND4_X1 port map( A1 => n2371, A2 => n2370, A3 => n2369, A4 => 
                           n2368, ZN => n2542);
   U1864 : AOI22_X1 port map( A1 => n1200, A2 => n199, B1 => n495, B2 => n4154,
                           ZN => n2372);
   U1865 : OAI221_X1 port map( B1 => n1207, B2 => n296, C1 => n255, C2 => n1202
                           , A => n2372, ZN => n2381);
   U1866 : AOI22_X1 port map( A1 => n998, A2 => n4218, B1 => n879, B2 => n4186,
                           ZN => n2373);
   U1867 : OAI221_X1 port map( B1 => n383, B2 => n6, C1 => n415, C2 => n1212, A
                           => n2373, ZN => n2380);
   U1868 : AOI22_X1 port map( A1 => n5113, A2 => n704, B1 => n5145, B2 => n1216
                           , ZN => n2374);
   U1869 : OAI221_X1 port map( B1 => n1223, B2 => n2376, C1 => n1219, C2 => 
                           n2375, A => n2374, ZN => n2379);
   U1870 : AOI22_X1 port map( A1 => n5177, A2 => n2, B1 => n5209, B2 => n750, 
                           ZN => n2377);
   U1871 : NOR4_X1 port map( A1 => n2381, A2 => n2380, A3 => n2379, A4 => n2378
                           , ZN => n2383);
   U1872 : OAI22_X1 port map( A1 => n498, A2 => n2386, B1 => n959, B2 => n1245,
                           ZN => n2387);
   U1873 : AOI221_X1 port map( B1 => n4793, B2 => n1253, C1 => n1250, C2 => 
                           n4334, A => n2387, ZN => n2395);
   U1874 : OAI222_X1 port map( A1 => n639, A2 => n1262, B1 => n1260, B2 => 
                           n2389, C1 => n590, C2 => n2388, ZN => n2390);
   U1875 : OAI22_X1 port map( A1 => n4697, A2 => n1277, B1 => n1388, B2 => 
                           n1271, ZN => n2391);
   U1876 : AOI221_X1 port map( B1 => n4953, B2 => n1281, C1 => n1278, C2 => 
                           n2392, A => n2391, ZN => n2393);
   U1877 : AOI22_X1 port map( A1 => n1200, A2 => n200, B1 => n9, B2 => n4153, 
                           ZN => n2397);
   U1878 : AOI22_X1 port map( A1 => n998, A2 => n4217, B1 => n879, B2 => n4185,
                           ZN => n2398);
   U1879 : OAI221_X1 port map( B1 => n382, B2 => n1213, C1 => n414, C2 => n8, A
                           => n2398, ZN => n2405);
   U1880 : AOI22_X1 port map( A1 => n5114, A2 => n704, B1 => n5146, B2 => n1216
                           , ZN => n2399);
   U1881 : OAI221_X1 port map( B1 => n1223, B2 => n2401, C1 => n1219, C2 => 
                           n2400, A => n2399, ZN => n2404);
   U1882 : AOI22_X1 port map( A1 => n5178, A2 => n932, B1 => n5210, B2 => n931,
                           ZN => n2402);
   U1883 : NOR4_X1 port map( A1 => n2406, A2 => n2405, A3 => n2403, A4 => n2404
                           , ZN => n2408);
   U1884 : OAI222_X1 port map( A1 => n830, A2 => n1237, B1 => n2408, B2 => 
                           n1234, C1 => n1231, C2 => n2407, ZN => n2409);
   U1885 : OAI22_X1 port map( A1 => n1248, A2 => n2411, B1 => n958, B2 => n480,
                           ZN => n2412);
   U1886 : AOI221_X1 port map( B1 => n4794, B2 => n1255, C1 => n1250, C2 => 
                           n4333, A => n2412, ZN => n2420);
   U1887 : OAI222_X1 port map( A1 => n638, A2 => n1262, B1 => n1260, B2 => 
                           n2414, C1 => n590, C2 => n2413, ZN => n2415);
   U1888 : AOI221_X1 port map( B1 => n1268, B2 => n4281, C1 => n1265, C2 => 
                           n4249, A => n2415, ZN => n2419);
   U1889 : OAI22_X1 port map( A1 => n4698, A2 => n1277, B1 => n1390, B2 => 
                           n1271, ZN => n2416);
   U1890 : AOI221_X1 port map( B1 => n4954, B2 => n1281, C1 => n1278, C2 => 
                           n2417, A => n2416, ZN => n2418);
   U1891 : NAND4_X1 port map( A1 => n2421, A2 => n2418, A3 => n2419, A4 => 
                           n2420, ZN => n2544);
   U1892 : AOI22_X1 port map( A1 => n66, A2 => n201, B1 => n496, B2 => n4152, 
                           ZN => n2422);
   U1893 : OAI221_X1 port map( B1 => n1206, B2 => n298, C1 => n253, C2 => n1202
                           , A => n2422, ZN => n2431);
   U1894 : AOI22_X1 port map( A1 => n998, A2 => n4216, B1 => n879, B2 => n4184,
                           ZN => n2423);
   U1895 : OAI221_X1 port map( B1 => n381, B2 => n1215, C1 => n413, C2 => n1212
                           , A => n2423, ZN => n2430);
   U1896 : AOI22_X1 port map( A1 => n5115, A2 => n589, B1 => n5147, B2 => n1216
                           , ZN => n2424);
   U1897 : OAI221_X1 port map( B1 => n1222, B2 => n2426, C1 => n1219, C2 => 
                           n2425, A => n2424, ZN => n2429);
   U1898 : AOI22_X1 port map( A1 => n5179, A2 => n932, B1 => n5211, B2 => n931,
                           ZN => n2427);
   U1899 : OAI221_X1 port map( B1 => n1230, B2 => n177, C1 => n1225, C2 => n326
                           , A => n2427, ZN => n2428);
   U1900 : NOR4_X1 port map( A1 => n2431, A2 => n2430, A3 => n2428, A4 => n2429
                           , ZN => n2433);
   U1901 : OAI222_X1 port map( A1 => n829, A2 => n1237, B1 => n2433, B2 => 
                           n1234, C1 => n1231, C2 => n2432, ZN => n2434);
   U1902 : OAI22_X1 port map( A1 => n498, A2 => n2436, B1 => n957, B2 => n1245,
                           ZN => n2437);
   U1903 : AOI221_X1 port map( B1 => n4795, B2 => n1253, C1 => n1250, C2 => 
                           n4332, A => n2437, ZN => n2445);
   U1904 : OAI222_X1 port map( A1 => n637, A2 => n1262, B1 => n1259, B2 => 
                           n2439, C1 => n1258, C2 => n2438, ZN => n2440);
   U1905 : OAI22_X1 port map( A1 => n4699, A2 => n1277, B1 => n1392, B2 => 
                           n1271, ZN => n2441);
   U1906 : AOI221_X1 port map( B1 => n4955, B2 => n1281, C1 => n1278, C2 => 
                           n2442, A => n2441, ZN => n2443);
   U1907 : AOI22_X1 port map( A1 => n1201, A2 => n202, B1 => n496, B2 => n4151,
                           ZN => n2447);
   U1908 : OAI221_X1 port map( B1 => n1207, B2 => n299, C1 => n252, C2 => n1202
                           , A => n2447, ZN => n2456);
   U1909 : AOI22_X1 port map( A1 => n998, A2 => n4215, B1 => n879, B2 => n4183,
                           ZN => n2448);
   U1910 : OAI221_X1 port map( B1 => n380, B2 => n1213, C1 => n412, C2 => n1210
                           , A => n2448, ZN => n2455);
   U1911 : AOI22_X1 port map( A1 => n5116, A2 => n987, B1 => n5148, B2 => n1216
                           , ZN => n2449);
   U1912 : OAI221_X1 port map( B1 => n1223, B2 => n2451, C1 => n1219, C2 => 
                           n2450, A => n2449, ZN => n2454);
   U1913 : AOI22_X1 port map( A1 => n5180, A2 => n932, B1 => n5212, B2 => n750,
                           ZN => n2452);
   U1914 : NOR4_X1 port map( A1 => n2456, A2 => n2455, A3 => n2453, A4 => n2454
                           , ZN => n2458);
   U1915 : OAI22_X1 port map( A1 => n498, A2 => n2461, B1 => n956, B2 => n1245,
                           ZN => n2462);
   U1916 : AOI221_X1 port map( B1 => n4796, B2 => n1253, C1 => n1250, C2 => 
                           n4331, A => n2462, ZN => n2470);
   U1917 : OAI222_X1 port map( A1 => n636, A2 => n1262, B1 => n1259, B2 => 
                           n2464, C1 => n1258, C2 => n2463, ZN => n2465);
   U1918 : OAI22_X1 port map( A1 => n4700, A2 => n1277, B1 => n1394, B2 => 
                           n1271, ZN => n2466);
   U1919 : AOI221_X1 port map( B1 => n4956, B2 => n1281, C1 => n1278, C2 => 
                           n2467, A => n2466, ZN => n2468);
   U1920 : AOI22_X1 port map( A1 => n66, A2 => n213, B1 => n9, B2 => n4150, ZN 
                           => n2472);
   U1921 : OAI221_X1 port map( B1 => n1206, B2 => n300, C1 => n251, C2 => n1202
                           , A => n2472, ZN => n2481);
   U1922 : AOI22_X1 port map( A1 => n689, A2 => n4214, B1 => n879, B2 => n4182,
                           ZN => n2473);
   U1923 : OAI221_X1 port map( B1 => n379, B2 => n6, C1 => n411, C2 => n8, A =>
                           n2473, ZN => n2480);
   U1924 : AOI22_X1 port map( A1 => n5117, A2 => n589, B1 => n5149, B2 => n1216
                           , ZN => n2474);
   U1925 : OAI221_X1 port map( B1 => n1222, B2 => n2476, C1 => n1219, C2 => 
                           n2475, A => n2474, ZN => n2479);
   U1926 : AOI22_X1 port map( A1 => n5181, A2 => n932, B1 => n5213, B2 => n40, 
                           ZN => n2477);
   U1927 : OAI221_X1 port map( B1 => n1228, B2 => n179, C1 => n1225, C2 => n328
                           , A => n2477, ZN => n2478);
   U1928 : NOR4_X1 port map( A1 => n2481, A2 => n2478, A3 => n2479, A4 => n2480
                           , ZN => n2483);
   U1929 : OAI222_X1 port map( A1 => n827, A2 => n1237, B1 => n2483, B2 => 
                           n1234, C1 => n1231, C2 => n2482, ZN => n2484);
   U1930 : OAI22_X1 port map( A1 => n498, A2 => n2486, B1 => n955, B2 => n1245,
                           ZN => n2487);
   U1931 : OAI22_X1 port map( A1 => n4701, A2 => n1277, B1 => n1396, B2 => 
                           n1271, ZN => n2491);
   U1932 : AOI221_X1 port map( B1 => n4957, B2 => n1281, C1 => n1278, C2 => 
                           n2492, A => n2491, ZN => n2493);
   U1933 : AOI22_X1 port map( A1 => n1200, A2 => n203, B1 => n1198, B2 => n4149
                           , ZN => n2497);
   U1934 : OAI221_X1 port map( B1 => n1206, B2 => n301, C1 => n250, C2 => n1202
                           , A => n2497, ZN => n3562);
   U1935 : AOI22_X1 port map( A1 => n689, A2 => n4213, B1 => n879, B2 => n4181,
                           ZN => n2498);
   U1936 : OAI221_X1 port map( B1 => n378, B2 => n1213, C1 => n410, C2 => n1210
                           , A => n2498, ZN => n2505);
   U1937 : AOI22_X1 port map( A1 => n5118, A2 => n589, B1 => n5150, B2 => n1216
                           , ZN => n2499);
   U1938 : OAI221_X1 port map( B1 => n1223, B2 => n2501, C1 => n1219, C2 => 
                           n2500, A => n2499, ZN => n2504);
   U1939 : AOI22_X1 port map( A1 => n5182, A2 => n2, B1 => n5214, B2 => n750, 
                           ZN => n2502);
   U1940 : OAI221_X1 port map( B1 => n1228, B2 => n180, C1 => n1225, C2 => n329
                           , A => n2502, ZN => n2503);
   U1941 : NOR4_X1 port map( A1 => n3562, A2 => n2503, A3 => n2505, A4 => n2504
                           , ZN => n3564);
   U1942 : OAI222_X1 port map( A1 => n826, A2 => n1237, B1 => n3564, B2 => 
                           n1234, C1 => n1231, C2 => n3563, ZN => n3565);
   U1943 : OAI22_X1 port map( A1 => n498, A2 => n3567, B1 => n954, B2 => n1245,
                           ZN => n3568);
   U1944 : AOI221_X1 port map( B1 => n4798, B2 => n1253, C1 => n1250, C2 => 
                           n4329, A => n3568, ZN => n3576);
   U1945 : OAI22_X1 port map( A1 => n4702, A2 => n1277, B1 => n1398, B2 => 
                           n1271, ZN => n3572);
   U1946 : AOI221_X1 port map( B1 => n4958, B2 => n1281, C1 => n1278, C2 => 
                           n3573, A => n3572, ZN => n3574);
   U1947 : AOI22_X1 port map( A1 => n697, A2 => n214, B1 => n688, B2 => n4148, 
                           ZN => n3578);
   U1948 : OAI221_X1 port map( B1 => n1206, B2 => n302, C1 => n249, C2 => n1202
                           , A => n3578, ZN => n3587);
   U1949 : AOI22_X1 port map( A1 => n689, A2 => n4212, B1 => n879, B2 => n4180,
                           ZN => n3579);
   U1950 : OAI221_X1 port map( B1 => n377, B2 => n1213, C1 => n409, C2 => n1210
                           , A => n3579, ZN => n3586);
   U1951 : AOI22_X1 port map( A1 => n987, A2 => n5119, B1 => n5151, B2 => n1216
                           , ZN => n3580);
   U1952 : OAI221_X1 port map( B1 => n1223, B2 => n3582, C1 => n1219, C2 => 
                           n3581, A => n3580, ZN => n3585);
   U1953 : AOI22_X1 port map( A1 => n5183, A2 => n1, B1 => n5215, B2 => n750, 
                           ZN => n3583);
   U1954 : NOR4_X1 port map( A1 => n3587, A2 => n3586, A3 => n3585, A4 => n3584
                           , ZN => n3589);
   U1955 : OAI222_X1 port map( A1 => n825, A2 => n1237, B1 => n3589, B2 => 
                           n1234, C1 => n1231, C2 => n3588, ZN => n3590);
   U1956 : OAI22_X1 port map( A1 => n509, A2 => n3592, B1 => n953, B2 => n480, 
                           ZN => n3593);
   U1957 : AOI221_X1 port map( B1 => n4799, B2 => n33, C1 => n1250, C2 => n4328
                           , A => n3593, ZN => n3601);
   U1958 : OAI222_X1 port map( A1 => n633, A2 => n1262, B1 => n1260, B2 => 
                           n3595, C1 => n1258, C2 => n3594, ZN => n3596);
   U1959 : AOI221_X1 port map( B1 => n1268, B2 => n4276, C1 => n1265, C2 => 
                           n4244, A => n3596, ZN => n3600);
   U1960 : OAI22_X1 port map( A1 => n4703, A2 => n1277, B1 => n1400, B2 => 
                           n1271, ZN => n3597);
   U1961 : AOI221_X1 port map( B1 => n4959, B2 => n1281, C1 => n1278, C2 => 
                           n3598, A => n3597, ZN => n3599);
   U1962 : NAND4_X1 port map( A1 => n3602, A2 => n3601, A3 => n3600, A4 => 
                           n3599, ZN => n2549);
   U1963 : AOI22_X1 port map( A1 => n1199, A2 => n215, B1 => n1197, B2 => n4147
                           , ZN => n3603);
   U1964 : AOI22_X1 port map( A1 => n87, A2 => n4211, B1 => n892, B2 => n4179, 
                           ZN => n3604);
   U1965 : AOI22_X1 port map( A1 => n5120, A2 => n589, B1 => n5152, B2 => n1217
                           , ZN => n3605);
   U1966 : OAI221_X1 port map( B1 => n1224, B2 => n3607, C1 => n1220, C2 => 
                           n3606, A => n3605, ZN => n3610);
   U1967 : AOI22_X1 port map( A1 => n2, A2 => n5184, B1 => n5216, B2 => n931, 
                           ZN => n3608);
   U1968 : OAI221_X1 port map( B1 => n1230, B2 => n181, C1 => n1226, C2 => n330
                           , A => n3608, ZN => n3609);
   U1969 : NOR4_X1 port map( A1 => n3611, A2 => n3612, A3 => n3609, A4 => n3610
                           , ZN => n3614);
   U1970 : OAI222_X1 port map( A1 => n824, A2 => n1238, B1 => n3614, B2 => 
                           n1235, C1 => n1232, C2 => n3613, ZN => n3615);
   U1971 : OAI22_X1 port map( A1 => n1249, A2 => n3617, B1 => n952, B2 => n1246
                           , ZN => n3618);
   U1972 : AOI221_X1 port map( B1 => n4800, B2 => n1255, C1 => n1251, C2 => 
                           n4327, A => n3618, ZN => n3626);
   U1973 : OAI222_X1 port map( A1 => n632, A2 => n1263, B1 => n1259, B2 => 
                           n3620, C1 => n590, C2 => n3619, ZN => n3621);
   U1974 : AOI221_X1 port map( B1 => n1269, B2 => n4275, C1 => n1266, C2 => 
                           n4243, A => n3621, ZN => n3625);
   U1975 : OAI22_X1 port map( A1 => n4704, A2 => n1277, B1 => n1402, B2 => 
                           n1272, ZN => n3622);
   U1976 : AOI221_X1 port map( B1 => n4960, B2 => n1282, C1 => n1279, C2 => 
                           n3623, A => n3622, ZN => n3624);
   U1977 : NAND4_X1 port map( A1 => n3627, A2 => n3626, A3 => n3625, A4 => 
                           n3624, ZN => n2550);
   U1978 : AOI22_X1 port map( A1 => n697, A2 => n216, B1 => n688, B2 => n4146, 
                           ZN => n3628);
   U1979 : AOI22_X1 port map( A1 => n998, A2 => n4210, B1 => n1208, B2 => n4178
                           , ZN => n3629);
   U1980 : OAI221_X1 port map( B1 => n375, B2 => n1215, C1 => n407, C2 => n1210
                           , A => n3629, ZN => n3636);
   U1981 : AOI22_X1 port map( A1 => n5121, A2 => n704, B1 => n5153, B2 => n1217
                           , ZN => n3630);
   U1982 : OAI221_X1 port map( B1 => n1222, B2 => n3632, C1 => n1220, C2 => 
                           n3631, A => n3630, ZN => n3635);
   U1983 : AOI22_X1 port map( A1 => n5185, A2 => n1, B1 => n5217, B2 => n750, 
                           ZN => n3633);
   U1984 : NOR4_X1 port map( A1 => n3637, A2 => n3636, A3 => n3634, A4 => n3635
                           , ZN => n3639);
   U1985 : OAI222_X1 port map( A1 => n823, A2 => n1238, B1 => n3639, B2 => 
                           n1235, C1 => n1232, C2 => n3638, ZN => n3640);
   U1986 : OAI22_X1 port map( A1 => n1248, A2 => n3642, B1 => n951, B2 => n480,
                           ZN => n3643);
   U1987 : AOI221_X1 port map( B1 => n4801, B2 => n33, C1 => n1251, C2 => n4326
                           , A => n3643, ZN => n3651);
   U1988 : OAI222_X1 port map( A1 => n631, A2 => n1263, B1 => n1259, B2 => 
                           n3645, C1 => n590, C2 => n3644, ZN => n3646);
   U1989 : AOI221_X1 port map( B1 => n1269, B2 => n4274, C1 => n1266, C2 => 
                           n4242, A => n3646, ZN => n3650);
   U1990 : OAI22_X1 port map( A1 => n4705, A2 => n1277, B1 => n1404, B2 => 
                           n1272, ZN => n3647);
   U1991 : AOI221_X1 port map( B1 => n4961, B2 => n1282, C1 => n1279, C2 => 
                           n3648, A => n3647, ZN => n3649);
   U1992 : NAND4_X1 port map( A1 => n3652, A2 => n3649, A3 => n3650, A4 => 
                           n3651, ZN => n2551);
   U1993 : AOI22_X1 port map( A1 => n697, A2 => n217, B1 => n496, B2 => n4145, 
                           ZN => n3653);
   U1994 : OAI221_X1 port map( B1 => n1206, B2 => n304, C1 => n246, C2 => n1203
                           , A => n3653, ZN => n3662);
   U1995 : AOI22_X1 port map( A1 => n689, A2 => n4209, B1 => n1209, B2 => n4177
                           , ZN => n3654);
   U1996 : OAI221_X1 port map( B1 => n374, B2 => n6, C1 => n406, C2 => n8, A =>
                           n3654, ZN => n3661);
   U1997 : AOI22_X1 port map( A1 => n5122, A2 => n987, B1 => n5154, B2 => n1217
                           , ZN => n3655);
   U1998 : OAI221_X1 port map( B1 => n1223, B2 => n3657, C1 => n1220, C2 => 
                           n3656, A => n3655, ZN => n3660);
   U1999 : AOI22_X1 port map( A1 => n5186, A2 => n932, B1 => n5218, B2 => n40, 
                           ZN => n3658);
   U2000 : NOR4_X1 port map( A1 => n3662, A2 => n3661, A3 => n3659, A4 => n3660
                           , ZN => n3664);
   U2001 : OAI222_X1 port map( A1 => n822, A2 => n1238, B1 => n3664, B2 => 
                           n1235, C1 => n1232, C2 => n3663, ZN => n3665);
   U2002 : OAI22_X1 port map( A1 => n509, A2 => n3667, B1 => n950, B2 => n1247,
                           ZN => n3668);
   U2003 : AOI221_X1 port map( B1 => n4802, B2 => n1254, C1 => n1251, C2 => 
                           n4325, A => n3668, ZN => n3676);
   U2004 : OAI222_X1 port map( A1 => n630, A2 => n1263, B1 => n1260, B2 => 
                           n3670, C1 => n1258, C2 => n3669, ZN => n3671);
   U2005 : AOI221_X1 port map( B1 => n1269, B2 => n4273, C1 => n1266, C2 => 
                           n4241, A => n3671, ZN => n3675);
   U2006 : OAI22_X1 port map( A1 => n4706, A2 => n1276, B1 => n1406, B2 => 
                           n1272, ZN => n3672);
   U2007 : AOI221_X1 port map( B1 => n4962, B2 => n1282, C1 => n1279, C2 => 
                           n3673, A => n3672, ZN => n3674);
   U2008 : NAND4_X1 port map( A1 => n3677, A2 => n3676, A3 => n3675, A4 => 
                           n3674, ZN => n2552);
   U2009 : AOI22_X1 port map( A1 => n1199, A2 => n204, B1 => n1198, B2 => n4144
                           , ZN => n3678);
   U2010 : OAI221_X1 port map( B1 => n1207, B2 => n305, C1 => n245, C2 => n1203
                           , A => n3678, ZN => n3687);
   U2011 : AOI22_X1 port map( A1 => n998, A2 => n4208, B1 => n1208, B2 => n4176
                           , ZN => n3679);
   U2012 : AOI22_X1 port map( A1 => n5123, A2 => n704, B1 => n5155, B2 => n1217
                           , ZN => n3680);
   U2013 : OAI221_X1 port map( B1 => n1224, B2 => n3682, C1 => n1220, C2 => 
                           n3681, A => n3680, ZN => n3685);
   U2014 : AOI22_X1 port map( A1 => n5187, A2 => n710, B1 => n5219, B2 => n40, 
                           ZN => n3683);
   U2015 : OAI221_X1 port map( B1 => n1229, B2 => n183, C1 => n1226, C2 => n332
                           , A => n3683, ZN => n3684);
   U2016 : NOR4_X1 port map( A1 => n3687, A2 => n3685, A3 => n3686, A4 => n3684
                           , ZN => n3689);
   U2017 : OAI22_X1 port map( A1 => n1249, A2 => n3692, B1 => n949, B2 => n1246
                           , ZN => n3693);
   U2018 : AOI221_X1 port map( B1 => n4803, B2 => n1255, C1 => n1251, C2 => 
                           n4324, A => n3693, ZN => n3701);
   U2019 : OAI222_X1 port map( A1 => n629, A2 => n1263, B1 => n1260, B2 => 
                           n3695, C1 => n1258, C2 => n3694, ZN => n3696);
   U2020 : AOI221_X1 port map( B1 => n1269, B2 => n4272, C1 => n1266, C2 => 
                           n4240, A => n3696, ZN => n3700);
   U2021 : OAI22_X1 port map( A1 => n4707, A2 => n1276, B1 => n1408, B2 => 
                           n1272, ZN => n3697);
   U2022 : AOI221_X1 port map( B1 => n4963, B2 => n1282, C1 => n1279, C2 => 
                           n3698, A => n3697, ZN => n3699);
   U2023 : NAND4_X1 port map( A1 => n3702, A2 => n3699, A3 => n3700, A4 => 
                           n3701, ZN => n2553);
   U2024 : AOI22_X1 port map( A1 => n1200, A2 => n205, B1 => n495, B2 => n4143,
                           ZN => n3703);
   U2025 : OAI221_X1 port map( B1 => n1207, B2 => n306, C1 => n244, C2 => n1203
                           , A => n3703, ZN => n3712);
   U2026 : AOI22_X1 port map( A1 => n998, A2 => n4207, B1 => n1208, B2 => n4175
                           , ZN => n3704);
   U2027 : OAI221_X1 port map( B1 => n372, B2 => n1213, C1 => n404, C2 => n8, A
                           => n3704, ZN => n3711);
   U2028 : AOI22_X1 port map( A1 => n5124, A2 => n704, B1 => n5156, B2 => n1217
                           , ZN => n3705);
   U2029 : OAI221_X1 port map( B1 => n1224, B2 => n3707, C1 => n1220, C2 => 
                           n3706, A => n3705, ZN => n3710);
   U2030 : AOI22_X1 port map( A1 => n5188, A2 => n1, B1 => n5220, B2 => n931, 
                           ZN => n3708);
   U2031 : NOR4_X1 port map( A1 => n3712, A2 => n3711, A3 => n3710, A4 => n3709
                           , ZN => n3714);
   U2032 : OAI222_X1 port map( A1 => n820, A2 => n1238, B1 => n3714, B2 => 
                           n1235, C1 => n1232, C2 => n3713, ZN => n3715);
   U2033 : OAI22_X1 port map( A1 => n509, A2 => n3717, B1 => n948, B2 => n1247,
                           ZN => n3718);
   U2034 : AOI221_X1 port map( B1 => n4804, B2 => n33, C1 => n1251, C2 => n4323
                           , A => n3718, ZN => n3726);
   U2035 : OAI222_X1 port map( A1 => n628, A2 => n1263, B1 => n1259, B2 => 
                           n3720, C1 => n1256, C2 => n3719, ZN => n3721);
   U2036 : AOI221_X1 port map( B1 => n1269, B2 => n4271, C1 => n1266, C2 => 
                           n4239, A => n3721, ZN => n3725);
   U2037 : OAI22_X1 port map( A1 => n4708, A2 => n1276, B1 => n1410, B2 => 
                           n1272, ZN => n3722);
   U2038 : AOI221_X1 port map( B1 => n4964, B2 => n1282, C1 => n1279, C2 => 
                           n3723, A => n3722, ZN => n3724);
   U2039 : NAND4_X1 port map( A1 => n3727, A2 => n3726, A3 => n3725, A4 => 
                           n3724, ZN => n2554);
   U2040 : AOI22_X1 port map( A1 => n697, A2 => n206, B1 => n495, B2 => n4142, 
                           ZN => n3728);
   U2041 : OAI221_X1 port map( B1 => n1206, B2 => n307, C1 => n243, C2 => n1203
                           , A => n3728, ZN => n3737);
   U2042 : AOI22_X1 port map( A1 => n998, A2 => n4206, B1 => n1209, B2 => n4174
                           , ZN => n3729);
   U2043 : OAI221_X1 port map( B1 => n371, B2 => n6, C1 => n403, C2 => n1210, A
                           => n3729, ZN => n3736);
   U2044 : AOI22_X1 port map( A1 => n5125, A2 => n987, B1 => n5157, B2 => n1217
                           , ZN => n3730);
   U2045 : OAI221_X1 port map( B1 => n1222, B2 => n3732, C1 => n1220, C2 => 
                           n3731, A => n3730, ZN => n3735);
   U2046 : AOI22_X1 port map( A1 => n5189, A2 => n2, B1 => n5221, B2 => n40, ZN
                           => n3733);
   U2047 : NOR4_X1 port map( A1 => n3737, A2 => n3736, A3 => n3735, A4 => n3734
                           , ZN => n3739);
   U2048 : OAI222_X1 port map( A1 => n819, A2 => n1238, B1 => n3739, B2 => 
                           n1235, C1 => n1232, C2 => n3738, ZN => n3740);
   U2049 : OAI22_X1 port map( A1 => n509, A2 => n3742, B1 => n947, B2 => n1246,
                           ZN => n3743);
   U2050 : AOI221_X1 port map( B1 => n4805, B2 => n33, C1 => n1251, C2 => n4322
                           , A => n3743, ZN => n3751);
   U2051 : OAI222_X1 port map( A1 => n627, A2 => n1263, B1 => n1260, B2 => 
                           n3745, C1 => n1258, C2 => n3744, ZN => n3746);
   U2052 : AOI221_X1 port map( B1 => n1269, B2 => n4270, C1 => n1266, C2 => 
                           n4238, A => n3746, ZN => n3750);
   U2053 : OAI22_X1 port map( A1 => n4709, A2 => n1276, B1 => n1412, B2 => 
                           n1272, ZN => n3747);
   U2054 : AOI221_X1 port map( B1 => n4965, B2 => n1282, C1 => n1279, C2 => 
                           n3748, A => n3747, ZN => n3749);
   U2055 : NAND4_X1 port map( A1 => n3752, A2 => n3751, A3 => n3750, A4 => 
                           n3749, ZN => n2555);
   U2056 : AOI22_X1 port map( A1 => n66, A2 => n207, B1 => n495, B2 => n4141, 
                           ZN => n3753);
   U2057 : AOI22_X1 port map( A1 => n998, A2 => n4205, B1 => n1208, B2 => n4173
                           , ZN => n3754);
   U2058 : OAI221_X1 port map( B1 => n370, B2 => n6, C1 => n402, C2 => n1212, A
                           => n3754, ZN => n3761);
   U2059 : AOI22_X1 port map( A1 => n589, A2 => n5126, B1 => n5158, B2 => n1217
                           , ZN => n3755);
   U2060 : OAI221_X1 port map( B1 => n1224, B2 => n3757, C1 => n1220, C2 => 
                           n3756, A => n3755, ZN => n3760);
   U2061 : AOI22_X1 port map( A1 => n5190, A2 => n932, B1 => n5222, B2 => n750,
                           ZN => n3758);
   U2062 : NOR4_X1 port map( A1 => n3762, A2 => n3761, A3 => n3759, A4 => n3760
                           , ZN => n3764);
   U2063 : OAI222_X1 port map( A1 => n818, A2 => n1238, B1 => n3764, B2 => 
                           n1235, C1 => n1232, C2 => n3763, ZN => n3765);
   U2064 : OAI22_X1 port map( A1 => n1248, A2 => n3767, B1 => n946, B2 => n1246
                           , ZN => n3768);
   U2065 : AOI221_X1 port map( B1 => n4806, B2 => n1254, C1 => n1251, C2 => 
                           n4321, A => n3768, ZN => n3776);
   U2066 : OAI222_X1 port map( A1 => n626, A2 => n1263, B1 => n1259, B2 => 
                           n3770, C1 => n1258, C2 => n3769, ZN => n3771);
   U2067 : AOI221_X1 port map( B1 => n1269, B2 => n4269, C1 => n1266, C2 => 
                           n4237, A => n3771, ZN => n3775);
   U2068 : OAI22_X1 port map( A1 => n4710, A2 => n1276, B1 => n1414, B2 => 
                           n1272, ZN => n3772);
   U2069 : AOI221_X1 port map( B1 => n4966, B2 => n1282, C1 => n1279, C2 => 
                           n3773, A => n3772, ZN => n3774);
   U2070 : NAND4_X1 port map( A1 => n3777, A2 => n3774, A3 => n3775, A4 => 
                           n3776, ZN => n2556);
   U2071 : AOI22_X1 port map( A1 => n1201, A2 => n208, B1 => n688, B2 => n4140,
                           ZN => n3778);
   U2072 : OAI221_X1 port map( B1 => n1206, B2 => n309, C1 => n241, C2 => n1203
                           , A => n3778, ZN => n3787);
   U2073 : AOI22_X1 port map( A1 => n689, A2 => n4204, B1 => n1208, B2 => n4172
                           , ZN => n3779);
   U2074 : OAI221_X1 port map( B1 => n369, B2 => n1213, C1 => n401, C2 => n8, A
                           => n3779, ZN => n3786);
   U2075 : AOI22_X1 port map( A1 => n5127, A2 => n987, B1 => n5159, B2 => n1217
                           , ZN => n3780);
   U2076 : OAI221_X1 port map( B1 => n1223, B2 => n3782, C1 => n1220, C2 => 
                           n3781, A => n3780, ZN => n3785);
   U2077 : AOI22_X1 port map( A1 => n5191, A2 => n2, B1 => n5223, B2 => n750, 
                           ZN => n3783);
   U2078 : NOR4_X1 port map( A1 => n3787, A2 => n3786, A3 => n3785, A4 => n3784
                           , ZN => n3789);
   U2079 : OAI222_X1 port map( A1 => n817, A2 => n1238, B1 => n3789, B2 => 
                           n1235, C1 => n1232, C2 => n3788, ZN => n3790);
   U2080 : OAI22_X1 port map( A1 => n509, A2 => n3792, B1 => n945, B2 => n480, 
                           ZN => n3793);
   U2081 : AOI221_X1 port map( B1 => n4807, B2 => n1255, C1 => n1251, C2 => 
                           n4320, A => n3793, ZN => n3801);
   U2082 : OAI222_X1 port map( A1 => n625, A2 => n1263, B1 => n1259, B2 => 
                           n3795, C1 => n590, C2 => n3794, ZN => n3796);
   U2083 : AOI221_X1 port map( B1 => n1269, B2 => n4268, C1 => n1266, C2 => 
                           n4236, A => n3796, ZN => n3800);
   U2084 : OAI22_X1 port map( A1 => n4711, A2 => n1276, B1 => n1416, B2 => 
                           n1272, ZN => n3797);
   U2085 : AOI221_X1 port map( B1 => n4967, B2 => n1282, C1 => n1279, C2 => 
                           n3798, A => n3797, ZN => n3799);
   U2086 : NAND4_X1 port map( A1 => n3802, A2 => n3801, A3 => n3800, A4 => 
                           n3799, ZN => n2557);
   U2087 : AOI22_X1 port map( A1 => n1200, A2 => n209, B1 => n1196, B2 => n4139
                           , ZN => n3803);
   U2088 : OAI221_X1 port map( B1 => n1206, B2 => n310, C1 => n240, C2 => n1203
                           , A => n3803, ZN => n3812);
   U2089 : AOI22_X1 port map( A1 => n689, A2 => n4203, B1 => n1209, B2 => n4171
                           , ZN => n3804);
   U2090 : OAI221_X1 port map( B1 => n368, B2 => n1215, C1 => n400, C2 => n1212
                           , A => n3804, ZN => n3811);
   U2091 : AOI22_X1 port map( A1 => n5128, A2 => n589, B1 => n5160, B2 => n1217
                           , ZN => n3805);
   U2092 : OAI221_X1 port map( B1 => n1224, B2 => n3807, C1 => n1220, C2 => 
                           n3806, A => n3805, ZN => n3810);
   U2093 : AOI22_X1 port map( A1 => n5192, A2 => n1, B1 => n5224, B2 => n750, 
                           ZN => n3808);
   U2094 : NOR4_X1 port map( A1 => n3812, A2 => n3811, A3 => n3810, A4 => n3809
                           , ZN => n3814);
   U2095 : OAI222_X1 port map( A1 => n816, A2 => n1238, B1 => n3814, B2 => 
                           n1235, C1 => n1232, C2 => n3813, ZN => n3815);
   U2096 : OAI22_X1 port map( A1 => n1249, A2 => n3817, B1 => n944, B2 => n480,
                           ZN => n3818);
   U2097 : AOI221_X1 port map( B1 => n4808, B2 => n33, C1 => n1251, C2 => n4319
                           , A => n3818, ZN => n3826);
   U2098 : OAI222_X1 port map( A1 => n624, A2 => n1263, B1 => n1259, B2 => 
                           n3820, C1 => n590, C2 => n3819, ZN => n3821);
   U2099 : AOI221_X1 port map( B1 => n1269, B2 => n4267, C1 => n1266, C2 => 
                           n4235, A => n3821, ZN => n3825);
   U2100 : OAI22_X1 port map( A1 => n4712, A2 => n1276, B1 => n1418, B2 => 
                           n1272, ZN => n3822);
   U2101 : AOI221_X1 port map( B1 => n4968, B2 => n1282, C1 => n1279, C2 => 
                           n3823, A => n3822, ZN => n3824);
   U2102 : NAND4_X1 port map( A1 => n3827, A2 => n3826, A3 => n3825, A4 => 
                           n3824, ZN => n2558);
   U2103 : AOI22_X1 port map( A1 => n66, A2 => n210, B1 => n688, B2 => n4138, 
                           ZN => n3828);
   U2104 : OAI221_X1 port map( B1 => n1207, B2 => n311, C1 => n239, C2 => n1203
                           , A => n3828, ZN => n3837);
   U2105 : AOI22_X1 port map( A1 => n998, A2 => n4202, B1 => n1208, B2 => n4170
                           , ZN => n3829);
   U2106 : OAI221_X1 port map( B1 => n367, B2 => n6, C1 => n399, C2 => n1210, A
                           => n3829, ZN => n3836);
   U2107 : AOI22_X1 port map( A1 => n5129, A2 => n589, B1 => n5161, B2 => n1217
                           , ZN => n3830);
   U2108 : OAI221_X1 port map( B1 => n1222, B2 => n3832, C1 => n1220, C2 => 
                           n3831, A => n3830, ZN => n3835);
   U2109 : AOI22_X1 port map( A1 => n5193, A2 => n932, B1 => n5225, B2 => n40, 
                           ZN => n3833);
   U2110 : NOR4_X1 port map( A1 => n3837, A2 => n3836, A3 => n3835, A4 => n3834
                           , ZN => n3839);
   U2111 : OAI222_X1 port map( A1 => n815, A2 => n1238, B1 => n3839, B2 => 
                           n1235, C1 => n1232, C2 => n3838, ZN => n3840);
   U2112 : OAI22_X1 port map( A1 => n1248, A2 => n3842, B1 => n943, B2 => n480,
                           ZN => n3843);
   U2113 : AOI221_X1 port map( B1 => n4809, B2 => n33, C1 => n1251, C2 => n4318
                           , A => n3843, ZN => n3851);
   U2114 : OAI222_X1 port map( A1 => n623, A2 => n1263, B1 => n1260, B2 => 
                           n3845, C1 => n1258, C2 => n3844, ZN => n3846);
   U2115 : AOI221_X1 port map( B1 => n1269, B2 => n4266, C1 => n1266, C2 => 
                           n4234, A => n3846, ZN => n3850);
   U2116 : OAI22_X1 port map( A1 => n4713, A2 => n1276, B1 => n1420, B2 => 
                           n1272, ZN => n3847);
   U2117 : AOI221_X1 port map( B1 => n4969, B2 => n1282, C1 => n1279, C2 => 
                           n3848, A => n3847, ZN => n3849);
   U2118 : NAND4_X1 port map( A1 => n3852, A2 => n3851, A3 => n3850, A4 => 
                           n3849, ZN => n2559);
   U2119 : AOI22_X1 port map( A1 => n66, A2 => n211, B1 => n496, B2 => n4137, 
                           ZN => n3853);
   U2120 : OAI221_X1 port map( B1 => n1207, B2 => n312, C1 => n238, C2 => n1203
                           , A => n3853, ZN => n3862);
   U2121 : AOI22_X1 port map( A1 => n998, A2 => n4201, B1 => n1209, B2 => n4169
                           , ZN => n3854);
   U2122 : OAI221_X1 port map( B1 => n366, B2 => n1215, C1 => n398, C2 => n8, A
                           => n3854, ZN => n3861);
   U2123 : AOI22_X1 port map( A1 => n5130, A2 => n704, B1 => n5162, B2 => n1217
                           , ZN => n3855);
   U2124 : OAI221_X1 port map( B1 => n1223, B2 => n3857, C1 => n1220, C2 => 
                           n3856, A => n3855, ZN => n3860);
   U2125 : AOI22_X1 port map( A1 => n5194, A2 => n932, B1 => n5226, B2 => n931,
                           ZN => n3858);
   U2126 : NOR4_X1 port map( A1 => n3862, A2 => n3861, A3 => n3860, A4 => n3859
                           , ZN => n3864);
   U2127 : OAI222_X1 port map( A1 => n814, A2 => n1238, B1 => n3864, B2 => 
                           n1235, C1 => n1232, C2 => n3863, ZN => n3865);
   U2128 : OAI22_X1 port map( A1 => n509, A2 => n3867, B1 => n942, B2 => n1246,
                           ZN => n3868);
   U2129 : AOI221_X1 port map( B1 => n4810, B2 => n33, C1 => n1251, C2 => n4317
                           , A => n3868, ZN => n3876);
   U2130 : OAI222_X1 port map( A1 => n622, A2 => n1263, B1 => n1260, B2 => 
                           n3870, C1 => n1258, C2 => n3869, ZN => n3871);
   U2131 : AOI221_X1 port map( B1 => n1269, B2 => n4265, C1 => n1266, C2 => 
                           n4233, A => n3871, ZN => n3875);
   U2132 : OAI22_X1 port map( A1 => n4714, A2 => n1276, B1 => n1422, B2 => 
                           n1272, ZN => n3872);
   U2133 : AOI221_X1 port map( B1 => n4970, B2 => n1282, C1 => n1279, C2 => 
                           n3873, A => n3872, ZN => n3874);
   U2134 : NAND4_X1 port map( A1 => n3877, A2 => n3876, A3 => n3875, A4 => 
                           n3874, ZN => n2560);
   U2135 : AOI22_X1 port map( A1 => n697, A2 => n212, B1 => n496, B2 => n4136, 
                           ZN => n3878);
   U2136 : AOI22_X1 port map( A1 => n998, A2 => n4200, B1 => n1209, B2 => n4168
                           , ZN => n3879);
   U2137 : OAI221_X1 port map( B1 => n365, B2 => n1213, C1 => n397, C2 => n1210
                           , A => n3879, ZN => n3886);
   U2138 : AOI22_X1 port map( A1 => n5131, A2 => n589, B1 => n5163, B2 => n1217
                           , ZN => n3880);
   U2139 : OAI221_X1 port map( B1 => n1222, B2 => n3882, C1 => n1220, C2 => 
                           n3881, A => n3880, ZN => n3885);
   U2140 : AOI22_X1 port map( A1 => n5195, A2 => n932, B1 => n5227, B2 => n40, 
                           ZN => n3883);
   U2141 : NOR4_X1 port map( A1 => n3887, A2 => n3886, A3 => n3884, A4 => n3885
                           , ZN => n3889);
   U2142 : OAI222_X1 port map( A1 => n813, A2 => n1238, B1 => n3889, B2 => 
                           n1235, C1 => n1232, C2 => n3888, ZN => n3890);
   U2143 : OAI22_X1 port map( A1 => n1248, A2 => n3892, B1 => n941, B2 => n1246
                           , ZN => n3893);
   U2144 : AOI221_X1 port map( B1 => n4811, B2 => n33, C1 => n1251, C2 => n4316
                           , A => n3893, ZN => n3901);
   U2145 : OAI222_X1 port map( A1 => n621, A2 => n1263, B1 => n1260, B2 => 
                           n3895, C1 => n1256, C2 => n3894, ZN => n3896);
   U2146 : AOI221_X1 port map( B1 => n1269, B2 => n4264, C1 => n1266, C2 => 
                           n4232, A => n3896, ZN => n3900);
   U2147 : OAI22_X1 port map( A1 => n4715, A2 => n1276, B1 => n1424, B2 => 
                           n1272, ZN => n3897);
   U2148 : AOI221_X1 port map( B1 => n4971, B2 => n1282, C1 => n1279, C2 => 
                           n3898, A => n3897, ZN => n3899);
   U2149 : NAND4_X1 port map( A1 => n3902, A2 => n3899, A3 => n3900, A4 => 
                           n3901, ZN => n2561);
   U2150 : AOI22_X1 port map( A1 => n66, A2 => n3903, B1 => n9, B2 => n4135, ZN
                           => n3904);
   U2151 : OAI221_X1 port map( B1 => n1207, B2 => n314, C1 => n236, C2 => n1204
                           , A => n3904, ZN => n3913);
   U2152 : AOI22_X1 port map( A1 => n998, A2 => n4199, B1 => n1209, B2 => n4167
                           , ZN => n3905);
   U2153 : OAI221_X1 port map( B1 => n364, B2 => n6, C1 => n396, C2 => n8, A =>
                           n3905, ZN => n3912);
   U2154 : AOI22_X1 port map( A1 => n5132, A2 => n704, B1 => n5164, B2 => n1218
                           , ZN => n3906);
   U2155 : OAI221_X1 port map( B1 => n1224, B2 => n3908, C1 => n1221, C2 => 
                           n3907, A => n3906, ZN => n3911);
   U2156 : AOI22_X1 port map( A1 => n5196, A2 => n2, B1 => n5228, B2 => n931, 
                           ZN => n3909);
   U2157 : NOR4_X1 port map( A1 => n3913, A2 => n3912, A3 => n3910, A4 => n3911
                           , ZN => n3915);
   U2158 : OAI22_X1 port map( A1 => n509, A2 => n3918, B1 => n940, B2 => n1247,
                           ZN => n3919);
   U2159 : AOI221_X1 port map( B1 => n4812, B2 => n1254, C1 => n1252, C2 => 
                           n4315, A => n3919, ZN => n3927);
   U2160 : OAI22_X1 port map( A1 => n4716, A2 => n1276, B1 => n1427, B2 => 
                           n1273, ZN => n3923);
   U2161 : AOI221_X1 port map( B1 => n4972, B2 => n1283, C1 => n1280, C2 => 
                           n3924, A => n3923, ZN => n3925);
   U2162 : AOI22_X1 port map( A1 => n1199, A2 => n3929, B1 => n1197, B2 => 
                           n4134, ZN => n3930);
   U2163 : OAI221_X1 port map( B1 => n1207, B2 => n315, C1 => n235, C2 => n1204
                           , A => n3930, ZN => n3939);
   U2164 : AOI22_X1 port map( A1 => n998, A2 => n4198, B1 => n1209, B2 => n4166
                           , ZN => n3931);
   U2165 : OAI221_X1 port map( B1 => n363, B2 => n6, C1 => n395, C2 => n1210, A
                           => n3931, ZN => n3938);
   U2166 : AOI22_X1 port map( A1 => n987, A2 => n5133, B1 => n5165, B2 => n1218
                           , ZN => n3932);
   U2167 : OAI221_X1 port map( B1 => n1223, B2 => n3934, C1 => n1221, C2 => 
                           n3933, A => n3932, ZN => n3937);
   U2168 : AOI22_X1 port map( A1 => n5197, A2 => n1, B1 => n5229, B2 => n40, ZN
                           => n3935);
   U2169 : NOR4_X1 port map( A1 => n3939, A2 => n3938, A3 => n3937, A4 => n3936
                           , ZN => n3941);
   U2170 : OAI222_X1 port map( A1 => n811, A2 => n1239, B1 => n3941, B2 => 
                           n1236, C1 => n1233, C2 => n3940, ZN => n3942);
   U2171 : OAI22_X1 port map( A1 => n1249, A2 => n3944, B1 => n939, B2 => n1247
                           , ZN => n3945);
   U2172 : AOI221_X1 port map( B1 => n4813, B2 => n1255, C1 => n1252, C2 => 
                           n4314, A => n3945, ZN => n3953);
   U2173 : OAI22_X1 port map( A1 => n4717, A2 => n1275, B1 => n1430, B2 => 
                           n1273, ZN => n3949);
   U2174 : AOI221_X1 port map( B1 => n4973, B2 => n1283, C1 => n1280, C2 => 
                           n3950, A => n3949, ZN => n3951);
   U2175 : AOI22_X1 port map( A1 => n697, A2 => n3955, B1 => n688, B2 => n4133,
                           ZN => n3956);
   U2176 : OAI221_X1 port map( B1 => n1206, B2 => n316, C1 => n234, C2 => n1204
                           , A => n3956, ZN => n3965);
   U2177 : AOI22_X1 port map( A1 => n689, A2 => n4197, B1 => n1208, B2 => n4165
                           , ZN => n3957);
   U2178 : OAI221_X1 port map( B1 => n362, B2 => n1213, C1 => n394, C2 => n8, A
                           => n3957, ZN => n3964);
   U2179 : AOI22_X1 port map( A1 => n5134, A2 => n987, B1 => n5166, B2 => n1218
                           , ZN => n3958);
   U2180 : OAI221_X1 port map( B1 => n1224, B2 => n3960, C1 => n1221, C2 => 
                           n3959, A => n3958, ZN => n3963);
   U2181 : AOI22_X1 port map( A1 => n5198, A2 => n2, B1 => n5230, B2 => n750, 
                           ZN => n3961);
   U2182 : OAI221_X1 port map( B1 => n1228, B2 => n188, C1 => n1227, C2 => n337
                           , A => n3961, ZN => n3962);
   U2183 : NOR4_X1 port map( A1 => n3965, A2 => n3962, A3 => n3964, A4 => n3963
                           , ZN => n3967);
   U2184 : OAI22_X1 port map( A1 => n1248, A2 => n3970, B1 => n938, B2 => n1246
                           , ZN => n3971);
   U2185 : AOI221_X1 port map( B1 => n4814, B2 => n33, C1 => n1252, C2 => n4313
                           , A => n3971, ZN => n3979);
   U2186 : OAI22_X1 port map( A1 => n4718, A2 => n1275, B1 => n1433, B2 => 
                           n1273, ZN => n3975);
   U2187 : AOI221_X1 port map( B1 => n4974, B2 => n1283, C1 => n1280, C2 => 
                           n3976, A => n3975, ZN => n3977);
   U2188 : AOI22_X1 port map( A1 => n1201, A2 => n3981, B1 => n9, B2 => n4132, 
                           ZN => n3982);
   U2189 : OAI221_X1 port map( B1 => n1207, B2 => n317, C1 => n233, C2 => n1204
                           , A => n3982, ZN => n3991);
   U2190 : AOI22_X1 port map( A1 => n998, A2 => n4196, B1 => n1209, B2 => n4164
                           , ZN => n3983);
   U2191 : OAI221_X1 port map( B1 => n361, B2 => n1213, C1 => n393, C2 => n1212
                           , A => n3983, ZN => n3990);
   U2192 : AOI22_X1 port map( A1 => n5135, A2 => n987, B1 => n5167, B2 => n1218
                           , ZN => n3984);
   U2193 : AOI22_X1 port map( A1 => n5199, A2 => n932, B1 => n5231, B2 => n40, 
                           ZN => n3987);
   U2194 : OAI221_X1 port map( B1 => n1229, B2 => n189, C1 => n1227, C2 => n338
                           , A => n3987, ZN => n3988);
   U2195 : NOR4_X1 port map( A1 => n3991, A2 => n3990, A3 => n3988, A4 => n3989
                           , ZN => n3993);
   U2196 : OAI222_X1 port map( A1 => n809, A2 => n1239, B1 => n3993, B2 => 
                           n1236, C1 => n1233, C2 => n3992, ZN => n3994);
   U2197 : OAI22_X1 port map( A1 => n509, A2 => n3996, B1 => n937, B2 => n480, 
                           ZN => n3997);
   U2198 : AOI221_X1 port map( B1 => n4815, B2 => n1254, C1 => n1252, C2 => 
                           n4312, A => n3997, ZN => n4005);
   U2199 : OAI22_X1 port map( A1 => n4719, A2 => n1275, B1 => n1436, B2 => 
                           n1273, ZN => n4001);
   U2200 : AOI221_X1 port map( B1 => n4975, B2 => n1283, C1 => n1280, C2 => 
                           n4002, A => n4001, ZN => n4003);
   U2201 : AOI22_X1 port map( A1 => n1199, A2 => n4007, B1 => n1196, B2 => 
                           n4131, ZN => n4008);
   U2202 : OAI221_X1 port map( B1 => n1207, B2 => n318, C1 => n232, C2 => n1204
                           , A => n4008, ZN => n4017);
   U2203 : AOI22_X1 port map( A1 => n998, A2 => n4195, B1 => n1208, B2 => n4163
                           , ZN => n4009);
   U2204 : OAI221_X1 port map( B1 => n360, B2 => n1215, C1 => n392, C2 => n8, A
                           => n4009, ZN => n4016);
   U2205 : AOI22_X1 port map( A1 => n5136, A2 => n589, B1 => n5168, B2 => n1218
                           , ZN => n4010);
   U2206 : OAI221_X1 port map( B1 => n1224, B2 => n4012, C1 => n1221, C2 => 
                           n4011, A => n4010, ZN => n4015);
   U2207 : AOI22_X1 port map( A1 => n5200, A2 => n710, B1 => n5232, B2 => n931,
                           ZN => n4013);
   U2208 : OAI221_X1 port map( B1 => n1228, B2 => n190, C1 => n1227, C2 => n339
                           , A => n4013, ZN => n4014);
   U2209 : NOR4_X1 port map( A1 => n4017, A2 => n4016, A3 => n4015, A4 => n4014
                           , ZN => n4019);
   U2210 : OAI222_X1 port map( A1 => n808, A2 => n1239, B1 => n4019, B2 => 
                           n1236, C1 => n1233, C2 => n4018, ZN => n4020);
   U2211 : OAI22_X1 port map( A1 => n1248, A2 => n4022, B1 => n936, B2 => n1247
                           , ZN => n4023);
   U2212 : AOI221_X1 port map( B1 => n4816, B2 => n1255, C1 => n1252, C2 => 
                           n4311, A => n4023, ZN => n4031);
   U2213 : OAI22_X1 port map( A1 => n4720, A2 => n1275, B1 => n1439, B2 => 
                           n1273, ZN => n4027);
   U2214 : AOI221_X1 port map( B1 => n4976, B2 => n1283, C1 => n1280, C2 => 
                           n4028, A => n4027, ZN => n4029);
   U2215 : AOI22_X1 port map( A1 => n1201, A2 => n4033, B1 => n1196, B2 => 
                           n4130, ZN => n4034);
   U2216 : AOI22_X1 port map( A1 => n689, A2 => n4194, B1 => n1208, B2 => n4162
                           , ZN => n4035);
   U2217 : OAI221_X1 port map( B1 => n359, B2 => n6, C1 => n391, C2 => n1210, A
                           => n4035, ZN => n4042);
   U2218 : AOI22_X1 port map( A1 => n5137, A2 => n987, B1 => n5169, B2 => n1218
                           , ZN => n4036);
   U2219 : OAI221_X1 port map( B1 => n1222, B2 => n4038, C1 => n1221, C2 => 
                           n4037, A => n4036, ZN => n4041);
   U2220 : AOI22_X1 port map( A1 => n5201, A2 => n710, B1 => n5233, B2 => n40, 
                           ZN => n4039);
   U2221 : OAI221_X1 port map( B1 => n1229, B2 => n191, C1 => n1227, C2 => n340
                           , A => n4039, ZN => n4040);
   U2222 : NOR4_X1 port map( A1 => n4043, A2 => n4042, A3 => n4041, A4 => n4040
                           , ZN => n4045);
   U2223 : OAI222_X1 port map( A1 => n807, A2 => n1239, B1 => n4045, B2 => 
                           n1236, C1 => n1233, C2 => n4044, ZN => n4046);
   U2224 : OAI22_X1 port map( A1 => n1249, A2 => n4048, B1 => n935, B2 => n1246
                           , ZN => n4049);
   U2225 : AOI221_X1 port map( B1 => n4817, B2 => n33, C1 => n1252, C2 => n4310
                           , A => n4049, ZN => n4057);
   U2226 : OAI222_X1 port map( A1 => n615, A2 => n1264, B1 => n1261, B2 => 
                           n4051, C1 => n1257, C2 => n4050, ZN => n4052);
   U2227 : AOI221_X1 port map( B1 => n1270, B2 => n4258, C1 => n1267, C2 => 
                           n4226, A => n4052, ZN => n4056);
   U2228 : OAI22_X1 port map( A1 => n4721, A2 => n1275, B1 => n1442, B2 => 
                           n1273, ZN => n4053);
   U2229 : AOI221_X1 port map( B1 => n4977, B2 => n1283, C1 => n1280, C2 => 
                           n4054, A => n4053, ZN => n4055);
   U2230 : AOI22_X1 port map( A1 => n1199, A2 => n4059, B1 => n1197, B2 => 
                           n4129, ZN => n4060);
   U2231 : OAI221_X1 port map( B1 => n1206, B2 => n320, C1 => n230, C2 => n1204
                           , A => n4060, ZN => n4069);
   U2232 : AOI22_X1 port map( A1 => n689, A2 => n4193, B1 => n1209, B2 => n4161
                           , ZN => n4061);
   U2233 : OAI221_X1 port map( B1 => n358, B2 => n6, C1 => n390, C2 => n1210, A
                           => n4061, ZN => n4068);
   U2234 : AOI22_X1 port map( A1 => n704, A2 => n5138, B1 => n5170, B2 => n1218
                           , ZN => n4062);
   U2235 : OAI221_X1 port map( B1 => n1222, B2 => n4064, C1 => n1221, C2 => 
                           n4063, A => n4062, ZN => n4067);
   U2236 : AOI22_X1 port map( A1 => n5202, A2 => n710, B1 => n5234, B2 => n40, 
                           ZN => n4065);
   U2237 : OAI221_X1 port map( B1 => n1229, B2 => n192, C1 => n1227, C2 => n341
                           , A => n4065, ZN => n4066);
   U2238 : NOR4_X1 port map( A1 => n4069, A2 => n4068, A3 => n4067, A4 => n4066
                           , ZN => n4071);
   U2239 : OAI222_X1 port map( A1 => n806, A2 => n1239, B1 => n4071, B2 => 
                           n1236, C1 => n1233, C2 => n4070, ZN => n4072);
   U2240 : OAI22_X1 port map( A1 => n1248, A2 => n4074, B1 => n934, B2 => n480,
                           ZN => n4075);
   U2241 : AOI221_X1 port map( B1 => n4818, B2 => n1254, C1 => n1252, C2 => 
                           n4309, A => n4075, ZN => n4083);
   U2242 : OAI222_X1 port map( A1 => n614, A2 => n1264, B1 => n1261, B2 => 
                           n4077, C1 => n1257, C2 => n4076, ZN => n4078);
   U2243 : AOI221_X1 port map( B1 => n1270, B2 => n4257, C1 => n1267, C2 => 
                           n4225, A => n4078, ZN => n4082);
   U2244 : OAI22_X1 port map( A1 => n4722, A2 => n1275, B1 => n1445, B2 => 
                           n1273, ZN => n4079);
   U2245 : AOI221_X1 port map( B1 => n4978, B2 => n1283, C1 => n1280, C2 => 
                           n4080, A => n4079, ZN => n4081);
   U2246 : AOI22_X1 port map( A1 => n1201, A2 => n4085, B1 => n1198, B2 => 
                           n4128, ZN => n4086);
   U2247 : OAI221_X1 port map( B1 => n1206, B2 => n321, C1 => n229, C2 => n1204
                           , A => n4086, ZN => n4103);
   U2248 : AOI22_X1 port map( A1 => n689, A2 => n4192, B1 => n1209, B2 => n4160
                           , ZN => n4089);
   U2249 : OAI221_X1 port map( B1 => n357, B2 => n1214, C1 => n389, C2 => n1211
                           , A => n4089, ZN => n4102);
   U2250 : AOI22_X1 port map( A1 => n589, A2 => n5139, B1 => n5171, B2 => n1218
                           , ZN => n4092);
   U2251 : OAI221_X1 port map( B1 => n1224, B2 => n4095, C1 => n1221, C2 => 
                           n4093, A => n4092, ZN => n4101);
   U2252 : AOI22_X1 port map( A1 => n5203, A2 => n2, B1 => n5235, B2 => n931, 
                           ZN => n4097);
   U2253 : OAI221_X1 port map( B1 => n1229, B2 => n193, C1 => n1227, C2 => n342
                           , A => n4097, ZN => n4100);
   U2254 : NOR4_X1 port map( A1 => n4103, A2 => n4100, A3 => n4102, A4 => n4101
                           , ZN => n4107);
   U2255 : OAI222_X1 port map( A1 => n805, A2 => n1239, B1 => n4107, B2 => 
                           n1236, C1 => n1233, C2 => n4104, ZN => n4109);
   U2256 : OAI22_X1 port map( A1 => n1248, A2 => n4112, B1 => n933, B2 => n480,
                           ZN => n4114);
   U2257 : AOI221_X1 port map( B1 => n4819, B2 => n1254, C1 => n1252, C2 => 
                           n4308, A => n4114, ZN => n4126);
   U2258 : OAI222_X1 port map( A1 => n613, A2 => n1264, B1 => n1260, B2 => 
                           n4117, C1 => n590, C2 => n4115, ZN => n4120);
   U2259 : AOI221_X1 port map( B1 => n1270, B2 => n4256, C1 => n1267, C2 => 
                           n4224, A => n4120, ZN => n4125);
   U2260 : OAI22_X1 port map( A1 => n4723, A2 => n1276, B1 => n1448, B2 => 
                           n1273, ZN => n4122);
   U2261 : AOI221_X1 port map( B1 => n4979, B2 => n1283, C1 => n1280, C2 => 
                           n4123, A => n4122, ZN => n4124);
   U2262 : NAND4_X1 port map( A1 => n4127, A2 => n4124, A3 => n4125, A4 => 
                           n4126, ZN => n2569);
   U2263 : MUX2_X1 port map( A => n4128, B => n1446, S => n1286, Z => n3561);
   U2264 : MUX2_X1 port map( A => n4129, B => n1443, S => n1286, Z => n3560);
   U2265 : MUX2_X1 port map( A => n4130, B => n1440, S => n1286, Z => n3559);
   U2266 : MUX2_X1 port map( A => n4131, B => n1437, S => n1286, Z => n3558);
   U2267 : MUX2_X1 port map( A => n4132, B => n1434, S => n1286, Z => n3557);
   U2268 : MUX2_X1 port map( A => n4133, B => n1431, S => n1286, Z => n3556);
   U2269 : MUX2_X1 port map( A => n4134, B => n1428, S => n1286, Z => n3555);
   U2270 : MUX2_X1 port map( A => n4135, B => n1425, S => n1286, Z => n3554);
   U2271 : MUX2_X1 port map( A => n4136, B => n1423, S => n1285, Z => n3553);
   U2272 : MUX2_X1 port map( A => n4137, B => n1421, S => n1285, Z => n3552);
   U2273 : MUX2_X1 port map( A => n4138, B => n1419, S => n1285, Z => n3551);
   U2274 : MUX2_X1 port map( A => n4139, B => n1417, S => n1285, Z => n3550);
   U2275 : MUX2_X1 port map( A => n4140, B => n1415, S => n1285, Z => n3549);
   U2276 : MUX2_X1 port map( A => n4141, B => n1413, S => n1285, Z => n3548);
   U2277 : MUX2_X1 port map( A => n4142, B => n1411, S => n1285, Z => n3547);
   U2278 : MUX2_X1 port map( A => n4143, B => n1409, S => n1285, Z => n3546);
   U2279 : MUX2_X1 port map( A => n4144, B => n1407, S => n1285, Z => n3545);
   U2280 : MUX2_X1 port map( A => n4145, B => n1405, S => n1285, Z => n3544);
   U2281 : MUX2_X1 port map( A => n4146, B => n1403, S => n1285, Z => n3543);
   U2282 : MUX2_X1 port map( A => n4147, B => n1401, S => n1285, Z => n3542);
   U2283 : MUX2_X1 port map( A => n4148, B => n1399, S => n1284, Z => n3541);
   U2284 : MUX2_X1 port map( A => n4149, B => n1397, S => n1284, Z => n3540);
   U2285 : MUX2_X1 port map( A => n4150, B => n1395, S => n1284, Z => n3539);
   U2286 : MUX2_X1 port map( A => n4151, B => n1393, S => n1284, Z => n3538);
   U2287 : MUX2_X1 port map( A => n4152, B => n1391, S => n1284, Z => n3537);
   U2288 : MUX2_X1 port map( A => n4153, B => n1389, S => n1284, Z => n3536);
   U2289 : MUX2_X1 port map( A => n4154, B => n1387, S => n1284, Z => n3535);
   U2290 : MUX2_X1 port map( A => n4155, B => n1385, S => n1284, Z => n3534);
   U2291 : MUX2_X1 port map( A => n4156, B => n1383, S => n1284, Z => n3533);
   U2292 : MUX2_X1 port map( A => n4157, B => n1381, S => n1284, Z => n3532);
   U2293 : MUX2_X1 port map( A => n4158, B => n1379, S => n1284, Z => n3531);
   U2294 : MUX2_X1 port map( A => n4159, B => n1377, S => n1284, Z => n3530);
   U2295 : AND2_X1 port map( A1 => n4341, A2 => n4342, ZN => n4340);
   U2296 : MUX2_X1 port map( A => n5235, B => n1446, S => n1289, Z => n3529);
   U2297 : MUX2_X1 port map( A => n5234, B => n1443, S => n1289, Z => n3528);
   U2298 : MUX2_X1 port map( A => n5233, B => n1440, S => n1289, Z => n3527);
   U2299 : MUX2_X1 port map( A => n5232, B => n1437, S => n1289, Z => n3526);
   U2300 : MUX2_X1 port map( A => n5231, B => n1434, S => n1289, Z => n3525);
   U2301 : MUX2_X1 port map( A => n5230, B => n1431, S => n1289, Z => n3524);
   U2302 : MUX2_X1 port map( A => n5229, B => n1428, S => n1289, Z => n3523);
   U2303 : MUX2_X1 port map( A => n5228, B => n1425, S => n1289, Z => n3522);
   U2304 : MUX2_X1 port map( A => n5227, B => n1423, S => n1288, Z => n3521);
   U2305 : MUX2_X1 port map( A => n5226, B => n1421, S => n1288, Z => n3520);
   U2306 : MUX2_X1 port map( A => n5225, B => n1419, S => n1288, Z => n3519);
   U2307 : MUX2_X1 port map( A => n5224, B => n1417, S => n1288, Z => n3518);
   U2308 : MUX2_X1 port map( A => n5223, B => n1415, S => n1288, Z => n3517);
   U2309 : MUX2_X1 port map( A => n5222, B => n1413, S => n1288, Z => n3516);
   U2310 : MUX2_X1 port map( A => n5221, B => n1411, S => n1288, Z => n3515);
   U2311 : MUX2_X1 port map( A => n5220, B => n1409, S => n1288, Z => n3514);
   U2312 : MUX2_X1 port map( A => n5219, B => n1407, S => n1288, Z => n3513);
   U2313 : MUX2_X1 port map( A => n5218, B => n1405, S => n1288, Z => n3512);
   U2314 : MUX2_X1 port map( A => n5217, B => n1403, S => n1288, Z => n3511);
   U2315 : MUX2_X1 port map( A => n5216, B => n1401, S => n1288, Z => n3510);
   U2316 : MUX2_X1 port map( A => n5215, B => n1399, S => n1287, Z => n3509);
   U2317 : MUX2_X1 port map( A => n5214, B => n1397, S => n1287, Z => n3508);
   U2318 : MUX2_X1 port map( A => n5213, B => n1395, S => n1287, Z => n3507);
   U2319 : MUX2_X1 port map( A => n5212, B => n1393, S => n1287, Z => n3506);
   U2320 : MUX2_X1 port map( A => n5211, B => n1391, S => n1287, Z => n3505);
   U2321 : MUX2_X1 port map( A => n5210, B => n1389, S => n1287, Z => n3504);
   U2322 : MUX2_X1 port map( A => n5209, B => n1387, S => n1287, Z => n3503);
   U2323 : MUX2_X1 port map( A => n5208, B => n1385, S => n1287, Z => n3502);
   U2324 : MUX2_X1 port map( A => n5207, B => n1383, S => n1287, Z => n3501);
   U2325 : MUX2_X1 port map( A => n5206, B => n1381, S => n1287, Z => n3500);
   U2326 : MUX2_X1 port map( A => n5205, B => n1379, S => n1287, Z => n3499);
   U2327 : MUX2_X1 port map( A => n5204, B => n1377, S => n1287, Z => n3498);
   U2328 : AND2_X1 port map( A1 => n4344, A2 => n4342, ZN => n4343);
   U2329 : MUX2_X1 port map( A => n5203, B => n1446, S => n1292, Z => n3497);
   U2330 : MUX2_X1 port map( A => n5202, B => n1443, S => n1292, Z => n3496);
   U2331 : MUX2_X1 port map( A => n5201, B => n1440, S => n1292, Z => n3495);
   U2332 : MUX2_X1 port map( A => n5200, B => n1437, S => n1292, Z => n3494);
   U2333 : MUX2_X1 port map( A => n5199, B => n1434, S => n1292, Z => n3493);
   U2334 : MUX2_X1 port map( A => n5198, B => n1431, S => n1292, Z => n3492);
   U2335 : MUX2_X1 port map( A => n5197, B => n1428, S => n1292, Z => n3491);
   U2336 : MUX2_X1 port map( A => n5196, B => n1425, S => n1292, Z => n3490);
   U2337 : MUX2_X1 port map( A => n5195, B => n1423, S => n1291, Z => n3489);
   U2338 : MUX2_X1 port map( A => n5194, B => n1421, S => n1291, Z => n3488);
   U2339 : MUX2_X1 port map( A => n5193, B => n1419, S => n1291, Z => n3487);
   U2340 : MUX2_X1 port map( A => n5192, B => n1417, S => n1291, Z => n3486);
   U2341 : MUX2_X1 port map( A => n5191, B => n1415, S => n1291, Z => n3485);
   U2342 : MUX2_X1 port map( A => n5190, B => n1413, S => n1291, Z => n3484);
   U2343 : MUX2_X1 port map( A => n5189, B => n1411, S => n1291, Z => n3483);
   U2344 : MUX2_X1 port map( A => n5188, B => n1409, S => n1291, Z => n3482);
   U2345 : MUX2_X1 port map( A => n5187, B => n1407, S => n1291, Z => n3481);
   U2346 : MUX2_X1 port map( A => n5186, B => n1405, S => n1291, Z => n3480);
   U2347 : MUX2_X1 port map( A => n5185, B => n1403, S => n1291, Z => n3479);
   U2348 : MUX2_X1 port map( A => n5184, B => n1401, S => n1291, Z => n3478);
   U2349 : MUX2_X1 port map( A => n5183, B => n1399, S => n1290, Z => n3477);
   U2350 : MUX2_X1 port map( A => n5182, B => n1397, S => n1290, Z => n3476);
   U2351 : MUX2_X1 port map( A => n5181, B => n1395, S => n1290, Z => n3475);
   U2352 : MUX2_X1 port map( A => n5180, B => n1393, S => n1290, Z => n3474);
   U2353 : MUX2_X1 port map( A => n5179, B => n1391, S => n1290, Z => n3473);
   U2354 : MUX2_X1 port map( A => n5178, B => n1389, S => n1290, Z => n3472);
   U2355 : MUX2_X1 port map( A => n5177, B => n1387, S => n1290, Z => n3471);
   U2356 : MUX2_X1 port map( A => n5176, B => n1385, S => n1290, Z => n3470);
   U2357 : MUX2_X1 port map( A => n5175, B => n1383, S => n1290, Z => n3469);
   U2358 : MUX2_X1 port map( A => n5174, B => n1381, S => n1290, Z => n3468);
   U2359 : MUX2_X1 port map( A => n5173, B => n1379, S => n1290, Z => n3467);
   U2360 : MUX2_X1 port map( A => n5172, B => n1377, S => n1290, Z => n3466);
   U2361 : AND2_X1 port map( A1 => n4346, A2 => n4342, ZN => n4345);
   U2362 : MUX2_X1 port map( A => n4160, B => n1446, S => n1295, Z => n3465);
   U2363 : MUX2_X1 port map( A => n4161, B => n1443, S => n1295, Z => n3464);
   U2364 : MUX2_X1 port map( A => n4162, B => n1440, S => n1295, Z => n3463);
   U2365 : MUX2_X1 port map( A => n4163, B => n1437, S => n1295, Z => n3462);
   U2366 : MUX2_X1 port map( A => n4164, B => n1434, S => n1295, Z => n3461);
   U2367 : MUX2_X1 port map( A => n4165, B => n1431, S => n1295, Z => n3460);
   U2368 : MUX2_X1 port map( A => n4166, B => n1428, S => n1295, Z => n3459);
   U2369 : MUX2_X1 port map( A => n4167, B => n1425, S => n1295, Z => n3458);
   U2370 : MUX2_X1 port map( A => n4168, B => n1423, S => n1294, Z => n3457);
   U2371 : MUX2_X1 port map( A => n4169, B => n1421, S => n1294, Z => n3456);
   U2372 : MUX2_X1 port map( A => n4170, B => n1419, S => n1294, Z => n3455);
   U2373 : MUX2_X1 port map( A => n4171, B => n1417, S => n1294, Z => n3454);
   U2374 : MUX2_X1 port map( A => n4172, B => n1415, S => n1294, Z => n3453);
   U2375 : MUX2_X1 port map( A => n4173, B => n1413, S => n1294, Z => n3452);
   U2376 : MUX2_X1 port map( A => n4174, B => n1411, S => n1294, Z => n3451);
   U2377 : MUX2_X1 port map( A => n4175, B => n1409, S => n1294, Z => n3450);
   U2378 : MUX2_X1 port map( A => n4176, B => n1407, S => n1294, Z => n3449);
   U2379 : MUX2_X1 port map( A => n4177, B => n1405, S => n1294, Z => n3448);
   U2380 : MUX2_X1 port map( A => n4178, B => n1403, S => n1294, Z => n3447);
   U2381 : MUX2_X1 port map( A => n4179, B => n1401, S => n1294, Z => n3446);
   U2382 : MUX2_X1 port map( A => n4180, B => n1399, S => n1293, Z => n3445);
   U2383 : MUX2_X1 port map( A => n4181, B => n1397, S => n1293, Z => n3444);
   U2384 : MUX2_X1 port map( A => n4182, B => n1395, S => n1293, Z => n3443);
   U2385 : MUX2_X1 port map( A => n4183, B => n1393, S => n1293, Z => n3442);
   U2386 : MUX2_X1 port map( A => n4184, B => n1391, S => n1293, Z => n3441);
   U2387 : MUX2_X1 port map( A => n4185, B => n1389, S => n1293, Z => n3440);
   U2388 : MUX2_X1 port map( A => n4186, B => n1387, S => n1293, Z => n3439);
   U2389 : MUX2_X1 port map( A => n4187, B => n1385, S => n1293, Z => n3438);
   U2390 : MUX2_X1 port map( A => n4188, B => n1383, S => n1293, Z => n3437);
   U2391 : MUX2_X1 port map( A => n4189, B => n1381, S => n1293, Z => n3436);
   U2392 : MUX2_X1 port map( A => n4190, B => n1379, S => n1293, Z => n3435);
   U2393 : MUX2_X1 port map( A => n4191, B => n1377, S => n1293, Z => n3434);
   U2394 : AND2_X1 port map( A1 => n4348, A2 => n4342, ZN => n4347);
   U2395 : MUX2_X1 port map( A => n4192, B => n1446, S => n1298, Z => n3433);
   U2396 : MUX2_X1 port map( A => n4193, B => n1443, S => n1298, Z => n3432);
   U2397 : MUX2_X1 port map( A => n4194, B => n1440, S => n1298, Z => n3431);
   U2398 : MUX2_X1 port map( A => n4195, B => n1437, S => n1298, Z => n3430);
   U2399 : MUX2_X1 port map( A => n4196, B => n1434, S => n1298, Z => n3429);
   U2400 : MUX2_X1 port map( A => n4197, B => n1431, S => n1298, Z => n3428);
   U2401 : MUX2_X1 port map( A => n4198, B => n1428, S => n1298, Z => n3427);
   U2402 : MUX2_X1 port map( A => n4199, B => n1425, S => n1298, Z => n3426);
   U2403 : MUX2_X1 port map( A => n4200, B => n1423, S => n1297, Z => n3425);
   U2404 : MUX2_X1 port map( A => n4201, B => n1421, S => n1297, Z => n3424);
   U2405 : MUX2_X1 port map( A => n4202, B => n1419, S => n1297, Z => n3423);
   U2406 : MUX2_X1 port map( A => n4203, B => n1417, S => n1297, Z => n3422);
   U2407 : MUX2_X1 port map( A => n4204, B => n1415, S => n1297, Z => n3421);
   U2408 : MUX2_X1 port map( A => n4205, B => n1413, S => n1297, Z => n3420);
   U2409 : MUX2_X1 port map( A => n4206, B => n1411, S => n1297, Z => n3419);
   U2410 : MUX2_X1 port map( A => n4207, B => n1409, S => n1297, Z => n3418);
   U2411 : MUX2_X1 port map( A => n4208, B => n1407, S => n1297, Z => n3417);
   U2412 : MUX2_X1 port map( A => n4209, B => n1405, S => n1297, Z => n3416);
   U2413 : MUX2_X1 port map( A => n4210, B => n1403, S => n1297, Z => n3415);
   U2414 : MUX2_X1 port map( A => n4211, B => n1401, S => n1297, Z => n3414);
   U2415 : MUX2_X1 port map( A => n4212, B => n1399, S => n1296, Z => n3413);
   U2416 : MUX2_X1 port map( A => n4213, B => n1397, S => n1296, Z => n3412);
   U2417 : MUX2_X1 port map( A => n4214, B => n1395, S => n1296, Z => n3411);
   U2418 : MUX2_X1 port map( A => n4215, B => n1393, S => n1296, Z => n3410);
   U2419 : MUX2_X1 port map( A => n4216, B => n1391, S => n1296, Z => n3409);
   U2420 : MUX2_X1 port map( A => n4217, B => n1389, S => n1296, Z => n3408);
   U2421 : MUX2_X1 port map( A => n4218, B => n1387, S => n1296, Z => n3407);
   U2422 : MUX2_X1 port map( A => n4219, B => n1385, S => n1296, Z => n3406);
   U2423 : MUX2_X1 port map( A => n4220, B => n1383, S => n1296, Z => n3405);
   U2424 : MUX2_X1 port map( A => n4221, B => n1381, S => n1296, Z => n3404);
   U2425 : MUX2_X1 port map( A => n4222, B => n1379, S => n1296, Z => n3403);
   U2426 : MUX2_X1 port map( A => n4223, B => n1377, S => n1296, Z => n3402);
   U2427 : AND2_X1 port map( A1 => n4350, A2 => n4342, ZN => n4349);
   U2428 : MUX2_X1 port map( A => n5171, B => n1446, S => n1301, Z => n3401);
   U2429 : MUX2_X1 port map( A => n5170, B => n1443, S => n1301, Z => n3400);
   U2430 : MUX2_X1 port map( A => n5169, B => n1440, S => n1301, Z => n3399);
   U2431 : MUX2_X1 port map( A => n5168, B => n1437, S => n1301, Z => n3398);
   U2432 : MUX2_X1 port map( A => n5167, B => n1434, S => n1301, Z => n3397);
   U2433 : MUX2_X1 port map( A => n5166, B => n1431, S => n1301, Z => n3396);
   U2434 : MUX2_X1 port map( A => n5165, B => n1428, S => n1301, Z => n3395);
   U2435 : MUX2_X1 port map( A => n5164, B => n1425, S => n1301, Z => n3394);
   U2436 : MUX2_X1 port map( A => n5163, B => n1423, S => n1300, Z => n3393);
   U2437 : MUX2_X1 port map( A => n5162, B => n1421, S => n1300, Z => n3392);
   U2438 : MUX2_X1 port map( A => n5161, B => n1419, S => n1300, Z => n3391);
   U2439 : MUX2_X1 port map( A => n5160, B => n1417, S => n1300, Z => n3390);
   U2440 : MUX2_X1 port map( A => n5159, B => n1415, S => n1300, Z => n3389);
   U2441 : MUX2_X1 port map( A => n5158, B => n1413, S => n1300, Z => n3388);
   U2442 : MUX2_X1 port map( A => n5157, B => n1411, S => n1300, Z => n3387);
   U2443 : MUX2_X1 port map( A => n5156, B => n1409, S => n1300, Z => n3386);
   U2444 : MUX2_X1 port map( A => n5155, B => n1407, S => n1300, Z => n3385);
   U2445 : MUX2_X1 port map( A => n5154, B => n1405, S => n1300, Z => n3384);
   U2446 : MUX2_X1 port map( A => n5153, B => n1403, S => n1300, Z => n3383);
   U2447 : MUX2_X1 port map( A => n5152, B => n1401, S => n1300, Z => n3382);
   U2448 : MUX2_X1 port map( A => n5151, B => n1399, S => n1299, Z => n3381);
   U2449 : MUX2_X1 port map( A => n5150, B => n1397, S => n1299, Z => n3380);
   U2450 : MUX2_X1 port map( A => n5149, B => n1395, S => n1299, Z => n3379);
   U2451 : MUX2_X1 port map( A => n5148, B => n1393, S => n1299, Z => n3378);
   U2452 : MUX2_X1 port map( A => n5147, B => n1391, S => n1299, Z => n3377);
   U2453 : MUX2_X1 port map( A => n5146, B => n1389, S => n1299, Z => n3376);
   U2454 : MUX2_X1 port map( A => n5145, B => n1387, S => n1299, Z => n3375);
   U2455 : MUX2_X1 port map( A => n5144, B => n1385, S => n1299, Z => n3374);
   U2456 : MUX2_X1 port map( A => n5143, B => n1383, S => n1299, Z => n3373);
   U2457 : MUX2_X1 port map( A => n5142, B => n1381, S => n1299, Z => n3372);
   U2458 : MUX2_X1 port map( A => n5141, B => n1379, S => n1299, Z => n3371);
   U2459 : MUX2_X1 port map( A => n5140, B => n1377, S => n1299, Z => n3370);
   U2460 : AND2_X1 port map( A1 => n4352, A2 => n4342, ZN => n4351);
   U2461 : MUX2_X1 port map( A => n5139, B => n1446, S => n1304, Z => n3369);
   U2462 : MUX2_X1 port map( A => n5138, B => n1443, S => n1304, Z => n3368);
   U2463 : MUX2_X1 port map( A => n5137, B => n1440, S => n1304, Z => n3367);
   U2464 : MUX2_X1 port map( A => n5136, B => n1437, S => n1304, Z => n3366);
   U2465 : MUX2_X1 port map( A => n5135, B => n1434, S => n1304, Z => n3365);
   U2466 : MUX2_X1 port map( A => n5134, B => n1431, S => n1304, Z => n3364);
   U2467 : MUX2_X1 port map( A => n5133, B => n1428, S => n1304, Z => n3363);
   U2468 : MUX2_X1 port map( A => n5132, B => n1425, S => n1304, Z => n3362);
   U2469 : MUX2_X1 port map( A => n5131, B => n1423, S => n1303, Z => n3361);
   U2470 : MUX2_X1 port map( A => n5130, B => n1421, S => n1303, Z => n3360);
   U2471 : MUX2_X1 port map( A => n5129, B => n1419, S => n1303, Z => n3359);
   U2472 : MUX2_X1 port map( A => n5128, B => n1417, S => n1303, Z => n3358);
   U2473 : MUX2_X1 port map( A => n5127, B => n1415, S => n1303, Z => n3357);
   U2474 : MUX2_X1 port map( A => n5126, B => n1413, S => n1303, Z => n3356);
   U2475 : MUX2_X1 port map( A => n5125, B => n1411, S => n1303, Z => n3355);
   U2476 : MUX2_X1 port map( A => n5124, B => n1409, S => n1303, Z => n3354);
   U2477 : MUX2_X1 port map( A => n5123, B => n1407, S => n1303, Z => n3353);
   U2478 : MUX2_X1 port map( A => n5122, B => n1405, S => n1303, Z => n3352);
   U2479 : MUX2_X1 port map( A => n5121, B => n1403, S => n1303, Z => n3351);
   U2480 : MUX2_X1 port map( A => n5120, B => n1401, S => n1303, Z => n3350);
   U2481 : MUX2_X1 port map( A => n5119, B => n1399, S => n1302, Z => n3349);
   U2482 : MUX2_X1 port map( A => n5118, B => n1397, S => n1302, Z => n3348);
   U2483 : MUX2_X1 port map( A => n5117, B => n1395, S => n1302, Z => n3347);
   U2484 : MUX2_X1 port map( A => n5116, B => n1393, S => n1302, Z => n3346);
   U2485 : MUX2_X1 port map( A => n5115, B => n1391, S => n1302, Z => n3345);
   U2486 : MUX2_X1 port map( A => n5114, B => n1389, S => n1302, Z => n3344);
   U2487 : MUX2_X1 port map( A => n5113, B => n1387, S => n1302, Z => n3343);
   U2488 : MUX2_X1 port map( A => n5112, B => n1385, S => n1302, Z => n3342);
   U2489 : MUX2_X1 port map( A => n5111, B => n1383, S => n1302, Z => n3341);
   U2490 : MUX2_X1 port map( A => n5110, B => n1381, S => n1302, Z => n3340);
   U2491 : MUX2_X1 port map( A => n5109, B => n1379, S => n1302, Z => n3339);
   U2492 : MUX2_X1 port map( A => n5108, B => n1377, S => n1302, Z => n3338);
   U2493 : AND2_X1 port map( A1 => n4354, A2 => n4342, ZN => n4353);
   U2494 : AND3_X1 port map( A1 => n4355, A2 => n4356, A3 => n4357, ZN => n4342
                           );
   U2495 : INV_X1 port map( A => n4358, ZN => n3337);
   U2496 : MUX2_X1 port map( A => n229, B => n1448, S => n1307, Z => n4358);
   U2497 : INV_X1 port map( A => n4360, ZN => n3336);
   U2498 : MUX2_X1 port map( A => n230, B => n1445, S => n1307, Z => n4360);
   U2499 : INV_X1 port map( A => n4361, ZN => n3335);
   U2500 : MUX2_X1 port map( A => n231, B => n1442, S => n1307, Z => n4361);
   U2501 : INV_X1 port map( A => n4362, ZN => n3334);
   U2502 : MUX2_X1 port map( A => n232, B => n1439, S => n1307, Z => n4362);
   U2503 : INV_X1 port map( A => n4363, ZN => n3333);
   U2504 : MUX2_X1 port map( A => n233, B => n1436, S => n1307, Z => n4363);
   U2505 : INV_X1 port map( A => n4364, ZN => n3332);
   U2506 : MUX2_X1 port map( A => n234, B => n1433, S => n1307, Z => n4364);
   U2507 : INV_X1 port map( A => n4365, ZN => n3331);
   U2508 : MUX2_X1 port map( A => n235, B => n1430, S => n1307, Z => n4365);
   U2509 : INV_X1 port map( A => n4366, ZN => n3330);
   U2510 : MUX2_X1 port map( A => n236, B => n1427, S => n1307, Z => n4366);
   U2511 : INV_X1 port map( A => n4367, ZN => n3329);
   U2512 : MUX2_X1 port map( A => n237, B => n1424, S => n1306, Z => n4367);
   U2513 : INV_X1 port map( A => n4368, ZN => n3328);
   U2514 : MUX2_X1 port map( A => n238, B => n1422, S => n1306, Z => n4368);
   U2515 : INV_X1 port map( A => n4369, ZN => n3327);
   U2516 : MUX2_X1 port map( A => n239, B => n1420, S => n1306, Z => n4369);
   U2517 : INV_X1 port map( A => n4370, ZN => n3326);
   U2518 : MUX2_X1 port map( A => n240, B => n1418, S => n1306, Z => n4370);
   U2519 : INV_X1 port map( A => n4371, ZN => n3325);
   U2520 : MUX2_X1 port map( A => n241, B => n1416, S => n1306, Z => n4371);
   U2521 : INV_X1 port map( A => n4372, ZN => n3324);
   U2522 : MUX2_X1 port map( A => n242, B => n1414, S => n1306, Z => n4372);
   U2523 : INV_X1 port map( A => n4373, ZN => n3323);
   U2524 : MUX2_X1 port map( A => n243, B => n1412, S => n1306, Z => n4373);
   U2525 : INV_X1 port map( A => n4374, ZN => n3322);
   U2526 : MUX2_X1 port map( A => n244, B => n1410, S => n1306, Z => n4374);
   U2527 : INV_X1 port map( A => n4375, ZN => n3321);
   U2528 : MUX2_X1 port map( A => n245, B => n1408, S => n1306, Z => n4375);
   U2529 : INV_X1 port map( A => n4376, ZN => n3320);
   U2530 : MUX2_X1 port map( A => n246, B => n1406, S => n1306, Z => n4376);
   U2531 : INV_X1 port map( A => n4377, ZN => n3319);
   U2532 : MUX2_X1 port map( A => n247, B => n1404, S => n1306, Z => n4377);
   U2533 : INV_X1 port map( A => n4378, ZN => n3318);
   U2534 : MUX2_X1 port map( A => n248, B => n1402, S => n1306, Z => n4378);
   U2535 : INV_X1 port map( A => n4379, ZN => n3317);
   U2536 : MUX2_X1 port map( A => n249, B => n1400, S => n1305, Z => n4379);
   U2537 : INV_X1 port map( A => n4380, ZN => n3316);
   U2538 : MUX2_X1 port map( A => n250, B => n1398, S => n1305, Z => n4380);
   U2539 : INV_X1 port map( A => n4381, ZN => n3315);
   U2540 : MUX2_X1 port map( A => n251, B => n1396, S => n1305, Z => n4381);
   U2541 : INV_X1 port map( A => n4382, ZN => n3314);
   U2542 : MUX2_X1 port map( A => n252, B => n1394, S => n1305, Z => n4382);
   U2543 : INV_X1 port map( A => n4383, ZN => n3313);
   U2544 : MUX2_X1 port map( A => n253, B => n1392, S => n1305, Z => n4383);
   U2545 : INV_X1 port map( A => n4384, ZN => n3312);
   U2546 : MUX2_X1 port map( A => n254, B => n1390, S => n1305, Z => n4384);
   U2547 : INV_X1 port map( A => n4385, ZN => n3311);
   U2548 : MUX2_X1 port map( A => n255, B => n1388, S => n1305, Z => n4385);
   U2549 : INV_X1 port map( A => n4386, ZN => n3310);
   U2550 : MUX2_X1 port map( A => n256, B => n1386, S => n1305, Z => n4386);
   U2551 : INV_X1 port map( A => n4387, ZN => n3309);
   U2552 : MUX2_X1 port map( A => n257, B => n1384, S => n1305, Z => n4387);
   U2553 : INV_X1 port map( A => n4388, ZN => n3308);
   U2554 : MUX2_X1 port map( A => n258, B => n1382, S => n1305, Z => n4388);
   U2555 : INV_X1 port map( A => n4389, ZN => n3307);
   U2556 : MUX2_X1 port map( A => n259, B => n1380, S => n1305, Z => n4389);
   U2557 : INV_X1 port map( A => n4390, ZN => n3306);
   U2558 : MUX2_X1 port map( A => n260, B => n1378, S => n1305, Z => n4390);
   U2559 : AND2_X1 port map( A1 => n4391, A2 => n4392, ZN => n4359);
   U2560 : INV_X1 port map( A => n4393, ZN => n3305);
   U2561 : MUX2_X1 port map( A => n261, B => n1448, S => n1310, Z => n4393);
   U2562 : INV_X1 port map( A => n4395, ZN => n3304);
   U2563 : MUX2_X1 port map( A => n262, B => n1445, S => n1310, Z => n4395);
   U2564 : INV_X1 port map( A => n4396, ZN => n3303);
   U2565 : MUX2_X1 port map( A => n263, B => n1442, S => n1310, Z => n4396);
   U2566 : INV_X1 port map( A => n4397, ZN => n3302);
   U2567 : MUX2_X1 port map( A => n264, B => n1439, S => n1310, Z => n4397);
   U2568 : INV_X1 port map( A => n4398, ZN => n3301);
   U2569 : MUX2_X1 port map( A => n265, B => n1436, S => n1310, Z => n4398);
   U2570 : INV_X1 port map( A => n4399, ZN => n3300);
   U2571 : MUX2_X1 port map( A => n266, B => n1433, S => n1310, Z => n4399);
   U2572 : INV_X1 port map( A => n4400, ZN => n3299);
   U2573 : MUX2_X1 port map( A => n267, B => n1430, S => n1310, Z => n4400);
   U2574 : INV_X1 port map( A => n4401, ZN => n3298);
   U2575 : MUX2_X1 port map( A => n268, B => n1427, S => n1310, Z => n4401);
   U2576 : INV_X1 port map( A => n4402, ZN => n3297);
   U2577 : MUX2_X1 port map( A => n269, B => n1424, S => n1309, Z => n4402);
   U2578 : INV_X1 port map( A => n4403, ZN => n3296);
   U2579 : MUX2_X1 port map( A => n270, B => n1422, S => n1309, Z => n4403);
   U2580 : INV_X1 port map( A => n4404, ZN => n3295);
   U2581 : MUX2_X1 port map( A => n271, B => n1420, S => n1309, Z => n4404);
   U2582 : INV_X1 port map( A => n4405, ZN => n3294);
   U2583 : MUX2_X1 port map( A => n272, B => n1418, S => n1309, Z => n4405);
   U2584 : INV_X1 port map( A => n4406, ZN => n3293);
   U2585 : MUX2_X1 port map( A => n273, B => n1416, S => n1309, Z => n4406);
   U2586 : INV_X1 port map( A => n4407, ZN => n3292);
   U2587 : MUX2_X1 port map( A => n274, B => n1414, S => n1309, Z => n4407);
   U2588 : INV_X1 port map( A => n4408, ZN => n3291);
   U2589 : MUX2_X1 port map( A => n275, B => n1412, S => n1309, Z => n4408);
   U2590 : INV_X1 port map( A => n4409, ZN => n3290);
   U2591 : MUX2_X1 port map( A => n276, B => n1410, S => n1309, Z => n4409);
   U2592 : INV_X1 port map( A => n4410, ZN => n3289);
   U2593 : MUX2_X1 port map( A => n277, B => n1408, S => n1309, Z => n4410);
   U2594 : INV_X1 port map( A => n4411, ZN => n3288);
   U2595 : MUX2_X1 port map( A => n278, B => n1406, S => n1309, Z => n4411);
   U2596 : INV_X1 port map( A => n4412, ZN => n3287);
   U2597 : MUX2_X1 port map( A => n279, B => n1404, S => n1309, Z => n4412);
   U2598 : INV_X1 port map( A => n4413, ZN => n3286);
   U2599 : MUX2_X1 port map( A => n280, B => n1402, S => n1309, Z => n4413);
   U2600 : INV_X1 port map( A => n4414, ZN => n3285);
   U2601 : MUX2_X1 port map( A => n281, B => n1400, S => n1308, Z => n4414);
   U2602 : INV_X1 port map( A => n4415, ZN => n3284);
   U2603 : MUX2_X1 port map( A => n282, B => n1398, S => n1308, Z => n4415);
   U2604 : INV_X1 port map( A => n4416, ZN => n3283);
   U2605 : MUX2_X1 port map( A => n283, B => n1396, S => n1308, Z => n4416);
   U2606 : INV_X1 port map( A => n4417, ZN => n3282);
   U2607 : MUX2_X1 port map( A => n284, B => n1394, S => n1308, Z => n4417);
   U2608 : INV_X1 port map( A => n4418, ZN => n3281);
   U2609 : MUX2_X1 port map( A => n285, B => n1392, S => n1308, Z => n4418);
   U2610 : INV_X1 port map( A => n4419, ZN => n3280);
   U2611 : MUX2_X1 port map( A => n286, B => n1390, S => n1308, Z => n4419);
   U2612 : INV_X1 port map( A => n4420, ZN => n3279);
   U2613 : MUX2_X1 port map( A => n287, B => n1388, S => n1308, Z => n4420);
   U2614 : INV_X1 port map( A => n4421, ZN => n3278);
   U2615 : MUX2_X1 port map( A => n288, B => n1386, S => n1308, Z => n4421);
   U2616 : INV_X1 port map( A => n4422, ZN => n3277);
   U2617 : MUX2_X1 port map( A => n289, B => n1384, S => n1308, Z => n4422);
   U2618 : INV_X1 port map( A => n4423, ZN => n3276);
   U2619 : MUX2_X1 port map( A => n290, B => n1382, S => n1308, Z => n4423);
   U2620 : INV_X1 port map( A => n4424, ZN => n3275);
   U2621 : MUX2_X1 port map( A => n291, B => n1380, S => n1308, Z => n4424);
   U2622 : INV_X1 port map( A => n4425, ZN => n3274);
   U2623 : MUX2_X1 port map( A => n292, B => n1378, S => n1308, Z => n4425);
   U2624 : AND2_X1 port map( A1 => n4391, A2 => n4341, ZN => n4394);
   U2625 : MUX2_X1 port map( A => n5107, B => n1446, S => n1313, Z => n3273);
   U2626 : MUX2_X1 port map( A => n5106, B => n1443, S => n1313, Z => n3272);
   U2627 : MUX2_X1 port map( A => n5105, B => n1440, S => n1313, Z => n3271);
   U2628 : MUX2_X1 port map( A => n5104, B => n1437, S => n1313, Z => n3270);
   U2629 : MUX2_X1 port map( A => n5103, B => n1434, S => n1313, Z => n3269);
   U2630 : MUX2_X1 port map( A => n5102, B => n1431, S => n1313, Z => n3268);
   U2631 : MUX2_X1 port map( A => n5101, B => n1428, S => n1313, Z => n3267);
   U2632 : MUX2_X1 port map( A => n5100, B => n1425, S => n1313, Z => n3266);
   U2633 : MUX2_X1 port map( A => n5099, B => n1423, S => n1312, Z => n3265);
   U2634 : MUX2_X1 port map( A => n5098, B => n1421, S => n1312, Z => n3264);
   U2635 : MUX2_X1 port map( A => n5097, B => n1419, S => n1312, Z => n3263);
   U2636 : MUX2_X1 port map( A => n5096, B => n1417, S => n1312, Z => n3262);
   U2637 : MUX2_X1 port map( A => n5095, B => n1415, S => n1312, Z => n3261);
   U2638 : MUX2_X1 port map( A => n5094, B => n1413, S => n1312, Z => n3260);
   U2639 : MUX2_X1 port map( A => n5093, B => n1411, S => n1312, Z => n3259);
   U2640 : MUX2_X1 port map( A => n5092, B => n1409, S => n1312, Z => n3258);
   U2641 : MUX2_X1 port map( A => n5091, B => n1407, S => n1312, Z => n3257);
   U2642 : MUX2_X1 port map( A => n5090, B => n1405, S => n1312, Z => n3256);
   U2643 : MUX2_X1 port map( A => n5089, B => n1403, S => n1312, Z => n3255);
   U2644 : MUX2_X1 port map( A => n5088, B => n1401, S => n1312, Z => n3254);
   U2645 : MUX2_X1 port map( A => n5087, B => n1399, S => n1311, Z => n3253);
   U2646 : MUX2_X1 port map( A => n5086, B => n1397, S => n1311, Z => n3252);
   U2647 : MUX2_X1 port map( A => n5085, B => n1395, S => n1311, Z => n3251);
   U2648 : MUX2_X1 port map( A => n5084, B => n1393, S => n1311, Z => n3250);
   U2649 : MUX2_X1 port map( A => n5083, B => n1391, S => n1311, Z => n3249);
   U2650 : MUX2_X1 port map( A => n5082, B => n1389, S => n1311, Z => n3248);
   U2651 : MUX2_X1 port map( A => n5081, B => n1387, S => n1311, Z => n3247);
   U2652 : MUX2_X1 port map( A => n5080, B => n1385, S => n1311, Z => n3246);
   U2653 : MUX2_X1 port map( A => n5079, B => n1383, S => n1311, Z => n3245);
   U2654 : MUX2_X1 port map( A => n5078, B => n1381, S => n1311, Z => n3244);
   U2655 : MUX2_X1 port map( A => n5077, B => n1379, S => n1311, Z => n3243);
   U2656 : MUX2_X1 port map( A => n5076, B => n1377, S => n1311, Z => n3242);
   U2657 : AND2_X1 port map( A1 => n4391, A2 => n4344, ZN => n4426);
   U2658 : MUX2_X1 port map( A => n5075, B => n1446, S => n1316, Z => n3241);
   U2659 : MUX2_X1 port map( A => n5074, B => n1443, S => n1316, Z => n3240);
   U2660 : MUX2_X1 port map( A => n5073, B => n1440, S => n1316, Z => n3239);
   U2661 : MUX2_X1 port map( A => n5072, B => n1437, S => n1316, Z => n3238);
   U2662 : MUX2_X1 port map( A => n5071, B => n1434, S => n1316, Z => n3237);
   U2663 : MUX2_X1 port map( A => n5070, B => n1431, S => n1316, Z => n3236);
   U2664 : MUX2_X1 port map( A => n5069, B => n1428, S => n1316, Z => n3235);
   U2665 : MUX2_X1 port map( A => n5068, B => n1425, S => n1316, Z => n3234);
   U2666 : MUX2_X1 port map( A => n5067, B => n1423, S => n1315, Z => n3233);
   U2667 : MUX2_X1 port map( A => n5066, B => n1421, S => n1315, Z => n3232);
   U2668 : MUX2_X1 port map( A => n5065, B => n1419, S => n1315, Z => n3231);
   U2669 : MUX2_X1 port map( A => n5064, B => n1417, S => n1315, Z => n3230);
   U2670 : MUX2_X1 port map( A => n5063, B => n1415, S => n1315, Z => n3229);
   U2671 : MUX2_X1 port map( A => n5062, B => n1413, S => n1315, Z => n3228);
   U2672 : MUX2_X1 port map( A => n5061, B => n1411, S => n1315, Z => n3227);
   U2673 : MUX2_X1 port map( A => n5060, B => n1409, S => n1315, Z => n3226);
   U2674 : MUX2_X1 port map( A => n5059, B => n1407, S => n1315, Z => n3225);
   U2675 : MUX2_X1 port map( A => n5058, B => n1405, S => n1315, Z => n3224);
   U2676 : MUX2_X1 port map( A => n5057, B => n1403, S => n1315, Z => n3223);
   U2677 : MUX2_X1 port map( A => n5056, B => n1401, S => n1315, Z => n3222);
   U2678 : MUX2_X1 port map( A => n5055, B => n1399, S => n1314, Z => n3221);
   U2679 : MUX2_X1 port map( A => n5054, B => n1397, S => n1314, Z => n3220);
   U2680 : MUX2_X1 port map( A => n5053, B => n1395, S => n1314, Z => n3219);
   U2681 : MUX2_X1 port map( A => n5052, B => n1393, S => n1314, Z => n3218);
   U2682 : MUX2_X1 port map( A => n5051, B => n1391, S => n1314, Z => n3217);
   U2683 : MUX2_X1 port map( A => n5050, B => n1389, S => n1314, Z => n3216);
   U2684 : MUX2_X1 port map( A => n5049, B => n1387, S => n1314, Z => n3215);
   U2685 : MUX2_X1 port map( A => n5048, B => n1385, S => n1314, Z => n3214);
   U2686 : MUX2_X1 port map( A => n5047, B => n1383, S => n1314, Z => n3213);
   U2687 : MUX2_X1 port map( A => n5046, B => n1381, S => n1314, Z => n3212);
   U2688 : MUX2_X1 port map( A => n5045, B => n1379, S => n1314, Z => n3211);
   U2689 : MUX2_X1 port map( A => n5044, B => n1377, S => n1314, Z => n3210);
   U2690 : AND2_X1 port map( A1 => n4391, A2 => n4346, ZN => n4427);
   U2691 : INV_X1 port map( A => n4428, ZN => n3209);
   U2692 : MUX2_X1 port map( A => n357, B => n1448, S => n1319, Z => n4428);
   U2693 : INV_X1 port map( A => n4430, ZN => n3208);
   U2694 : MUX2_X1 port map( A => n358, B => n1445, S => n1319, Z => n4430);
   U2695 : INV_X1 port map( A => n4431, ZN => n3207);
   U2696 : MUX2_X1 port map( A => n359, B => n1442, S => n1319, Z => n4431);
   U2697 : INV_X1 port map( A => n4432, ZN => n3206);
   U2698 : MUX2_X1 port map( A => n360, B => n1439, S => n1319, Z => n4432);
   U2699 : INV_X1 port map( A => n4433, ZN => n3205);
   U2700 : MUX2_X1 port map( A => n361, B => n1436, S => n1319, Z => n4433);
   U2701 : INV_X1 port map( A => n4434, ZN => n3204);
   U2702 : MUX2_X1 port map( A => n362, B => n1433, S => n1319, Z => n4434);
   U2703 : INV_X1 port map( A => n4435, ZN => n3203);
   U2704 : MUX2_X1 port map( A => n363, B => n1430, S => n1319, Z => n4435);
   U2705 : INV_X1 port map( A => n4436, ZN => n3202);
   U2706 : MUX2_X1 port map( A => n364, B => n1427, S => n1319, Z => n4436);
   U2707 : INV_X1 port map( A => n4437, ZN => n3201);
   U2708 : MUX2_X1 port map( A => n365, B => n1424, S => n1318, Z => n4437);
   U2709 : INV_X1 port map( A => n4438, ZN => n3200);
   U2710 : MUX2_X1 port map( A => n366, B => n1422, S => n1318, Z => n4438);
   U2711 : INV_X1 port map( A => n4439, ZN => n3199);
   U2712 : MUX2_X1 port map( A => n367, B => n1420, S => n1318, Z => n4439);
   U2713 : INV_X1 port map( A => n4440, ZN => n3198);
   U2714 : MUX2_X1 port map( A => n368, B => n1418, S => n1318, Z => n4440);
   U2715 : INV_X1 port map( A => n4441, ZN => n3197);
   U2716 : MUX2_X1 port map( A => n369, B => n1416, S => n1318, Z => n4441);
   U2717 : INV_X1 port map( A => n4442, ZN => n3196);
   U2718 : MUX2_X1 port map( A => n370, B => n1414, S => n1318, Z => n4442);
   U2719 : INV_X1 port map( A => n4443, ZN => n3195);
   U2720 : MUX2_X1 port map( A => n371, B => n1412, S => n1318, Z => n4443);
   U2721 : INV_X1 port map( A => n4444, ZN => n3194);
   U2722 : MUX2_X1 port map( A => n372, B => n1410, S => n1318, Z => n4444);
   U2723 : INV_X1 port map( A => n4445, ZN => n3193);
   U2724 : MUX2_X1 port map( A => n373, B => n1408, S => n1318, Z => n4445);
   U2725 : INV_X1 port map( A => n4446, ZN => n3192);
   U2726 : MUX2_X1 port map( A => n374, B => n1406, S => n1318, Z => n4446);
   U2727 : INV_X1 port map( A => n4447, ZN => n3191);
   U2728 : MUX2_X1 port map( A => n375, B => n1404, S => n1318, Z => n4447);
   U2729 : INV_X1 port map( A => n4448, ZN => n3190);
   U2730 : MUX2_X1 port map( A => n376, B => n1402, S => n1318, Z => n4448);
   U2731 : INV_X1 port map( A => n4449, ZN => n3189);
   U2732 : MUX2_X1 port map( A => n377, B => n1400, S => n1317, Z => n4449);
   U2733 : INV_X1 port map( A => n4450, ZN => n3188);
   U2734 : MUX2_X1 port map( A => n378, B => n1398, S => n1317, Z => n4450);
   U2735 : INV_X1 port map( A => n4451, ZN => n3187);
   U2736 : MUX2_X1 port map( A => n379, B => n1396, S => n1317, Z => n4451);
   U2737 : INV_X1 port map( A => n4452, ZN => n3186);
   U2738 : MUX2_X1 port map( A => n380, B => n1394, S => n1317, Z => n4452);
   U2739 : INV_X1 port map( A => n4453, ZN => n3185);
   U2740 : MUX2_X1 port map( A => n381, B => n1392, S => n1317, Z => n4453);
   U2741 : INV_X1 port map( A => n4454, ZN => n3184);
   U2742 : MUX2_X1 port map( A => n382, B => n1390, S => n1317, Z => n4454);
   U2743 : INV_X1 port map( A => n4455, ZN => n3183);
   U2744 : MUX2_X1 port map( A => n383, B => n1388, S => n1317, Z => n4455);
   U2745 : INV_X1 port map( A => n4456, ZN => n3182);
   U2746 : MUX2_X1 port map( A => n384, B => n1386, S => n1317, Z => n4456);
   U2747 : INV_X1 port map( A => n4457, ZN => n3181);
   U2748 : MUX2_X1 port map( A => n385, B => n1384, S => n1317, Z => n4457);
   U2749 : INV_X1 port map( A => n4458, ZN => n3180);
   U2750 : MUX2_X1 port map( A => n386, B => n1382, S => n1317, Z => n4458);
   U2751 : INV_X1 port map( A => n4459, ZN => n3179);
   U2752 : MUX2_X1 port map( A => n387, B => n1380, S => n1317, Z => n4459);
   U2753 : INV_X1 port map( A => n4460, ZN => n3178);
   U2754 : MUX2_X1 port map( A => n388, B => n1378, S => n1317, Z => n4460);
   U2755 : AND2_X1 port map( A1 => n4391, A2 => n4348, ZN => n4429);
   U2756 : INV_X1 port map( A => n4461, ZN => n3177);
   U2757 : MUX2_X1 port map( A => n389, B => n1448, S => n1322, Z => n4461);
   U2758 : INV_X1 port map( A => n4463, ZN => n3176);
   U2759 : MUX2_X1 port map( A => n390, B => n1445, S => n1322, Z => n4463);
   U2760 : INV_X1 port map( A => n4464, ZN => n3175);
   U2761 : MUX2_X1 port map( A => n391, B => n1442, S => n1322, Z => n4464);
   U2762 : INV_X1 port map( A => n4465, ZN => n3174);
   U2763 : MUX2_X1 port map( A => n392, B => n1439, S => n1322, Z => n4465);
   U2764 : INV_X1 port map( A => n4466, ZN => n3173);
   U2765 : MUX2_X1 port map( A => n393, B => n1436, S => n1322, Z => n4466);
   U2766 : INV_X1 port map( A => n4467, ZN => n3172);
   U2767 : MUX2_X1 port map( A => n394, B => n1433, S => n1322, Z => n4467);
   U2768 : INV_X1 port map( A => n4468, ZN => n3171);
   U2769 : MUX2_X1 port map( A => n395, B => n1430, S => n1322, Z => n4468);
   U2770 : INV_X1 port map( A => n4469, ZN => n3170);
   U2771 : MUX2_X1 port map( A => n396, B => n1427, S => n1322, Z => n4469);
   U2772 : INV_X1 port map( A => n4470, ZN => n3169);
   U2773 : MUX2_X1 port map( A => n397, B => n1424, S => n1321, Z => n4470);
   U2774 : INV_X1 port map( A => n4471, ZN => n3168);
   U2775 : MUX2_X1 port map( A => n398, B => n1422, S => n1321, Z => n4471);
   U2776 : INV_X1 port map( A => n4472, ZN => n3167);
   U2777 : MUX2_X1 port map( A => n399, B => n1420, S => n1321, Z => n4472);
   U2778 : INV_X1 port map( A => n4473, ZN => n3166);
   U2779 : MUX2_X1 port map( A => n400, B => n1418, S => n1321, Z => n4473);
   U2780 : INV_X1 port map( A => n4474, ZN => n3165);
   U2781 : MUX2_X1 port map( A => n401, B => n1416, S => n1321, Z => n4474);
   U2782 : INV_X1 port map( A => n4475, ZN => n3164);
   U2783 : MUX2_X1 port map( A => n402, B => n1414, S => n1321, Z => n4475);
   U2784 : INV_X1 port map( A => n4476, ZN => n3163);
   U2785 : MUX2_X1 port map( A => n403, B => n1412, S => n1321, Z => n4476);
   U2786 : INV_X1 port map( A => n4477, ZN => n3162);
   U2787 : MUX2_X1 port map( A => n404, B => n1410, S => n1321, Z => n4477);
   U2788 : INV_X1 port map( A => n4478, ZN => n3161);
   U2789 : MUX2_X1 port map( A => n405, B => n1408, S => n1321, Z => n4478);
   U2790 : INV_X1 port map( A => n4479, ZN => n3160);
   U2791 : MUX2_X1 port map( A => n406, B => n1406, S => n1321, Z => n4479);
   U2792 : INV_X1 port map( A => n4480, ZN => n3159);
   U2793 : MUX2_X1 port map( A => n407, B => n1404, S => n1321, Z => n4480);
   U2794 : INV_X1 port map( A => n4481, ZN => n3158);
   U2795 : MUX2_X1 port map( A => n408, B => n1402, S => n1321, Z => n4481);
   U2796 : INV_X1 port map( A => n4482, ZN => n3157);
   U2797 : MUX2_X1 port map( A => n409, B => n1400, S => n1320, Z => n4482);
   U2798 : INV_X1 port map( A => n4483, ZN => n3156);
   U2799 : MUX2_X1 port map( A => n410, B => n1398, S => n1320, Z => n4483);
   U2800 : INV_X1 port map( A => n4484, ZN => n3155);
   U2801 : MUX2_X1 port map( A => n411, B => n1396, S => n1320, Z => n4484);
   U2802 : INV_X1 port map( A => n4485, ZN => n3154);
   U2803 : MUX2_X1 port map( A => n412, B => n1394, S => n1320, Z => n4485);
   U2804 : INV_X1 port map( A => n4486, ZN => n3153);
   U2805 : MUX2_X1 port map( A => n413, B => n1392, S => n1320, Z => n4486);
   U2806 : INV_X1 port map( A => n4487, ZN => n3152);
   U2807 : MUX2_X1 port map( A => n414, B => n1390, S => n1320, Z => n4487);
   U2808 : INV_X1 port map( A => n4488, ZN => n3151);
   U2809 : MUX2_X1 port map( A => n415, B => n1388, S => n1320, Z => n4488);
   U2810 : INV_X1 port map( A => n4489, ZN => n3150);
   U2811 : MUX2_X1 port map( A => n416, B => n1386, S => n1320, Z => n4489);
   U2812 : INV_X1 port map( A => n4490, ZN => n3149);
   U2813 : MUX2_X1 port map( A => n417, B => n1384, S => n1320, Z => n4490);
   U2814 : INV_X1 port map( A => n4491, ZN => n3148);
   U2815 : MUX2_X1 port map( A => n418, B => n1382, S => n1320, Z => n4491);
   U2816 : INV_X1 port map( A => n4492, ZN => n3147);
   U2817 : MUX2_X1 port map( A => n419, B => n1380, S => n1320, Z => n4492);
   U2818 : INV_X1 port map( A => n4493, ZN => n3146);
   U2819 : MUX2_X1 port map( A => n420, B => n1378, S => n1320, Z => n4493);
   U2820 : AND2_X1 port map( A1 => n4391, A2 => n4350, ZN => n4462);
   U2821 : MUX2_X1 port map( A => n5043, B => n1446, S => n1325, Z => n3145);
   U2822 : MUX2_X1 port map( A => n5042, B => n1443, S => n1325, Z => n3144);
   U2823 : MUX2_X1 port map( A => n5041, B => n1440, S => n1325, Z => n3143);
   U2824 : MUX2_X1 port map( A => n5040, B => n1437, S => n1325, Z => n3142);
   U2825 : MUX2_X1 port map( A => n5039, B => n1434, S => n1325, Z => n3141);
   U2826 : MUX2_X1 port map( A => n5038, B => n1431, S => n1325, Z => n3140);
   U2827 : MUX2_X1 port map( A => n5037, B => n1428, S => n1325, Z => n3139);
   U2828 : MUX2_X1 port map( A => n5036, B => n1425, S => n1325, Z => n3138);
   U2829 : MUX2_X1 port map( A => n5035, B => n1423, S => n1324, Z => n3137);
   U2830 : MUX2_X1 port map( A => n5034, B => n1421, S => n1324, Z => n3136);
   U2831 : MUX2_X1 port map( A => n5033, B => n1419, S => n1324, Z => n3135);
   U2832 : MUX2_X1 port map( A => n5032, B => n1417, S => n1324, Z => n3134);
   U2833 : MUX2_X1 port map( A => n5031, B => n1415, S => n1324, Z => n3133);
   U2834 : MUX2_X1 port map( A => n5030, B => n1413, S => n1324, Z => n3132);
   U2835 : MUX2_X1 port map( A => n5029, B => n1411, S => n1324, Z => n3131);
   U2836 : MUX2_X1 port map( A => n5028, B => n1409, S => n1324, Z => n3130);
   U2837 : MUX2_X1 port map( A => n5027, B => n1407, S => n1324, Z => n3129);
   U2838 : MUX2_X1 port map( A => n5026, B => n1405, S => n1324, Z => n3128);
   U2839 : MUX2_X1 port map( A => n5025, B => n1403, S => n1324, Z => n3127);
   U2840 : MUX2_X1 port map( A => n5024, B => n1401, S => n1324, Z => n3126);
   U2841 : MUX2_X1 port map( A => n5023, B => n1399, S => n1323, Z => n3125);
   U2842 : MUX2_X1 port map( A => n5022, B => n1397, S => n1323, Z => n3124);
   U2843 : MUX2_X1 port map( A => n5021, B => n1395, S => n1323, Z => n3123);
   U2844 : MUX2_X1 port map( A => n5020, B => n1393, S => n1323, Z => n3122);
   U2845 : MUX2_X1 port map( A => n5019, B => n1391, S => n1323, Z => n3121);
   U2846 : MUX2_X1 port map( A => n5018, B => n1389, S => n1323, Z => n3120);
   U2847 : MUX2_X1 port map( A => n5017, B => n1387, S => n1323, Z => n3119);
   U2848 : MUX2_X1 port map( A => n5016, B => n1385, S => n1323, Z => n3118);
   U2849 : MUX2_X1 port map( A => n5015, B => n1383, S => n1323, Z => n3117);
   U2850 : MUX2_X1 port map( A => n5014, B => n1381, S => n1323, Z => n3116);
   U2851 : MUX2_X1 port map( A => n5013, B => n1379, S => n1323, Z => n3115);
   U2852 : MUX2_X1 port map( A => n5012, B => n1377, S => n1323, Z => n3114);
   U2853 : AND2_X1 port map( A1 => n4391, A2 => n4352, ZN => n4494);
   U2854 : MUX2_X1 port map( A => n5011, B => n1446, S => n1328, Z => n3113);
   U2855 : MUX2_X1 port map( A => n5010, B => n1443, S => n1328, Z => n3112);
   U2856 : MUX2_X1 port map( A => n5009, B => n1440, S => n1328, Z => n3111);
   U2857 : MUX2_X1 port map( A => n5008, B => n1437, S => n1328, Z => n3110);
   U2858 : MUX2_X1 port map( A => n5007, B => n1434, S => n1328, Z => n3109);
   U2859 : MUX2_X1 port map( A => n5006, B => n1431, S => n1328, Z => n3108);
   U2860 : MUX2_X1 port map( A => n5005, B => n1428, S => n1328, Z => n3107);
   U2861 : MUX2_X1 port map( A => n5004, B => n1425, S => n1328, Z => n3106);
   U2862 : MUX2_X1 port map( A => n5003, B => n1423, S => n1327, Z => n3105);
   U2863 : MUX2_X1 port map( A => n5002, B => n1421, S => n1327, Z => n3104);
   U2864 : MUX2_X1 port map( A => n5001, B => n1419, S => n1327, Z => n3103);
   U2865 : MUX2_X1 port map( A => n5000, B => n1417, S => n1327, Z => n3102);
   U2866 : MUX2_X1 port map( A => n4999, B => n1415, S => n1327, Z => n3101);
   U2867 : MUX2_X1 port map( A => n4998, B => n1413, S => n1327, Z => n3100);
   U2868 : MUX2_X1 port map( A => n4997, B => n1411, S => n1327, Z => n3099);
   U2869 : MUX2_X1 port map( A => n4996, B => n1409, S => n1327, Z => n3098);
   U2870 : MUX2_X1 port map( A => n4995, B => n1407, S => n1327, Z => n3097);
   U2871 : MUX2_X1 port map( A => n4994, B => n1405, S => n1327, Z => n3096);
   U2872 : MUX2_X1 port map( A => n4993, B => n1403, S => n1327, Z => n3095);
   U2873 : MUX2_X1 port map( A => n4992, B => n1401, S => n1327, Z => n3094);
   U2874 : MUX2_X1 port map( A => n4991, B => n1399, S => n1326, Z => n3093);
   U2875 : MUX2_X1 port map( A => n4990, B => n1397, S => n1326, Z => n3092);
   U2876 : MUX2_X1 port map( A => n4989, B => n1395, S => n1326, Z => n3091);
   U2877 : MUX2_X1 port map( A => n4988, B => n1393, S => n1326, Z => n3090);
   U2878 : MUX2_X1 port map( A => n4987, B => n1391, S => n1326, Z => n3089);
   U2879 : MUX2_X1 port map( A => n4986, B => n1389, S => n1326, Z => n3088);
   U2880 : MUX2_X1 port map( A => n4985, B => n1387, S => n1326, Z => n3087);
   U2881 : MUX2_X1 port map( A => n4984, B => n1385, S => n1326, Z => n3086);
   U2882 : MUX2_X1 port map( A => n4983, B => n1383, S => n1326, Z => n3085);
   U2883 : MUX2_X1 port map( A => n4982, B => n1381, S => n1326, Z => n3084);
   U2884 : MUX2_X1 port map( A => n4981, B => n1379, S => n1326, Z => n3083);
   U2885 : MUX2_X1 port map( A => n4980, B => n1377, S => n1326, Z => n3082);
   U2886 : AND2_X1 port map( A1 => n4391, A2 => n4354, ZN => n4495);
   U2887 : AND3_X1 port map( A1 => n4357, A2 => n4356, A3 => ADD_WR(3), ZN => 
                           n4391);
   U2888 : MUX2_X1 port map( A => n4224, B => n1447, S => n1331, Z => n3081);
   U2889 : MUX2_X1 port map( A => n4225, B => n1444, S => n1331, Z => n3080);
   U2890 : MUX2_X1 port map( A => n4226, B => n1441, S => n1331, Z => n3079);
   U2891 : MUX2_X1 port map( A => n4227, B => n1438, S => n1331, Z => n3078);
   U2892 : MUX2_X1 port map( A => n4228, B => n1435, S => n1331, Z => n3077);
   U2893 : MUX2_X1 port map( A => n4229, B => n1432, S => n1331, Z => n3076);
   U2894 : MUX2_X1 port map( A => n4230, B => n1429, S => n1331, Z => n3075);
   U2895 : MUX2_X1 port map( A => n4231, B => n1426, S => n1331, Z => n3074);
   U2896 : MUX2_X1 port map( A => n4232, B => n1423, S => n1330, Z => n3073);
   U2897 : MUX2_X1 port map( A => n4233, B => n1421, S => n1330, Z => n3072);
   U2898 : MUX2_X1 port map( A => n4234, B => n1419, S => n1330, Z => n3071);
   U2899 : MUX2_X1 port map( A => n4235, B => n1417, S => n1330, Z => n3070);
   U2900 : MUX2_X1 port map( A => n4236, B => n1415, S => n1330, Z => n3069);
   U2901 : MUX2_X1 port map( A => n4237, B => n1413, S => n1330, Z => n3068);
   U2902 : MUX2_X1 port map( A => n4238, B => n1411, S => n1330, Z => n3067);
   U2903 : MUX2_X1 port map( A => n4239, B => n1409, S => n1330, Z => n3066);
   U2904 : MUX2_X1 port map( A => n4240, B => n1407, S => n1330, Z => n3065);
   U2905 : MUX2_X1 port map( A => n4241, B => n1405, S => n1330, Z => n3064);
   U2906 : MUX2_X1 port map( A => n4242, B => n1403, S => n1330, Z => n3063);
   U2907 : MUX2_X1 port map( A => n4243, B => n1401, S => n1330, Z => n3062);
   U2908 : MUX2_X1 port map( A => n4244, B => n1399, S => n1329, Z => n3061);
   U2909 : MUX2_X1 port map( A => n4245, B => n1397, S => n1329, Z => n3060);
   U2910 : MUX2_X1 port map( A => n4246, B => n1395, S => n1329, Z => n3059);
   U2911 : MUX2_X1 port map( A => n4247, B => n1393, S => n1329, Z => n3058);
   U2912 : MUX2_X1 port map( A => n4248, B => n1391, S => n1329, Z => n3057);
   U2913 : MUX2_X1 port map( A => n4249, B => n1389, S => n1329, Z => n3056);
   U2914 : MUX2_X1 port map( A => n4250, B => n1387, S => n1329, Z => n3055);
   U2915 : MUX2_X1 port map( A => n4251, B => n1385, S => n1329, Z => n3054);
   U2916 : MUX2_X1 port map( A => n4252, B => n1383, S => n1329, Z => n3053);
   U2917 : MUX2_X1 port map( A => n4253, B => n1381, S => n1329, Z => n3052);
   U2918 : MUX2_X1 port map( A => n4254, B => n1379, S => n1329, Z => n3051);
   U2919 : MUX2_X1 port map( A => n4255, B => n1377, S => n1329, Z => n3050);
   U2920 : AND2_X1 port map( A1 => n4497, A2 => n4392, ZN => n4496);
   U2921 : INV_X1 port map( A => n4498, ZN => n3049);
   U2922 : MUX2_X1 port map( A => n517, B => n1448, S => n1334, Z => n4498);
   U2923 : INV_X1 port map( A => n4500, ZN => n3048);
   U2924 : MUX2_X1 port map( A => n518, B => n1445, S => n1334, Z => n4500);
   U2925 : INV_X1 port map( A => n4501, ZN => n3047);
   U2926 : MUX2_X1 port map( A => n519, B => n1442, S => n1334, Z => n4501);
   U2927 : INV_X1 port map( A => n4502, ZN => n3046);
   U2928 : MUX2_X1 port map( A => n520, B => n1439, S => n1334, Z => n4502);
   U2929 : INV_X1 port map( A => n4503, ZN => n3045);
   U2930 : MUX2_X1 port map( A => n521, B => n1436, S => n1334, Z => n4503);
   U2931 : INV_X1 port map( A => n4504, ZN => n3044);
   U2932 : MUX2_X1 port map( A => n522, B => n1433, S => n1334, Z => n4504);
   U2933 : INV_X1 port map( A => n4505, ZN => n3043);
   U2934 : MUX2_X1 port map( A => n523, B => n1430, S => n1334, Z => n4505);
   U2935 : INV_X1 port map( A => n4506, ZN => n3042);
   U2936 : MUX2_X1 port map( A => n524, B => n1427, S => n1334, Z => n4506);
   U2937 : INV_X1 port map( A => n4507, ZN => n3041);
   U2938 : MUX2_X1 port map( A => n525, B => n1424, S => n1333, Z => n4507);
   U2939 : INV_X1 port map( A => n4508, ZN => n3040);
   U2940 : MUX2_X1 port map( A => n526, B => n1422, S => n1333, Z => n4508);
   U2941 : INV_X1 port map( A => n4509, ZN => n3039);
   U2942 : MUX2_X1 port map( A => n527, B => n1420, S => n1333, Z => n4509);
   U2943 : INV_X1 port map( A => n4510, ZN => n3038);
   U2944 : MUX2_X1 port map( A => n528, B => n1418, S => n1333, Z => n4510);
   U2945 : INV_X1 port map( A => n4511, ZN => n3037);
   U2946 : MUX2_X1 port map( A => n529, B => n1416, S => n1333, Z => n4511);
   U2947 : INV_X1 port map( A => n4512, ZN => n3036);
   U2948 : MUX2_X1 port map( A => n530, B => n1414, S => n1333, Z => n4512);
   U2949 : INV_X1 port map( A => n4513, ZN => n3035);
   U2950 : MUX2_X1 port map( A => n531, B => n1412, S => n1333, Z => n4513);
   U2951 : INV_X1 port map( A => n4514, ZN => n3034);
   U2952 : MUX2_X1 port map( A => n532, B => n1410, S => n1333, Z => n4514);
   U2953 : INV_X1 port map( A => n4515, ZN => n3033);
   U2954 : MUX2_X1 port map( A => n533, B => n1408, S => n1333, Z => n4515);
   U2955 : INV_X1 port map( A => n4516, ZN => n3032);
   U2956 : MUX2_X1 port map( A => n534, B => n1406, S => n1333, Z => n4516);
   U2957 : INV_X1 port map( A => n4517, ZN => n3031);
   U2958 : MUX2_X1 port map( A => n535, B => n1404, S => n1333, Z => n4517);
   U2959 : INV_X1 port map( A => n4518, ZN => n3030);
   U2960 : MUX2_X1 port map( A => n536, B => n1402, S => n1333, Z => n4518);
   U2961 : INV_X1 port map( A => n4519, ZN => n3029);
   U2962 : MUX2_X1 port map( A => n537, B => n1400, S => n1332, Z => n4519);
   U2963 : INV_X1 port map( A => n4520, ZN => n3028);
   U2964 : MUX2_X1 port map( A => n538, B => n1398, S => n1332, Z => n4520);
   U2965 : INV_X1 port map( A => n4521, ZN => n3027);
   U2966 : MUX2_X1 port map( A => n539, B => n1396, S => n1332, Z => n4521);
   U2967 : INV_X1 port map( A => n4522, ZN => n3026);
   U2968 : MUX2_X1 port map( A => n540, B => n1394, S => n1332, Z => n4522);
   U2969 : INV_X1 port map( A => n4523, ZN => n3025);
   U2970 : MUX2_X1 port map( A => n541, B => n1392, S => n1332, Z => n4523);
   U2971 : INV_X1 port map( A => n4524, ZN => n3024);
   U2972 : MUX2_X1 port map( A => n542, B => n1390, S => n1332, Z => n4524);
   U2973 : INV_X1 port map( A => n4525, ZN => n3023);
   U2974 : MUX2_X1 port map( A => n543, B => n1388, S => n1332, Z => n4525);
   U2975 : INV_X1 port map( A => n4526, ZN => n3022);
   U2976 : MUX2_X1 port map( A => n544, B => n1386, S => n1332, Z => n4526);
   U2977 : INV_X1 port map( A => n4527, ZN => n3021);
   U2978 : MUX2_X1 port map( A => n545, B => n1384, S => n1332, Z => n4527);
   U2979 : INV_X1 port map( A => n4528, ZN => n3020);
   U2980 : MUX2_X1 port map( A => n546, B => n1382, S => n1332, Z => n4528);
   U2981 : INV_X1 port map( A => n4529, ZN => n3019);
   U2982 : MUX2_X1 port map( A => n547, B => n1380, S => n1332, Z => n4529);
   U2983 : INV_X1 port map( A => n4530, ZN => n3018);
   U2984 : MUX2_X1 port map( A => n548, B => n1378, S => n1332, Z => n4530);
   U2985 : AND2_X1 port map( A1 => n4497, A2 => n4341, ZN => n4499);
   U2986 : MUX2_X1 port map( A => n4979, B => n1447, S => n1337, Z => n3017);
   U2987 : MUX2_X1 port map( A => n4978, B => n1444, S => n1337, Z => n3016);
   U2988 : MUX2_X1 port map( A => n4977, B => n1441, S => n1337, Z => n3015);
   U2989 : MUX2_X1 port map( A => n4976, B => n1438, S => n1337, Z => n3014);
   U2990 : MUX2_X1 port map( A => n4975, B => n1435, S => n1337, Z => n3013);
   U2991 : MUX2_X1 port map( A => n4974, B => n1432, S => n1337, Z => n3012);
   U2992 : MUX2_X1 port map( A => n4973, B => n1429, S => n1337, Z => n3011);
   U2993 : MUX2_X1 port map( A => n4972, B => n1426, S => n1337, Z => n3010);
   U2994 : MUX2_X1 port map( A => n4971, B => n1423, S => n1336, Z => n3009);
   U2995 : MUX2_X1 port map( A => n4970, B => n1421, S => n1336, Z => n3008);
   U2996 : MUX2_X1 port map( A => n4969, B => n1419, S => n1336, Z => n3007);
   U2997 : MUX2_X1 port map( A => n4968, B => n1417, S => n1336, Z => n3006);
   U2998 : MUX2_X1 port map( A => n4967, B => n1415, S => n1336, Z => n3005);
   U2999 : MUX2_X1 port map( A => n4966, B => n1413, S => n1336, Z => n3004);
   U3000 : MUX2_X1 port map( A => n4965, B => n1411, S => n1336, Z => n3003);
   U3001 : MUX2_X1 port map( A => n4964, B => n1409, S => n1336, Z => n3002);
   U3002 : MUX2_X1 port map( A => n4963, B => n1407, S => n1336, Z => n3001);
   U3003 : MUX2_X1 port map( A => n4962, B => n1405, S => n1336, Z => n3000);
   U3004 : MUX2_X1 port map( A => n4961, B => n1403, S => n1336, Z => n2999);
   U3005 : MUX2_X1 port map( A => n4960, B => n1401, S => n1336, Z => n2998);
   U3006 : MUX2_X1 port map( A => n4959, B => n1399, S => n1335, Z => n2997);
   U3007 : MUX2_X1 port map( A => n4958, B => n1397, S => n1335, Z => n2996);
   U3008 : MUX2_X1 port map( A => n4957, B => n1395, S => n1335, Z => n2995);
   U3009 : MUX2_X1 port map( A => n4956, B => n1393, S => n1335, Z => n2994);
   U3010 : MUX2_X1 port map( A => n4955, B => n1391, S => n1335, Z => n2993);
   U3011 : MUX2_X1 port map( A => n4954, B => n1389, S => n1335, Z => n2992);
   U3012 : MUX2_X1 port map( A => n4953, B => n1387, S => n1335, Z => n2991);
   U3013 : MUX2_X1 port map( A => n4952, B => n1385, S => n1335, Z => n2990);
   U3014 : MUX2_X1 port map( A => n4951, B => n1383, S => n1335, Z => n2989);
   U3015 : MUX2_X1 port map( A => n4950, B => n1381, S => n1335, Z => n2988);
   U3016 : MUX2_X1 port map( A => n4949, B => n1379, S => n1335, Z => n2987);
   U3017 : MUX2_X1 port map( A => n4948, B => n1377, S => n1335, Z => n2986);
   U3018 : AND2_X1 port map( A1 => n4497, A2 => n4344, ZN => n4531);
   U3019 : MUX2_X1 port map( A => n4947, B => n1447, S => n1340, Z => n2985);
   U3020 : MUX2_X1 port map( A => n4946, B => n1444, S => n1340, Z => n2984);
   U3021 : MUX2_X1 port map( A => n4945, B => n1441, S => n1340, Z => n2983);
   U3022 : MUX2_X1 port map( A => n4944, B => n1438, S => n1340, Z => n2982);
   U3023 : MUX2_X1 port map( A => n4943, B => n1435, S => n1340, Z => n2981);
   U3024 : MUX2_X1 port map( A => n4942, B => n1432, S => n1340, Z => n2980);
   U3025 : MUX2_X1 port map( A => n4941, B => n1429, S => n1340, Z => n2979);
   U3026 : MUX2_X1 port map( A => n4940, B => n1426, S => n1340, Z => n2978);
   U3027 : MUX2_X1 port map( A => n4939, B => n1423, S => n1339, Z => n2977);
   U3028 : MUX2_X1 port map( A => n4938, B => n1421, S => n1339, Z => n2976);
   U3029 : MUX2_X1 port map( A => n4937, B => n1419, S => n1339, Z => n2975);
   U3030 : MUX2_X1 port map( A => n4936, B => n1417, S => n1339, Z => n2974);
   U3031 : MUX2_X1 port map( A => n4935, B => n1415, S => n1339, Z => n2973);
   U3032 : MUX2_X1 port map( A => n4934, B => n1413, S => n1339, Z => n2972);
   U3033 : MUX2_X1 port map( A => n4933, B => n1411, S => n1339, Z => n2971);
   U3034 : MUX2_X1 port map( A => n4932, B => n1409, S => n1339, Z => n2970);
   U3035 : MUX2_X1 port map( A => n4931, B => n1407, S => n1339, Z => n2969);
   U3036 : MUX2_X1 port map( A => n4930, B => n1405, S => n1339, Z => n2968);
   U3037 : MUX2_X1 port map( A => n4929, B => n1403, S => n1339, Z => n2967);
   U3038 : MUX2_X1 port map( A => n4928, B => n1401, S => n1339, Z => n2966);
   U3039 : MUX2_X1 port map( A => n4927, B => n1399, S => n1338, Z => n2965);
   U3040 : MUX2_X1 port map( A => n4926, B => n1397, S => n1338, Z => n2964);
   U3041 : MUX2_X1 port map( A => n4925, B => n1395, S => n1338, Z => n2963);
   U3042 : MUX2_X1 port map( A => n4924, B => n1393, S => n1338, Z => n2962);
   U3043 : MUX2_X1 port map( A => n4923, B => n1391, S => n1338, Z => n2961);
   U3044 : MUX2_X1 port map( A => n4922, B => n1389, S => n1338, Z => n2960);
   U3045 : MUX2_X1 port map( A => n4921, B => n1387, S => n1338, Z => n2959);
   U3046 : MUX2_X1 port map( A => n4920, B => n1385, S => n1338, Z => n2958);
   U3047 : MUX2_X1 port map( A => n4919, B => n1383, S => n1338, Z => n2957);
   U3048 : MUX2_X1 port map( A => n4918, B => n1381, S => n1338, Z => n2956);
   U3049 : MUX2_X1 port map( A => n4917, B => n1379, S => n1338, Z => n2955);
   U3050 : MUX2_X1 port map( A => n4916, B => n1377, S => n1338, Z => n2954);
   U3051 : AND2_X1 port map( A1 => n4497, A2 => n4346, ZN => n4532);
   U3052 : INV_X1 port map( A => n4533, ZN => n2953);
   U3053 : MUX2_X1 port map( A => n613, B => n1448, S => n1343, Z => n4533);
   U3054 : INV_X1 port map( A => n4535, ZN => n2952);
   U3055 : MUX2_X1 port map( A => n614, B => n1445, S => n1343, Z => n4535);
   U3056 : INV_X1 port map( A => n4536, ZN => n2951);
   U3057 : MUX2_X1 port map( A => n615, B => n1442, S => n1343, Z => n4536);
   U3058 : INV_X1 port map( A => n4537, ZN => n2950);
   U3059 : MUX2_X1 port map( A => n616, B => n1439, S => n1343, Z => n4537);
   U3060 : INV_X1 port map( A => n4538, ZN => n2949);
   U3061 : MUX2_X1 port map( A => n617, B => n1436, S => n1343, Z => n4538);
   U3062 : INV_X1 port map( A => n4539, ZN => n2948);
   U3063 : MUX2_X1 port map( A => n618, B => n1433, S => n1343, Z => n4539);
   U3064 : INV_X1 port map( A => n4540, ZN => n2947);
   U3065 : MUX2_X1 port map( A => n619, B => n1430, S => n1343, Z => n4540);
   U3066 : INV_X1 port map( A => n4541, ZN => n2946);
   U3067 : MUX2_X1 port map( A => n620, B => n1427, S => n1343, Z => n4541);
   U3068 : INV_X1 port map( A => n4542, ZN => n2945);
   U3069 : MUX2_X1 port map( A => n621, B => n1424, S => n1342, Z => n4542);
   U3070 : INV_X1 port map( A => n4543, ZN => n2944);
   U3071 : MUX2_X1 port map( A => n622, B => n1422, S => n1342, Z => n4543);
   U3072 : INV_X1 port map( A => n4544, ZN => n2943);
   U3073 : MUX2_X1 port map( A => n623, B => n1420, S => n1342, Z => n4544);
   U3074 : INV_X1 port map( A => n4545, ZN => n2942);
   U3075 : MUX2_X1 port map( A => n624, B => n1418, S => n1342, Z => n4545);
   U3076 : INV_X1 port map( A => n4546, ZN => n2941);
   U3077 : MUX2_X1 port map( A => n625, B => n1416, S => n1342, Z => n4546);
   U3078 : INV_X1 port map( A => n4547, ZN => n2940);
   U3079 : MUX2_X1 port map( A => n626, B => n1414, S => n1342, Z => n4547);
   U3080 : INV_X1 port map( A => n4548, ZN => n2939);
   U3081 : MUX2_X1 port map( A => n627, B => n1412, S => n1342, Z => n4548);
   U3082 : INV_X1 port map( A => n4549, ZN => n2938);
   U3083 : MUX2_X1 port map( A => n628, B => n1410, S => n1342, Z => n4549);
   U3084 : INV_X1 port map( A => n4550, ZN => n2937);
   U3085 : MUX2_X1 port map( A => n629, B => n1408, S => n1342, Z => n4550);
   U3086 : INV_X1 port map( A => n4551, ZN => n2936);
   U3087 : MUX2_X1 port map( A => n630, B => n1406, S => n1342, Z => n4551);
   U3088 : INV_X1 port map( A => n4552, ZN => n2935);
   U3089 : MUX2_X1 port map( A => n631, B => n1404, S => n1342, Z => n4552);
   U3090 : INV_X1 port map( A => n4553, ZN => n2934);
   U3091 : MUX2_X1 port map( A => n632, B => n1402, S => n1342, Z => n4553);
   U3092 : INV_X1 port map( A => n4554, ZN => n2933);
   U3093 : MUX2_X1 port map( A => n633, B => n1400, S => n1341, Z => n4554);
   U3094 : INV_X1 port map( A => n4555, ZN => n2932);
   U3095 : MUX2_X1 port map( A => n634, B => n1398, S => n1341, Z => n4555);
   U3096 : INV_X1 port map( A => n4556, ZN => n2931);
   U3097 : MUX2_X1 port map( A => n635, B => n1396, S => n1341, Z => n4556);
   U3098 : INV_X1 port map( A => n4557, ZN => n2930);
   U3099 : MUX2_X1 port map( A => n636, B => n1394, S => n1341, Z => n4557);
   U3100 : INV_X1 port map( A => n4558, ZN => n2929);
   U3101 : MUX2_X1 port map( A => n637, B => n1392, S => n1341, Z => n4558);
   U3102 : INV_X1 port map( A => n4559, ZN => n2928);
   U3103 : MUX2_X1 port map( A => n638, B => n1390, S => n1341, Z => n4559);
   U3104 : INV_X1 port map( A => n4560, ZN => n2927);
   U3105 : MUX2_X1 port map( A => n639, B => n1388, S => n1341, Z => n4560);
   U3106 : INV_X1 port map( A => n4561, ZN => n2926);
   U3107 : MUX2_X1 port map( A => n640, B => n1386, S => n1341, Z => n4561);
   U3108 : INV_X1 port map( A => n4562, ZN => n2925);
   U3109 : MUX2_X1 port map( A => n641, B => n1384, S => n1341, Z => n4562);
   U3110 : INV_X1 port map( A => n4563, ZN => n2924);
   U3111 : MUX2_X1 port map( A => n642, B => n1382, S => n1341, Z => n4563);
   U3112 : INV_X1 port map( A => n4564, ZN => n2923);
   U3113 : MUX2_X1 port map( A => n643, B => n1380, S => n1341, Z => n4564);
   U3114 : INV_X1 port map( A => n4565, ZN => n2922);
   U3115 : MUX2_X1 port map( A => n644, B => n1378, S => n1341, Z => n4565);
   U3116 : AND2_X1 port map( A1 => n4497, A2 => n4348, ZN => n4534);
   U3117 : MUX2_X1 port map( A => n4256, B => n1447, S => n1346, Z => n2921);
   U3118 : MUX2_X1 port map( A => n4257, B => n1444, S => n1346, Z => n2920);
   U3119 : MUX2_X1 port map( A => n4258, B => n1441, S => n1346, Z => n2919);
   U3120 : MUX2_X1 port map( A => n4259, B => n1438, S => n1346, Z => n2918);
   U3121 : MUX2_X1 port map( A => n4260, B => n1435, S => n1346, Z => n2917);
   U3122 : MUX2_X1 port map( A => n4261, B => n1432, S => n1346, Z => n2916);
   U3123 : MUX2_X1 port map( A => n4262, B => n1429, S => n1346, Z => n2915);
   U3124 : MUX2_X1 port map( A => n4263, B => n1426, S => n1346, Z => n2914);
   U3125 : MUX2_X1 port map( A => n4264, B => n1423, S => n1345, Z => n2913);
   U3126 : MUX2_X1 port map( A => n4265, B => n1421, S => n1345, Z => n2912);
   U3127 : MUX2_X1 port map( A => n4266, B => n1419, S => n1345, Z => n2911);
   U3128 : MUX2_X1 port map( A => n4267, B => n1417, S => n1345, Z => n2910);
   U3129 : MUX2_X1 port map( A => n4268, B => n1415, S => n1345, Z => n2909);
   U3130 : MUX2_X1 port map( A => n4269, B => n1413, S => n1345, Z => n2908);
   U3131 : MUX2_X1 port map( A => n4270, B => n1411, S => n1345, Z => n2907);
   U3132 : MUX2_X1 port map( A => n4271, B => n1409, S => n1345, Z => n2906);
   U3133 : MUX2_X1 port map( A => n4272, B => n1407, S => n1345, Z => n2905);
   U3134 : MUX2_X1 port map( A => n4273, B => n1405, S => n1345, Z => n2904);
   U3135 : MUX2_X1 port map( A => n4274, B => n1403, S => n1345, Z => n2903);
   U3136 : MUX2_X1 port map( A => n4275, B => n1401, S => n1345, Z => n2902);
   U3137 : MUX2_X1 port map( A => n4276, B => n1399, S => n1344, Z => n2901);
   U3138 : MUX2_X1 port map( A => n4277, B => n1397, S => n1344, Z => n2900);
   U3139 : MUX2_X1 port map( A => n4278, B => n1395, S => n1344, Z => n2899);
   U3140 : MUX2_X1 port map( A => n4279, B => n1393, S => n1344, Z => n2898);
   U3141 : MUX2_X1 port map( A => n4280, B => n1391, S => n1344, Z => n2897);
   U3142 : MUX2_X1 port map( A => n4281, B => n1389, S => n1344, Z => n2896);
   U3143 : MUX2_X1 port map( A => n4282, B => n1387, S => n1344, Z => n2895);
   U3144 : MUX2_X1 port map( A => n4283, B => n1385, S => n1344, Z => n2894);
   U3145 : MUX2_X1 port map( A => n4284, B => n1383, S => n1344, Z => n2893);
   U3146 : MUX2_X1 port map( A => n4285, B => n1381, S => n1344, Z => n2892);
   U3147 : MUX2_X1 port map( A => n4286, B => n1379, S => n1344, Z => n2891);
   U3148 : MUX2_X1 port map( A => n4287, B => n1377, S => n1344, Z => n2890);
   U3149 : AND2_X1 port map( A1 => n4497, A2 => n4350, ZN => n4566);
   U3150 : MUX2_X1 port map( A => n4915, B => n1447, S => n1349, Z => n2889);
   U3151 : MUX2_X1 port map( A => n4914, B => n1444, S => n1349, Z => n2888);
   U3152 : MUX2_X1 port map( A => n4913, B => n1441, S => n1349, Z => n2887);
   U3153 : MUX2_X1 port map( A => n4912, B => n1438, S => n1349, Z => n2886);
   U3154 : MUX2_X1 port map( A => n4911, B => n1435, S => n1349, Z => n2885);
   U3155 : MUX2_X1 port map( A => n4910, B => n1432, S => n1349, Z => n2884);
   U3156 : MUX2_X1 port map( A => n4909, B => n1429, S => n1349, Z => n2883);
   U3157 : MUX2_X1 port map( A => n4908, B => n1426, S => n1349, Z => n2882);
   U3158 : MUX2_X1 port map( A => n4907, B => n1423, S => n1348, Z => n2881);
   U3159 : MUX2_X1 port map( A => n4906, B => n1421, S => n1348, Z => n2880);
   U3160 : MUX2_X1 port map( A => n4905, B => n1419, S => n1348, Z => n2879);
   U3161 : MUX2_X1 port map( A => n4904, B => n1417, S => n1348, Z => n2878);
   U3162 : MUX2_X1 port map( A => n4903, B => n1415, S => n1348, Z => n2877);
   U3163 : MUX2_X1 port map( A => n4902, B => n1413, S => n1348, Z => n2876);
   U3164 : MUX2_X1 port map( A => n4901, B => n1411, S => n1348, Z => n2875);
   U3165 : MUX2_X1 port map( A => n4900, B => n1409, S => n1348, Z => n2874);
   U3166 : MUX2_X1 port map( A => n4899, B => n1407, S => n1348, Z => n2873);
   U3167 : MUX2_X1 port map( A => n4898, B => n1405, S => n1348, Z => n2872);
   U3168 : MUX2_X1 port map( A => n4897, B => n1403, S => n1348, Z => n2871);
   U3169 : MUX2_X1 port map( A => n4896, B => n1401, S => n1348, Z => n2870);
   U3170 : MUX2_X1 port map( A => n4895, B => n1399, S => n1347, Z => n2869);
   U3171 : MUX2_X1 port map( A => n4894, B => n1397, S => n1347, Z => n2868);
   U3172 : MUX2_X1 port map( A => n4893, B => n1395, S => n1347, Z => n2867);
   U3173 : MUX2_X1 port map( A => n4892, B => n1393, S => n1347, Z => n2866);
   U3174 : MUX2_X1 port map( A => n4891, B => n1391, S => n1347, Z => n2865);
   U3175 : MUX2_X1 port map( A => n4890, B => n1389, S => n1347, Z => n2864);
   U3176 : MUX2_X1 port map( A => n4889, B => n1387, S => n1347, Z => n2863);
   U3177 : MUX2_X1 port map( A => n4888, B => n1385, S => n1347, Z => n2862);
   U3178 : MUX2_X1 port map( A => n4887, B => n1383, S => n1347, Z => n2861);
   U3179 : MUX2_X1 port map( A => n4886, B => n1381, S => n1347, Z => n2860);
   U3180 : MUX2_X1 port map( A => n4885, B => n1379, S => n1347, Z => n2859);
   U3181 : MUX2_X1 port map( A => n4884, B => n1377, S => n1347, Z => n2858);
   U3182 : AND2_X1 port map( A1 => n4497, A2 => n4352, ZN => n4567);
   U3183 : MUX2_X1 port map( A => n4883, B => n1447, S => n1352, Z => n2857);
   U3184 : MUX2_X1 port map( A => n4882, B => n1444, S => n1352, Z => n2856);
   U3185 : MUX2_X1 port map( A => n4881, B => n1441, S => n1352, Z => n2855);
   U3186 : MUX2_X1 port map( A => n4880, B => n1438, S => n1352, Z => n2854);
   U3187 : MUX2_X1 port map( A => n4879, B => n1435, S => n1352, Z => n2853);
   U3188 : MUX2_X1 port map( A => n4878, B => n1432, S => n1352, Z => n2852);
   U3189 : MUX2_X1 port map( A => n4877, B => n1429, S => n1352, Z => n2851);
   U3190 : MUX2_X1 port map( A => n4876, B => n1426, S => n1352, Z => n2850);
   U3191 : MUX2_X1 port map( A => n4875, B => n1423, S => n1351, Z => n2849);
   U3192 : MUX2_X1 port map( A => n4874, B => n1421, S => n1351, Z => n2848);
   U3193 : MUX2_X1 port map( A => n4873, B => n1419, S => n1351, Z => n2847);
   U3194 : MUX2_X1 port map( A => n4872, B => n1417, S => n1351, Z => n2846);
   U3195 : MUX2_X1 port map( A => n4871, B => n1415, S => n1351, Z => n2845);
   U3196 : MUX2_X1 port map( A => n4870, B => n1413, S => n1351, Z => n2844);
   U3197 : MUX2_X1 port map( A => n4869, B => n1411, S => n1351, Z => n2843);
   U3198 : MUX2_X1 port map( A => n4868, B => n1409, S => n1351, Z => n2842);
   U3199 : MUX2_X1 port map( A => n4867, B => n1407, S => n1351, Z => n2841);
   U3200 : MUX2_X1 port map( A => n4866, B => n1405, S => n1351, Z => n2840);
   U3201 : MUX2_X1 port map( A => n4865, B => n1403, S => n1351, Z => n2839);
   U3202 : MUX2_X1 port map( A => n4864, B => n1401, S => n1351, Z => n2838);
   U3203 : MUX2_X1 port map( A => n4863, B => n1399, S => n1350, Z => n2837);
   U3204 : MUX2_X1 port map( A => n4862, B => n1397, S => n1350, Z => n2836);
   U3205 : MUX2_X1 port map( A => n4861, B => n1395, S => n1350, Z => n2835);
   U3206 : MUX2_X1 port map( A => n4860, B => n1393, S => n1350, Z => n2834);
   U3207 : MUX2_X1 port map( A => n4859, B => n1391, S => n1350, Z => n2833);
   U3208 : MUX2_X1 port map( A => n4858, B => n1389, S => n1350, Z => n2832);
   U3209 : MUX2_X1 port map( A => n4857, B => n1387, S => n1350, Z => n2831);
   U3210 : MUX2_X1 port map( A => n4856, B => n1385, S => n1350, Z => n2830);
   U3211 : MUX2_X1 port map( A => n4855, B => n1383, S => n1350, Z => n2829);
   U3212 : MUX2_X1 port map( A => n4854, B => n1381, S => n1350, Z => n2828);
   U3213 : MUX2_X1 port map( A => n4853, B => n1379, S => n1350, Z => n2827);
   U3214 : MUX2_X1 port map( A => n4852, B => n1377, S => n1350, Z => n2826);
   U3215 : AND2_X1 port map( A1 => n4497, A2 => n4354, ZN => n4568);
   U3216 : AND3_X1 port map( A1 => n4357, A2 => n4355, A3 => ADD_WR(4), ZN => 
                           n4497);
   U3217 : MUX2_X1 port map( A => n4851, B => n1447, S => n1355, Z => n2825);
   U3218 : MUX2_X1 port map( A => n4850, B => n1444, S => n1355, Z => n2824);
   U3219 : MUX2_X1 port map( A => n4849, B => n1441, S => n1355, Z => n2823);
   U3220 : MUX2_X1 port map( A => n4848, B => n1438, S => n1355, Z => n2822);
   U3221 : MUX2_X1 port map( A => n4847, B => n1435, S => n1355, Z => n2821);
   U3222 : MUX2_X1 port map( A => n4846, B => n1432, S => n1355, Z => n2820);
   U3223 : MUX2_X1 port map( A => n4845, B => n1429, S => n1355, Z => n2819);
   U3224 : MUX2_X1 port map( A => n4844, B => n1426, S => n1355, Z => n2818);
   U3225 : MUX2_X1 port map( A => n4843, B => n1423, S => n1354, Z => n2817);
   U3226 : MUX2_X1 port map( A => n4842, B => n1421, S => n1354, Z => n2816);
   U3227 : MUX2_X1 port map( A => n4841, B => n1419, S => n1354, Z => n2815);
   U3228 : MUX2_X1 port map( A => n4840, B => n1417, S => n1354, Z => n2814);
   U3229 : MUX2_X1 port map( A => n4839, B => n1415, S => n1354, Z => n2813);
   U3230 : MUX2_X1 port map( A => n4838, B => n1413, S => n1354, Z => n2812);
   U3231 : MUX2_X1 port map( A => n4837, B => n1411, S => n1354, Z => n2811);
   U3232 : MUX2_X1 port map( A => n4836, B => n1409, S => n1354, Z => n2810);
   U3233 : MUX2_X1 port map( A => n4835, B => n1407, S => n1354, Z => n2809);
   U3234 : MUX2_X1 port map( A => n4834, B => n1405, S => n1354, Z => n2808);
   U3235 : MUX2_X1 port map( A => n4833, B => n1403, S => n1354, Z => n2807);
   U3236 : MUX2_X1 port map( A => n4832, B => n1401, S => n1354, Z => n2806);
   U3237 : MUX2_X1 port map( A => n4831, B => n1399, S => n1353, Z => n2805);
   U3238 : MUX2_X1 port map( A => n4830, B => n1397, S => n1353, Z => n2804);
   U3239 : MUX2_X1 port map( A => n4829, B => n1395, S => n1353, Z => n2803);
   U3240 : MUX2_X1 port map( A => n4828, B => n1393, S => n1353, Z => n2802);
   U3241 : MUX2_X1 port map( A => n4827, B => n1391, S => n1353, Z => n2801);
   U3242 : MUX2_X1 port map( A => n4826, B => n1389, S => n1353, Z => n2800);
   U3243 : MUX2_X1 port map( A => n4825, B => n1387, S => n1353, Z => n2799);
   U3244 : MUX2_X1 port map( A => n4824, B => n1385, S => n1353, Z => n2798);
   U3245 : MUX2_X1 port map( A => n4823, B => n1383, S => n1353, Z => n2797);
   U3246 : MUX2_X1 port map( A => n4822, B => n1381, S => n1353, Z => n2796);
   U3247 : MUX2_X1 port map( A => n4821, B => n1379, S => n1353, Z => n2795);
   U3248 : MUX2_X1 port map( A => n4820, B => n1377, S => n1353, Z => n2794);
   U3249 : AND2_X1 port map( A1 => n4570, A2 => n4392, ZN => n4569);
   U3250 : MUX2_X1 port map( A => n4819, B => n1447, S => n1358, Z => n2793);
   U3251 : MUX2_X1 port map( A => n4818, B => n1444, S => n1358, Z => n2792);
   U3252 : MUX2_X1 port map( A => n4817, B => n1441, S => n1358, Z => n2791);
   U3253 : MUX2_X1 port map( A => n4816, B => n1438, S => n1358, Z => n2790);
   U3254 : MUX2_X1 port map( A => n4815, B => n1435, S => n1358, Z => n2789);
   U3255 : MUX2_X1 port map( A => n4814, B => n1432, S => n1358, Z => n2788);
   U3256 : MUX2_X1 port map( A => n4813, B => n1429, S => n1358, Z => n2787);
   U3257 : MUX2_X1 port map( A => n4812, B => n1426, S => n1358, Z => n2786);
   U3258 : MUX2_X1 port map( A => n4811, B => n1423, S => n1357, Z => n2785);
   U3259 : MUX2_X1 port map( A => n4810, B => n1421, S => n1357, Z => n2784);
   U3260 : MUX2_X1 port map( A => n4809, B => n1419, S => n1357, Z => n2783);
   U3261 : MUX2_X1 port map( A => n4808, B => n1417, S => n1357, Z => n2782);
   U3262 : MUX2_X1 port map( A => n4807, B => n1415, S => n1357, Z => n2781);
   U3263 : MUX2_X1 port map( A => n4806, B => n1413, S => n1357, Z => n2780);
   U3264 : MUX2_X1 port map( A => n4805, B => n1411, S => n1357, Z => n2779);
   U3265 : MUX2_X1 port map( A => n4804, B => n1409, S => n1357, Z => n2778);
   U3266 : MUX2_X1 port map( A => n4803, B => n1407, S => n1357, Z => n2777);
   U3267 : MUX2_X1 port map( A => n4802, B => n1405, S => n1357, Z => n2776);
   U3268 : MUX2_X1 port map( A => n4801, B => n1403, S => n1357, Z => n2775);
   U3269 : MUX2_X1 port map( A => n4800, B => n1401, S => n1357, Z => n2774);
   U3270 : MUX2_X1 port map( A => n4799, B => n1399, S => n1356, Z => n2773);
   U3271 : MUX2_X1 port map( A => n4798, B => n1397, S => n1356, Z => n2772);
   U3272 : MUX2_X1 port map( A => n4797, B => n1395, S => n1356, Z => n2771);
   U3273 : MUX2_X1 port map( A => n4796, B => n1393, S => n1356, Z => n2770);
   U3274 : MUX2_X1 port map( A => n4795, B => n1391, S => n1356, Z => n2769);
   U3275 : MUX2_X1 port map( A => n4794, B => n1389, S => n1356, Z => n2768);
   U3276 : MUX2_X1 port map( A => n4793, B => n1387, S => n1356, Z => n2767);
   U3277 : MUX2_X1 port map( A => n4792, B => n1385, S => n1356, Z => n2766);
   U3278 : MUX2_X1 port map( A => n4791, B => n1383, S => n1356, Z => n2765);
   U3279 : MUX2_X1 port map( A => n4790, B => n1381, S => n1356, Z => n2764);
   U3280 : MUX2_X1 port map( A => n4789, B => n1379, S => n1356, Z => n2763);
   U3281 : MUX2_X1 port map( A => n4788, B => n1377, S => n1356, Z => n2762);
   U3282 : AND2_X1 port map( A1 => n4570, A2 => n4341, ZN => n4571);
   U3283 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => n4572, ZN 
                           => n4341);
   U3284 : MUX2_X1 port map( A => n4288, B => n1447, S => n1361, Z => n2761);
   U3285 : MUX2_X1 port map( A => n4289, B => n1444, S => n1361, Z => n2760);
   U3286 : MUX2_X1 port map( A => n4290, B => n1441, S => n1361, Z => n2759);
   U3287 : MUX2_X1 port map( A => n4291, B => n1438, S => n1361, Z => n2758);
   U3288 : MUX2_X1 port map( A => n4292, B => n1435, S => n1361, Z => n2757);
   U3289 : MUX2_X1 port map( A => n4293, B => n1432, S => n1361, Z => n2756);
   U3290 : MUX2_X1 port map( A => n4294, B => n1429, S => n1361, Z => n2755);
   U3291 : MUX2_X1 port map( A => n4295, B => n1426, S => n1361, Z => n2754);
   U3292 : MUX2_X1 port map( A => n4296, B => n1423, S => n1360, Z => n2753);
   U3293 : MUX2_X1 port map( A => n4297, B => n1421, S => n1360, Z => n2752);
   U3294 : MUX2_X1 port map( A => n224, B => n1419, S => n1360, Z => n2751);
   U3295 : MUX2_X1 port map( A => n4298, B => n1417, S => n1360, Z => n2750);
   U3296 : MUX2_X1 port map( A => n343, B => n1415, S => n1360, Z => n2749);
   U3297 : MUX2_X1 port map( A => n344, B => n1413, S => n1360, Z => n2748);
   U3298 : MUX2_X1 port map( A => n225, B => n1411, S => n1360, Z => n2747);
   U3299 : MUX2_X1 port map( A => n4299, B => n1409, S => n1360, Z => n2746);
   U3300 : MUX2_X1 port map( A => n345, B => n1407, S => n1360, Z => n2745);
   U3301 : MUX2_X1 port map( A => n4300, B => n1405, S => n1360, Z => n2744);
   U3302 : MUX2_X1 port map( A => n4301, B => n1403, S => n1360, Z => n2743);
   U3303 : MUX2_X1 port map( A => n346, B => n1401, S => n1360, Z => n2742);
   U3304 : MUX2_X1 port map( A => n4302, B => n1399, S => n1359, Z => n2741);
   U3305 : MUX2_X1 port map( A => n226, B => n1397, S => n1359, Z => n2740);
   U3306 : MUX2_X1 port map( A => n4303, B => n1395, S => n1359, Z => n2739);
   U3307 : MUX2_X1 port map( A => n347, B => n1393, S => n1359, Z => n2738);
   U3308 : MUX2_X1 port map( A => n4304, B => n1391, S => n1359, Z => n2737);
   U3309 : MUX2_X1 port map( A => n4305, B => n1389, S => n1359, Z => n2736);
   U3310 : MUX2_X1 port map( A => n351, B => n1387, S => n1359, Z => n2735);
   U3311 : MUX2_X1 port map( A => n348, B => n1385, S => n1359, Z => n2734);
   U3312 : MUX2_X1 port map( A => n349, B => n1383, S => n1359, Z => n2733);
   U3313 : MUX2_X1 port map( A => n4306, B => n1381, S => n1359, Z => n2732);
   U3314 : MUX2_X1 port map( A => n350, B => n1379, S => n1359, Z => n2731);
   U3315 : MUX2_X1 port map( A => n4307, B => n1377, S => n1359, Z => n2730);
   U3316 : AND2_X1 port map( A1 => n4570, A2 => n4344, ZN => n4573);
   U3317 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(2), A3 => n4574, ZN 
                           => n4344);
   U3318 : INV_X1 port map( A => n4575, ZN => n2729);
   U3319 : MUX2_X1 port map( A => n837, B => n1448, S => n1364, Z => n4575);
   U3320 : INV_X1 port map( A => n4577, ZN => n2728);
   U3321 : MUX2_X1 port map( A => n838, B => n1445, S => n1364, Z => n4577);
   U3322 : INV_X1 port map( A => n4578, ZN => n2727);
   U3323 : MUX2_X1 port map( A => n839, B => n1442, S => n1364, Z => n4578);
   U3324 : INV_X1 port map( A => n4579, ZN => n2726);
   U3325 : MUX2_X1 port map( A => n840, B => n1439, S => n1364, Z => n4579);
   U3326 : INV_X1 port map( A => n4580, ZN => n2725);
   U3327 : MUX2_X1 port map( A => n841, B => n1436, S => n1364, Z => n4580);
   U3328 : INV_X1 port map( A => n4581, ZN => n2724);
   U3329 : MUX2_X1 port map( A => n842, B => n1433, S => n1364, Z => n4581);
   U3330 : INV_X1 port map( A => n4582, ZN => n2723);
   U3331 : MUX2_X1 port map( A => n843, B => n1430, S => n1364, Z => n4582);
   U3332 : INV_X1 port map( A => n4583, ZN => n2722);
   U3333 : MUX2_X1 port map( A => n844, B => n1427, S => n1364, Z => n4583);
   U3334 : INV_X1 port map( A => n4584, ZN => n2721);
   U3335 : MUX2_X1 port map( A => n845, B => n1424, S => n1363, Z => n4584);
   U3336 : INV_X1 port map( A => n4585, ZN => n2720);
   U3337 : MUX2_X1 port map( A => n846, B => n1422, S => n1363, Z => n4585);
   U3338 : INV_X1 port map( A => n4586, ZN => n2719);
   U3339 : MUX2_X1 port map( A => n847, B => n1420, S => n1363, Z => n4586);
   U3340 : INV_X1 port map( A => n4587, ZN => n2718);
   U3341 : MUX2_X1 port map( A => n848, B => n1418, S => n1363, Z => n4587);
   U3342 : INV_X1 port map( A => n4588, ZN => n2717);
   U3343 : MUX2_X1 port map( A => n849, B => n1416, S => n1363, Z => n4588);
   U3344 : INV_X1 port map( A => n4589, ZN => n2716);
   U3345 : MUX2_X1 port map( A => n850, B => n1414, S => n1363, Z => n4589);
   U3346 : INV_X1 port map( A => n4590, ZN => n2715);
   U3347 : MUX2_X1 port map( A => n851, B => n1412, S => n1363, Z => n4590);
   U3348 : INV_X1 port map( A => n4591, ZN => n2714);
   U3349 : MUX2_X1 port map( A => n852, B => n1410, S => n1363, Z => n4591);
   U3350 : INV_X1 port map( A => n4592, ZN => n2713);
   U3351 : MUX2_X1 port map( A => n853, B => n1408, S => n1363, Z => n4592);
   U3352 : INV_X1 port map( A => n4593, ZN => n2712);
   U3353 : MUX2_X1 port map( A => n854, B => n1406, S => n1363, Z => n4593);
   U3354 : INV_X1 port map( A => n4594, ZN => n2711);
   U3355 : MUX2_X1 port map( A => n855, B => n1404, S => n1363, Z => n4594);
   U3356 : INV_X1 port map( A => n4595, ZN => n2710);
   U3357 : MUX2_X1 port map( A => n856, B => n1402, S => n1363, Z => n4595);
   U3358 : INV_X1 port map( A => n4596, ZN => n2709);
   U3359 : MUX2_X1 port map( A => n857, B => n1400, S => n1362, Z => n4596);
   U3360 : INV_X1 port map( A => n4597, ZN => n2708);
   U3361 : MUX2_X1 port map( A => n858, B => n1398, S => n1362, Z => n4597);
   U3362 : INV_X1 port map( A => n4598, ZN => n2707);
   U3363 : MUX2_X1 port map( A => n859, B => n1396, S => n1362, Z => n4598);
   U3364 : INV_X1 port map( A => n4599, ZN => n2706);
   U3365 : MUX2_X1 port map( A => n860, B => n1394, S => n1362, Z => n4599);
   U3366 : INV_X1 port map( A => n4600, ZN => n2705);
   U3367 : MUX2_X1 port map( A => n861, B => n1392, S => n1362, Z => n4600);
   U3368 : INV_X1 port map( A => n4601, ZN => n2704);
   U3369 : MUX2_X1 port map( A => n862, B => n1390, S => n1362, Z => n4601);
   U3370 : INV_X1 port map( A => n4602, ZN => n2703);
   U3371 : MUX2_X1 port map( A => n863, B => n1388, S => n1362, Z => n4602);
   U3372 : INV_X1 port map( A => n4603, ZN => n2702);
   U3373 : MUX2_X1 port map( A => n864, B => n1386, S => n1362, Z => n4603);
   U3374 : INV_X1 port map( A => n4604, ZN => n2701);
   U3375 : MUX2_X1 port map( A => n865, B => n1384, S => n1362, Z => n4604);
   U3376 : INV_X1 port map( A => n4605, ZN => n2700);
   U3377 : MUX2_X1 port map( A => n866, B => n1382, S => n1362, Z => n4605);
   U3378 : INV_X1 port map( A => n4606, ZN => n2699);
   U3379 : MUX2_X1 port map( A => n867, B => n1380, S => n1362, Z => n4606);
   U3380 : INV_X1 port map( A => n4607, ZN => n2698);
   U3381 : MUX2_X1 port map( A => n868, B => n1378, S => n1362, Z => n4607);
   U3382 : AND2_X1 port map( A1 => n4570, A2 => n4346, ZN => n4576);
   U3383 : NOR3_X1 port map( A1 => n4572, A2 => ADD_WR(2), A3 => n4574, ZN => 
                           n4346);
   U3384 : MUX2_X1 port map( A => n4787, B => n1447, S => n1367, Z => n2697);
   U3385 : MUX2_X1 port map( A => n4786, B => n1444, S => n1367, Z => n2696);
   U3386 : MUX2_X1 port map( A => n4785, B => n1441, S => n1367, Z => n2695);
   U3387 : MUX2_X1 port map( A => n4784, B => n1438, S => n1367, Z => n2694);
   U3388 : MUX2_X1 port map( A => n4783, B => n1435, S => n1367, Z => n2693);
   U3389 : MUX2_X1 port map( A => n4782, B => n1432, S => n1367, Z => n2692);
   U3390 : MUX2_X1 port map( A => n4781, B => n1429, S => n1367, Z => n2691);
   U3391 : MUX2_X1 port map( A => n4780, B => n1426, S => n1367, Z => n2690);
   U3392 : MUX2_X1 port map( A => n4779, B => n1423, S => n1366, Z => n2689);
   U3393 : MUX2_X1 port map( A => n4778, B => n1421, S => n1366, Z => n2688);
   U3394 : MUX2_X1 port map( A => n4777, B => n1419, S => n1366, Z => n2687);
   U3395 : MUX2_X1 port map( A => n4776, B => n1417, S => n1366, Z => n2686);
   U3396 : MUX2_X1 port map( A => n4775, B => n1415, S => n1366, Z => n2685);
   U3397 : MUX2_X1 port map( A => n4774, B => n1413, S => n1366, Z => n2684);
   U3398 : MUX2_X1 port map( A => n4773, B => n1411, S => n1366, Z => n2683);
   U3399 : MUX2_X1 port map( A => n4772, B => n1409, S => n1366, Z => n2682);
   U3400 : MUX2_X1 port map( A => n4771, B => n1407, S => n1366, Z => n2681);
   U3401 : MUX2_X1 port map( A => n4770, B => n1405, S => n1366, Z => n2680);
   U3402 : MUX2_X1 port map( A => n4769, B => n1403, S => n1366, Z => n2679);
   U3403 : MUX2_X1 port map( A => n4768, B => n1401, S => n1366, Z => n2678);
   U3404 : MUX2_X1 port map( A => n4767, B => n1399, S => n1365, Z => n2677);
   U3405 : MUX2_X1 port map( A => n4766, B => n1397, S => n1365, Z => n2676);
   U3406 : MUX2_X1 port map( A => n4765, B => n1395, S => n1365, Z => n2675);
   U3407 : MUX2_X1 port map( A => n4764, B => n1393, S => n1365, Z => n2674);
   U3408 : MUX2_X1 port map( A => n4763, B => n1391, S => n1365, Z => n2673);
   U3409 : MUX2_X1 port map( A => n4762, B => n1389, S => n1365, Z => n2672);
   U3410 : MUX2_X1 port map( A => n4761, B => n1387, S => n1365, Z => n2671);
   U3411 : MUX2_X1 port map( A => n4760, B => n1385, S => n1365, Z => n2670);
   U3412 : MUX2_X1 port map( A => n4759, B => n1383, S => n1365, Z => n2669);
   U3413 : MUX2_X1 port map( A => n4758, B => n1381, S => n1365, Z => n2668);
   U3414 : MUX2_X1 port map( A => n4757, B => n1379, S => n1365, Z => n2667);
   U3415 : MUX2_X1 port map( A => n4756, B => n1377, S => n1365, Z => n2666);
   U3416 : AND2_X1 port map( A1 => n4570, A2 => n4348, ZN => n4608);
   U3417 : AND3_X1 port map( A1 => n4572, A2 => n4574, A3 => ADD_WR(2), ZN => 
                           n4348);
   U3418 : MUX2_X1 port map( A => n4755, B => n1447, S => n1370, Z => n2665);
   U3419 : MUX2_X1 port map( A => n4754, B => n1444, S => n1370, Z => n2664);
   U3420 : MUX2_X1 port map( A => n4753, B => n1441, S => n1370, Z => n2663);
   U3421 : MUX2_X1 port map( A => n4752, B => n1438, S => n1370, Z => n2662);
   U3422 : MUX2_X1 port map( A => n4751, B => n1435, S => n1370, Z => n2661);
   U3423 : MUX2_X1 port map( A => n4750, B => n1432, S => n1370, Z => n2660);
   U3424 : MUX2_X1 port map( A => n4749, B => n1429, S => n1370, Z => n2659);
   U3425 : MUX2_X1 port map( A => n4748, B => n1426, S => n1370, Z => n2658);
   U3426 : MUX2_X1 port map( A => n4747, B => n1423, S => n1369, Z => n2657);
   U3427 : MUX2_X1 port map( A => n4746, B => n1421, S => n1369, Z => n2656);
   U3428 : MUX2_X1 port map( A => n4745, B => n1419, S => n1369, Z => n2655);
   U3429 : MUX2_X1 port map( A => n4744, B => n1417, S => n1369, Z => n2654);
   U3430 : MUX2_X1 port map( A => n4743, B => n1415, S => n1369, Z => n2653);
   U3431 : MUX2_X1 port map( A => n4742, B => n1413, S => n1369, Z => n2652);
   U3432 : MUX2_X1 port map( A => n4741, B => n1411, S => n1369, Z => n2651);
   U3433 : MUX2_X1 port map( A => n4740, B => n1409, S => n1369, Z => n2650);
   U3434 : MUX2_X1 port map( A => n4739, B => n1407, S => n1369, Z => n2649);
   U3435 : MUX2_X1 port map( A => n4738, B => n1405, S => n1369, Z => n2648);
   U3436 : MUX2_X1 port map( A => n4737, B => n1403, S => n1369, Z => n2647);
   U3437 : MUX2_X1 port map( A => n4736, B => n1401, S => n1369, Z => n2646);
   U3438 : MUX2_X1 port map( A => n4735, B => n1399, S => n1368, Z => n2645);
   U3439 : MUX2_X1 port map( A => n4734, B => n1397, S => n1368, Z => n2644);
   U3440 : MUX2_X1 port map( A => n4733, B => n1395, S => n1368, Z => n2643);
   U3441 : MUX2_X1 port map( A => n4732, B => n1393, S => n1368, Z => n2642);
   U3442 : MUX2_X1 port map( A => n4731, B => n1391, S => n1368, Z => n2641);
   U3443 : MUX2_X1 port map( A => n4730, B => n1389, S => n1368, Z => n2640);
   U3444 : MUX2_X1 port map( A => n4729, B => n1387, S => n1368, Z => n2639);
   U3445 : MUX2_X1 port map( A => n4728, B => n1385, S => n1368, Z => n2638);
   U3446 : MUX2_X1 port map( A => n4727, B => n1383, S => n1368, Z => n2637);
   U3447 : MUX2_X1 port map( A => n4726, B => n1381, S => n1368, Z => n2636);
   U3448 : MUX2_X1 port map( A => n4725, B => n1379, S => n1368, Z => n2635);
   U3449 : MUX2_X1 port map( A => n4724, B => n1377, S => n1368, Z => n2634);
   U3450 : AND2_X1 port map( A1 => n4570, A2 => n4350, ZN => n4609);
   U3451 : AND3_X1 port map( A1 => ADD_WR(0), A2 => n4574, A3 => ADD_WR(2), ZN 
                           => n4350);
   U3452 : INV_X1 port map( A => n4610, ZN => n2633);
   U3453 : MUX2_X1 port map( A => n933, B => n1448, S => n1373, Z => n4610);
   U3454 : INV_X1 port map( A => n4612, ZN => n2632);
   U3455 : MUX2_X1 port map( A => n934, B => n1445, S => n1373, Z => n4612);
   U3456 : INV_X1 port map( A => n4613, ZN => n2631);
   U3457 : MUX2_X1 port map( A => n935, B => n1442, S => n1373, Z => n4613);
   U3458 : INV_X1 port map( A => n4614, ZN => n2630);
   U3459 : MUX2_X1 port map( A => n936, B => n1439, S => n1373, Z => n4614);
   U3460 : INV_X1 port map( A => n4615, ZN => n2629);
   U3461 : MUX2_X1 port map( A => n937, B => n1436, S => n1373, Z => n4615);
   U3462 : INV_X1 port map( A => n4616, ZN => n2628);
   U3463 : MUX2_X1 port map( A => n938, B => n1433, S => n1373, Z => n4616);
   U3464 : INV_X1 port map( A => n4617, ZN => n2627);
   U3465 : MUX2_X1 port map( A => n939, B => n1430, S => n1373, Z => n4617);
   U3466 : INV_X1 port map( A => n4618, ZN => n2626);
   U3467 : MUX2_X1 port map( A => n940, B => n1427, S => n1373, Z => n4618);
   U3468 : INV_X1 port map( A => n4619, ZN => n2625);
   U3469 : MUX2_X1 port map( A => n941, B => n1424, S => n1372, Z => n4619);
   U3470 : INV_X1 port map( A => n4620, ZN => n2624);
   U3471 : MUX2_X1 port map( A => n942, B => n1422, S => n1372, Z => n4620);
   U3472 : INV_X1 port map( A => n4621, ZN => n2623);
   U3473 : MUX2_X1 port map( A => n943, B => n1420, S => n1372, Z => n4621);
   U3474 : INV_X1 port map( A => n4622, ZN => n2622);
   U3475 : MUX2_X1 port map( A => n944, B => n1418, S => n1372, Z => n4622);
   U3476 : INV_X1 port map( A => n4623, ZN => n2621);
   U3477 : MUX2_X1 port map( A => n945, B => n1416, S => n1372, Z => n4623);
   U3478 : INV_X1 port map( A => n4624, ZN => n2620);
   U3479 : MUX2_X1 port map( A => n946, B => n1414, S => n1372, Z => n4624);
   U3480 : INV_X1 port map( A => n4625, ZN => n2619);
   U3481 : MUX2_X1 port map( A => n947, B => n1412, S => n1372, Z => n4625);
   U3482 : INV_X1 port map( A => n4626, ZN => n2618);
   U3483 : MUX2_X1 port map( A => n948, B => n1410, S => n1372, Z => n4626);
   U3484 : INV_X1 port map( A => n4627, ZN => n2617);
   U3485 : MUX2_X1 port map( A => n949, B => n1408, S => n1372, Z => n4627);
   U3486 : INV_X1 port map( A => n4628, ZN => n2616);
   U3487 : MUX2_X1 port map( A => n950, B => n1406, S => n1372, Z => n4628);
   U3488 : INV_X1 port map( A => n4629, ZN => n2615);
   U3489 : MUX2_X1 port map( A => n951, B => n1404, S => n1372, Z => n4629);
   U3490 : INV_X1 port map( A => n4630, ZN => n2614);
   U3491 : MUX2_X1 port map( A => n952, B => n1402, S => n1372, Z => n4630);
   U3492 : INV_X1 port map( A => n4631, ZN => n2613);
   U3493 : MUX2_X1 port map( A => n953, B => n1400, S => n1371, Z => n4631);
   U3494 : INV_X1 port map( A => n4632, ZN => n2612);
   U3495 : MUX2_X1 port map( A => n954, B => n1398, S => n1371, Z => n4632);
   U3496 : INV_X1 port map( A => n4633, ZN => n2611);
   U3497 : MUX2_X1 port map( A => n955, B => n1396, S => n1371, Z => n4633);
   U3498 : INV_X1 port map( A => n4634, ZN => n2610);
   U3499 : MUX2_X1 port map( A => n956, B => n1394, S => n1371, Z => n4634);
   U3500 : INV_X1 port map( A => n4635, ZN => n2609);
   U3501 : MUX2_X1 port map( A => n957, B => n1392, S => n1371, Z => n4635);
   U3502 : INV_X1 port map( A => n4636, ZN => n2608);
   U3503 : MUX2_X1 port map( A => n958, B => n1390, S => n1371, Z => n4636);
   U3504 : INV_X1 port map( A => n4637, ZN => n2607);
   U3505 : MUX2_X1 port map( A => n959, B => n1388, S => n1371, Z => n4637);
   U3506 : INV_X1 port map( A => n4638, ZN => n2606);
   U3507 : MUX2_X1 port map( A => n960, B => n1386, S => n1371, Z => n4638);
   U3508 : INV_X1 port map( A => n4639, ZN => n2605);
   U3509 : MUX2_X1 port map( A => n961, B => n1384, S => n1371, Z => n4639);
   U3510 : INV_X1 port map( A => n4640, ZN => n2604);
   U3511 : MUX2_X1 port map( A => n962, B => n1382, S => n1371, Z => n4640);
   U3512 : INV_X1 port map( A => n4641, ZN => n2603);
   U3513 : MUX2_X1 port map( A => n963, B => n1380, S => n1371, Z => n4641);
   U3514 : INV_X1 port map( A => n4642, ZN => n2602);
   U3515 : MUX2_X1 port map( A => n964, B => n1378, S => n1371, Z => n4642);
   U3516 : AND2_X1 port map( A1 => n4570, A2 => n4352, ZN => n4611);
   U3517 : AND3_X1 port map( A1 => ADD_WR(1), A2 => n4572, A3 => ADD_WR(2), ZN 
                           => n4352);
   U3518 : MUX2_X1 port map( A => n4308, B => n1446, S => n1376, Z => n2601);
   U3519 : MUX2_X1 port map( A => n4309, B => n1443, S => n1376, Z => n2600);
   U3520 : MUX2_X1 port map( A => n4310, B => n1440, S => n1376, Z => n2599);
   U3521 : MUX2_X1 port map( A => n4311, B => n1437, S => n1376, Z => n2598);
   U3522 : MUX2_X1 port map( A => n4312, B => n1434, S => n1376, Z => n2597);
   U3523 : MUX2_X1 port map( A => n4313, B => n1431, S => n1376, Z => n2596);
   U3524 : MUX2_X1 port map( A => n4314, B => n1428, S => n1376, Z => n2595);
   U3525 : MUX2_X1 port map( A => n4315, B => n1425, S => n1376, Z => n2594);
   U3526 : MUX2_X1 port map( A => n4316, B => n1423, S => n1375, Z => n2593);
   U3527 : MUX2_X1 port map( A => n4317, B => n1421, S => n1375, Z => n2592);
   U3528 : MUX2_X1 port map( A => n4318, B => n1419, S => n1375, Z => n2591);
   U3529 : MUX2_X1 port map( A => n4319, B => n1417, S => n1375, Z => n2590);
   U3530 : MUX2_X1 port map( A => n4320, B => n1415, S => n1375, Z => n2589);
   U3531 : MUX2_X1 port map( A => n4321, B => n1413, S => n1375, Z => n2588);
   U3532 : MUX2_X1 port map( A => n4322, B => n1411, S => n1375, Z => n2587);
   U3533 : MUX2_X1 port map( A => n4323, B => n1409, S => n1375, Z => n2586);
   U3534 : MUX2_X1 port map( A => n4324, B => n1407, S => n1375, Z => n2585);
   U3535 : MUX2_X1 port map( A => n4325, B => n1405, S => n1375, Z => n2584);
   U3536 : MUX2_X1 port map( A => n4326, B => n1403, S => n1375, Z => n2583);
   U3537 : MUX2_X1 port map( A => n4327, B => n1401, S => n1375, Z => n2582);
   U3538 : MUX2_X1 port map( A => n4328, B => n1399, S => n1374, Z => n2581);
   U3539 : MUX2_X1 port map( A => n4329, B => n1397, S => n1374, Z => n2580);
   U3540 : MUX2_X1 port map( A => n4330, B => n1395, S => n1374, Z => n2579);
   U3541 : MUX2_X1 port map( A => n4331, B => n1393, S => n1374, Z => n2578);
   U3542 : MUX2_X1 port map( A => n4332, B => n1391, S => n1374, Z => n2577);
   U3543 : MUX2_X1 port map( A => n4333, B => n1389, S => n1374, Z => n2576);
   U3544 : MUX2_X1 port map( A => n4334, B => n1387, S => n1374, Z => n2575);
   U3545 : MUX2_X1 port map( A => n4335, B => n1385, S => n1374, Z => n2574);
   U3546 : MUX2_X1 port map( A => n4336, B => n1383, S => n1374, Z => n2573);
   U3547 : MUX2_X1 port map( A => n4337, B => n1381, S => n1374, Z => n2572);
   U3548 : MUX2_X1 port map( A => n4338, B => n1379, S => n1374, Z => n2571);
   U3549 : MUX2_X1 port map( A => n4339, B => n1377, S => n1374, Z => n2570);
   U3550 : AND2_X1 port map( A1 => n4570, A2 => n4354, ZN => n4643);
   U3551 : AND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2),
                           ZN => n4354);
   U3552 : AND3_X1 port map( A1 => ADD_WR(3), A2 => n4357, A3 => ADD_WR(4), ZN 
                           => n4570);
   U3553 : NOR2_X1 port map( A1 => n4644, A2 => n4645, ZN => n4357);
   U3554 : INV_X1 port map( A => ENABLE, ZN => n4644);
   U3555 : XNOR2_X1 port map( A => ADD_RS2(1), B => n4574, ZN => n4651);
   U3556 : XNOR2_X1 port map( A => ADD_RS2(0), B => n4572, ZN => n4650);
   U3557 : XNOR2_X1 port map( A => ADD_RS2(3), B => ADD_WR(3), ZN => n4648);
   U3558 : XNOR2_X1 port map( A => ADD_RS2(4), B => ADD_WR(4), ZN => n4647);
   U3559 : XNOR2_X1 port map( A => ADD_RS2(2), B => ADD_WR(2), ZN => n4646);
   U3560 : XNOR2_X1 port map( A => n4574, B => n784, ZN => n4657);
   U3561 : INV_X1 port map( A => ADD_WR(1), ZN => n4574);
   U3562 : OAI21_X1 port map( B1 => n4658, B2 => n4659, A => WR, ZN => n4645);
   U3563 : NAND2_X1 port map( A1 => n4355, A2 => n4356, ZN => n4659);
   U3564 : INV_X1 port map( A => ADD_WR(4), ZN => n4356);
   U3565 : INV_X1 port map( A => ADD_WR(3), ZN => n4355);
   U3566 : INV_X1 port map( A => n4392, ZN => n4658);
   U3567 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => ADD_WR(0),
                           ZN => n4392);
   U3568 : XNOR2_X1 port map( A => ADD_RS1(0), B => n4572, ZN => n4656);
   U3569 : INV_X1 port map( A => ADD_WR(0), ZN => n4572);
   U3570 : XNOR2_X1 port map( A => n84, B => ADD_WR(3), ZN => n4654);
   U3571 : XNOR2_X1 port map( A => n1092, B => ADD_WR(4), ZN => n4653);
   U3572 : XNOR2_X1 port map( A => n764, B => ADD_WR(2), ZN => n4652);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT5_0 is

   port( A, B : in std_logic_vector (4 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (4 downto 0));

end mux21_NBIT5_0;

architecture SYN_bhv of mux21_NBIT5_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8, n9, n10, n11, n1, n2 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => S, Z => n1);
   U2 : INV_X1 port map( A => n10, ZN => Z(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n2, B1 => B(1), B2 => n1, ZN => 
                           n10);
   U4 : INV_X1 port map( A => n9, ZN => Z(2));
   U5 : INV_X1 port map( A => n7, ZN => Z(4));
   U6 : INV_X1 port map( A => n11, ZN => Z(0));
   U7 : INV_X1 port map( A => n8, ZN => Z(3));
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n2, B1 => B(3), B2 => n1, ZN => n8
                           );
   U9 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => n1, ZN => n9
                           );
   U10 : AOI22_X1 port map( A1 => A(4), A2 => n2, B1 => S, B2 => B(4), ZN => n7
                           );
   U11 : AOI22_X1 port map( A1 => A(0), A2 => n2, B1 => B(0), B2 => n1, ZN => 
                           n11);
   U12 : INV_X1 port map( A => S, ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_0 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_0;

architecture SYN_bhv of regn_N5_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15 : 
      std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n15, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n10);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n14, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n9);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n13, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n8);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n12, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n7);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n11, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n6);
   U2 : OAI21_X1 port map( B1 => n7, B2 => EN, A => n2, ZN => n12);
   U3 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n2);
   U4 : OAI21_X1 port map( B1 => n8, B2 => EN, A => n3, ZN => n13);
   U5 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n3);
   U6 : OAI21_X1 port map( B1 => n9, B2 => EN, A => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n4);
   U8 : OAI21_X1 port map( B1 => n10, B2 => EN, A => n5, ZN => n15);
   U9 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n5);
   U10 : OAI21_X1 port map( B1 => n6, B2 => EN, A => n1, ZN => n11);
   U11 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n1);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity instruction_decomposition is

   port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype : in
         std_logic;  ADD_RS1, ADD_RS2, ADD_WR : out std_logic_vector (4 downto 
         0);  IMM : out std_logic_vector (31 downto 0);  RD1, RD2 : out 
         std_logic);

end instruction_decomposition;

architecture SYN_bhv of instruction_decomposition is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal IMM_24_port, IMM_23_port, IMM_22_port, IMM_21_port, IMM_20_port, 
      IMM_19_port, IMM_18_port, IMM_17_port, IMM_16_port, IMM_15_port, 
      IMM_14_port, IMM_13_port, IMM_12_port, IMM_11_port, IMM_10_port, 
      IMM_9_port, IMM_8_port, IMM_7_port, IMM_6_port, IMM_5_port, IMM_4_port, 
      IMM_3_port, IMM_2_port, IMM_1_port, IMM_0_port, n56, RD2_port, n33, n1, 
      RD1_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      IMM_31_port, n50, n51, n52, n53, n54, n55 : std_logic;

begin
   IMM <= ( IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, 
      IMM_31_port, IMM_31_port, IMM_24_port, IMM_23_port, IMM_22_port, 
      IMM_21_port, IMM_20_port, IMM_19_port, IMM_18_port, IMM_17_port, 
      IMM_16_port, IMM_15_port, IMM_14_port, IMM_13_port, IMM_12_port, 
      IMM_11_port, IMM_10_port, IMM_9_port, IMM_8_port, IMM_7_port, IMM_6_port,
      IMM_5_port, IMM_4_port, IMM_3_port, IMM_2_port, IMM_1_port, IMM_0_port );
   RD1 <= RD1_port;
   RD2 <= RD2_port;
   
   U3 : INV_X1 port map( A => RD1_port, ZN => n1);
   U4 : CLKBUF_X1 port map( A => n7, Z => RD1_port);
   U5 : CLKBUF_X1 port map( A => n1, Z => n3);
   U6 : BUF_X1 port map( A => n56, Z => n7);
   U7 : AND2_X1 port map( A1 => n56, A2 => INST_IN(23), ZN => ADD_RS1(2));
   U8 : NOR2_X1 port map( A1 => n17, A2 => n18, ZN => n4);
   U9 : NOR2_X1 port map( A1 => n19, A2 => n5, ZN => n20);
   U10 : INV_X1 port map( A => n4, ZN => n5);
   U11 : BUF_X1 port map( A => n31, Z => n8);
   U12 : AND2_X2 port map( A1 => n7, A2 => INST_IN(21), ZN => ADD_RS1(0));
   U13 : AND2_X2 port map( A1 => n41, A2 => n13, ZN => n14);
   U14 : AND2_X1 port map( A1 => n31, A2 => n12, ZN => n6);
   U15 : AND2_X1 port map( A1 => n31, A2 => n12, ZN => n15);
   U16 : INV_X1 port map( A => n16, ZN => n9);
   U17 : AOI211_X4 port map( C1 => n16, C2 => n13, A => n34, B => n15, ZN => 
                           ADD_RS2(1));
   U18 : CLKBUF_X1 port map( A => n13, Z => n10);
   U19 : NAND2_X1 port map( A1 => INST_IN(15), A2 => n24, ZN => n25);
   U20 : AND2_X1 port map( A1 => n29, A2 => n28, ZN => n11);
   U21 : INV_X1 port map( A => INST_IN(15), ZN => n51);
   U22 : INV_X1 port map( A => INST_IN(11), ZN => n55);
   U23 : INV_X1 port map( A => INST_IN(12), ZN => n54);
   U24 : INV_X1 port map( A => INST_IN(13), ZN => n53);
   U25 : INV_X1 port map( A => INST_IN(14), ZN => n52);
   U26 : CLKBUF_X1 port map( A => n40, Z => n12);
   U27 : BUF_X2 port map( A => n40, Z => n13);
   U28 : NAND2_X1 port map( A1 => n3, A2 => Jtype, ZN => n28);
   U29 : INV_X1 port map( A => n56, ZN => n45);
   U30 : NOR2_X1 port map( A1 => n43, A2 => n14, ZN => ADD_RS1(3));
   U31 : AND2_X2 port map( A1 => RD2_port, A2 => INST_IN(18), ZN => ADD_RS2(2))
                           ;
   U32 : INV_X1 port map( A => Itype, ZN => n16);
   U33 : NOR3_X1 port map( A1 => n14, A2 => n6, A3 => n36, ZN => ADD_RS2(3));
   U34 : OR4_X1 port map( A1 => n50, A2 => INST_IN(28), A3 => INST_IN(29), A4 
                           => INST_IN(31), ZN => n33);
   U35 : NOR3_X2 port map( A1 => n14, A2 => n6, A3 => n32, ZN => ADD_RS2(0));
   U36 : INV_X1 port map( A => INST_IN(28), ZN => n21);
   U37 : INV_X1 port map( A => INST_IN(30), ZN => n26);
   U38 : XOR2_X1 port map( A => INST_IN(26), B => INST_IN(27), Z => n19);
   U39 : INV_X1 port map( A => INST_IN(31), ZN => n18);
   U40 : INV_X1 port map( A => INST_IN(29), ZN => n17);
   U41 : NAND3_X1 port map( A1 => n20, A2 => n26, A3 => n21, ZN => n31);
   U42 : INV_X1 port map( A => Itype, ZN => n41);
   U43 : INV_X1 port map( A => Rtype, ZN => n40);
   U44 : OAI21_X1 port map( B1 => n8, B2 => n16, A => n13, ZN => RD2_port);
   U45 : NAND2_X1 port map( A1 => n41, A2 => n13, ZN => n56);
   U46 : OAI21_X1 port map( B1 => Jtype, B2 => n9, A => n10, ZN => n23);
   U47 : INV_X1 port map( A => n23, ZN => n22);
   U48 : AND2_X1 port map( A1 => INST_IN(0), A2 => n22, ZN => IMM_0_port);
   U49 : AND2_X1 port map( A1 => INST_IN(1), A2 => n22, ZN => IMM_1_port);
   U50 : AND2_X1 port map( A1 => INST_IN(2), A2 => n22, ZN => IMM_2_port);
   U51 : AND2_X1 port map( A1 => INST_IN(3), A2 => n22, ZN => IMM_3_port);
   U52 : AND2_X1 port map( A1 => INST_IN(4), A2 => n22, ZN => IMM_4_port);
   U53 : AND2_X1 port map( A1 => INST_IN(5), A2 => n22, ZN => IMM_5_port);
   U54 : AND2_X1 port map( A1 => INST_IN(6), A2 => n22, ZN => IMM_6_port);
   U55 : AND2_X1 port map( A1 => INST_IN(7), A2 => n22, ZN => IMM_7_port);
   U56 : AND2_X1 port map( A1 => INST_IN(8), A2 => n22, ZN => IMM_8_port);
   U57 : AND2_X1 port map( A1 => INST_IN(9), A2 => n22, ZN => IMM_9_port);
   U58 : AND2_X1 port map( A1 => INST_IN(10), A2 => n22, ZN => IMM_10_port);
   U59 : NOR2_X1 port map( A1 => n55, A2 => n23, ZN => IMM_11_port);
   U60 : NOR2_X1 port map( A1 => n54, A2 => n23, ZN => IMM_12_port);
   U61 : NOR2_X1 port map( A1 => n53, A2 => n23, ZN => IMM_13_port);
   U62 : NOR2_X1 port map( A1 => n52, A2 => n23, ZN => IMM_14_port);
   U63 : NOR2_X1 port map( A1 => n51, A2 => n23, ZN => IMM_15_port);
   U64 : INV_X1 port map( A => INST_IN(16), ZN => n32);
   U65 : NAND2_X1 port map( A1 => n9, A2 => n13, ZN => n30);
   U66 : INV_X1 port map( A => n30, ZN => n24);
   U67 : OAI21_X1 port map( B1 => n32, B2 => n28, A => n25, ZN => IMM_16_port);
   U68 : INV_X1 port map( A => INST_IN(17), ZN => n34);
   U69 : OAI21_X1 port map( B1 => n34, B2 => n28, A => n25, ZN => IMM_17_port);
   U70 : INV_X1 port map( A => INST_IN(18), ZN => n35);
   U71 : OAI21_X1 port map( B1 => n35, B2 => n28, A => n25, ZN => IMM_18_port);
   U72 : INV_X1 port map( A => INST_IN(19), ZN => n36);
   U73 : OAI21_X1 port map( B1 => n36, B2 => n28, A => n25, ZN => IMM_19_port);
   U74 : INV_X1 port map( A => INST_IN(20), ZN => n37);
   U75 : OAI21_X1 port map( B1 => n37, B2 => n28, A => n25, ZN => IMM_20_port);
   U76 : INV_X1 port map( A => INST_IN(21), ZN => n38);
   U77 : OAI21_X1 port map( B1 => n38, B2 => n28, A => n25, ZN => IMM_21_port);
   U78 : INV_X1 port map( A => INST_IN(22), ZN => n39);
   U79 : OAI21_X1 port map( B1 => n39, B2 => n28, A => n25, ZN => IMM_22_port);
   U80 : INV_X1 port map( A => INST_IN(23), ZN => n42);
   U81 : OAI21_X1 port map( B1 => n42, B2 => n28, A => n25, ZN => IMM_23_port);
   U82 : INV_X1 port map( A => INST_IN(24), ZN => n43);
   U83 : OAI21_X1 port map( B1 => n43, B2 => n28, A => n25, ZN => IMM_24_port);
   U84 : INV_X1 port map( A => INST_IN(25), ZN => n44);
   U85 : OAI22_X1 port map( A1 => n51, A2 => n30, B1 => n44, B2 => n28, ZN => 
                           IMM_31_port);
   U86 : INV_X1 port map( A => INST_IN(26), ZN => n27);
   U87 : OR4_X1 port map( A1 => n27, A2 => n26, A3 => n33, A4 => n30, ZN => n29
                           );
   U88 : OAI221_X1 port map( B1 => n32, B2 => n30, C1 => n55, C2 => n10, A => 
                           n11, ZN => ADD_WR(0));
   U89 : OAI221_X1 port map( B1 => n34, B2 => n30, C1 => n54, C2 => n10, A => 
                           n11, ZN => ADD_WR(1));
   U90 : OAI221_X1 port map( B1 => n35, B2 => n30, C1 => n53, C2 => n10, A => 
                           n11, ZN => ADD_WR(2));
   U91 : OAI221_X1 port map( B1 => n36, B2 => n30, C1 => n52, C2 => n10, A => 
                           n11, ZN => ADD_WR(3));
   U92 : OAI221_X1 port map( B1 => n37, B2 => n30, C1 => n51, C2 => n10, A => 
                           n11, ZN => ADD_WR(4));
   U93 : NOR3_X1 port map( A1 => n14, A2 => n6, A3 => n37, ZN => ADD_RS2(4));
   U94 : AOI21_X1 port map( B1 => n16, B2 => n13, A => n39, ZN => ADD_RS1(1));
   U95 : NOR2_X1 port map( A1 => n45, A2 => n44, ZN => ADD_RS1(4));
   U96 : INV_X1 port map( A => INST_IN(27), ZN => n50);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity instruction_type is

   port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype : 
         out std_logic);

end instruction_type;

architecture SYN_bhv of instruction_type is

   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => INST_IN(30), Z => n5);
   U2 : CLKBUF_X1 port map( A => n9, Z => n1);
   U3 : BUF_X1 port map( A => INST_IN(26), Z => n9);
   U4 : INV_X1 port map( A => INST_IN(30), ZN => n2);
   U5 : INV_X1 port map( A => INST_IN(30), ZN => n3);
   U6 : CLKBUF_X1 port map( A => INST_IN(27), Z => n4);
   U7 : INV_X1 port map( A => n15, ZN => n6);
   U8 : INV_X1 port map( A => INST_IN(27), ZN => n7);
   U9 : NAND4_X1 port map( A1 => n13, A2 => n11, A3 => n2, A4 => n18, ZN => n8)
                           ;
   U10 : INV_X1 port map( A => INST_IN(31), ZN => n10);
   U11 : INV_X1 port map( A => INST_IN(28), ZN => n13);
   U12 : INV_X1 port map( A => INST_IN(29), ZN => n11);
   U13 : INV_X1 port map( A => INST_IN(30), ZN => n24);
   U14 : INV_X1 port map( A => INST_IN(31), ZN => n18);
   U15 : NAND4_X1 port map( A1 => n13, A2 => n11, A3 => n24, A4 => n18, ZN => 
                           n28);
   U16 : INV_X1 port map( A => INST_IN(27), ZN => n15);
   U17 : NOR2_X1 port map( A1 => n15, A2 => n8, ZN => Jtype);
   U18 : MUX2_X1 port map( A => n2, B => n10, S => INST_IN(29), Z => n12);
   U19 : NAND3_X1 port map( A1 => n15, A2 => INST_IN(28), A3 => n12, ZN => n27)
                           ;
   U20 : OAI211_X1 port map( C1 => n13, C2 => n24, A => INST_IN(29), B => n10, 
                           ZN => n26);
   U21 : NAND3_X1 port map( A1 => n9, A2 => n7, A3 => INST_IN(28), ZN => n14);
   U22 : OAI211_X1 port map( C1 => INST_IN(28), C2 => n15, A => n14, B => 
                           INST_IN(29), ZN => n23);
   U23 : XOR2_X1 port map( A => INST_IN(27), B => INST_IN(26), Z => n16);
   U24 : NOR3_X1 port map( A1 => n16, A2 => INST_IN(28), A3 => n10, ZN => n22);
   U25 : INV_X1 port map( A => INST_IN(26), ZN => n17);
   U26 : NAND3_X1 port map( A1 => INST_IN(28), A2 => n18, A3 => n17, ZN => n20)
                           ;
   U27 : AOI21_X1 port map( B1 => n4, B2 => n18, A => INST_IN(29), ZN => n19);
   U28 : NAND3_X1 port map( A1 => n19, A2 => n20, A3 => n5, ZN => n21);
   U29 : OAI221_X1 port map( B1 => n23, B2 => n3, C1 => n22, C2 => n5, A => n21
                           , ZN => n25);
   U30 : NAND3_X1 port map( A1 => n25, A2 => n26, A3 => n27, ZN => Itype);
   U31 : NOR3_X1 port map( A1 => n28, A2 => n1, A3 => n6, ZN => Rtype);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_0 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_0;

architecture SYN_bhv of regn_N32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DOUT_18_port, DOUT_17_port, DOUT_16_port, DOUT_15_port, DOUT_14_port,
      DOUT_13_port, DOUT_12_port, DOUT_10_port, DOUT_9_port, DOUT_8_port, 
      DOUT_7_port, DOUT_6_port, DOUT_5_port, DOUT_4_port, DOUT_3_port, 
      DOUT_2_port, DOUT_1_port, DOUT_0_port, n1, n2, n3, n4, n5, n6, n7, n8, 
      n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48
      , n49, n50, n51, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, n93, n94, n95, n96, n9, n10, n11, n12, n13, n14, DOUT_11_port
      , n16, n17, n18, n19, n20, n21, n22, DOUT_19_port, DOUT_20_port, 
      DOUT_21_port, DOUT_22_port, DOUT_23_port, DOUT_24_port, DOUT_25_port, 
      DOUT_26_port, DOUT_27_port, DOUT_28_port, DOUT_29_port, DOUT_30_port, 
      DOUT_31_port, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, 
      n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594 : std_logic;

begin
   DOUT <= ( DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, 
      DOUT_27_port, DOUT_26_port, DOUT_25_port, DOUT_24_port, DOUT_23_port, 
      DOUT_22_port, DOUT_21_port, DOUT_20_port, DOUT_19_port, DOUT_18_port, 
      DOUT_17_port, DOUT_16_port, DOUT_15_port, DOUT_14_port, DOUT_13_port, 
      DOUT_12_port, DOUT_11_port, DOUT_10_port, DOUT_9_port, DOUT_8_port, 
      DOUT_7_port, DOUT_6_port, DOUT_5_port, DOUT_4_port, DOUT_3_port, 
      DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n96, CK => CLK, RN => n11, Q => 
                           DOUT_31_port, QN => n_1581);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n95, CK => CLK, RN => n11, Q => 
                           DOUT_30_port, QN => n_1582);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n94, CK => CLK, RN => n11, Q => 
                           DOUT_29_port, QN => n_1583);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n93, CK => CLK, RN => n11, Q => 
                           DOUT_28_port, QN => n_1584);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n92, CK => CLK, RN => n11, Q => 
                           DOUT_27_port, QN => n_1585);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n91, CK => CLK, RN => n11, Q => 
                           DOUT_26_port, QN => n_1586);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n90, CK => CLK, RN => n11, Q => 
                           DOUT_25_port, QN => n_1587);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n89, CK => CLK, RN => n11, Q => 
                           DOUT_24_port, QN => n_1588);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n88, CK => CLK, RN => n10, Q => 
                           DOUT_23_port, QN => n_1589);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n87, CK => CLK, RN => n10, Q => 
                           DOUT_22_port, QN => n_1590);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n86, CK => CLK, RN => n10, Q => 
                           DOUT_21_port, QN => n_1591);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n85, CK => CLK, RN => n10, Q => 
                           DOUT_20_port, QN => n_1592);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n84, CK => CLK, RN => n10, Q => 
                           DOUT_19_port, QN => n_1593);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n83, CK => CLK, RN => n10, Q => 
                           DOUT_18_port, QN => n51);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n82, CK => CLK, RN => n10, Q => 
                           DOUT_17_port, QN => n50);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n81, CK => CLK, RN => n10, Q => 
                           DOUT_16_port, QN => n49);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n80, CK => CLK, RN => n10, Q => 
                           DOUT_15_port, QN => n48);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n79, CK => CLK, RN => n10, Q => 
                           DOUT_14_port, QN => n47);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n78, CK => CLK, RN => n10, Q => 
                           DOUT_13_port, QN => n46);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n77, CK => CLK, RN => n10, Q => 
                           DOUT_12_port, QN => n45);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n76, CK => CLK, RN => n9, Q => 
                           DOUT_11_port, QN => n_1594);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n75, CK => CLK, RN => n9, Q => 
                           DOUT_10_port, QN => n43);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n74, CK => CLK, RN => n9, Q => 
                           DOUT_9_port, QN => n42);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n73, CK => CLK, RN => n9, Q => 
                           DOUT_8_port, QN => n41);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n72, CK => CLK, RN => n9, Q => 
                           DOUT_7_port, QN => n40);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n71, CK => CLK, RN => n9, Q => 
                           DOUT_6_port, QN => n39);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n70, CK => CLK, RN => n9, Q => 
                           DOUT_5_port, QN => n38);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n69, CK => CLK, RN => n9, Q => 
                           DOUT_4_port, QN => n37);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n68, CK => CLK, RN => n9, Q => 
                           DOUT_3_port, QN => n36);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n67, CK => CLK, RN => n9, Q => 
                           DOUT_2_port, QN => n35);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n66, CK => CLK, RN => n9, Q => 
                           DOUT_1_port, QN => n34);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n65, CK => CLK, RN => n9, Q => 
                           DOUT_0_port, QN => n33);
   U2 : BUF_X1 port map( A => RST, Z => n9);
   U3 : BUF_X1 port map( A => RST, Z => n10);
   U4 : BUF_X1 port map( A => RST, Z => n11);
   U5 : OAI21_X1 port map( B1 => n34, B2 => EN, A => n2, ZN => n66);
   U6 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n35, B2 => EN, A => n3, ZN => n67);
   U8 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n3);
   U9 : OAI21_X1 port map( B1 => n36, B2 => EN, A => n4, ZN => n68);
   U10 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n4);
   U11 : OAI21_X1 port map( B1 => n40, B2 => EN, A => n8, ZN => n72);
   U12 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n8);
   U13 : OAI21_X1 port map( B1 => n39, B2 => EN, A => n7, ZN => n71);
   U14 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n38, B2 => EN, A => n6, ZN => n70);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n6);
   U17 : OAI21_X1 port map( B1 => n37, B2 => EN, A => n5, ZN => n69);
   U18 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n5);
   U19 : OAI21_X1 port map( B1 => n33, B2 => EN, A => n1, ZN => n65);
   U20 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n1);
   U21 : INV_X1 port map( A => n41, ZN => n12);
   U22 : MUX2_X1 port map( A => n12, B => DIN(8), S => EN, Z => n73);
   U23 : INV_X1 port map( A => n42, ZN => n13);
   U24 : MUX2_X1 port map( A => n13, B => DIN(9), S => EN, Z => n74);
   U25 : INV_X1 port map( A => n43, ZN => n14);
   U26 : MUX2_X1 port map( A => n14, B => DIN(10), S => EN, Z => n75);
   U27 : MUX2_X1 port map( A => DOUT_11_port, B => DIN(11), S => EN, Z => n76);
   U28 : INV_X1 port map( A => n45, ZN => n16);
   U29 : MUX2_X1 port map( A => n16, B => DIN(12), S => EN, Z => n77);
   U30 : INV_X1 port map( A => n46, ZN => n17);
   U31 : MUX2_X1 port map( A => n17, B => DIN(13), S => EN, Z => n78);
   U32 : INV_X1 port map( A => n47, ZN => n18);
   U33 : MUX2_X1 port map( A => n18, B => DIN(14), S => EN, Z => n79);
   U34 : INV_X1 port map( A => n48, ZN => n19);
   U35 : MUX2_X1 port map( A => n19, B => DIN(15), S => EN, Z => n80);
   U36 : INV_X1 port map( A => n49, ZN => n20);
   U37 : MUX2_X1 port map( A => n20, B => DIN(16), S => EN, Z => n81);
   U38 : INV_X1 port map( A => n50, ZN => n21);
   U39 : MUX2_X1 port map( A => n21, B => DIN(17), S => EN, Z => n82);
   U40 : INV_X1 port map( A => n51, ZN => n22);
   U41 : MUX2_X1 port map( A => n22, B => DIN(18), S => EN, Z => n83);
   U42 : MUX2_X1 port map( A => DOUT_19_port, B => DIN(19), S => EN, Z => n84);
   U43 : MUX2_X1 port map( A => DOUT_20_port, B => DIN(20), S => EN, Z => n85);
   U44 : MUX2_X1 port map( A => DOUT_21_port, B => DIN(21), S => EN, Z => n86);
   U45 : MUX2_X1 port map( A => DOUT_22_port, B => DIN(22), S => EN, Z => n87);
   U46 : MUX2_X1 port map( A => DOUT_23_port, B => DIN(23), S => EN, Z => n88);
   U47 : MUX2_X1 port map( A => DOUT_24_port, B => DIN(24), S => EN, Z => n89);
   U48 : MUX2_X1 port map( A => DOUT_25_port, B => DIN(25), S => EN, Z => n90);
   U49 : MUX2_X1 port map( A => DOUT_26_port, B => DIN(26), S => EN, Z => n91);
   U50 : MUX2_X1 port map( A => DOUT_27_port, B => DIN(27), S => EN, Z => n92);
   U51 : MUX2_X1 port map( A => DOUT_28_port, B => DIN(28), S => EN, Z => n93);
   U52 : MUX2_X1 port map( A => DOUT_29_port, B => DIN(29), S => EN, Z => n94);
   U53 : MUX2_X1 port map( A => DOUT_30_port, B => DIN(30), S => EN, Z => n95);
   U54 : MUX2_X1 port map( A => DOUT_31_port, B => DIN(31), S => EN, Z => n96);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_0;

architecture SYN_bhv of mux21_NBIT32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n43, n54, n65, n1, n2, n3 : std_logic;

begin
   
   U1 : INV_X2 port map( A => n2, ZN => n1);
   U2 : INV_X1 port map( A => n54, ZN => Z(1));
   U3 : AOI22_X1 port map( A1 => A(1), A2 => n2, B1 => B(1), B2 => S, ZN => n54
                           );
   U4 : INV_X1 port map( A => n43, ZN => Z(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => n3, B1 => B(2), B2 => S, ZN => n43
                           );
   U6 : INV_X1 port map( A => n40, ZN => Z(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n2, B1 => B(3), B2 => S, ZN => n40
                           );
   U8 : INV_X1 port map( A => n36, ZN => Z(7));
   U9 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => S, ZN => n36
                           );
   U10 : INV_X1 port map( A => n37, ZN => Z(6));
   U11 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => S, ZN => 
                           n37);
   U12 : INV_X1 port map( A => n38, ZN => Z(5));
   U13 : AOI22_X1 port map( A1 => A(5), A2 => n2, B1 => B(5), B2 => S, ZN => 
                           n38);
   U14 : INV_X1 port map( A => n39, ZN => Z(4));
   U15 : AOI22_X1 port map( A1 => A(4), A2 => n2, B1 => B(4), B2 => S, ZN => 
                           n39);
   U16 : INV_X1 port map( A => n65, ZN => Z(0));
   U17 : AOI22_X1 port map( A1 => A(0), A2 => n3, B1 => B(0), B2 => S, ZN => 
                           n65);
   U18 : INV_X1 port map( A => S, ZN => n2);
   U19 : INV_X1 port map( A => S, ZN => n3);
   U20 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Z(8));
   U21 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Z(9));
   U22 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Z(10));
   U23 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Z(11));
   U24 : MUX2_X1 port map( A => A(12), B => B(12), S => n1, Z => Z(12));
   U25 : MUX2_X1 port map( A => A(13), B => B(13), S => n1, Z => Z(13));
   U26 : MUX2_X1 port map( A => A(14), B => B(14), S => n1, Z => Z(14));
   U27 : MUX2_X1 port map( A => A(15), B => B(15), S => n1, Z => Z(15));
   U28 : MUX2_X1 port map( A => A(16), B => B(16), S => n1, Z => Z(16));
   U29 : MUX2_X1 port map( A => A(17), B => B(17), S => n1, Z => Z(17));
   U30 : MUX2_X1 port map( A => A(18), B => B(18), S => n1, Z => Z(18));
   U31 : MUX2_X1 port map( A => A(19), B => B(19), S => n1, Z => Z(19));
   U32 : MUX2_X1 port map( A => A(20), B => B(20), S => n1, Z => Z(20));
   U33 : MUX2_X1 port map( A => A(21), B => B(21), S => n1, Z => Z(21));
   U34 : MUX2_X1 port map( A => A(22), B => B(22), S => n1, Z => Z(22));
   U35 : MUX2_X1 port map( A => A(23), B => B(23), S => n1, Z => Z(23));
   U36 : MUX2_X1 port map( A => A(24), B => B(24), S => n1, Z => Z(24));
   U37 : MUX2_X1 port map( A => A(25), B => B(25), S => n1, Z => Z(25));
   U38 : MUX2_X1 port map( A => A(26), B => B(26), S => n1, Z => Z(26));
   U39 : MUX2_X1 port map( A => A(27), B => B(27), S => n1, Z => Z(27));
   U40 : MUX2_X1 port map( A => A(28), B => B(28), S => n1, Z => Z(28));
   U41 : MUX2_X1 port map( A => A(29), B => B(29), S => n1, Z => Z(29));
   U42 : MUX2_X1 port map( A => A(30), B => B(30), S => n1, Z => Z(30));
   U43 : MUX2_X1 port map( A => A(31), B => B(31), S => n1, Z => Z(31));

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HazardDetection is

   port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : in std_logic_vector (4
         downto 0);  DRAM_R : in std_logic;  INS_IN, PC_IN : in 
         std_logic_vector (31 downto 0);  Bubble : out std_logic;  HDU_INS_OUT,
         HDU_PC_OUT, HDU_NPC_OUT : out std_logic_vector (31 downto 0));

end HazardDetection;

architecture SYN_arch of HazardDetection is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component HazardDetection_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n7, n8, n11, n1, n2, n3, n4, n5, n6, n9, n10, n12, n13, n14, n15, n16
      , n_1595 : std_logic;

begin
   HDU_INS_OUT <= ( INS_IN(31), INS_IN(30), INS_IN(29), INS_IN(28), INS_IN(27),
      INS_IN(26), INS_IN(25), INS_IN(24), INS_IN(23), INS_IN(22), INS_IN(21), 
      INS_IN(20), INS_IN(19), INS_IN(18), INS_IN(17), INS_IN(16), INS_IN(15), 
      INS_IN(14), INS_IN(13), INS_IN(12), INS_IN(11), INS_IN(10), INS_IN(9), 
      INS_IN(8), INS_IN(7), INS_IN(6), INS_IN(5), INS_IN(4), INS_IN(3), 
      INS_IN(2), INS_IN(1), INS_IN(0) );
   HDU_PC_OUT <= ( PC_IN(31), PC_IN(30), PC_IN(29), PC_IN(28), PC_IN(27), 
      PC_IN(26), PC_IN(25), PC_IN(24), PC_IN(23), PC_IN(22), PC_IN(21), 
      PC_IN(20), PC_IN(19), PC_IN(18), PC_IN(17), PC_IN(16), PC_IN(15), 
      PC_IN(14), PC_IN(13), PC_IN(12), PC_IN(11), PC_IN(10), PC_IN(9), PC_IN(8)
      , PC_IN(7), PC_IN(6), PC_IN(5), PC_IN(4), PC_IN(3), PC_IN(2), PC_IN(1), 
      PC_IN(0) );
   
   n7 <= '0';
   n8 <= '1';
   n11 <= '0';
   add_32 : HazardDetection_DW01_add_0 port map( A(31) => PC_IN(31), A(30) => 
                           PC_IN(30), A(29) => PC_IN(29), A(28) => PC_IN(28), 
                           A(27) => PC_IN(27), A(26) => PC_IN(26), A(25) => 
                           PC_IN(25), A(24) => PC_IN(24), A(23) => PC_IN(23), 
                           A(22) => PC_IN(22), A(21) => PC_IN(21), A(20) => 
                           PC_IN(20), A(19) => PC_IN(19), A(18) => PC_IN(18), 
                           A(17) => PC_IN(17), A(16) => PC_IN(16), A(15) => 
                           PC_IN(15), A(14) => PC_IN(14), A(13) => PC_IN(13), 
                           A(12) => PC_IN(12), A(11) => PC_IN(11), A(10) => 
                           PC_IN(10), A(9) => PC_IN(9), A(8) => PC_IN(8), A(7) 
                           => PC_IN(7), A(6) => PC_IN(6), A(5) => PC_IN(5), 
                           A(4) => PC_IN(4), A(3) => PC_IN(3), A(2) => PC_IN(2)
                           , A(1) => PC_IN(1), A(0) => PC_IN(0), B(31) => n7, 
                           B(30) => n7, B(29) => n7, B(28) => n7, B(27) => n7, 
                           B(26) => n7, B(25) => n7, B(24) => n7, B(23) => n7, 
                           B(22) => n7, B(21) => n7, B(20) => n7, B(19) => n7, 
                           B(18) => n7, B(17) => n7, B(16) => n7, B(15) => n7, 
                           B(14) => n7, B(13) => n7, B(12) => n7, B(11) => n7, 
                           B(10) => n7, B(9) => n7, B(8) => n7, B(7) => n7, 
                           B(6) => n7, B(5) => n7, B(4) => n7, B(3) => n7, B(2)
                           => n8, B(1) => n7, B(0) => n7, CI => n11, SUM(31) =>
                           HDU_NPC_OUT(31), SUM(30) => HDU_NPC_OUT(30), SUM(29)
                           => HDU_NPC_OUT(29), SUM(28) => HDU_NPC_OUT(28), 
                           SUM(27) => HDU_NPC_OUT(27), SUM(26) => 
                           HDU_NPC_OUT(26), SUM(25) => HDU_NPC_OUT(25), SUM(24)
                           => HDU_NPC_OUT(24), SUM(23) => HDU_NPC_OUT(23), 
                           SUM(22) => HDU_NPC_OUT(22), SUM(21) => 
                           HDU_NPC_OUT(21), SUM(20) => HDU_NPC_OUT(20), SUM(19)
                           => HDU_NPC_OUT(19), SUM(18) => HDU_NPC_OUT(18), 
                           SUM(17) => HDU_NPC_OUT(17), SUM(16) => 
                           HDU_NPC_OUT(16), SUM(15) => HDU_NPC_OUT(15), SUM(14)
                           => HDU_NPC_OUT(14), SUM(13) => HDU_NPC_OUT(13), 
                           SUM(12) => HDU_NPC_OUT(12), SUM(11) => 
                           HDU_NPC_OUT(11), SUM(10) => HDU_NPC_OUT(10), SUM(9) 
                           => HDU_NPC_OUT(9), SUM(8) => HDU_NPC_OUT(8), SUM(7) 
                           => HDU_NPC_OUT(7), SUM(6) => HDU_NPC_OUT(6), SUM(5) 
                           => HDU_NPC_OUT(5), SUM(4) => HDU_NPC_OUT(4), SUM(3) 
                           => HDU_NPC_OUT(3), SUM(2) => HDU_NPC_OUT(2), SUM(1) 
                           => HDU_NPC_OUT(1), SUM(0) => HDU_NPC_OUT(0), CO => 
                           n_1595);
   U4 : AND3_X1 port map( A1 => DRAM_R, A2 => n1, A3 => RST, ZN => Bubble);
   U5 : OAI33_X1 port map( A1 => n2, A2 => n3, A3 => n4, B1 => n5, B2 => n6, B3
                           => n9, ZN => n1);
   U6 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RS2(4), Z => n9);
   U8 : XOR2_X1 port map( A => ADD_WR(2), B => ADD_RS2(2), Z => n6);
   U9 : NAND3_X1 port map( A1 => n10, A2 => n12, A3 => n13, ZN => n5);
   U11 : XNOR2_X1 port map( A => ADD_WR(0), B => ADD_RS2(0), ZN => n13);
   U12 : XNOR2_X1 port map( A => ADD_WR(1), B => ADD_RS2(1), ZN => n12);
   U13 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS2(3), ZN => n10);
   U14 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RS1(4), Z => n4);
   U15 : XOR2_X1 port map( A => ADD_WR(2), B => ADD_RS1(2), Z => n3);
   U16 : NAND3_X1 port map( A1 => n14, A2 => n15, A3 => n16, ZN => n2);
   U17 : XNOR2_X1 port map( A => ADD_WR(0), B => ADD_RS1(0), ZN => n16);
   U18 : XNOR2_X1 port map( A => ADD_WR(1), B => ADD_RS1(1), ZN => n15);
   U19 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS1(3), ZN => n14);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Writeback is

   port( WB_MUX_SEL : in std_logic;  DATA_IN, ALU_RES_IN : in std_logic_vector 
         (31 downto 0);  ADD_WR_IN : in std_logic_vector (4 downto 0);  
         DATA_OUT : out std_logic_vector (31 downto 0);  ADD_WR_OUT : out 
         std_logic_vector (4 downto 0));

end Writeback;

architecture SYN_struct of Writeback is

   component mux21_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;

begin
   ADD_WR_OUT <= ( ADD_WR_IN(4), ADD_WR_IN(3), ADD_WR_IN(2), ADD_WR_IN(1), 
      ADD_WR_IN(0) );
   
   WBmux : mux21_NBIT32_3 port map( A(31) => ALU_RES_IN(31), A(30) => 
                           ALU_RES_IN(30), A(29) => ALU_RES_IN(29), A(28) => 
                           ALU_RES_IN(28), A(27) => ALU_RES_IN(27), A(26) => 
                           ALU_RES_IN(26), A(25) => ALU_RES_IN(25), A(24) => 
                           ALU_RES_IN(24), A(23) => ALU_RES_IN(23), A(22) => 
                           ALU_RES_IN(22), A(21) => ALU_RES_IN(21), A(20) => 
                           ALU_RES_IN(20), A(19) => ALU_RES_IN(19), A(18) => 
                           ALU_RES_IN(18), A(17) => ALU_RES_IN(17), A(16) => 
                           ALU_RES_IN(16), A(15) => ALU_RES_IN(15), A(14) => 
                           ALU_RES_IN(14), A(13) => ALU_RES_IN(13), A(12) => 
                           ALU_RES_IN(12), A(11) => ALU_RES_IN(11), A(10) => 
                           ALU_RES_IN(10), A(9) => ALU_RES_IN(9), A(8) => 
                           ALU_RES_IN(8), A(7) => ALU_RES_IN(7), A(6) => 
                           ALU_RES_IN(6), A(5) => ALU_RES_IN(5), A(4) => 
                           ALU_RES_IN(4), A(3) => ALU_RES_IN(3), A(2) => 
                           ALU_RES_IN(2), A(1) => ALU_RES_IN(1), A(0) => 
                           ALU_RES_IN(0), B(31) => DATA_IN(31), B(30) => 
                           DATA_IN(30), B(29) => DATA_IN(29), B(28) => 
                           DATA_IN(28), B(27) => DATA_IN(27), B(26) => 
                           DATA_IN(26), B(25) => DATA_IN(25), B(24) => 
                           DATA_IN(24), B(23) => DATA_IN(23), B(22) => 
                           DATA_IN(22), B(21) => DATA_IN(21), B(20) => 
                           DATA_IN(20), B(19) => DATA_IN(19), B(18) => 
                           DATA_IN(18), B(17) => DATA_IN(17), B(16) => 
                           DATA_IN(16), B(15) => DATA_IN(15), B(14) => 
                           DATA_IN(14), B(13) => DATA_IN(13), B(12) => 
                           DATA_IN(12), B(11) => DATA_IN(11), B(10) => 
                           DATA_IN(10), B(9) => DATA_IN(9), B(8) => DATA_IN(8),
                           B(7) => DATA_IN(7), B(6) => DATA_IN(6), B(5) => 
                           DATA_IN(5), B(4) => DATA_IN(4), B(3) => DATA_IN(3), 
                           B(2) => DATA_IN(2), B(1) => DATA_IN(1), B(0) => 
                           DATA_IN(0), S => WB_MUX_SEL, Z(31) => DATA_OUT(31), 
                           Z(30) => DATA_OUT(30), Z(29) => DATA_OUT(29), Z(28) 
                           => DATA_OUT(28), Z(27) => DATA_OUT(27), Z(26) => 
                           DATA_OUT(26), Z(25) => DATA_OUT(25), Z(24) => 
                           DATA_OUT(24), Z(23) => DATA_OUT(23), Z(22) => 
                           DATA_OUT(22), Z(21) => DATA_OUT(21), Z(20) => 
                           DATA_OUT(20), Z(19) => DATA_OUT(19), Z(18) => 
                           DATA_OUT(18), Z(17) => DATA_OUT(17), Z(16) => 
                           DATA_OUT(16), Z(15) => DATA_OUT(15), Z(14) => 
                           DATA_OUT(14), Z(13) => DATA_OUT(13), Z(12) => 
                           DATA_OUT(12), Z(11) => DATA_OUT(11), Z(10) => 
                           DATA_OUT(10), Z(9) => DATA_OUT(9), Z(8) => 
                           DATA_OUT(8), Z(7) => DATA_OUT(7), Z(6) => 
                           DATA_OUT(6), Z(5) => DATA_OUT(5), Z(4) => 
                           DATA_OUT(4), Z(3) => DATA_OUT(3), Z(2) => 
                           DATA_OUT(2), Z(1) => DATA_OUT(1), Z(0) => 
                           DATA_OUT(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Memory is

   port( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN : in std_logic;  PC_SEL : in
         std_logic_vector (1 downto 0);  NPC_IN, NPC_ABS, NPC_REL, ALU_RES_IN, 
         B_IN : in std_logic_vector (31 downto 0);  ADD_WR_IN : in 
         std_logic_vector (4 downto 0);  DRAM_DATA_IN : in std_logic_vector (31
         downto 0);  LOAD_TYPE_IN : in std_logic_vector (1 downto 0);  
         STORE_TYPE_IN : in std_logic;  PC_OUT : out std_logic_vector (31 
         downto 0);  DRAM_R_OUT, DRAM_W_OUT : out std_logic;  DRAM_ADDR_OUT, 
         DRAM_DATA_OUT, DATA_OUT, ALU_RES_OUT, OP_MEM : out std_logic_vector 
         (31 downto 0);  ADD_WR_MEM, ADD_WR_OUT : out std_logic_vector (4 
         downto 0);  LOAD_TYPE_OUT : out std_logic_vector (1 downto 0);  
         STORE_TYPE_OUT : out std_logic);

end Memory;

architecture SYN_struct of Memory is

   component mux41_NBIT32_2
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component regn_N32_1
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N5_1
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   signal X_Logic0_port : std_logic;

begin
   DRAM_R_OUT <= DRAM_R_IN;
   DRAM_W_OUT <= DRAM_W_IN;
   DRAM_ADDR_OUT <= ( ALU_RES_IN(31), ALU_RES_IN(30), ALU_RES_IN(29), 
      ALU_RES_IN(28), ALU_RES_IN(27), ALU_RES_IN(26), ALU_RES_IN(25), 
      ALU_RES_IN(24), ALU_RES_IN(23), ALU_RES_IN(22), ALU_RES_IN(21), 
      ALU_RES_IN(20), ALU_RES_IN(19), ALU_RES_IN(18), ALU_RES_IN(17), 
      ALU_RES_IN(16), ALU_RES_IN(15), ALU_RES_IN(14), ALU_RES_IN(13), 
      ALU_RES_IN(12), ALU_RES_IN(11), ALU_RES_IN(10), ALU_RES_IN(9), 
      ALU_RES_IN(8), ALU_RES_IN(7), ALU_RES_IN(6), ALU_RES_IN(5), ALU_RES_IN(4)
      , ALU_RES_IN(3), ALU_RES_IN(2), ALU_RES_IN(1), ALU_RES_IN(0) );
   DRAM_DATA_OUT <= ( B_IN(31), B_IN(30), B_IN(29), B_IN(28), B_IN(27), 
      B_IN(26), B_IN(25), B_IN(24), B_IN(23), B_IN(22), B_IN(21), B_IN(20), 
      B_IN(19), B_IN(18), B_IN(17), B_IN(16), B_IN(15), B_IN(14), B_IN(13), 
      B_IN(12), B_IN(11), B_IN(10), B_IN(9), B_IN(8), B_IN(7), B_IN(6), B_IN(5)
      , B_IN(4), B_IN(3), B_IN(2), B_IN(1), B_IN(0) );
   DATA_OUT <= ( DRAM_DATA_IN(31), DRAM_DATA_IN(30), DRAM_DATA_IN(29), 
      DRAM_DATA_IN(28), DRAM_DATA_IN(27), DRAM_DATA_IN(26), DRAM_DATA_IN(25), 
      DRAM_DATA_IN(24), DRAM_DATA_IN(23), DRAM_DATA_IN(22), DRAM_DATA_IN(21), 
      DRAM_DATA_IN(20), DRAM_DATA_IN(19), DRAM_DATA_IN(18), DRAM_DATA_IN(17), 
      DRAM_DATA_IN(16), DRAM_DATA_IN(15), DRAM_DATA_IN(14), DRAM_DATA_IN(13), 
      DRAM_DATA_IN(12), DRAM_DATA_IN(11), DRAM_DATA_IN(10), DRAM_DATA_IN(9), 
      DRAM_DATA_IN(8), DRAM_DATA_IN(7), DRAM_DATA_IN(6), DRAM_DATA_IN(5), 
      DRAM_DATA_IN(4), DRAM_DATA_IN(3), DRAM_DATA_IN(2), DRAM_DATA_IN(1), 
      DRAM_DATA_IN(0) );
   OP_MEM <= ( ALU_RES_IN(31), ALU_RES_IN(30), ALU_RES_IN(29), ALU_RES_IN(28), 
      ALU_RES_IN(27), ALU_RES_IN(26), ALU_RES_IN(25), ALU_RES_IN(24), 
      ALU_RES_IN(23), ALU_RES_IN(22), ALU_RES_IN(21), ALU_RES_IN(20), 
      ALU_RES_IN(19), ALU_RES_IN(18), ALU_RES_IN(17), ALU_RES_IN(16), 
      ALU_RES_IN(15), ALU_RES_IN(14), ALU_RES_IN(13), ALU_RES_IN(12), 
      ALU_RES_IN(11), ALU_RES_IN(10), ALU_RES_IN(9), ALU_RES_IN(8), 
      ALU_RES_IN(7), ALU_RES_IN(6), ALU_RES_IN(5), ALU_RES_IN(4), ALU_RES_IN(3)
      , ALU_RES_IN(2), ALU_RES_IN(1), ALU_RES_IN(0) );
   ADD_WR_MEM <= ( ADD_WR_IN(4), ADD_WR_IN(3), ADD_WR_IN(2), ADD_WR_IN(1), 
      ADD_WR_IN(0) );
   LOAD_TYPE_OUT <= ( LOAD_TYPE_IN(1), LOAD_TYPE_IN(0) );
   STORE_TYPE_OUT <= STORE_TYPE_IN;
   
   X_Logic0_port <= '0';
   reg0 : regn_N5_1 port map( DIN(4) => ADD_WR_IN(4), DIN(3) => ADD_WR_IN(3), 
                           DIN(2) => ADD_WR_IN(2), DIN(1) => ADD_WR_IN(1), 
                           DIN(0) => ADD_WR_IN(0), CLK => CLK, EN => MEM_EN_IN,
                           RST => RST, DOUT(4) => ADD_WR_OUT(4), DOUT(3) => 
                           ADD_WR_OUT(3), DOUT(2) => ADD_WR_OUT(2), DOUT(1) => 
                           ADD_WR_OUT(1), DOUT(0) => ADD_WR_OUT(0));
   reg1 : regn_N32_1 port map( DIN(31) => ALU_RES_IN(31), DIN(30) => 
                           ALU_RES_IN(30), DIN(29) => ALU_RES_IN(29), DIN(28) 
                           => ALU_RES_IN(28), DIN(27) => ALU_RES_IN(27), 
                           DIN(26) => ALU_RES_IN(26), DIN(25) => ALU_RES_IN(25)
                           , DIN(24) => ALU_RES_IN(24), DIN(23) => 
                           ALU_RES_IN(23), DIN(22) => ALU_RES_IN(22), DIN(21) 
                           => ALU_RES_IN(21), DIN(20) => ALU_RES_IN(20), 
                           DIN(19) => ALU_RES_IN(19), DIN(18) => ALU_RES_IN(18)
                           , DIN(17) => ALU_RES_IN(17), DIN(16) => 
                           ALU_RES_IN(16), DIN(15) => ALU_RES_IN(15), DIN(14) 
                           => ALU_RES_IN(14), DIN(13) => ALU_RES_IN(13), 
                           DIN(12) => ALU_RES_IN(12), DIN(11) => ALU_RES_IN(11)
                           , DIN(10) => ALU_RES_IN(10), DIN(9) => ALU_RES_IN(9)
                           , DIN(8) => ALU_RES_IN(8), DIN(7) => ALU_RES_IN(7), 
                           DIN(6) => ALU_RES_IN(6), DIN(5) => ALU_RES_IN(5), 
                           DIN(4) => ALU_RES_IN(4), DIN(3) => ALU_RES_IN(3), 
                           DIN(2) => ALU_RES_IN(2), DIN(1) => ALU_RES_IN(1), 
                           DIN(0) => ALU_RES_IN(0), CLK => CLK, EN => MEM_EN_IN
                           , RST => RST, DOUT(31) => ALU_RES_OUT(31), DOUT(30) 
                           => ALU_RES_OUT(30), DOUT(29) => ALU_RES_OUT(29), 
                           DOUT(28) => ALU_RES_OUT(28), DOUT(27) => 
                           ALU_RES_OUT(27), DOUT(26) => ALU_RES_OUT(26), 
                           DOUT(25) => ALU_RES_OUT(25), DOUT(24) => 
                           ALU_RES_OUT(24), DOUT(23) => ALU_RES_OUT(23), 
                           DOUT(22) => ALU_RES_OUT(22), DOUT(21) => 
                           ALU_RES_OUT(21), DOUT(20) => ALU_RES_OUT(20), 
                           DOUT(19) => ALU_RES_OUT(19), DOUT(18) => 
                           ALU_RES_OUT(18), DOUT(17) => ALU_RES_OUT(17), 
                           DOUT(16) => ALU_RES_OUT(16), DOUT(15) => 
                           ALU_RES_OUT(15), DOUT(14) => ALU_RES_OUT(14), 
                           DOUT(13) => ALU_RES_OUT(13), DOUT(12) => 
                           ALU_RES_OUT(12), DOUT(11) => ALU_RES_OUT(11), 
                           DOUT(10) => ALU_RES_OUT(10), DOUT(9) => 
                           ALU_RES_OUT(9), DOUT(8) => ALU_RES_OUT(8), DOUT(7) 
                           => ALU_RES_OUT(7), DOUT(6) => ALU_RES_OUT(6), 
                           DOUT(5) => ALU_RES_OUT(5), DOUT(4) => ALU_RES_OUT(4)
                           , DOUT(3) => ALU_RES_OUT(3), DOUT(2) => 
                           ALU_RES_OUT(2), DOUT(1) => ALU_RES_OUT(1), DOUT(0) 
                           => ALU_RES_OUT(0));
   PCsel : mux41_NBIT32_2 port map( A(31) => NPC_IN(31), A(30) => NPC_IN(30), 
                           A(29) => NPC_IN(29), A(28) => NPC_IN(28), A(27) => 
                           NPC_IN(27), A(26) => NPC_IN(26), A(25) => NPC_IN(25)
                           , A(24) => NPC_IN(24), A(23) => NPC_IN(23), A(22) =>
                           NPC_IN(22), A(21) => NPC_IN(21), A(20) => NPC_IN(20)
                           , A(19) => NPC_IN(19), A(18) => NPC_IN(18), A(17) =>
                           NPC_IN(17), A(16) => NPC_IN(16), A(15) => NPC_IN(15)
                           , A(14) => NPC_IN(14), A(13) => NPC_IN(13), A(12) =>
                           NPC_IN(12), A(11) => NPC_IN(11), A(10) => NPC_IN(10)
                           , A(9) => NPC_IN(9), A(8) => NPC_IN(8), A(7) => 
                           NPC_IN(7), A(6) => NPC_IN(6), A(5) => NPC_IN(5), 
                           A(4) => NPC_IN(4), A(3) => NPC_IN(3), A(2) => 
                           NPC_IN(2), A(1) => NPC_IN(1), A(0) => NPC_IN(0), 
                           B(31) => NPC_REL(31), B(30) => NPC_REL(30), B(29) =>
                           NPC_REL(29), B(28) => NPC_REL(28), B(27) => 
                           NPC_REL(27), B(26) => NPC_REL(26), B(25) => 
                           NPC_REL(25), B(24) => NPC_REL(24), B(23) => 
                           NPC_REL(23), B(22) => NPC_REL(22), B(21) => 
                           NPC_REL(21), B(20) => NPC_REL(20), B(19) => 
                           NPC_REL(19), B(18) => NPC_REL(18), B(17) => 
                           NPC_REL(17), B(16) => NPC_REL(16), B(15) => 
                           NPC_REL(15), B(14) => NPC_REL(14), B(13) => 
                           NPC_REL(13), B(12) => NPC_REL(12), B(11) => 
                           NPC_REL(11), B(10) => NPC_REL(10), B(9) => 
                           NPC_REL(9), B(8) => NPC_REL(8), B(7) => NPC_REL(7), 
                           B(6) => NPC_REL(6), B(5) => NPC_REL(5), B(4) => 
                           NPC_REL(4), B(3) => NPC_REL(3), B(2) => NPC_REL(2), 
                           B(1) => NPC_REL(1), B(0) => NPC_REL(0), C(31) => 
                           NPC_ABS(31), C(30) => NPC_ABS(30), C(29) => 
                           NPC_ABS(29), C(28) => NPC_ABS(28), C(27) => 
                           NPC_ABS(27), C(26) => NPC_ABS(26), C(25) => 
                           NPC_ABS(25), C(24) => NPC_ABS(24), C(23) => 
                           NPC_ABS(23), C(22) => NPC_ABS(22), C(21) => 
                           NPC_ABS(21), C(20) => NPC_ABS(20), C(19) => 
                           NPC_ABS(19), C(18) => NPC_ABS(18), C(17) => 
                           NPC_ABS(17), C(16) => NPC_ABS(16), C(15) => 
                           NPC_ABS(15), C(14) => NPC_ABS(14), C(13) => 
                           NPC_ABS(13), C(12) => NPC_ABS(12), C(11) => 
                           NPC_ABS(11), C(10) => NPC_ABS(10), C(9) => 
                           NPC_ABS(9), C(8) => NPC_ABS(8), C(7) => NPC_ABS(7), 
                           C(6) => NPC_ABS(6), C(5) => NPC_ABS(5), C(4) => 
                           NPC_ABS(4), C(3) => NPC_ABS(3), C(2) => NPC_ABS(2), 
                           C(1) => NPC_ABS(1), C(0) => NPC_ABS(0), D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => X_Logic0_port, D(25) => 
                           X_Logic0_port, D(24) => X_Logic0_port, D(23) => 
                           X_Logic0_port, D(22) => X_Logic0_port, D(21) => 
                           X_Logic0_port, D(20) => X_Logic0_port, D(19) => 
                           X_Logic0_port, D(18) => X_Logic0_port, D(17) => 
                           X_Logic0_port, D(16) => X_Logic0_port, D(15) => 
                           X_Logic0_port, D(14) => X_Logic0_port, D(13) => 
                           X_Logic0_port, D(12) => X_Logic0_port, D(11) => 
                           X_Logic0_port, D(10) => X_Logic0_port, D(9) => 
                           X_Logic0_port, D(8) => X_Logic0_port, D(7) => 
                           X_Logic0_port, D(6) => X_Logic0_port, D(5) => 
                           X_Logic0_port, D(4) => X_Logic0_port, D(3) => 
                           X_Logic0_port, D(2) => X_Logic0_port, D(1) => 
                           X_Logic0_port, D(0) => X_Logic0_port, S(1) => 
                           PC_SEL(1), S(0) => PC_SEL(0), Z(31) => PC_OUT(31), 
                           Z(30) => PC_OUT(30), Z(29) => PC_OUT(29), Z(28) => 
                           PC_OUT(28), Z(27) => PC_OUT(27), Z(26) => PC_OUT(26)
                           , Z(25) => PC_OUT(25), Z(24) => PC_OUT(24), Z(23) =>
                           PC_OUT(23), Z(22) => PC_OUT(22), Z(21) => PC_OUT(21)
                           , Z(20) => PC_OUT(20), Z(19) => PC_OUT(19), Z(18) =>
                           PC_OUT(18), Z(17) => PC_OUT(17), Z(16) => PC_OUT(16)
                           , Z(15) => PC_OUT(15), Z(14) => PC_OUT(14), Z(13) =>
                           PC_OUT(13), Z(12) => PC_OUT(12), Z(11) => PC_OUT(11)
                           , Z(10) => PC_OUT(10), Z(9) => PC_OUT(9), Z(8) => 
                           PC_OUT(8), Z(7) => PC_OUT(7), Z(6) => PC_OUT(6), 
                           Z(5) => PC_OUT(5), Z(4) => PC_OUT(4), Z(3) => 
                           PC_OUT(3), Z(2) => PC_OUT(2), Z(1) => PC_OUT(1), 
                           Z(0) => PC_OUT(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ff_0 is

   port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);

end ff_0;

architecture SYN_bhv of ff_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n3, CK => CLK, RN => RST, Q => Q, QN => n2);
   U2 : OAI21_X1 port map( B1 => n2, B2 => EN, A => n1, ZN => n3);
   U3 : NAND2_X1 port map( A1 => EN, A2 => D, ZN => n1);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute is

   port( CLK, RST, MUX_A_SEL : in std_logic;  MUX_B_SEL : in std_logic_vector 
         (1 downto 0);  ALU_OPC : in std_logic_vector (0 to 4);  ALU_OUTREG_EN 
         : in std_logic;  JUMP_TYPE : in std_logic_vector (1 downto 0);  PC_IN,
         A_IN, B_IN, IMM_IN : in std_logic_vector (31 downto 0);  ADD_WR_IN, 
         ADD_RS1_IN, ADD_RS2_IN, ADD_WR_MEM, ADD_WR_WB : in std_logic_vector (4
         downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;  OP_MEM, OP_WB : in 
         std_logic_vector (31 downto 0);  PC_SEL : out std_logic_vector (1 
         downto 0);  ZERO_FLAG : out std_logic;  NPC_ABS, NPC_REL, ALU_RES, 
         B_OUT : out std_logic_vector (31 downto 0);  ADD_WR_OUT : out 
         std_logic_vector (4 downto 0));

end Execute;

architecture SYN_struct of Execute is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component Execute_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component Execute_DW01_add_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component regn_N32_2
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_3
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N5_2
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N32_4
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_5
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component ALU_NBIT32
      port( OP1, OP2 : in std_logic_vector (31 downto 0);  ALU_OPC : in 
            std_logic_vector (0 to 4);  ALU_RES : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux41_NBIT32_3
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux21_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux41_NBIT32_4
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux41_NBIT32_0
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component FWD_Unit
      port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB : in 
            std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;
            FWDA, FWDB : out std_logic_vector (1 downto 0));
   end component;
   
   component regn_N2
      port( DIN : in std_logic_vector (1 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (1 downto 0));
   end component;
   
   component ff_1
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Branch_Cond_Unit_NBIT32
      port( RST : in std_logic;  A : in std_logic_vector (31 downto 0);  
            ALU_OPC : in std_logic_vector (0 to 4);  JUMP_TYPE : in 
            std_logic_vector (1 downto 0);  PC_SEL : out std_logic_vector (1 
            downto 0);  ZERO : out std_logic);
   end component;
   
   signal ZERO_FLAG_port, sig_RST, sig_NPC_ABS_31_port, sig_NPC_ABS_30_port, 
      sig_NPC_ABS_29_port, sig_NPC_ABS_28_port, sig_NPC_ABS_27_port, 
      sig_NPC_ABS_26_port, sig_NPC_ABS_25_port, sig_NPC_ABS_24_port, 
      sig_NPC_ABS_23_port, sig_NPC_ABS_22_port, sig_NPC_ABS_21_port, 
      sig_NPC_ABS_20_port, sig_NPC_ABS_19_port, sig_NPC_ABS_18_port, 
      sig_NPC_ABS_17_port, sig_NPC_ABS_16_port, sig_NPC_ABS_15_port, 
      sig_NPC_ABS_14_port, sig_NPC_ABS_13_port, sig_NPC_ABS_12_port, 
      sig_NPC_ABS_11_port, sig_NPC_ABS_10_port, sig_NPC_ABS_9_port, 
      sig_NPC_ABS_8_port, sig_NPC_ABS_7_port, sig_NPC_ABS_6_port, 
      sig_NPC_ABS_5_port, sig_NPC_ABS_4_port, sig_NPC_ABS_3_port, 
      sig_NPC_ABS_2_port, sig_NPC_ABS_1_port, sig_NPC_ABS_0_port, 
      sig_NPC_REL_31_port, sig_NPC_REL_30_port, sig_NPC_REL_29_port, 
      sig_NPC_REL_28_port, sig_NPC_REL_27_port, sig_NPC_REL_26_port, 
      sig_NPC_REL_25_port, sig_NPC_REL_24_port, sig_NPC_REL_23_port, 
      sig_NPC_REL_22_port, sig_NPC_REL_21_port, sig_NPC_REL_20_port, 
      sig_NPC_REL_19_port, sig_NPC_REL_18_port, sig_NPC_REL_17_port, 
      sig_NPC_REL_16_port, sig_NPC_REL_15_port, sig_NPC_REL_14_port, 
      sig_NPC_REL_13_port, sig_NPC_REL_12_port, sig_NPC_REL_11_port, 
      sig_NPC_REL_10_port, sig_NPC_REL_9_port, sig_NPC_REL_8_port, 
      sig_NPC_REL_7_port, sig_NPC_REL_6_port, sig_NPC_REL_5_port, 
      sig_NPC_REL_4_port, sig_NPC_REL_3_port, sig_NPC_REL_2_port, 
      sig_NPC_REL_1_port, sig_NPC_REL_0_port, sig_PC_SEL_1_port, 
      sig_PC_SEL_0_port, sig_ZERO_FLAG, FWDA_1_port, FWDA_0_port, FWDB_1_port, 
      FWDB_0_port, OP2_FW_31_port, OP2_FW_30_port, OP2_FW_29_port, 
      OP2_FW_28_port, OP2_FW_27_port, OP2_FW_26_port, OP2_FW_25_port, 
      OP2_FW_24_port, OP2_FW_23_port, OP2_FW_22_port, OP2_FW_21_port, 
      OP2_FW_20_port, OP2_FW_19_port, OP2_FW_18_port, OP2_FW_17_port, 
      OP2_FW_16_port, OP2_FW_15_port, OP2_FW_14_port, OP2_FW_13_port, 
      OP2_FW_12_port, OP2_FW_11_port, OP2_FW_10_port, OP2_FW_9_port, 
      OP2_FW_8_port, OP2_FW_7_port, OP2_FW_6_port, OP2_FW_5_port, OP2_FW_4_port
      , OP2_FW_3_port, OP2_FW_2_port, OP2_FW_1_port, OP2_FW_0_port, 
      sig_OP1_31_port, sig_OP1_30_port, sig_OP1_29_port, sig_OP1_28_port, 
      sig_OP1_27_port, sig_OP1_26_port, sig_OP1_25_port, sig_OP1_24_port, 
      sig_OP1_23_port, sig_OP1_22_port, sig_OP1_21_port, sig_OP1_20_port, 
      sig_OP1_19_port, sig_OP1_18_port, sig_OP1_17_port, sig_OP1_16_port, 
      sig_OP1_15_port, sig_OP1_14_port, sig_OP1_13_port, sig_OP1_12_port, 
      sig_OP1_11_port, sig_OP1_10_port, sig_OP1_9_port, sig_OP1_8_port, 
      sig_OP1_7_port, sig_OP1_6_port, sig_OP1_5_port, sig_OP1_4_port, 
      sig_OP1_3_port, sig_OP1_2_port, sig_OP1_1_port, sig_OP1_0_port, 
      sig_OP2_31_port, sig_OP2_30_port, sig_OP2_29_port, sig_OP2_28_port, 
      sig_OP2_27_port, sig_OP2_26_port, sig_OP2_25_port, sig_OP2_24_port, 
      sig_OP2_23_port, sig_OP2_22_port, sig_OP2_21_port, sig_OP2_20_port, 
      sig_OP2_19_port, sig_OP2_18_port, sig_OP2_17_port, sig_OP2_16_port, 
      sig_OP2_15_port, sig_OP2_14_port, sig_OP2_13_port, sig_OP2_12_port, 
      sig_OP2_11_port, sig_OP2_10_port, sig_OP2_9_port, sig_OP2_8_port, 
      sig_OP2_7_port, sig_OP2_6_port, sig_OP2_5_port, sig_OP2_4_port, 
      sig_OP2_3_port, sig_OP2_2_port, sig_OP2_1_port, sig_OP2_0_port, 
      sig_ALU_RES_31_port, sig_ALU_RES_30_port, sig_ALU_RES_29_port, 
      sig_ALU_RES_28_port, sig_ALU_RES_27_port, sig_ALU_RES_26_port, 
      sig_ALU_RES_25_port, sig_ALU_RES_24_port, sig_ALU_RES_23_port, 
      sig_ALU_RES_22_port, sig_ALU_RES_21_port, sig_ALU_RES_20_port, 
      sig_ALU_RES_19_port, sig_ALU_RES_18_port, sig_ALU_RES_17_port, 
      sig_ALU_RES_16_port, sig_ALU_RES_15_port, sig_ALU_RES_14_port, 
      sig_ALU_RES_13_port, sig_ALU_RES_12_port, sig_ALU_RES_11_port, 
      sig_ALU_RES_10_port, sig_ALU_RES_9_port, sig_ALU_RES_8_port, 
      sig_ALU_RES_7_port, sig_ALU_RES_6_port, sig_ALU_RES_5_port, 
      sig_ALU_RES_4_port, sig_ALU_RES_3_port, sig_ALU_RES_2_port, 
      sig_ALU_RES_1_port, sig_ALU_RES_0_port, N9, N8, N7, N6, N5, N4, N31, N30,
      N3, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N2, N19, N18, N17, 
      N16, N15, N14, N13, N12, N11, N10, N1, N0, n1_port, n2_port, n3_port, 
      n4_port, n5_port, n6_port, n7_port, n_1596, n_1597 : std_logic;

begin
   ZERO_FLAG <= ZERO_FLAG_port;
   
   n7_port <= '1';
   n6_port <= '0';
   Branch_Cond : Branch_Cond_Unit_NBIT32 port map( RST => sig_RST, A(31) => 
                           sig_NPC_ABS_31_port, A(30) => sig_NPC_ABS_30_port, 
                           A(29) => sig_NPC_ABS_29_port, A(28) => 
                           sig_NPC_ABS_28_port, A(27) => sig_NPC_ABS_27_port, 
                           A(26) => sig_NPC_ABS_26_port, A(25) => 
                           sig_NPC_ABS_25_port, A(24) => sig_NPC_ABS_24_port, 
                           A(23) => sig_NPC_ABS_23_port, A(22) => 
                           sig_NPC_ABS_22_port, A(21) => sig_NPC_ABS_21_port, 
                           A(20) => sig_NPC_ABS_20_port, A(19) => 
                           sig_NPC_ABS_19_port, A(18) => sig_NPC_ABS_18_port, 
                           A(17) => sig_NPC_ABS_17_port, A(16) => 
                           sig_NPC_ABS_16_port, A(15) => sig_NPC_ABS_15_port, 
                           A(14) => sig_NPC_ABS_14_port, A(13) => 
                           sig_NPC_ABS_13_port, A(12) => sig_NPC_ABS_12_port, 
                           A(11) => sig_NPC_ABS_11_port, A(10) => 
                           sig_NPC_ABS_10_port, A(9) => sig_NPC_ABS_9_port, 
                           A(8) => sig_NPC_ABS_8_port, A(7) => 
                           sig_NPC_ABS_7_port, A(6) => sig_NPC_ABS_6_port, A(5)
                           => sig_NPC_ABS_5_port, A(4) => sig_NPC_ABS_4_port, 
                           A(3) => sig_NPC_ABS_3_port, A(2) => 
                           sig_NPC_ABS_2_port, A(1) => sig_NPC_ABS_1_port, A(0)
                           => sig_NPC_ABS_0_port, ALU_OPC(0) => ALU_OPC(0), 
                           ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => ALU_OPC(2), 
                           ALU_OPC(3) => ALU_OPC(3), ALU_OPC(4) => ALU_OPC(4), 
                           JUMP_TYPE(1) => JUMP_TYPE(1), JUMP_TYPE(0) => 
                           JUMP_TYPE(0), PC_SEL(1) => sig_PC_SEL_1_port, 
                           PC_SEL(0) => sig_PC_SEL_0_port, ZERO => 
                           sig_ZERO_FLAG);
   ff0 : ff_1 port map( D => sig_ZERO_FLAG, CLK => CLK, EN => n7_port, RST => 
                           RST, Q => ZERO_FLAG_port);
   reg0 : regn_N2 port map( DIN(1) => sig_PC_SEL_1_port, DIN(0) => 
                           sig_PC_SEL_0_port, CLK => CLK, EN => n7_port, RST =>
                           RST, DOUT(1) => PC_SEL(1), DOUT(0) => PC_SEL(0));
   FWD : FWD_Unit port map( RST => sig_RST, ADD_RS1(4) => ADD_RS1_IN(4), 
                           ADD_RS1(3) => ADD_RS1_IN(3), ADD_RS1(2) => 
                           ADD_RS1_IN(2), ADD_RS1(1) => ADD_RS1_IN(1), 
                           ADD_RS1(0) => ADD_RS1_IN(0), ADD_RS2(4) => 
                           ADD_RS2_IN(4), ADD_RS2(3) => ADD_RS2_IN(3), 
                           ADD_RS2(2) => ADD_RS2_IN(2), ADD_RS2(1) => 
                           ADD_RS2_IN(1), ADD_RS2(0) => ADD_RS2_IN(0), 
                           ADD_WR_MEM(4) => ADD_WR_MEM(4), ADD_WR_MEM(3) => 
                           ADD_WR_MEM(3), ADD_WR_MEM(2) => ADD_WR_MEM(2), 
                           ADD_WR_MEM(1) => ADD_WR_MEM(1), ADD_WR_MEM(0) => 
                           ADD_WR_MEM(0), ADD_WR_WB(4) => ADD_WR_WB(4), 
                           ADD_WR_WB(3) => ADD_WR_WB(3), ADD_WR_WB(2) => 
                           ADD_WR_WB(2), ADD_WR_WB(1) => ADD_WR_WB(1), 
                           ADD_WR_WB(0) => ADD_WR_WB(0), RF_WE_MEM => RF_WE_MEM
                           , RF_WE_WB => RF_WE_WB, FWDA(1) => FWDA_1_port, 
                           FWDA(0) => FWDA_0_port, FWDB(1) => FWDB_1_port, 
                           FWDB(0) => FWDB_0_port);
   FW1 : mux41_NBIT32_0 port map( A(31) => A_IN(31), A(30) => A_IN(30), A(29) 
                           => A_IN(29), A(28) => A_IN(28), A(27) => A_IN(27), 
                           A(26) => A_IN(26), A(25) => A_IN(25), A(24) => 
                           A_IN(24), A(23) => A_IN(23), A(22) => A_IN(22), 
                           A(21) => A_IN(21), A(20) => A_IN(20), A(19) => 
                           A_IN(19), A(18) => A_IN(18), A(17) => A_IN(17), 
                           A(16) => A_IN(16), A(15) => A_IN(15), A(14) => 
                           A_IN(14), A(13) => A_IN(13), A(12) => A_IN(12), 
                           A(11) => A_IN(11), A(10) => A_IN(10), A(9) => 
                           A_IN(9), A(8) => A_IN(8), A(7) => A_IN(7), A(6) => 
                           A_IN(6), A(5) => A_IN(5), A(4) => A_IN(4), A(3) => 
                           A_IN(3), A(2) => A_IN(2), A(1) => A_IN(1), A(0) => 
                           A_IN(0), B(31) => OP_WB(31), B(30) => OP_WB(30), 
                           B(29) => OP_WB(29), B(28) => OP_WB(28), B(27) => 
                           OP_WB(27), B(26) => OP_WB(26), B(25) => OP_WB(25), 
                           B(24) => OP_WB(24), B(23) => OP_WB(23), B(22) => 
                           OP_WB(22), B(21) => OP_WB(21), B(20) => OP_WB(20), 
                           B(19) => OP_WB(19), B(18) => OP_WB(18), B(17) => 
                           OP_WB(17), B(16) => OP_WB(16), B(15) => OP_WB(15), 
                           B(14) => OP_WB(14), B(13) => OP_WB(13), B(12) => 
                           OP_WB(12), B(11) => OP_WB(11), B(10) => OP_WB(10), 
                           B(9) => OP_WB(9), B(8) => OP_WB(8), B(7) => OP_WB(7)
                           , B(6) => OP_WB(6), B(5) => OP_WB(5), B(4) => 
                           OP_WB(4), B(3) => OP_WB(3), B(2) => OP_WB(2), B(1) 
                           => OP_WB(1), B(0) => OP_WB(0), C(31) => OP_MEM(31), 
                           C(30) => OP_MEM(30), C(29) => OP_MEM(29), C(28) => 
                           OP_MEM(28), C(27) => OP_MEM(27), C(26) => OP_MEM(26)
                           , C(25) => OP_MEM(25), C(24) => OP_MEM(24), C(23) =>
                           OP_MEM(23), C(22) => OP_MEM(22), C(21) => OP_MEM(21)
                           , C(20) => OP_MEM(20), C(19) => OP_MEM(19), C(18) =>
                           OP_MEM(18), C(17) => OP_MEM(17), C(16) => OP_MEM(16)
                           , C(15) => OP_MEM(15), C(14) => OP_MEM(14), C(13) =>
                           OP_MEM(13), C(12) => OP_MEM(12), C(11) => OP_MEM(11)
                           , C(10) => OP_MEM(10), C(9) => OP_MEM(9), C(8) => 
                           OP_MEM(8), C(7) => OP_MEM(7), C(6) => OP_MEM(6), 
                           C(5) => OP_MEM(5), C(4) => OP_MEM(4), C(3) => 
                           OP_MEM(3), C(2) => OP_MEM(2), C(1) => OP_MEM(1), 
                           C(0) => OP_MEM(0), D(31) => A_IN(31), D(30) => 
                           A_IN(30), D(29) => A_IN(29), D(28) => A_IN(28), 
                           D(27) => A_IN(27), D(26) => A_IN(26), D(25) => 
                           A_IN(25), D(24) => A_IN(24), D(23) => A_IN(23), 
                           D(22) => A_IN(22), D(21) => A_IN(21), D(20) => 
                           A_IN(20), D(19) => A_IN(19), D(18) => A_IN(18), 
                           D(17) => A_IN(17), D(16) => A_IN(16), D(15) => 
                           A_IN(15), D(14) => A_IN(14), D(13) => A_IN(13), 
                           D(12) => A_IN(12), D(11) => A_IN(11), D(10) => 
                           A_IN(10), D(9) => A_IN(9), D(8) => A_IN(8), D(7) => 
                           A_IN(7), D(6) => A_IN(6), D(5) => A_IN(5), D(4) => 
                           A_IN(4), D(3) => A_IN(3), D(2) => A_IN(2), D(1) => 
                           A_IN(1), D(0) => A_IN(0), S(1) => FWDA_1_port, S(0) 
                           => FWDA_0_port, Z(31) => sig_NPC_ABS_31_port, Z(30) 
                           => sig_NPC_ABS_30_port, Z(29) => sig_NPC_ABS_29_port
                           , Z(28) => sig_NPC_ABS_28_port, Z(27) => 
                           sig_NPC_ABS_27_port, Z(26) => sig_NPC_ABS_26_port, 
                           Z(25) => sig_NPC_ABS_25_port, Z(24) => 
                           sig_NPC_ABS_24_port, Z(23) => sig_NPC_ABS_23_port, 
                           Z(22) => sig_NPC_ABS_22_port, Z(21) => 
                           sig_NPC_ABS_21_port, Z(20) => sig_NPC_ABS_20_port, 
                           Z(19) => sig_NPC_ABS_19_port, Z(18) => 
                           sig_NPC_ABS_18_port, Z(17) => sig_NPC_ABS_17_port, 
                           Z(16) => sig_NPC_ABS_16_port, Z(15) => 
                           sig_NPC_ABS_15_port, Z(14) => sig_NPC_ABS_14_port, 
                           Z(13) => sig_NPC_ABS_13_port, Z(12) => 
                           sig_NPC_ABS_12_port, Z(11) => sig_NPC_ABS_11_port, 
                           Z(10) => sig_NPC_ABS_10_port, Z(9) => 
                           sig_NPC_ABS_9_port, Z(8) => sig_NPC_ABS_8_port, Z(7)
                           => sig_NPC_ABS_7_port, Z(6) => sig_NPC_ABS_6_port, 
                           Z(5) => sig_NPC_ABS_5_port, Z(4) => 
                           sig_NPC_ABS_4_port, Z(3) => sig_NPC_ABS_3_port, Z(2)
                           => sig_NPC_ABS_2_port, Z(1) => sig_NPC_ABS_1_port, 
                           Z(0) => sig_NPC_ABS_0_port);
   FW2 : mux41_NBIT32_4 port map( A(31) => B_IN(31), A(30) => B_IN(30), A(29) 
                           => B_IN(29), A(28) => B_IN(28), A(27) => B_IN(27), 
                           A(26) => B_IN(26), A(25) => B_IN(25), A(24) => 
                           B_IN(24), A(23) => B_IN(23), A(22) => B_IN(22), 
                           A(21) => B_IN(21), A(20) => B_IN(20), A(19) => 
                           B_IN(19), A(18) => B_IN(18), A(17) => B_IN(17), 
                           A(16) => B_IN(16), A(15) => B_IN(15), A(14) => 
                           B_IN(14), A(13) => B_IN(13), A(12) => B_IN(12), 
                           A(11) => B_IN(11), A(10) => B_IN(10), A(9) => 
                           B_IN(9), A(8) => B_IN(8), A(7) => B_IN(7), A(6) => 
                           B_IN(6), A(5) => B_IN(5), A(4) => B_IN(4), A(3) => 
                           B_IN(3), A(2) => B_IN(2), A(1) => B_IN(1), A(0) => 
                           B_IN(0), B(31) => OP_WB(31), B(30) => OP_WB(30), 
                           B(29) => OP_WB(29), B(28) => OP_WB(28), B(27) => 
                           OP_WB(27), B(26) => OP_WB(26), B(25) => OP_WB(25), 
                           B(24) => OP_WB(24), B(23) => OP_WB(23), B(22) => 
                           OP_WB(22), B(21) => OP_WB(21), B(20) => OP_WB(20), 
                           B(19) => OP_WB(19), B(18) => OP_WB(18), B(17) => 
                           OP_WB(17), B(16) => OP_WB(16), B(15) => OP_WB(15), 
                           B(14) => OP_WB(14), B(13) => OP_WB(13), B(12) => 
                           OP_WB(12), B(11) => OP_WB(11), B(10) => OP_WB(10), 
                           B(9) => OP_WB(9), B(8) => OP_WB(8), B(7) => OP_WB(7)
                           , B(6) => OP_WB(6), B(5) => OP_WB(5), B(4) => 
                           OP_WB(4), B(3) => OP_WB(3), B(2) => OP_WB(2), B(1) 
                           => OP_WB(1), B(0) => OP_WB(0), C(31) => OP_MEM(31), 
                           C(30) => OP_MEM(30), C(29) => OP_MEM(29), C(28) => 
                           OP_MEM(28), C(27) => OP_MEM(27), C(26) => OP_MEM(26)
                           , C(25) => OP_MEM(25), C(24) => OP_MEM(24), C(23) =>
                           OP_MEM(23), C(22) => OP_MEM(22), C(21) => OP_MEM(21)
                           , C(20) => OP_MEM(20), C(19) => OP_MEM(19), C(18) =>
                           OP_MEM(18), C(17) => OP_MEM(17), C(16) => OP_MEM(16)
                           , C(15) => OP_MEM(15), C(14) => OP_MEM(14), C(13) =>
                           OP_MEM(13), C(12) => OP_MEM(12), C(11) => OP_MEM(11)
                           , C(10) => OP_MEM(10), C(9) => OP_MEM(9), C(8) => 
                           OP_MEM(8), C(7) => OP_MEM(7), C(6) => OP_MEM(6), 
                           C(5) => OP_MEM(5), C(4) => OP_MEM(4), C(3) => 
                           OP_MEM(3), C(2) => OP_MEM(2), C(1) => OP_MEM(1), 
                           C(0) => OP_MEM(0), D(31) => B_IN(31), D(30) => 
                           B_IN(30), D(29) => B_IN(29), D(28) => B_IN(28), 
                           D(27) => B_IN(27), D(26) => B_IN(26), D(25) => 
                           B_IN(25), D(24) => B_IN(24), D(23) => B_IN(23), 
                           D(22) => B_IN(22), D(21) => B_IN(21), D(20) => 
                           B_IN(20), D(19) => B_IN(19), D(18) => B_IN(18), 
                           D(17) => B_IN(17), D(16) => B_IN(16), D(15) => 
                           B_IN(15), D(14) => B_IN(14), D(13) => B_IN(13), 
                           D(12) => B_IN(12), D(11) => B_IN(11), D(10) => 
                           B_IN(10), D(9) => B_IN(9), D(8) => B_IN(8), D(7) => 
                           B_IN(7), D(6) => B_IN(6), D(5) => B_IN(5), D(4) => 
                           B_IN(4), D(3) => B_IN(3), D(2) => B_IN(2), D(1) => 
                           B_IN(1), D(0) => B_IN(0), S(1) => FWDB_1_port, S(0) 
                           => FWDB_0_port, Z(31) => OP2_FW_31_port, Z(30) => 
                           OP2_FW_30_port, Z(29) => OP2_FW_29_port, Z(28) => 
                           OP2_FW_28_port, Z(27) => OP2_FW_27_port, Z(26) => 
                           OP2_FW_26_port, Z(25) => OP2_FW_25_port, Z(24) => 
                           OP2_FW_24_port, Z(23) => OP2_FW_23_port, Z(22) => 
                           OP2_FW_22_port, Z(21) => OP2_FW_21_port, Z(20) => 
                           OP2_FW_20_port, Z(19) => OP2_FW_19_port, Z(18) => 
                           OP2_FW_18_port, Z(17) => OP2_FW_17_port, Z(16) => 
                           OP2_FW_16_port, Z(15) => OP2_FW_15_port, Z(14) => 
                           OP2_FW_14_port, Z(13) => OP2_FW_13_port, Z(12) => 
                           OP2_FW_12_port, Z(11) => OP2_FW_11_port, Z(10) => 
                           OP2_FW_10_port, Z(9) => OP2_FW_9_port, Z(8) => 
                           OP2_FW_8_port, Z(7) => OP2_FW_7_port, Z(6) => 
                           OP2_FW_6_port, Z(5) => OP2_FW_5_port, Z(4) => 
                           OP2_FW_4_port, Z(3) => OP2_FW_3_port, Z(2) => 
                           OP2_FW_2_port, Z(1) => OP2_FW_1_port, Z(0) => 
                           OP2_FW_0_port);
   muxA : mux21_NBIT32_4 port map( A(31) => sig_NPC_ABS_31_port, A(30) => 
                           sig_NPC_ABS_30_port, A(29) => sig_NPC_ABS_29_port, 
                           A(28) => sig_NPC_ABS_28_port, A(27) => 
                           sig_NPC_ABS_27_port, A(26) => sig_NPC_ABS_26_port, 
                           A(25) => sig_NPC_ABS_25_port, A(24) => 
                           sig_NPC_ABS_24_port, A(23) => sig_NPC_ABS_23_port, 
                           A(22) => sig_NPC_ABS_22_port, A(21) => 
                           sig_NPC_ABS_21_port, A(20) => sig_NPC_ABS_20_port, 
                           A(19) => sig_NPC_ABS_19_port, A(18) => 
                           sig_NPC_ABS_18_port, A(17) => sig_NPC_ABS_17_port, 
                           A(16) => sig_NPC_ABS_16_port, A(15) => 
                           sig_NPC_ABS_15_port, A(14) => sig_NPC_ABS_14_port, 
                           A(13) => sig_NPC_ABS_13_port, A(12) => 
                           sig_NPC_ABS_12_port, A(11) => sig_NPC_ABS_11_port, 
                           A(10) => sig_NPC_ABS_10_port, A(9) => 
                           sig_NPC_ABS_9_port, A(8) => sig_NPC_ABS_8_port, A(7)
                           => sig_NPC_ABS_7_port, A(6) => sig_NPC_ABS_6_port, 
                           A(5) => sig_NPC_ABS_5_port, A(4) => 
                           sig_NPC_ABS_4_port, A(3) => sig_NPC_ABS_3_port, A(2)
                           => sig_NPC_ABS_2_port, A(1) => sig_NPC_ABS_1_port, 
                           A(0) => sig_NPC_ABS_0_port, B(31) => PC_IN(31), 
                           B(30) => PC_IN(30), B(29) => PC_IN(29), B(28) => 
                           PC_IN(28), B(27) => PC_IN(27), B(26) => PC_IN(26), 
                           B(25) => PC_IN(25), B(24) => PC_IN(24), B(23) => 
                           PC_IN(23), B(22) => PC_IN(22), B(21) => PC_IN(21), 
                           B(20) => PC_IN(20), B(19) => PC_IN(19), B(18) => 
                           PC_IN(18), B(17) => PC_IN(17), B(16) => PC_IN(16), 
                           B(15) => PC_IN(15), B(14) => PC_IN(14), B(13) => 
                           PC_IN(13), B(12) => PC_IN(12), B(11) => PC_IN(11), 
                           B(10) => PC_IN(10), B(9) => PC_IN(9), B(8) => 
                           PC_IN(8), B(7) => PC_IN(7), B(6) => PC_IN(6), B(5) 
                           => PC_IN(5), B(4) => PC_IN(4), B(3) => PC_IN(3), 
                           B(2) => PC_IN(2), B(1) => PC_IN(1), B(0) => PC_IN(0)
                           , S => MUX_A_SEL, Z(31) => sig_OP1_31_port, Z(30) =>
                           sig_OP1_30_port, Z(29) => sig_OP1_29_port, Z(28) => 
                           sig_OP1_28_port, Z(27) => sig_OP1_27_port, Z(26) => 
                           sig_OP1_26_port, Z(25) => sig_OP1_25_port, Z(24) => 
                           sig_OP1_24_port, Z(23) => sig_OP1_23_port, Z(22) => 
                           sig_OP1_22_port, Z(21) => sig_OP1_21_port, Z(20) => 
                           sig_OP1_20_port, Z(19) => sig_OP1_19_port, Z(18) => 
                           sig_OP1_18_port, Z(17) => sig_OP1_17_port, Z(16) => 
                           sig_OP1_16_port, Z(15) => sig_OP1_15_port, Z(14) => 
                           sig_OP1_14_port, Z(13) => sig_OP1_13_port, Z(12) => 
                           sig_OP1_12_port, Z(11) => sig_OP1_11_port, Z(10) => 
                           sig_OP1_10_port, Z(9) => sig_OP1_9_port, Z(8) => 
                           sig_OP1_8_port, Z(7) => sig_OP1_7_port, Z(6) => 
                           sig_OP1_6_port, Z(5) => sig_OP1_5_port, Z(4) => 
                           sig_OP1_4_port, Z(3) => sig_OP1_3_port, Z(2) => 
                           sig_OP1_2_port, Z(1) => sig_OP1_1_port, Z(0) => 
                           sig_OP1_0_port);
   muxB : mux41_NBIT32_3 port map( A(31) => OP2_FW_31_port, A(30) => 
                           OP2_FW_30_port, A(29) => OP2_FW_29_port, A(28) => 
                           OP2_FW_28_port, A(27) => OP2_FW_27_port, A(26) => 
                           OP2_FW_26_port, A(25) => OP2_FW_25_port, A(24) => 
                           OP2_FW_24_port, A(23) => OP2_FW_23_port, A(22) => 
                           OP2_FW_22_port, A(21) => OP2_FW_21_port, A(20) => 
                           OP2_FW_20_port, A(19) => OP2_FW_19_port, A(18) => 
                           OP2_FW_18_port, A(17) => OP2_FW_17_port, A(16) => 
                           OP2_FW_16_port, A(15) => OP2_FW_15_port, A(14) => 
                           OP2_FW_14_port, A(13) => OP2_FW_13_port, A(12) => 
                           OP2_FW_12_port, A(11) => OP2_FW_11_port, A(10) => 
                           OP2_FW_10_port, A(9) => OP2_FW_9_port, A(8) => 
                           OP2_FW_8_port, A(7) => OP2_FW_7_port, A(6) => 
                           OP2_FW_6_port, A(5) => OP2_FW_5_port, A(4) => 
                           OP2_FW_4_port, A(3) => OP2_FW_3_port, A(2) => 
                           OP2_FW_2_port, A(1) => OP2_FW_1_port, A(0) => 
                           OP2_FW_0_port, B(31) => IMM_IN(31), B(30) => 
                           IMM_IN(30), B(29) => IMM_IN(29), B(28) => IMM_IN(28)
                           , B(27) => IMM_IN(27), B(26) => IMM_IN(26), B(25) =>
                           IMM_IN(25), B(24) => IMM_IN(24), B(23) => IMM_IN(23)
                           , B(22) => IMM_IN(22), B(21) => IMM_IN(21), B(20) =>
                           IMM_IN(20), B(19) => IMM_IN(19), B(18) => IMM_IN(18)
                           , B(17) => IMM_IN(17), B(16) => IMM_IN(16), B(15) =>
                           IMM_IN(15), B(14) => IMM_IN(14), B(13) => IMM_IN(13)
                           , B(12) => IMM_IN(12), B(11) => IMM_IN(11), B(10) =>
                           IMM_IN(10), B(9) => IMM_IN(9), B(8) => IMM_IN(8), 
                           B(7) => IMM_IN(7), B(6) => IMM_IN(6), B(5) => 
                           IMM_IN(5), B(4) => IMM_IN(4), B(3) => IMM_IN(3), 
                           B(2) => IMM_IN(2), B(1) => IMM_IN(1), B(0) => 
                           IMM_IN(0), C(31) => n6_port, C(30) => n6_port, C(29)
                           => n6_port, C(28) => n6_port, C(27) => n6_port, 
                           C(26) => n6_port, C(25) => n6_port, C(24) => n6_port
                           , C(23) => n6_port, C(22) => n6_port, C(21) => 
                           n6_port, C(20) => n6_port, C(19) => n6_port, C(18) 
                           => n6_port, C(17) => n6_port, C(16) => n6_port, 
                           C(15) => n6_port, C(14) => n6_port, C(13) => n6_port
                           , C(12) => n6_port, C(11) => n6_port, C(10) => 
                           n6_port, C(9) => n6_port, C(8) => n6_port, C(7) => 
                           n6_port, C(6) => n6_port, C(5) => n6_port, C(4) => 
                           n6_port, C(3) => n6_port, C(2) => n7_port, C(1) => 
                           n6_port, C(0) => n6_port, D(31) => n6_port, D(30) =>
                           n6_port, D(29) => n6_port, D(28) => n6_port, D(27) 
                           => n6_port, D(26) => n6_port, D(25) => n6_port, 
                           D(24) => n6_port, D(23) => n6_port, D(22) => n6_port
                           , D(21) => n6_port, D(20) => n6_port, D(19) => 
                           n6_port, D(18) => n6_port, D(17) => n6_port, D(16) 
                           => n6_port, D(15) => n6_port, D(14) => n6_port, 
                           D(13) => n6_port, D(12) => n6_port, D(11) => n6_port
                           , D(10) => n6_port, D(9) => n6_port, D(8) => n6_port
                           , D(7) => n6_port, D(6) => n6_port, D(5) => n6_port,
                           D(4) => n6_port, D(3) => n6_port, D(2) => n6_port, 
                           D(1) => n6_port, D(0) => n6_port, S(1) => 
                           MUX_B_SEL(1), S(0) => MUX_B_SEL(0), Z(31) => 
                           sig_OP2_31_port, Z(30) => sig_OP2_30_port, Z(29) => 
                           sig_OP2_29_port, Z(28) => sig_OP2_28_port, Z(27) => 
                           sig_OP2_27_port, Z(26) => sig_OP2_26_port, Z(25) => 
                           sig_OP2_25_port, Z(24) => sig_OP2_24_port, Z(23) => 
                           sig_OP2_23_port, Z(22) => sig_OP2_22_port, Z(21) => 
                           sig_OP2_21_port, Z(20) => sig_OP2_20_port, Z(19) => 
                           sig_OP2_19_port, Z(18) => sig_OP2_18_port, Z(17) => 
                           sig_OP2_17_port, Z(16) => sig_OP2_16_port, Z(15) => 
                           sig_OP2_15_port, Z(14) => sig_OP2_14_port, Z(13) => 
                           sig_OP2_13_port, Z(12) => sig_OP2_12_port, Z(11) => 
                           sig_OP2_11_port, Z(10) => sig_OP2_10_port, Z(9) => 
                           sig_OP2_9_port, Z(8) => sig_OP2_8_port, Z(7) => 
                           sig_OP2_7_port, Z(6) => sig_OP2_6_port, Z(5) => 
                           sig_OP2_5_port, Z(4) => sig_OP2_4_port, Z(3) => 
                           sig_OP2_3_port, Z(2) => sig_OP2_2_port, Z(1) => 
                           sig_OP2_1_port, Z(0) => sig_OP2_0_port);
   alu0 : ALU_NBIT32 port map( OP1(31) => sig_OP1_31_port, OP1(30) => 
                           sig_OP1_30_port, OP1(29) => sig_OP1_29_port, OP1(28)
                           => sig_OP1_28_port, OP1(27) => sig_OP1_27_port, 
                           OP1(26) => sig_OP1_26_port, OP1(25) => 
                           sig_OP1_25_port, OP1(24) => sig_OP1_24_port, OP1(23)
                           => sig_OP1_23_port, OP1(22) => sig_OP1_22_port, 
                           OP1(21) => sig_OP1_21_port, OP1(20) => 
                           sig_OP1_20_port, OP1(19) => sig_OP1_19_port, OP1(18)
                           => sig_OP1_18_port, OP1(17) => sig_OP1_17_port, 
                           OP1(16) => sig_OP1_16_port, OP1(15) => 
                           sig_OP1_15_port, OP1(14) => sig_OP1_14_port, OP1(13)
                           => sig_OP1_13_port, OP1(12) => sig_OP1_12_port, 
                           OP1(11) => sig_OP1_11_port, OP1(10) => 
                           sig_OP1_10_port, OP1(9) => sig_OP1_9_port, OP1(8) =>
                           sig_OP1_8_port, OP1(7) => sig_OP1_7_port, OP1(6) => 
                           sig_OP1_6_port, OP1(5) => sig_OP1_5_port, OP1(4) => 
                           sig_OP1_4_port, OP1(3) => sig_OP1_3_port, OP1(2) => 
                           sig_OP1_2_port, OP1(1) => sig_OP1_1_port, OP1(0) => 
                           sig_OP1_0_port, OP2(31) => sig_OP2_31_port, OP2(30) 
                           => sig_OP2_30_port, OP2(29) => sig_OP2_29_port, 
                           OP2(28) => sig_OP2_28_port, OP2(27) => 
                           sig_OP2_27_port, OP2(26) => sig_OP2_26_port, OP2(25)
                           => sig_OP2_25_port, OP2(24) => sig_OP2_24_port, 
                           OP2(23) => sig_OP2_23_port, OP2(22) => 
                           sig_OP2_22_port, OP2(21) => sig_OP2_21_port, OP2(20)
                           => sig_OP2_20_port, OP2(19) => sig_OP2_19_port, 
                           OP2(18) => sig_OP2_18_port, OP2(17) => 
                           sig_OP2_17_port, OP2(16) => sig_OP2_16_port, OP2(15)
                           => sig_OP2_15_port, OP2(14) => sig_OP2_14_port, 
                           OP2(13) => sig_OP2_13_port, OP2(12) => 
                           sig_OP2_12_port, OP2(11) => sig_OP2_11_port, OP2(10)
                           => sig_OP2_10_port, OP2(9) => sig_OP2_9_port, OP2(8)
                           => sig_OP2_8_port, OP2(7) => sig_OP2_7_port, OP2(6) 
                           => sig_OP2_6_port, OP2(5) => sig_OP2_5_port, OP2(4) 
                           => sig_OP2_4_port, OP2(3) => sig_OP2_3_port, OP2(2) 
                           => sig_OP2_2_port, OP2(1) => sig_OP2_1_port, OP2(0) 
                           => sig_OP2_0_port, ALU_OPC(0) => ALU_OPC(0), 
                           ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => ALU_OPC(2), 
                           ALU_OPC(3) => ALU_OPC(3), ALU_OPC(4) => ALU_OPC(4), 
                           ALU_RES(31) => sig_ALU_RES_31_port, ALU_RES(30) => 
                           sig_ALU_RES_30_port, ALU_RES(29) => 
                           sig_ALU_RES_29_port, ALU_RES(28) => 
                           sig_ALU_RES_28_port, ALU_RES(27) => 
                           sig_ALU_RES_27_port, ALU_RES(26) => 
                           sig_ALU_RES_26_port, ALU_RES(25) => 
                           sig_ALU_RES_25_port, ALU_RES(24) => 
                           sig_ALU_RES_24_port, ALU_RES(23) => 
                           sig_ALU_RES_23_port, ALU_RES(22) => 
                           sig_ALU_RES_22_port, ALU_RES(21) => 
                           sig_ALU_RES_21_port, ALU_RES(20) => 
                           sig_ALU_RES_20_port, ALU_RES(19) => 
                           sig_ALU_RES_19_port, ALU_RES(18) => 
                           sig_ALU_RES_18_port, ALU_RES(17) => 
                           sig_ALU_RES_17_port, ALU_RES(16) => 
                           sig_ALU_RES_16_port, ALU_RES(15) => 
                           sig_ALU_RES_15_port, ALU_RES(14) => 
                           sig_ALU_RES_14_port, ALU_RES(13) => 
                           sig_ALU_RES_13_port, ALU_RES(12) => 
                           sig_ALU_RES_12_port, ALU_RES(11) => 
                           sig_ALU_RES_11_port, ALU_RES(10) => 
                           sig_ALU_RES_10_port, ALU_RES(9) => 
                           sig_ALU_RES_9_port, ALU_RES(8) => sig_ALU_RES_8_port
                           , ALU_RES(7) => sig_ALU_RES_7_port, ALU_RES(6) => 
                           sig_ALU_RES_6_port, ALU_RES(5) => sig_ALU_RES_5_port
                           , ALU_RES(4) => sig_ALU_RES_4_port, ALU_RES(3) => 
                           sig_ALU_RES_3_port, ALU_RES(2) => sig_ALU_RES_2_port
                           , ALU_RES(1) => sig_ALU_RES_1_port, ALU_RES(0) => 
                           sig_ALU_RES_0_port);
   alureg : regn_N32_5 port map( DIN(31) => sig_ALU_RES_31_port, DIN(30) => 
                           sig_ALU_RES_30_port, DIN(29) => sig_ALU_RES_29_port,
                           DIN(28) => sig_ALU_RES_28_port, DIN(27) => 
                           sig_ALU_RES_27_port, DIN(26) => sig_ALU_RES_26_port,
                           DIN(25) => sig_ALU_RES_25_port, DIN(24) => 
                           sig_ALU_RES_24_port, DIN(23) => sig_ALU_RES_23_port,
                           DIN(22) => sig_ALU_RES_22_port, DIN(21) => 
                           sig_ALU_RES_21_port, DIN(20) => sig_ALU_RES_20_port,
                           DIN(19) => sig_ALU_RES_19_port, DIN(18) => 
                           sig_ALU_RES_18_port, DIN(17) => sig_ALU_RES_17_port,
                           DIN(16) => sig_ALU_RES_16_port, DIN(15) => 
                           sig_ALU_RES_15_port, DIN(14) => sig_ALU_RES_14_port,
                           DIN(13) => sig_ALU_RES_13_port, DIN(12) => 
                           sig_ALU_RES_12_port, DIN(11) => sig_ALU_RES_11_port,
                           DIN(10) => sig_ALU_RES_10_port, DIN(9) => 
                           sig_ALU_RES_9_port, DIN(8) => sig_ALU_RES_8_port, 
                           DIN(7) => sig_ALU_RES_7_port, DIN(6) => 
                           sig_ALU_RES_6_port, DIN(5) => sig_ALU_RES_5_port, 
                           DIN(4) => sig_ALU_RES_4_port, DIN(3) => 
                           sig_ALU_RES_3_port, DIN(2) => sig_ALU_RES_2_port, 
                           DIN(1) => sig_ALU_RES_1_port, DIN(0) => 
                           sig_ALU_RES_0_port, CLK => CLK, EN => ALU_OUTREG_EN,
                           RST => RST, DOUT(31) => ALU_RES(31), DOUT(30) => 
                           ALU_RES(30), DOUT(29) => ALU_RES(29), DOUT(28) => 
                           ALU_RES(28), DOUT(27) => ALU_RES(27), DOUT(26) => 
                           ALU_RES(26), DOUT(25) => ALU_RES(25), DOUT(24) => 
                           ALU_RES(24), DOUT(23) => ALU_RES(23), DOUT(22) => 
                           ALU_RES(22), DOUT(21) => ALU_RES(21), DOUT(20) => 
                           ALU_RES(20), DOUT(19) => ALU_RES(19), DOUT(18) => 
                           ALU_RES(18), DOUT(17) => ALU_RES(17), DOUT(16) => 
                           ALU_RES(16), DOUT(15) => ALU_RES(15), DOUT(14) => 
                           ALU_RES(14), DOUT(13) => ALU_RES(13), DOUT(12) => 
                           ALU_RES(12), DOUT(11) => ALU_RES(11), DOUT(10) => 
                           ALU_RES(10), DOUT(9) => ALU_RES(9), DOUT(8) => 
                           ALU_RES(8), DOUT(7) => ALU_RES(7), DOUT(6) => 
                           ALU_RES(6), DOUT(5) => ALU_RES(5), DOUT(4) => 
                           ALU_RES(4), DOUT(3) => ALU_RES(3), DOUT(2) => 
                           ALU_RES(2), DOUT(1) => ALU_RES(1), DOUT(0) => 
                           ALU_RES(0));
   B_reg : regn_N32_4 port map( DIN(31) => OP2_FW_31_port, DIN(30) => 
                           OP2_FW_30_port, DIN(29) => OP2_FW_29_port, DIN(28) 
                           => OP2_FW_28_port, DIN(27) => OP2_FW_27_port, 
                           DIN(26) => OP2_FW_26_port, DIN(25) => OP2_FW_25_port
                           , DIN(24) => OP2_FW_24_port, DIN(23) => 
                           OP2_FW_23_port, DIN(22) => OP2_FW_22_port, DIN(21) 
                           => OP2_FW_21_port, DIN(20) => OP2_FW_20_port, 
                           DIN(19) => OP2_FW_19_port, DIN(18) => OP2_FW_18_port
                           , DIN(17) => OP2_FW_17_port, DIN(16) => 
                           OP2_FW_16_port, DIN(15) => OP2_FW_15_port, DIN(14) 
                           => OP2_FW_14_port, DIN(13) => OP2_FW_13_port, 
                           DIN(12) => OP2_FW_12_port, DIN(11) => OP2_FW_11_port
                           , DIN(10) => OP2_FW_10_port, DIN(9) => OP2_FW_9_port
                           , DIN(8) => OP2_FW_8_port, DIN(7) => OP2_FW_7_port, 
                           DIN(6) => OP2_FW_6_port, DIN(5) => OP2_FW_5_port, 
                           DIN(4) => OP2_FW_4_port, DIN(3) => OP2_FW_3_port, 
                           DIN(2) => OP2_FW_2_port, DIN(1) => OP2_FW_1_port, 
                           DIN(0) => OP2_FW_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => B_OUT(31), 
                           DOUT(30) => B_OUT(30), DOUT(29) => B_OUT(29), 
                           DOUT(28) => B_OUT(28), DOUT(27) => B_OUT(27), 
                           DOUT(26) => B_OUT(26), DOUT(25) => B_OUT(25), 
                           DOUT(24) => B_OUT(24), DOUT(23) => B_OUT(23), 
                           DOUT(22) => B_OUT(22), DOUT(21) => B_OUT(21), 
                           DOUT(20) => B_OUT(20), DOUT(19) => B_OUT(19), 
                           DOUT(18) => B_OUT(18), DOUT(17) => B_OUT(17), 
                           DOUT(16) => B_OUT(16), DOUT(15) => B_OUT(15), 
                           DOUT(14) => B_OUT(14), DOUT(13) => B_OUT(13), 
                           DOUT(12) => B_OUT(12), DOUT(11) => B_OUT(11), 
                           DOUT(10) => B_OUT(10), DOUT(9) => B_OUT(9), DOUT(8) 
                           => B_OUT(8), DOUT(7) => B_OUT(7), DOUT(6) => 
                           B_OUT(6), DOUT(5) => B_OUT(5), DOUT(4) => B_OUT(4), 
                           DOUT(3) => B_OUT(3), DOUT(2) => B_OUT(2), DOUT(1) =>
                           B_OUT(1), DOUT(0) => B_OUT(0));
   ADD_WR_reg : regn_N5_2 port map( DIN(4) => ADD_WR_IN(4), DIN(3) => 
                           ADD_WR_IN(3), DIN(2) => ADD_WR_IN(2), DIN(1) => 
                           ADD_WR_IN(1), DIN(0) => ADD_WR_IN(0), CLK => CLK, EN
                           => n7_port, RST => RST, DOUT(4) => ADD_WR_OUT(4), 
                           DOUT(3) => ADD_WR_OUT(3), DOUT(2) => ADD_WR_OUT(2), 
                           DOUT(1) => ADD_WR_OUT(1), DOUT(0) => ADD_WR_OUT(0));
   NPC_ABS_reg : regn_N32_3 port map( DIN(31) => sig_NPC_ABS_31_port, DIN(30) 
                           => sig_NPC_ABS_30_port, DIN(29) => 
                           sig_NPC_ABS_29_port, DIN(28) => sig_NPC_ABS_28_port,
                           DIN(27) => sig_NPC_ABS_27_port, DIN(26) => 
                           sig_NPC_ABS_26_port, DIN(25) => sig_NPC_ABS_25_port,
                           DIN(24) => sig_NPC_ABS_24_port, DIN(23) => 
                           sig_NPC_ABS_23_port, DIN(22) => sig_NPC_ABS_22_port,
                           DIN(21) => sig_NPC_ABS_21_port, DIN(20) => 
                           sig_NPC_ABS_20_port, DIN(19) => sig_NPC_ABS_19_port,
                           DIN(18) => sig_NPC_ABS_18_port, DIN(17) => 
                           sig_NPC_ABS_17_port, DIN(16) => sig_NPC_ABS_16_port,
                           DIN(15) => sig_NPC_ABS_15_port, DIN(14) => 
                           sig_NPC_ABS_14_port, DIN(13) => sig_NPC_ABS_13_port,
                           DIN(12) => sig_NPC_ABS_12_port, DIN(11) => 
                           sig_NPC_ABS_11_port, DIN(10) => sig_NPC_ABS_10_port,
                           DIN(9) => sig_NPC_ABS_9_port, DIN(8) => 
                           sig_NPC_ABS_8_port, DIN(7) => sig_NPC_ABS_7_port, 
                           DIN(6) => sig_NPC_ABS_6_port, DIN(5) => 
                           sig_NPC_ABS_5_port, DIN(4) => sig_NPC_ABS_4_port, 
                           DIN(3) => sig_NPC_ABS_3_port, DIN(2) => 
                           sig_NPC_ABS_2_port, DIN(1) => sig_NPC_ABS_1_port, 
                           DIN(0) => sig_NPC_ABS_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => NPC_ABS(31), 
                           DOUT(30) => NPC_ABS(30), DOUT(29) => NPC_ABS(29), 
                           DOUT(28) => NPC_ABS(28), DOUT(27) => NPC_ABS(27), 
                           DOUT(26) => NPC_ABS(26), DOUT(25) => NPC_ABS(25), 
                           DOUT(24) => NPC_ABS(24), DOUT(23) => NPC_ABS(23), 
                           DOUT(22) => NPC_ABS(22), DOUT(21) => NPC_ABS(21), 
                           DOUT(20) => NPC_ABS(20), DOUT(19) => NPC_ABS(19), 
                           DOUT(18) => NPC_ABS(18), DOUT(17) => NPC_ABS(17), 
                           DOUT(16) => NPC_ABS(16), DOUT(15) => NPC_ABS(15), 
                           DOUT(14) => NPC_ABS(14), DOUT(13) => NPC_ABS(13), 
                           DOUT(12) => NPC_ABS(12), DOUT(11) => NPC_ABS(11), 
                           DOUT(10) => NPC_ABS(10), DOUT(9) => NPC_ABS(9), 
                           DOUT(8) => NPC_ABS(8), DOUT(7) => NPC_ABS(7), 
                           DOUT(6) => NPC_ABS(6), DOUT(5) => NPC_ABS(5), 
                           DOUT(4) => NPC_ABS(4), DOUT(3) => NPC_ABS(3), 
                           DOUT(2) => NPC_ABS(2), DOUT(1) => NPC_ABS(1), 
                           DOUT(0) => NPC_ABS(0));
   NPC_REL_reg : regn_N32_2 port map( DIN(31) => sig_NPC_REL_31_port, DIN(30) 
                           => sig_NPC_REL_30_port, DIN(29) => 
                           sig_NPC_REL_29_port, DIN(28) => sig_NPC_REL_28_port,
                           DIN(27) => sig_NPC_REL_27_port, DIN(26) => 
                           sig_NPC_REL_26_port, DIN(25) => sig_NPC_REL_25_port,
                           DIN(24) => sig_NPC_REL_24_port, DIN(23) => 
                           sig_NPC_REL_23_port, DIN(22) => sig_NPC_REL_22_port,
                           DIN(21) => sig_NPC_REL_21_port, DIN(20) => 
                           sig_NPC_REL_20_port, DIN(19) => sig_NPC_REL_19_port,
                           DIN(18) => sig_NPC_REL_18_port, DIN(17) => 
                           sig_NPC_REL_17_port, DIN(16) => sig_NPC_REL_16_port,
                           DIN(15) => sig_NPC_REL_15_port, DIN(14) => 
                           sig_NPC_REL_14_port, DIN(13) => sig_NPC_REL_13_port,
                           DIN(12) => sig_NPC_REL_12_port, DIN(11) => 
                           sig_NPC_REL_11_port, DIN(10) => sig_NPC_REL_10_port,
                           DIN(9) => sig_NPC_REL_9_port, DIN(8) => 
                           sig_NPC_REL_8_port, DIN(7) => sig_NPC_REL_7_port, 
                           DIN(6) => sig_NPC_REL_6_port, DIN(5) => 
                           sig_NPC_REL_5_port, DIN(4) => sig_NPC_REL_4_port, 
                           DIN(3) => sig_NPC_REL_3_port, DIN(2) => 
                           sig_NPC_REL_2_port, DIN(1) => sig_NPC_REL_1_port, 
                           DIN(0) => sig_NPC_REL_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => NPC_REL(31), 
                           DOUT(30) => NPC_REL(30), DOUT(29) => NPC_REL(29), 
                           DOUT(28) => NPC_REL(28), DOUT(27) => NPC_REL(27), 
                           DOUT(26) => NPC_REL(26), DOUT(25) => NPC_REL(25), 
                           DOUT(24) => NPC_REL(24), DOUT(23) => NPC_REL(23), 
                           DOUT(22) => NPC_REL(22), DOUT(21) => NPC_REL(21), 
                           DOUT(20) => NPC_REL(20), DOUT(19) => NPC_REL(19), 
                           DOUT(18) => NPC_REL(18), DOUT(17) => NPC_REL(17), 
                           DOUT(16) => NPC_REL(16), DOUT(15) => NPC_REL(15), 
                           DOUT(14) => NPC_REL(14), DOUT(13) => NPC_REL(13), 
                           DOUT(12) => NPC_REL(12), DOUT(11) => NPC_REL(11), 
                           DOUT(10) => NPC_REL(10), DOUT(9) => NPC_REL(9), 
                           DOUT(8) => NPC_REL(8), DOUT(7) => NPC_REL(7), 
                           DOUT(6) => NPC_REL(6), DOUT(5) => NPC_REL(5), 
                           DOUT(4) => NPC_REL(4), DOUT(3) => NPC_REL(3), 
                           DOUT(2) => NPC_REL(2), DOUT(1) => NPC_REL(1), 
                           DOUT(0) => NPC_REL(0));
   add_1_root_add_0_root_add_122_2 : Execute_DW01_add_1 port map( A(31) => 
                           n2_port, A(30) => n2_port, A(29) => n2_port, A(28) 
                           => n2_port, A(27) => n2_port, A(26) => n2_port, 
                           A(25) => n2_port, A(24) => n2_port, A(23) => n2_port
                           , A(22) => n2_port, A(21) => n2_port, A(20) => 
                           n2_port, A(19) => n2_port, A(18) => n2_port, A(17) 
                           => n2_port, A(16) => n2_port, A(15) => n2_port, 
                           A(14) => n2_port, A(13) => n2_port, A(12) => n2_port
                           , A(11) => n2_port, A(10) => n2_port, A(9) => 
                           n2_port, A(8) => n2_port, A(7) => n2_port, A(6) => 
                           n2_port, A(5) => n2_port, A(4) => n2_port, A(3) => 
                           n2_port, A(2) => n3_port, A(1) => n2_port, A(0) => 
                           n2_port, B(31) => IMM_IN(31), B(30) => IMM_IN(30), 
                           B(29) => IMM_IN(29), B(28) => IMM_IN(28), B(27) => 
                           IMM_IN(27), B(26) => IMM_IN(26), B(25) => IMM_IN(25)
                           , B(24) => IMM_IN(24), B(23) => IMM_IN(23), B(22) =>
                           IMM_IN(22), B(21) => IMM_IN(21), B(20) => IMM_IN(20)
                           , B(19) => IMM_IN(19), B(18) => IMM_IN(18), B(17) =>
                           IMM_IN(17), B(16) => IMM_IN(16), B(15) => IMM_IN(15)
                           , B(14) => IMM_IN(14), B(13) => IMM_IN(13), B(12) =>
                           IMM_IN(12), B(11) => IMM_IN(11), B(10) => IMM_IN(10)
                           , B(9) => IMM_IN(9), B(8) => IMM_IN(8), B(7) => 
                           IMM_IN(7), B(6) => IMM_IN(6), B(5) => IMM_IN(5), 
                           B(4) => IMM_IN(4), B(3) => IMM_IN(3), B(2) => 
                           IMM_IN(2), B(1) => IMM_IN(1), B(0) => IMM_IN(0), CI 
                           => n4_port, SUM(31) => N31, SUM(30) => N30, SUM(29) 
                           => N29, SUM(28) => N28, SUM(27) => N27, SUM(26) => 
                           N26, SUM(25) => N25, SUM(24) => N24, SUM(23) => N23,
                           SUM(22) => N22, SUM(21) => N21, SUM(20) => N20, 
                           SUM(19) => N19, SUM(18) => N18, SUM(17) => N17, 
                           SUM(16) => N16, SUM(15) => N15, SUM(14) => N14, 
                           SUM(13) => N13, SUM(12) => N12, SUM(11) => N11, 
                           SUM(10) => N10, SUM(9) => N9, SUM(8) => N8, SUM(7) 
                           => N7, SUM(6) => N6, SUM(5) => N5, SUM(4) => N4, 
                           SUM(3) => N3, SUM(2) => N2, SUM(1) => N1, SUM(0) => 
                           N0, CO => n_1596);
   add_0_root_add_0_root_add_122_2 : Execute_DW01_add_0 port map( A(31) => 
                           PC_IN(31), A(30) => PC_IN(30), A(29) => PC_IN(29), 
                           A(28) => PC_IN(28), A(27) => PC_IN(27), A(26) => 
                           PC_IN(26), A(25) => PC_IN(25), A(24) => PC_IN(24), 
                           A(23) => PC_IN(23), A(22) => PC_IN(22), A(21) => 
                           PC_IN(21), A(20) => PC_IN(20), A(19) => PC_IN(19), 
                           A(18) => PC_IN(18), A(17) => PC_IN(17), A(16) => 
                           PC_IN(16), A(15) => PC_IN(15), A(14) => PC_IN(14), 
                           A(13) => PC_IN(13), A(12) => PC_IN(12), A(11) => 
                           PC_IN(11), A(10) => PC_IN(10), A(9) => PC_IN(9), 
                           A(8) => PC_IN(8), A(7) => PC_IN(7), A(6) => PC_IN(6)
                           , A(5) => PC_IN(5), A(4) => PC_IN(4), A(3) => 
                           PC_IN(3), A(2) => PC_IN(2), A(1) => PC_IN(1), A(0) 
                           => PC_IN(0), B(31) => N31, B(30) => N30, B(29) => 
                           N29, B(28) => N28, B(27) => N27, B(26) => N26, B(25)
                           => N25, B(24) => N24, B(23) => N23, B(22) => N22, 
                           B(21) => N21, B(20) => N20, B(19) => N19, B(18) => 
                           N18, B(17) => N17, B(16) => N16, B(15) => N15, B(14)
                           => N14, B(13) => N13, B(12) => N12, B(11) => N11, 
                           B(10) => N10, B(9) => N9, B(8) => N8, B(7) => N7, 
                           B(6) => N6, B(5) => N5, B(4) => N4, B(3) => N3, B(2)
                           => N2, B(1) => N1, B(0) => N0, CI => n5_port, 
                           SUM(31) => sig_NPC_REL_31_port, SUM(30) => 
                           sig_NPC_REL_30_port, SUM(29) => sig_NPC_REL_29_port,
                           SUM(28) => sig_NPC_REL_28_port, SUM(27) => 
                           sig_NPC_REL_27_port, SUM(26) => sig_NPC_REL_26_port,
                           SUM(25) => sig_NPC_REL_25_port, SUM(24) => 
                           sig_NPC_REL_24_port, SUM(23) => sig_NPC_REL_23_port,
                           SUM(22) => sig_NPC_REL_22_port, SUM(21) => 
                           sig_NPC_REL_21_port, SUM(20) => sig_NPC_REL_20_port,
                           SUM(19) => sig_NPC_REL_19_port, SUM(18) => 
                           sig_NPC_REL_18_port, SUM(17) => sig_NPC_REL_17_port,
                           SUM(16) => sig_NPC_REL_16_port, SUM(15) => 
                           sig_NPC_REL_15_port, SUM(14) => sig_NPC_REL_14_port,
                           SUM(13) => sig_NPC_REL_13_port, SUM(12) => 
                           sig_NPC_REL_12_port, SUM(11) => sig_NPC_REL_11_port,
                           SUM(10) => sig_NPC_REL_10_port, SUM(9) => 
                           sig_NPC_REL_9_port, SUM(8) => sig_NPC_REL_8_port, 
                           SUM(7) => sig_NPC_REL_7_port, SUM(6) => 
                           sig_NPC_REL_6_port, SUM(5) => sig_NPC_REL_5_port, 
                           SUM(4) => sig_NPC_REL_4_port, SUM(3) => 
                           sig_NPC_REL_3_port, SUM(2) => sig_NPC_REL_2_port, 
                           SUM(1) => sig_NPC_REL_1_port, SUM(0) => 
                           sig_NPC_REL_0_port, CO => n_1597);
   U3 : NOR2_X1 port map( A1 => ZERO_FLAG_port, A2 => n1_port, ZN => sig_RST);
   U4 : INV_X1 port map( A => RST, ZN => n1_port);
   n2_port <= '0';
   n3_port <= '1';
   n4_port <= '0';
   n5_port <= '0';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Decode is

   port( CLK, RST, Bubble, RF_WE, ZERO_FLAG : in std_logic;  PC_IN, INS_IN : in
         std_logic_vector (31 downto 0);  ADD_WR : in std_logic_vector (4 
         downto 0);  DATA_WR_IN : in std_logic_vector (31 downto 0);  PC_OUT, 
         A_OUT, B_OUT, IMM_OUT : out std_logic_vector (31 downto 0);  
         ADD_RS1_HDU, ADD_RS2_HDU, ADD_WR_OUT, ADD_RS1_OUT, ADD_RS2_OUT : out 
         std_logic_vector (4 downto 0));

end Decode;

architecture SYN_struct of Decode is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component register_file_NBIT_ADD5_NBIT_DATA32
      port( CLK, RST, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RS1, 
            ADD_RS2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component mux21_NBIT5_1
      port( A, B : in std_logic_vector (4 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component mux21_NBIT5_2
      port( A, B : in std_logic_vector (4 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component mux21_NBIT5_0
      port( A, B : in std_logic_vector (4 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N5_3
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N5_4
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N5_0
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N32_6
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_7
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component instruction_decomposition
      port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype :
            in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : out std_logic_vector (4 
            downto 0);  IMM : out std_logic_vector (31 downto 0);  RD1, RD2 : 
            out std_logic);
   end component;
   
   component instruction_type
      port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype :
            out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, n21, n22, n23, n24, n25, n26, n27, n28,
      n29, n30, sig_RST, sig_Rtype, sig_Itype, sig_Jtype, sig_ADD_WR_4_port, 
      sig_ADD_WR_3_port, sig_ADD_WR_2_port, sig_ADD_WR_1_port, 
      sig_ADD_WR_0_port, sig_IMM_31_port, sig_IMM_30_port, sig_IMM_29_port, 
      sig_IMM_28_port, sig_IMM_27_port, sig_IMM_26_port, sig_IMM_25_port, 
      sig_IMM_24_port, sig_IMM_23_port, sig_IMM_22_port, sig_IMM_21_port, 
      sig_IMM_20_port, sig_IMM_19_port, sig_IMM_18_port, sig_IMM_17_port, 
      sig_IMM_16_port, sig_IMM_15_port, sig_IMM_14_port, sig_IMM_13_port, 
      sig_IMM_12_port, sig_IMM_11_port, sig_IMM_10_port, sig_IMM_9_port, 
      sig_IMM_8_port, sig_IMM_7_port, sig_IMM_6_port, sig_IMM_5_port, 
      sig_IMM_4_port, sig_IMM_3_port, sig_IMM_2_port, sig_IMM_1_port, 
      sig_IMM_0_port, RD1, RD2, sig_ADD_WRHAZ_4_port, sig_ADD_WRHAZ_3_port, 
      sig_ADD_WRHAZ_2_port, sig_ADD_WRHAZ_1_port, sig_ADD_WRHAZ_0_port, 
      sig_ADD_RS1HAZ_4_port, sig_ADD_RS1HAZ_3_port, sig_ADD_RS1HAZ_2_port, 
      sig_ADD_RS1HAZ_1_port, sig_ADD_RS1HAZ_0_port, sig_ADD_RS2HAZ_4_port, 
      sig_ADD_RS2HAZ_3_port, sig_ADD_RS2HAZ_2_port, sig_ADD_RS2HAZ_1_port, 
      sig_ADD_RS2HAZ_0_port, n1, ADD_RS1_HDU_1_port, n3, n4, ADD_RS1_HDU_0_port
      , n6, ADD_RS2_HDU_1_port, ADD_RS2_HDU_3_port, ADD_RS2_HDU_4_port, n10, 
      n11, n12, ADD_RS1_HDU_2_port, ADD_RS2_HDU_0_port, ADD_RS2_HDU_2_port, 
      ADD_RS1_HDU_3_port, ADD_RS1_HDU_4_port, n18, n19, n20 : std_logic;

begin
   ADD_RS1_HDU <= ( ADD_RS1_HDU_4_port, ADD_RS1_HDU_3_port, ADD_RS1_HDU_2_port,
      ADD_RS1_HDU_1_port, ADD_RS1_HDU_0_port );
   ADD_RS2_HDU <= ( ADD_RS2_HDU_4_port, ADD_RS2_HDU_3_port, ADD_RS2_HDU_2_port,
      ADD_RS2_HDU_1_port, ADD_RS2_HDU_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   U3 : NOR2_X2 port map( A1 => ZERO_FLAG, A2 => n20, ZN => sig_RST);
   ins_type : instruction_type port map( INST_IN(31) => INS_IN(31), INST_IN(30)
                           => INS_IN(30), INST_IN(29) => INS_IN(29), 
                           INST_IN(28) => INS_IN(28), INST_IN(27) => INS_IN(27)
                           , INST_IN(26) => INS_IN(26), INST_IN(25) => 
                           INS_IN(25), INST_IN(24) => INS_IN(24), INST_IN(23) 
                           => INS_IN(23), INST_IN(22) => INS_IN(22), 
                           INST_IN(21) => INS_IN(21), INST_IN(20) => INS_IN(20)
                           , INST_IN(19) => INS_IN(19), INST_IN(18) => 
                           INS_IN(18), INST_IN(17) => INS_IN(17), INST_IN(16) 
                           => INS_IN(16), INST_IN(15) => INS_IN(15), 
                           INST_IN(14) => INS_IN(14), INST_IN(13) => INS_IN(13)
                           , INST_IN(12) => INS_IN(12), INST_IN(11) => 
                           INS_IN(11), INST_IN(10) => INS_IN(10), INST_IN(9) =>
                           INS_IN(9), INST_IN(8) => INS_IN(8), INST_IN(7) => 
                           INS_IN(7), INST_IN(6) => INS_IN(6), INST_IN(5) => 
                           INS_IN(5), INST_IN(4) => INS_IN(4), INST_IN(3) => 
                           INS_IN(3), INST_IN(2) => INS_IN(2), INST_IN(1) => 
                           INS_IN(1), INST_IN(0) => INS_IN(0), Rtype => 
                           sig_Rtype, Itype => sig_Itype, Jtype => sig_Jtype);
   ins_dec : instruction_decomposition port map( INST_IN(31) => INS_IN(31), 
                           INST_IN(30) => INS_IN(30), INST_IN(29) => INS_IN(29)
                           , INST_IN(28) => INS_IN(28), INST_IN(27) => n12, 
                           INST_IN(26) => n11, INST_IN(25) => INS_IN(25), 
                           INST_IN(24) => INS_IN(24), INST_IN(23) => INS_IN(23)
                           , INST_IN(22) => INS_IN(22), INST_IN(21) => 
                           INS_IN(21), INST_IN(20) => INS_IN(20), INST_IN(19) 
                           => INS_IN(19), INST_IN(18) => INS_IN(18), 
                           INST_IN(17) => INS_IN(17), INST_IN(16) => INS_IN(16)
                           , INST_IN(15) => INS_IN(15), INST_IN(14) => 
                           INS_IN(14), INST_IN(13) => INS_IN(13), INST_IN(12) 
                           => INS_IN(12), INST_IN(11) => INS_IN(11), 
                           INST_IN(10) => INS_IN(10), INST_IN(9) => INS_IN(9), 
                           INST_IN(8) => INS_IN(8), INST_IN(7) => INS_IN(7), 
                           INST_IN(6) => INS_IN(6), INST_IN(5) => INS_IN(5), 
                           INST_IN(4) => INS_IN(4), INST_IN(3) => INS_IN(3), 
                           INST_IN(2) => INS_IN(2), INST_IN(1) => INS_IN(1), 
                           INST_IN(0) => INS_IN(0), Rtype => sig_Rtype, Itype 
                           => sig_Itype, Jtype => sig_Jtype, ADD_RS1(4) => n21,
                           ADD_RS1(3) => n22, ADD_RS1(2) => n23, ADD_RS1(1) => 
                           n24, ADD_RS1(0) => n25, ADD_RS2(4) => n26, 
                           ADD_RS2(3) => n27, ADD_RS2(2) => n28, ADD_RS2(1) => 
                           n29, ADD_RS2(0) => n30, ADD_WR(4) => 
                           sig_ADD_WR_4_port, ADD_WR(3) => sig_ADD_WR_3_port, 
                           ADD_WR(2) => sig_ADD_WR_2_port, ADD_WR(1) => 
                           sig_ADD_WR_1_port, ADD_WR(0) => sig_ADD_WR_0_port, 
                           IMM(31) => sig_IMM_31_port, IMM(30) => 
                           sig_IMM_30_port, IMM(29) => sig_IMM_29_port, IMM(28)
                           => sig_IMM_28_port, IMM(27) => sig_IMM_27_port, 
                           IMM(26) => sig_IMM_26_port, IMM(25) => 
                           sig_IMM_25_port, IMM(24) => sig_IMM_24_port, IMM(23)
                           => sig_IMM_23_port, IMM(22) => sig_IMM_22_port, 
                           IMM(21) => sig_IMM_21_port, IMM(20) => 
                           sig_IMM_20_port, IMM(19) => sig_IMM_19_port, IMM(18)
                           => sig_IMM_18_port, IMM(17) => sig_IMM_17_port, 
                           IMM(16) => sig_IMM_16_port, IMM(15) => 
                           sig_IMM_15_port, IMM(14) => sig_IMM_14_port, IMM(13)
                           => sig_IMM_13_port, IMM(12) => sig_IMM_12_port, 
                           IMM(11) => sig_IMM_11_port, IMM(10) => 
                           sig_IMM_10_port, IMM(9) => sig_IMM_9_port, IMM(8) =>
                           sig_IMM_8_port, IMM(7) => sig_IMM_7_port, IMM(6) => 
                           sig_IMM_6_port, IMM(5) => sig_IMM_5_port, IMM(4) => 
                           sig_IMM_4_port, IMM(3) => sig_IMM_3_port, IMM(2) => 
                           sig_IMM_2_port, IMM(1) => sig_IMM_1_port, IMM(0) => 
                           sig_IMM_0_port, RD1 => RD1, RD2 => RD2);
   regPC : regn_N32_7 port map( DIN(31) => PC_IN(31), DIN(30) => PC_IN(30), 
                           DIN(29) => PC_IN(29), DIN(28) => PC_IN(28), DIN(27) 
                           => PC_IN(27), DIN(26) => PC_IN(26), DIN(25) => 
                           PC_IN(25), DIN(24) => PC_IN(24), DIN(23) => 
                           PC_IN(23), DIN(22) => PC_IN(22), DIN(21) => 
                           PC_IN(21), DIN(20) => PC_IN(20), DIN(19) => 
                           PC_IN(19), DIN(18) => PC_IN(18), DIN(17) => 
                           PC_IN(17), DIN(16) => PC_IN(16), DIN(15) => 
                           PC_IN(15), DIN(14) => PC_IN(14), DIN(13) => 
                           PC_IN(13), DIN(12) => PC_IN(12), DIN(11) => 
                           PC_IN(11), DIN(10) => PC_IN(10), DIN(9) => PC_IN(9),
                           DIN(8) => PC_IN(8), DIN(7) => PC_IN(7), DIN(6) => 
                           PC_IN(6), DIN(5) => PC_IN(5), DIN(4) => PC_IN(4), 
                           DIN(3) => PC_IN(3), DIN(2) => PC_IN(2), DIN(1) => 
                           PC_IN(1), DIN(0) => PC_IN(0), CLK => CLK, EN => 
                           X_Logic1_port, RST => sig_RST, DOUT(31) => 
                           PC_OUT(31), DOUT(30) => PC_OUT(30), DOUT(29) => 
                           PC_OUT(29), DOUT(28) => PC_OUT(28), DOUT(27) => 
                           PC_OUT(27), DOUT(26) => PC_OUT(26), DOUT(25) => 
                           PC_OUT(25), DOUT(24) => PC_OUT(24), DOUT(23) => 
                           PC_OUT(23), DOUT(22) => PC_OUT(22), DOUT(21) => 
                           PC_OUT(21), DOUT(20) => PC_OUT(20), DOUT(19) => 
                           PC_OUT(19), DOUT(18) => PC_OUT(18), DOUT(17) => 
                           PC_OUT(17), DOUT(16) => PC_OUT(16), DOUT(15) => 
                           PC_OUT(15), DOUT(14) => PC_OUT(14), DOUT(13) => 
                           PC_OUT(13), DOUT(12) => PC_OUT(12), DOUT(11) => 
                           PC_OUT(11), DOUT(10) => PC_OUT(10), DOUT(9) => 
                           PC_OUT(9), DOUT(8) => PC_OUT(8), DOUT(7) => 
                           PC_OUT(7), DOUT(6) => PC_OUT(6), DOUT(5) => 
                           PC_OUT(5), DOUT(4) => PC_OUT(4), DOUT(3) => 
                           PC_OUT(3), DOUT(2) => PC_OUT(2), DOUT(1) => 
                           PC_OUT(1), DOUT(0) => PC_OUT(0));
   regIMM : regn_N32_6 port map( DIN(31) => sig_IMM_31_port, DIN(30) => 
                           sig_IMM_30_port, DIN(29) => sig_IMM_29_port, DIN(28)
                           => sig_IMM_28_port, DIN(27) => sig_IMM_27_port, 
                           DIN(26) => sig_IMM_26_port, DIN(25) => 
                           sig_IMM_25_port, DIN(24) => sig_IMM_24_port, DIN(23)
                           => sig_IMM_23_port, DIN(22) => sig_IMM_22_port, 
                           DIN(21) => sig_IMM_21_port, DIN(20) => 
                           sig_IMM_20_port, DIN(19) => sig_IMM_19_port, DIN(18)
                           => sig_IMM_18_port, DIN(17) => sig_IMM_17_port, 
                           DIN(16) => sig_IMM_16_port, DIN(15) => 
                           sig_IMM_15_port, DIN(14) => sig_IMM_14_port, DIN(13)
                           => sig_IMM_13_port, DIN(12) => sig_IMM_12_port, 
                           DIN(11) => sig_IMM_11_port, DIN(10) => 
                           sig_IMM_10_port, DIN(9) => sig_IMM_9_port, DIN(8) =>
                           sig_IMM_8_port, DIN(7) => sig_IMM_7_port, DIN(6) => 
                           sig_IMM_6_port, DIN(5) => sig_IMM_5_port, DIN(4) => 
                           sig_IMM_4_port, DIN(3) => sig_IMM_3_port, DIN(2) => 
                           sig_IMM_2_port, DIN(1) => sig_IMM_1_port, DIN(0) => 
                           sig_IMM_0_port, CLK => CLK, EN => X_Logic1_port, RST
                           => sig_RST, DOUT(31) => IMM_OUT(31), DOUT(30) => 
                           IMM_OUT(30), DOUT(29) => IMM_OUT(29), DOUT(28) => 
                           IMM_OUT(28), DOUT(27) => IMM_OUT(27), DOUT(26) => 
                           IMM_OUT(26), DOUT(25) => IMM_OUT(25), DOUT(24) => 
                           IMM_OUT(24), DOUT(23) => IMM_OUT(23), DOUT(22) => 
                           IMM_OUT(22), DOUT(21) => IMM_OUT(21), DOUT(20) => 
                           IMM_OUT(20), DOUT(19) => IMM_OUT(19), DOUT(18) => 
                           IMM_OUT(18), DOUT(17) => IMM_OUT(17), DOUT(16) => 
                           IMM_OUT(16), DOUT(15) => IMM_OUT(15), DOUT(14) => 
                           IMM_OUT(14), DOUT(13) => IMM_OUT(13), DOUT(12) => 
                           IMM_OUT(12), DOUT(11) => IMM_OUT(11), DOUT(10) => 
                           IMM_OUT(10), DOUT(9) => IMM_OUT(9), DOUT(8) => 
                           IMM_OUT(8), DOUT(7) => IMM_OUT(7), DOUT(6) => 
                           IMM_OUT(6), DOUT(5) => IMM_OUT(5), DOUT(4) => 
                           IMM_OUT(4), DOUT(3) => IMM_OUT(3), DOUT(2) => 
                           IMM_OUT(2), DOUT(1) => IMM_OUT(1), DOUT(0) => 
                           IMM_OUT(0));
   regWR : regn_N5_0 port map( DIN(4) => sig_ADD_WRHAZ_4_port, DIN(3) => 
                           sig_ADD_WRHAZ_3_port, DIN(2) => sig_ADD_WRHAZ_2_port
                           , DIN(1) => sig_ADD_WRHAZ_1_port, DIN(0) => 
                           sig_ADD_WRHAZ_0_port, CLK => CLK, EN => 
                           X_Logic1_port, RST => sig_RST, DOUT(4) => 
                           ADD_WR_OUT(4), DOUT(3) => ADD_WR_OUT(3), DOUT(2) => 
                           ADD_WR_OUT(2), DOUT(1) => ADD_WR_OUT(1), DOUT(0) => 
                           ADD_WR_OUT(0));
   regRS1 : regn_N5_4 port map( DIN(4) => sig_ADD_RS1HAZ_4_port, DIN(3) => 
                           sig_ADD_RS1HAZ_3_port, DIN(2) => 
                           sig_ADD_RS1HAZ_2_port, DIN(1) => 
                           sig_ADD_RS1HAZ_1_port, DIN(0) => 
                           sig_ADD_RS1HAZ_0_port, CLK => CLK, EN => 
                           X_Logic1_port, RST => sig_RST, DOUT(4) => 
                           ADD_RS1_OUT(4), DOUT(3) => ADD_RS1_OUT(3), DOUT(2) 
                           => ADD_RS1_OUT(2), DOUT(1) => ADD_RS1_OUT(1), 
                           DOUT(0) => ADD_RS1_OUT(0));
   regRS2 : regn_N5_3 port map( DIN(4) => sig_ADD_RS2HAZ_4_port, DIN(3) => 
                           sig_ADD_RS2HAZ_3_port, DIN(2) => 
                           sig_ADD_RS2HAZ_2_port, DIN(1) => 
                           sig_ADD_RS2HAZ_1_port, DIN(0) => 
                           sig_ADD_RS2HAZ_0_port, CLK => CLK, EN => 
                           X_Logic1_port, RST => sig_RST, DOUT(4) => 
                           ADD_RS2_OUT(4), DOUT(3) => ADD_RS2_OUT(3), DOUT(2) 
                           => ADD_RS2_OUT(2), DOUT(1) => ADD_RS2_OUT(1), 
                           DOUT(0) => ADD_RS2_OUT(0));
   muxRS1 : mux21_NBIT5_0 port map( A(4) => ADD_RS1_HDU_4_port, A(3) => 
                           ADD_RS1_HDU_3_port, A(2) => n10, A(1) => 
                           ADD_RS1_HDU_1_port, A(0) => n4, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, S => Bubble, Z(4) => 
                           sig_ADD_RS1HAZ_4_port, Z(3) => sig_ADD_RS1HAZ_3_port
                           , Z(2) => sig_ADD_RS1HAZ_2_port, Z(1) => 
                           sig_ADD_RS1HAZ_1_port, Z(0) => sig_ADD_RS1HAZ_0_port
                           );
   muxRS2 : mux21_NBIT5_2 port map( A(4) => n3, A(3) => n1, A(2) => n6, A(1) =>
                           n29, A(0) => ADD_RS2_HDU_0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, S => Bubble, Z(4) => 
                           sig_ADD_RS2HAZ_4_port, Z(3) => sig_ADD_RS2HAZ_3_port
                           , Z(2) => sig_ADD_RS2HAZ_2_port, Z(1) => 
                           sig_ADD_RS2HAZ_1_port, Z(0) => sig_ADD_RS2HAZ_0_port
                           );
   muxWR : mux21_NBIT5_1 port map( A(4) => sig_ADD_WR_4_port, A(3) => 
                           sig_ADD_WR_3_port, A(2) => sig_ADD_WR_2_port, A(1) 
                           => sig_ADD_WR_1_port, A(0) => sig_ADD_WR_0_port, 
                           B(4) => X_Logic0_port, B(3) => X_Logic0_port, B(2) 
                           => X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, S => Bubble, Z(4) => 
                           sig_ADD_WRHAZ_4_port, Z(3) => sig_ADD_WRHAZ_3_port, 
                           Z(2) => sig_ADD_WRHAZ_2_port, Z(1) => 
                           sig_ADD_WRHAZ_1_port, Z(0) => sig_ADD_WRHAZ_0_port);
   rf : register_file_NBIT_ADD5_NBIT_DATA32 port map( CLK => CLK, RST => RST, 
                           ENABLE => X_Logic1_port, RD1 => RD1, RD2 => RD2, WR 
                           => RF_WE, ADD_WR(4) => ADD_WR(4), ADD_WR(3) => 
                           ADD_WR(3), ADD_WR(2) => ADD_WR(2), ADD_WR(1) => 
                           ADD_WR(1), ADD_WR(0) => ADD_WR(0), ADD_RS1(4) => n21
                           , ADD_RS1(3) => n22, ADD_RS1(2) => n23, ADD_RS1(1) 
                           => n24, ADD_RS1(0) => n25, ADD_RS2(4) => n19, 
                           ADD_RS2(3) => n18, ADD_RS2(2) => n28, ADD_RS2(1) => 
                           n29, ADD_RS2(0) => n30, DATAIN(31) => DATA_WR_IN(31)
                           , DATAIN(30) => DATA_WR_IN(30), DATAIN(29) => 
                           DATA_WR_IN(29), DATAIN(28) => DATA_WR_IN(28), 
                           DATAIN(27) => DATA_WR_IN(27), DATAIN(26) => 
                           DATA_WR_IN(26), DATAIN(25) => DATA_WR_IN(25), 
                           DATAIN(24) => DATA_WR_IN(24), DATAIN(23) => 
                           DATA_WR_IN(23), DATAIN(22) => DATA_WR_IN(22), 
                           DATAIN(21) => DATA_WR_IN(21), DATAIN(20) => 
                           DATA_WR_IN(20), DATAIN(19) => DATA_WR_IN(19), 
                           DATAIN(18) => DATA_WR_IN(18), DATAIN(17) => 
                           DATA_WR_IN(17), DATAIN(16) => DATA_WR_IN(16), 
                           DATAIN(15) => DATA_WR_IN(15), DATAIN(14) => 
                           DATA_WR_IN(14), DATAIN(13) => DATA_WR_IN(13), 
                           DATAIN(12) => DATA_WR_IN(12), DATAIN(11) => 
                           DATA_WR_IN(11), DATAIN(10) => DATA_WR_IN(10), 
                           DATAIN(9) => DATA_WR_IN(9), DATAIN(8) => 
                           DATA_WR_IN(8), DATAIN(7) => DATA_WR_IN(7), DATAIN(6)
                           => DATA_WR_IN(6), DATAIN(5) => DATA_WR_IN(5), 
                           DATAIN(4) => DATA_WR_IN(4), DATAIN(3) => 
                           DATA_WR_IN(3), DATAIN(2) => DATA_WR_IN(2), DATAIN(1)
                           => DATA_WR_IN(1), DATAIN(0) => DATA_WR_IN(0), 
                           OUT1(31) => A_OUT(31), OUT1(30) => A_OUT(30), 
                           OUT1(29) => A_OUT(29), OUT1(28) => A_OUT(28), 
                           OUT1(27) => A_OUT(27), OUT1(26) => A_OUT(26), 
                           OUT1(25) => A_OUT(25), OUT1(24) => A_OUT(24), 
                           OUT1(23) => A_OUT(23), OUT1(22) => A_OUT(22), 
                           OUT1(21) => A_OUT(21), OUT1(20) => A_OUT(20), 
                           OUT1(19) => A_OUT(19), OUT1(18) => A_OUT(18), 
                           OUT1(17) => A_OUT(17), OUT1(16) => A_OUT(16), 
                           OUT1(15) => A_OUT(15), OUT1(14) => A_OUT(14), 
                           OUT1(13) => A_OUT(13), OUT1(12) => A_OUT(12), 
                           OUT1(11) => A_OUT(11), OUT1(10) => A_OUT(10), 
                           OUT1(9) => A_OUT(9), OUT1(8) => A_OUT(8), OUT1(7) =>
                           A_OUT(7), OUT1(6) => A_OUT(6), OUT1(5) => A_OUT(5), 
                           OUT1(4) => A_OUT(4), OUT1(3) => A_OUT(3), OUT1(2) =>
                           A_OUT(2), OUT1(1) => A_OUT(1), OUT1(0) => A_OUT(0), 
                           OUT2(31) => B_OUT(31), OUT2(30) => B_OUT(30), 
                           OUT2(29) => B_OUT(29), OUT2(28) => B_OUT(28), 
                           OUT2(27) => B_OUT(27), OUT2(26) => B_OUT(26), 
                           OUT2(25) => B_OUT(25), OUT2(24) => B_OUT(24), 
                           OUT2(23) => B_OUT(23), OUT2(22) => B_OUT(22), 
                           OUT2(21) => B_OUT(21), OUT2(20) => B_OUT(20), 
                           OUT2(19) => B_OUT(19), OUT2(18) => B_OUT(18), 
                           OUT2(17) => B_OUT(17), OUT2(16) => B_OUT(16), 
                           OUT2(15) => B_OUT(15), OUT2(14) => B_OUT(14), 
                           OUT2(13) => B_OUT(13), OUT2(12) => B_OUT(12), 
                           OUT2(11) => B_OUT(11), OUT2(10) => B_OUT(10), 
                           OUT2(9) => B_OUT(9), OUT2(8) => B_OUT(8), OUT2(7) =>
                           B_OUT(7), OUT2(6) => B_OUT(6), OUT2(5) => B_OUT(5), 
                           OUT2(4) => B_OUT(4), OUT2(3) => B_OUT(3), OUT2(2) =>
                           B_OUT(2), OUT2(1) => B_OUT(1), OUT2(0) => B_OUT(0));
   U4 : CLKBUF_X1 port map( A => n30, Z => ADD_RS2_HDU_0_port);
   U5 : BUF_X1 port map( A => n22, Z => ADD_RS1_HDU_3_port);
   U6 : CLKBUF_X1 port map( A => INS_IN(27), Z => n12);
   U7 : CLKBUF_X1 port map( A => n18, Z => n1);
   U8 : CLKBUF_X1 port map( A => n24, Z => ADD_RS1_HDU_1_port);
   U9 : CLKBUF_X1 port map( A => n19, Z => n3);
   U10 : BUF_X2 port map( A => n26, Z => n19);
   U11 : CLKBUF_X1 port map( A => n25, Z => n4);
   U12 : CLKBUF_X1 port map( A => n4, Z => ADD_RS1_HDU_0_port);
   U13 : CLKBUF_X1 port map( A => n28, Z => n6);
   U14 : CLKBUF_X1 port map( A => n29, Z => ADD_RS2_HDU_1_port);
   U15 : CLKBUF_X1 port map( A => n1, Z => ADD_RS2_HDU_3_port);
   U16 : CLKBUF_X1 port map( A => n3, Z => ADD_RS2_HDU_4_port);
   U17 : CLKBUF_X1 port map( A => n21, Z => ADD_RS1_HDU_4_port);
   U18 : CLKBUF_X3 port map( A => n27, Z => n18);
   U19 : CLKBUF_X1 port map( A => n23, Z => n10);
   U20 : CLKBUF_X1 port map( A => INS_IN(26), Z => n11);
   U21 : CLKBUF_X1 port map( A => n10, Z => ADD_RS1_HDU_2_port);
   U22 : CLKBUF_X1 port map( A => n6, Z => ADD_RS2_HDU_2_port);
   U23 : INV_X1 port map( A => RST, ZN => n20);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Fetch is

   port( CLK, RST, ZERO_FLAG : in std_logic;  PC_EXT, INS_IN : in 
         std_logic_vector (31 downto 0);  Bubble_in : in std_logic;  HDU_INS_IN
         , HDU_PC_IN, HDU_NPC_IN : in std_logic_vector (31 downto 0);  PC_OUT, 
         ADDR_OUT, NPC_OUT, INS_OUT : out std_logic_vector (31 downto 0));

end Fetch;

architecture SYN_struct of Fetch is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component Fetch_DW01_add_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component regn_N32_8
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_9
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_0
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_6
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, ADDR_OUT_31_port, ADDR_OUT_30_port, ADDR_OUT_29_port, 
      ADDR_OUT_28_port, ADDR_OUT_27_port, ADDR_OUT_26_port, ADDR_OUT_25_port, 
      ADDR_OUT_24_port, ADDR_OUT_23_port, ADDR_OUT_22_port, ADDR_OUT_21_port, 
      ADDR_OUT_20_port, ADDR_OUT_19_port, ADDR_OUT_18_port, ADDR_OUT_17_port, 
      ADDR_OUT_16_port, ADDR_OUT_15_port, ADDR_OUT_14_port, ADDR_OUT_13_port, 
      ADDR_OUT_12_port, ADDR_OUT_11_port, ADDR_OUT_10_port, ADDR_OUT_9_port, 
      ADDR_OUT_8_port, ADDR_OUT_7_port, ADDR_OUT_6_port, ADDR_OUT_5_port, 
      ADDR_OUT_4_port, ADDR_OUT_3_port, ADDR_OUT_2_port, ADDR_OUT_1_port, 
      ADDR_OUT_0_port, sig_RST, sig_NPC_31_port, sig_NPC_30_port, 
      sig_NPC_29_port, sig_NPC_28_port, sig_NPC_27_port, sig_NPC_26_port, 
      sig_NPC_25_port, sig_NPC_24_port, sig_NPC_23_port, sig_NPC_22_port, 
      sig_NPC_21_port, sig_NPC_20_port, sig_NPC_19_port, sig_NPC_18_port, 
      sig_NPC_17_port, sig_NPC_16_port, sig_NPC_15_port, sig_NPC_14_port, 
      sig_NPC_13_port, sig_NPC_12_port, sig_NPC_11_port, sig_NPC_10_port, 
      sig_NPC_9_port, sig_NPC_8_port, sig_NPC_7_port, sig_NPC_6_port, 
      sig_NPC_5_port, sig_NPC_4_port, sig_NPC_3_port, sig_NPC_2_port, 
      sig_NPC_1_port, sig_NPC_0_port, PC_MUX_OUT_31_port, PC_MUX_OUT_30_port, 
      PC_MUX_OUT_29_port, PC_MUX_OUT_28_port, PC_MUX_OUT_27_port, 
      PC_MUX_OUT_26_port, PC_MUX_OUT_25_port, PC_MUX_OUT_24_port, 
      PC_MUX_OUT_23_port, PC_MUX_OUT_22_port, PC_MUX_OUT_21_port, 
      PC_MUX_OUT_20_port, PC_MUX_OUT_19_port, PC_MUX_OUT_18_port, 
      PC_MUX_OUT_17_port, PC_MUX_OUT_16_port, PC_MUX_OUT_15_port, 
      PC_MUX_OUT_14_port, PC_MUX_OUT_13_port, PC_MUX_OUT_12_port, 
      PC_MUX_OUT_11_port, PC_MUX_OUT_10_port, PC_MUX_OUT_9_port, 
      PC_MUX_OUT_8_port, PC_MUX_OUT_7_port, PC_MUX_OUT_6_port, 
      PC_MUX_OUT_5_port, PC_MUX_OUT_4_port, PC_MUX_OUT_3_port, 
      PC_MUX_OUT_2_port, PC_MUX_OUT_1_port, PC_MUX_OUT_0_port, sig_INS_31_port,
      sig_INS_30_port, sig_INS_29_port, sig_INS_28_port, sig_INS_27_port, 
      sig_INS_26_port, sig_INS_25_port, sig_INS_24_port, sig_INS_23_port, 
      sig_INS_22_port, sig_INS_21_port, sig_INS_20_port, sig_INS_19_port, 
      sig_INS_18_port, sig_INS_17_port, sig_INS_16_port, sig_INS_15_port, 
      sig_INS_14_port, sig_INS_13_port, sig_INS_12_port, sig_INS_11_port, 
      sig_INS_10_port, sig_INS_9_port, sig_INS_8_port, sig_INS_7_port, 
      sig_INS_6_port, sig_INS_5_port, sig_INS_4_port, sig_INS_3_port, 
      sig_INS_2_port, sig_INS_1_port, sig_INS_0_port, n1, n2, n3, n4, n_1598 : 
      std_logic;

begin
   ADDR_OUT <= ( ADDR_OUT_31_port, ADDR_OUT_30_port, ADDR_OUT_29_port, 
      ADDR_OUT_28_port, ADDR_OUT_27_port, ADDR_OUT_26_port, ADDR_OUT_25_port, 
      ADDR_OUT_24_port, ADDR_OUT_23_port, ADDR_OUT_22_port, ADDR_OUT_21_port, 
      ADDR_OUT_20_port, ADDR_OUT_19_port, ADDR_OUT_18_port, ADDR_OUT_17_port, 
      ADDR_OUT_16_port, ADDR_OUT_15_port, ADDR_OUT_14_port, ADDR_OUT_13_port, 
      ADDR_OUT_12_port, ADDR_OUT_11_port, ADDR_OUT_10_port, ADDR_OUT_9_port, 
      ADDR_OUT_8_port, ADDR_OUT_7_port, ADDR_OUT_6_port, ADDR_OUT_5_port, 
      ADDR_OUT_4_port, ADDR_OUT_3_port, ADDR_OUT_2_port, ADDR_OUT_1_port, 
      ADDR_OUT_0_port );
   
   X_Logic1_port <= '1';
   n1 <= '0';
   n2 <= '1';
   n3 <= '0';
   NPC_or_NPC_HDU : mux21_NBIT32_0 port map( A(31) => PC_EXT(31), A(30) => 
                           PC_EXT(30), A(29) => PC_EXT(29), A(28) => PC_EXT(28)
                           , A(27) => PC_EXT(27), A(26) => PC_EXT(26), A(25) =>
                           PC_EXT(25), A(24) => PC_EXT(24), A(23) => PC_EXT(23)
                           , A(22) => PC_EXT(22), A(21) => PC_EXT(21), A(20) =>
                           PC_EXT(20), A(19) => PC_EXT(19), A(18) => PC_EXT(18)
                           , A(17) => PC_EXT(17), A(16) => PC_EXT(16), A(15) =>
                           PC_EXT(15), A(14) => PC_EXT(14), A(13) => PC_EXT(13)
                           , A(12) => PC_EXT(12), A(11) => PC_EXT(11), A(10) =>
                           PC_EXT(10), A(9) => PC_EXT(9), A(8) => PC_EXT(8), 
                           A(7) => PC_EXT(7), A(6) => PC_EXT(6), A(5) => 
                           PC_EXT(5), A(4) => PC_EXT(4), A(3) => PC_EXT(3), 
                           A(2) => PC_EXT(2), A(1) => PC_EXT(1), A(0) => 
                           PC_EXT(0), B(31) => HDU_NPC_IN(31), B(30) => 
                           HDU_NPC_IN(30), B(29) => HDU_NPC_IN(29), B(28) => 
                           HDU_NPC_IN(28), B(27) => HDU_NPC_IN(27), B(26) => 
                           HDU_NPC_IN(26), B(25) => HDU_NPC_IN(25), B(24) => 
                           HDU_NPC_IN(24), B(23) => HDU_NPC_IN(23), B(22) => 
                           HDU_NPC_IN(22), B(21) => HDU_NPC_IN(21), B(20) => 
                           HDU_NPC_IN(20), B(19) => HDU_NPC_IN(19), B(18) => 
                           HDU_NPC_IN(18), B(17) => HDU_NPC_IN(17), B(16) => 
                           HDU_NPC_IN(16), B(15) => HDU_NPC_IN(15), B(14) => 
                           HDU_NPC_IN(14), B(13) => HDU_NPC_IN(13), B(12) => 
                           HDU_NPC_IN(12), B(11) => HDU_NPC_IN(11), B(10) => 
                           HDU_NPC_IN(10), B(9) => HDU_NPC_IN(9), B(8) => 
                           HDU_NPC_IN(8), B(7) => HDU_NPC_IN(7), B(6) => 
                           HDU_NPC_IN(6), B(5) => HDU_NPC_IN(5), B(4) => 
                           HDU_NPC_IN(4), B(3) => HDU_NPC_IN(3), B(2) => 
                           HDU_NPC_IN(2), B(1) => HDU_NPC_IN(1), B(0) => 
                           HDU_NPC_IN(0), S => Bubble_in, Z(31) => 
                           sig_NPC_31_port, Z(30) => sig_NPC_30_port, Z(29) => 
                           sig_NPC_29_port, Z(28) => sig_NPC_28_port, Z(27) => 
                           sig_NPC_27_port, Z(26) => sig_NPC_26_port, Z(25) => 
                           sig_NPC_25_port, Z(24) => sig_NPC_24_port, Z(23) => 
                           sig_NPC_23_port, Z(22) => sig_NPC_22_port, Z(21) => 
                           sig_NPC_21_port, Z(20) => sig_NPC_20_port, Z(19) => 
                           sig_NPC_19_port, Z(18) => sig_NPC_18_port, Z(17) => 
                           sig_NPC_17_port, Z(16) => sig_NPC_16_port, Z(15) => 
                           sig_NPC_15_port, Z(14) => sig_NPC_14_port, Z(13) => 
                           sig_NPC_13_port, Z(12) => sig_NPC_12_port, Z(11) => 
                           sig_NPC_11_port, Z(10) => sig_NPC_10_port, Z(9) => 
                           sig_NPC_9_port, Z(8) => sig_NPC_8_port, Z(7) => 
                           sig_NPC_7_port, Z(6) => sig_NPC_6_port, Z(5) => 
                           sig_NPC_5_port, Z(4) => sig_NPC_4_port, Z(3) => 
                           sig_NPC_3_port, Z(2) => sig_NPC_2_port, Z(1) => 
                           sig_NPC_1_port, Z(0) => sig_NPC_0_port);
   PC_or_PC_HDU : mux21_NBIT32_6 port map( A(31) => ADDR_OUT_31_port, A(30) => 
                           ADDR_OUT_30_port, A(29) => ADDR_OUT_29_port, A(28) 
                           => ADDR_OUT_28_port, A(27) => ADDR_OUT_27_port, 
                           A(26) => ADDR_OUT_26_port, A(25) => ADDR_OUT_25_port
                           , A(24) => ADDR_OUT_24_port, A(23) => 
                           ADDR_OUT_23_port, A(22) => ADDR_OUT_22_port, A(21) 
                           => ADDR_OUT_21_port, A(20) => ADDR_OUT_20_port, 
                           A(19) => ADDR_OUT_19_port, A(18) => ADDR_OUT_18_port
                           , A(17) => ADDR_OUT_17_port, A(16) => 
                           ADDR_OUT_16_port, A(15) => ADDR_OUT_15_port, A(14) 
                           => ADDR_OUT_14_port, A(13) => ADDR_OUT_13_port, 
                           A(12) => ADDR_OUT_12_port, A(11) => ADDR_OUT_11_port
                           , A(10) => ADDR_OUT_10_port, A(9) => ADDR_OUT_9_port
                           , A(8) => ADDR_OUT_8_port, A(7) => ADDR_OUT_7_port, 
                           A(6) => ADDR_OUT_6_port, A(5) => ADDR_OUT_5_port, 
                           A(4) => ADDR_OUT_4_port, A(3) => ADDR_OUT_3_port, 
                           A(2) => ADDR_OUT_2_port, A(1) => ADDR_OUT_1_port, 
                           A(0) => ADDR_OUT_0_port, B(31) => HDU_PC_IN(31), 
                           B(30) => HDU_PC_IN(30), B(29) => HDU_PC_IN(29), 
                           B(28) => HDU_PC_IN(28), B(27) => HDU_PC_IN(27), 
                           B(26) => HDU_PC_IN(26), B(25) => HDU_PC_IN(25), 
                           B(24) => HDU_PC_IN(24), B(23) => HDU_PC_IN(23), 
                           B(22) => HDU_PC_IN(22), B(21) => HDU_PC_IN(21), 
                           B(20) => HDU_PC_IN(20), B(19) => HDU_PC_IN(19), 
                           B(18) => HDU_PC_IN(18), B(17) => HDU_PC_IN(17), 
                           B(16) => HDU_PC_IN(16), B(15) => HDU_PC_IN(15), 
                           B(14) => HDU_PC_IN(14), B(13) => HDU_PC_IN(13), 
                           B(12) => HDU_PC_IN(12), B(11) => HDU_PC_IN(11), 
                           B(10) => HDU_PC_IN(10), B(9) => HDU_PC_IN(9), B(8) 
                           => HDU_PC_IN(8), B(7) => HDU_PC_IN(7), B(6) => 
                           HDU_PC_IN(6), B(5) => HDU_PC_IN(5), B(4) => 
                           HDU_PC_IN(4), B(3) => HDU_PC_IN(3), B(2) => 
                           HDU_PC_IN(2), B(1) => HDU_PC_IN(1), B(0) => 
                           HDU_PC_IN(0), S => Bubble_in, Z(31) => 
                           PC_MUX_OUT_31_port, Z(30) => PC_MUX_OUT_30_port, 
                           Z(29) => PC_MUX_OUT_29_port, Z(28) => 
                           PC_MUX_OUT_28_port, Z(27) => PC_MUX_OUT_27_port, 
                           Z(26) => PC_MUX_OUT_26_port, Z(25) => 
                           PC_MUX_OUT_25_port, Z(24) => PC_MUX_OUT_24_port, 
                           Z(23) => PC_MUX_OUT_23_port, Z(22) => 
                           PC_MUX_OUT_22_port, Z(21) => PC_MUX_OUT_21_port, 
                           Z(20) => PC_MUX_OUT_20_port, Z(19) => 
                           PC_MUX_OUT_19_port, Z(18) => PC_MUX_OUT_18_port, 
                           Z(17) => PC_MUX_OUT_17_port, Z(16) => 
                           PC_MUX_OUT_16_port, Z(15) => PC_MUX_OUT_15_port, 
                           Z(14) => PC_MUX_OUT_14_port, Z(13) => 
                           PC_MUX_OUT_13_port, Z(12) => PC_MUX_OUT_12_port, 
                           Z(11) => PC_MUX_OUT_11_port, Z(10) => 
                           PC_MUX_OUT_10_port, Z(9) => PC_MUX_OUT_9_port, Z(8) 
                           => PC_MUX_OUT_8_port, Z(7) => PC_MUX_OUT_7_port, 
                           Z(6) => PC_MUX_OUT_6_port, Z(5) => PC_MUX_OUT_5_port
                           , Z(4) => PC_MUX_OUT_4_port, Z(3) => 
                           PC_MUX_OUT_3_port, Z(2) => PC_MUX_OUT_2_port, Z(1) 
                           => PC_MUX_OUT_1_port, Z(0) => PC_MUX_OUT_0_port);
   INS_or_HDU_INS : mux21_NBIT32_5 port map( A(31) => INS_IN(31), A(30) => 
                           INS_IN(30), A(29) => INS_IN(29), A(28) => INS_IN(28)
                           , A(27) => INS_IN(27), A(26) => INS_IN(26), A(25) =>
                           INS_IN(25), A(24) => INS_IN(24), A(23) => INS_IN(23)
                           , A(22) => INS_IN(22), A(21) => INS_IN(21), A(20) =>
                           INS_IN(20), A(19) => INS_IN(19), A(18) => INS_IN(18)
                           , A(17) => INS_IN(17), A(16) => INS_IN(16), A(15) =>
                           INS_IN(15), A(14) => INS_IN(14), A(13) => INS_IN(13)
                           , A(12) => INS_IN(12), A(11) => INS_IN(11), A(10) =>
                           INS_IN(10), A(9) => INS_IN(9), A(8) => INS_IN(8), 
                           A(7) => INS_IN(7), A(6) => INS_IN(6), A(5) => 
                           INS_IN(5), A(4) => INS_IN(4), A(3) => INS_IN(3), 
                           A(2) => INS_IN(2), A(1) => INS_IN(1), A(0) => 
                           INS_IN(0), B(31) => HDU_INS_IN(31), B(30) => 
                           HDU_INS_IN(30), B(29) => HDU_INS_IN(29), B(28) => 
                           HDU_INS_IN(28), B(27) => HDU_INS_IN(27), B(26) => 
                           HDU_INS_IN(26), B(25) => HDU_INS_IN(25), B(24) => 
                           HDU_INS_IN(24), B(23) => HDU_INS_IN(23), B(22) => 
                           HDU_INS_IN(22), B(21) => HDU_INS_IN(21), B(20) => 
                           HDU_INS_IN(20), B(19) => HDU_INS_IN(19), B(18) => 
                           HDU_INS_IN(18), B(17) => HDU_INS_IN(17), B(16) => 
                           HDU_INS_IN(16), B(15) => HDU_INS_IN(15), B(14) => 
                           HDU_INS_IN(14), B(13) => HDU_INS_IN(13), B(12) => 
                           HDU_INS_IN(12), B(11) => HDU_INS_IN(11), B(10) => 
                           HDU_INS_IN(10), B(9) => HDU_INS_IN(9), B(8) => 
                           HDU_INS_IN(8), B(7) => HDU_INS_IN(7), B(6) => 
                           HDU_INS_IN(6), B(5) => HDU_INS_IN(5), B(4) => 
                           HDU_INS_IN(4), B(3) => HDU_INS_IN(3), B(2) => 
                           HDU_INS_IN(2), B(1) => HDU_INS_IN(1), B(0) => 
                           HDU_INS_IN(0), S => Bubble_in, Z(31) => 
                           sig_INS_31_port, Z(30) => sig_INS_30_port, Z(29) => 
                           sig_INS_29_port, Z(28) => sig_INS_28_port, Z(27) => 
                           sig_INS_27_port, Z(26) => sig_INS_26_port, Z(25) => 
                           sig_INS_25_port, Z(24) => sig_INS_24_port, Z(23) => 
                           sig_INS_23_port, Z(22) => sig_INS_22_port, Z(21) => 
                           sig_INS_21_port, Z(20) => sig_INS_20_port, Z(19) => 
                           sig_INS_19_port, Z(18) => sig_INS_18_port, Z(17) => 
                           sig_INS_17_port, Z(16) => sig_INS_16_port, Z(15) => 
                           sig_INS_15_port, Z(14) => sig_INS_14_port, Z(13) => 
                           sig_INS_13_port, Z(12) => sig_INS_12_port, Z(11) => 
                           sig_INS_11_port, Z(10) => sig_INS_10_port, Z(9) => 
                           sig_INS_9_port, Z(8) => sig_INS_8_port, Z(7) => 
                           sig_INS_7_port, Z(6) => sig_INS_6_port, Z(5) => 
                           sig_INS_5_port, Z(4) => sig_INS_4_port, Z(3) => 
                           sig_INS_3_port, Z(2) => sig_INS_2_port, Z(1) => 
                           sig_INS_1_port, Z(0) => sig_INS_0_port);
   PC : regn_N32_0 port map( DIN(31) => sig_NPC_31_port, DIN(30) => 
                           sig_NPC_30_port, DIN(29) => sig_NPC_29_port, DIN(28)
                           => sig_NPC_28_port, DIN(27) => sig_NPC_27_port, 
                           DIN(26) => sig_NPC_26_port, DIN(25) => 
                           sig_NPC_25_port, DIN(24) => sig_NPC_24_port, DIN(23)
                           => sig_NPC_23_port, DIN(22) => sig_NPC_22_port, 
                           DIN(21) => sig_NPC_21_port, DIN(20) => 
                           sig_NPC_20_port, DIN(19) => sig_NPC_19_port, DIN(18)
                           => sig_NPC_18_port, DIN(17) => sig_NPC_17_port, 
                           DIN(16) => sig_NPC_16_port, DIN(15) => 
                           sig_NPC_15_port, DIN(14) => sig_NPC_14_port, DIN(13)
                           => sig_NPC_13_port, DIN(12) => sig_NPC_12_port, 
                           DIN(11) => sig_NPC_11_port, DIN(10) => 
                           sig_NPC_10_port, DIN(9) => sig_NPC_9_port, DIN(8) =>
                           sig_NPC_8_port, DIN(7) => sig_NPC_7_port, DIN(6) => 
                           sig_NPC_6_port, DIN(5) => sig_NPC_5_port, DIN(4) => 
                           sig_NPC_4_port, DIN(3) => sig_NPC_3_port, DIN(2) => 
                           sig_NPC_2_port, DIN(1) => sig_NPC_1_port, DIN(0) => 
                           sig_NPC_0_port, CLK => CLK, EN => X_Logic1_port, RST
                           => RST, DOUT(31) => ADDR_OUT_31_port, DOUT(30) => 
                           ADDR_OUT_30_port, DOUT(29) => ADDR_OUT_29_port, 
                           DOUT(28) => ADDR_OUT_28_port, DOUT(27) => 
                           ADDR_OUT_27_port, DOUT(26) => ADDR_OUT_26_port, 
                           DOUT(25) => ADDR_OUT_25_port, DOUT(24) => 
                           ADDR_OUT_24_port, DOUT(23) => ADDR_OUT_23_port, 
                           DOUT(22) => ADDR_OUT_22_port, DOUT(21) => 
                           ADDR_OUT_21_port, DOUT(20) => ADDR_OUT_20_port, 
                           DOUT(19) => ADDR_OUT_19_port, DOUT(18) => 
                           ADDR_OUT_18_port, DOUT(17) => ADDR_OUT_17_port, 
                           DOUT(16) => ADDR_OUT_16_port, DOUT(15) => 
                           ADDR_OUT_15_port, DOUT(14) => ADDR_OUT_14_port, 
                           DOUT(13) => ADDR_OUT_13_port, DOUT(12) => 
                           ADDR_OUT_12_port, DOUT(11) => ADDR_OUT_11_port, 
                           DOUT(10) => ADDR_OUT_10_port, DOUT(9) => 
                           ADDR_OUT_9_port, DOUT(8) => ADDR_OUT_8_port, DOUT(7)
                           => ADDR_OUT_7_port, DOUT(6) => ADDR_OUT_6_port, 
                           DOUT(5) => ADDR_OUT_5_port, DOUT(4) => 
                           ADDR_OUT_4_port, DOUT(3) => ADDR_OUT_3_port, DOUT(2)
                           => ADDR_OUT_2_port, DOUT(1) => ADDR_OUT_1_port, 
                           DOUT(0) => ADDR_OUT_0_port);
   PC_reg : regn_N32_9 port map( DIN(31) => PC_MUX_OUT_31_port, DIN(30) => 
                           PC_MUX_OUT_30_port, DIN(29) => PC_MUX_OUT_29_port, 
                           DIN(28) => PC_MUX_OUT_28_port, DIN(27) => 
                           PC_MUX_OUT_27_port, DIN(26) => PC_MUX_OUT_26_port, 
                           DIN(25) => PC_MUX_OUT_25_port, DIN(24) => 
                           PC_MUX_OUT_24_port, DIN(23) => PC_MUX_OUT_23_port, 
                           DIN(22) => PC_MUX_OUT_22_port, DIN(21) => 
                           PC_MUX_OUT_21_port, DIN(20) => PC_MUX_OUT_20_port, 
                           DIN(19) => PC_MUX_OUT_19_port, DIN(18) => 
                           PC_MUX_OUT_18_port, DIN(17) => PC_MUX_OUT_17_port, 
                           DIN(16) => PC_MUX_OUT_16_port, DIN(15) => 
                           PC_MUX_OUT_15_port, DIN(14) => PC_MUX_OUT_14_port, 
                           DIN(13) => PC_MUX_OUT_13_port, DIN(12) => 
                           PC_MUX_OUT_12_port, DIN(11) => PC_MUX_OUT_11_port, 
                           DIN(10) => PC_MUX_OUT_10_port, DIN(9) => 
                           PC_MUX_OUT_9_port, DIN(8) => PC_MUX_OUT_8_port, 
                           DIN(7) => PC_MUX_OUT_7_port, DIN(6) => 
                           PC_MUX_OUT_6_port, DIN(5) => PC_MUX_OUT_5_port, 
                           DIN(4) => PC_MUX_OUT_4_port, DIN(3) => 
                           PC_MUX_OUT_3_port, DIN(2) => PC_MUX_OUT_2_port, 
                           DIN(1) => PC_MUX_OUT_1_port, DIN(0) => 
                           PC_MUX_OUT_0_port, CLK => CLK, EN => X_Logic1_port, 
                           RST => sig_RST, DOUT(31) => PC_OUT(31), DOUT(30) => 
                           PC_OUT(30), DOUT(29) => PC_OUT(29), DOUT(28) => 
                           PC_OUT(28), DOUT(27) => PC_OUT(27), DOUT(26) => 
                           PC_OUT(26), DOUT(25) => PC_OUT(25), DOUT(24) => 
                           PC_OUT(24), DOUT(23) => PC_OUT(23), DOUT(22) => 
                           PC_OUT(22), DOUT(21) => PC_OUT(21), DOUT(20) => 
                           PC_OUT(20), DOUT(19) => PC_OUT(19), DOUT(18) => 
                           PC_OUT(18), DOUT(17) => PC_OUT(17), DOUT(16) => 
                           PC_OUT(16), DOUT(15) => PC_OUT(15), DOUT(14) => 
                           PC_OUT(14), DOUT(13) => PC_OUT(13), DOUT(12) => 
                           PC_OUT(12), DOUT(11) => PC_OUT(11), DOUT(10) => 
                           PC_OUT(10), DOUT(9) => PC_OUT(9), DOUT(8) => 
                           PC_OUT(8), DOUT(7) => PC_OUT(7), DOUT(6) => 
                           PC_OUT(6), DOUT(5) => PC_OUT(5), DOUT(4) => 
                           PC_OUT(4), DOUT(3) => PC_OUT(3), DOUT(2) => 
                           PC_OUT(2), DOUT(1) => PC_OUT(1), DOUT(0) => 
                           PC_OUT(0));
   IR : regn_N32_8 port map( DIN(31) => sig_INS_31_port, DIN(30) => 
                           sig_INS_30_port, DIN(29) => sig_INS_29_port, DIN(28)
                           => sig_INS_28_port, DIN(27) => sig_INS_27_port, 
                           DIN(26) => sig_INS_26_port, DIN(25) => 
                           sig_INS_25_port, DIN(24) => sig_INS_24_port, DIN(23)
                           => sig_INS_23_port, DIN(22) => sig_INS_22_port, 
                           DIN(21) => sig_INS_21_port, DIN(20) => 
                           sig_INS_20_port, DIN(19) => sig_INS_19_port, DIN(18)
                           => sig_INS_18_port, DIN(17) => sig_INS_17_port, 
                           DIN(16) => sig_INS_16_port, DIN(15) => 
                           sig_INS_15_port, DIN(14) => sig_INS_14_port, DIN(13)
                           => sig_INS_13_port, DIN(12) => sig_INS_12_port, 
                           DIN(11) => sig_INS_11_port, DIN(10) => 
                           sig_INS_10_port, DIN(9) => sig_INS_9_port, DIN(8) =>
                           sig_INS_8_port, DIN(7) => sig_INS_7_port, DIN(6) => 
                           sig_INS_6_port, DIN(5) => sig_INS_5_port, DIN(4) => 
                           sig_INS_4_port, DIN(3) => sig_INS_3_port, DIN(2) => 
                           sig_INS_2_port, DIN(1) => sig_INS_1_port, DIN(0) => 
                           sig_INS_0_port, CLK => CLK, EN => X_Logic1_port, RST
                           => sig_RST, DOUT(31) => INS_OUT(31), DOUT(30) => 
                           INS_OUT(30), DOUT(29) => INS_OUT(29), DOUT(28) => 
                           INS_OUT(28), DOUT(27) => INS_OUT(27), DOUT(26) => 
                           INS_OUT(26), DOUT(25) => INS_OUT(25), DOUT(24) => 
                           INS_OUT(24), DOUT(23) => INS_OUT(23), DOUT(22) => 
                           INS_OUT(22), DOUT(21) => INS_OUT(21), DOUT(20) => 
                           INS_OUT(20), DOUT(19) => INS_OUT(19), DOUT(18) => 
                           INS_OUT(18), DOUT(17) => INS_OUT(17), DOUT(16) => 
                           INS_OUT(16), DOUT(15) => INS_OUT(15), DOUT(14) => 
                           INS_OUT(14), DOUT(13) => INS_OUT(13), DOUT(12) => 
                           INS_OUT(12), DOUT(11) => INS_OUT(11), DOUT(10) => 
                           INS_OUT(10), DOUT(9) => INS_OUT(9), DOUT(8) => 
                           INS_OUT(8), DOUT(7) => INS_OUT(7), DOUT(6) => 
                           INS_OUT(6), DOUT(5) => INS_OUT(5), DOUT(4) => 
                           INS_OUT(4), DOUT(3) => INS_OUT(3), DOUT(2) => 
                           INS_OUT(2), DOUT(1) => INS_OUT(1), DOUT(0) => 
                           INS_OUT(0));
   add_54 : Fetch_DW01_add_1 port map( A(31) => ADDR_OUT_31_port, A(30) => 
                           ADDR_OUT_30_port, A(29) => ADDR_OUT_29_port, A(28) 
                           => ADDR_OUT_28_port, A(27) => ADDR_OUT_27_port, 
                           A(26) => ADDR_OUT_26_port, A(25) => ADDR_OUT_25_port
                           , A(24) => ADDR_OUT_24_port, A(23) => 
                           ADDR_OUT_23_port, A(22) => ADDR_OUT_22_port, A(21) 
                           => ADDR_OUT_21_port, A(20) => ADDR_OUT_20_port, 
                           A(19) => ADDR_OUT_19_port, A(18) => ADDR_OUT_18_port
                           , A(17) => ADDR_OUT_17_port, A(16) => 
                           ADDR_OUT_16_port, A(15) => ADDR_OUT_15_port, A(14) 
                           => ADDR_OUT_14_port, A(13) => ADDR_OUT_13_port, 
                           A(12) => ADDR_OUT_12_port, A(11) => ADDR_OUT_11_port
                           , A(10) => ADDR_OUT_10_port, A(9) => ADDR_OUT_9_port
                           , A(8) => ADDR_OUT_8_port, A(7) => ADDR_OUT_7_port, 
                           A(6) => ADDR_OUT_6_port, A(5) => ADDR_OUT_5_port, 
                           A(4) => ADDR_OUT_4_port, A(3) => ADDR_OUT_3_port, 
                           A(2) => ADDR_OUT_2_port, A(1) => ADDR_OUT_1_port, 
                           A(0) => ADDR_OUT_0_port, B(31) => n1, B(30) => n1, 
                           B(29) => n1, B(28) => n1, B(27) => n1, B(26) => n1, 
                           B(25) => n1, B(24) => n1, B(23) => n1, B(22) => n1, 
                           B(21) => n1, B(20) => n1, B(19) => n1, B(18) => n1, 
                           B(17) => n1, B(16) => n1, B(15) => n1, B(14) => n1, 
                           B(13) => n1, B(12) => n1, B(11) => n1, B(10) => n1, 
                           B(9) => n1, B(8) => n1, B(7) => n1, B(6) => n1, B(5)
                           => n1, B(4) => n1, B(3) => n1, B(2) => n2, B(1) => 
                           n1, B(0) => n1, CI => n3, SUM(31) => NPC_OUT(31), 
                           SUM(30) => NPC_OUT(30), SUM(29) => NPC_OUT(29), 
                           SUM(28) => NPC_OUT(28), SUM(27) => NPC_OUT(27), 
                           SUM(26) => NPC_OUT(26), SUM(25) => NPC_OUT(25), 
                           SUM(24) => NPC_OUT(24), SUM(23) => NPC_OUT(23), 
                           SUM(22) => NPC_OUT(22), SUM(21) => NPC_OUT(21), 
                           SUM(20) => NPC_OUT(20), SUM(19) => NPC_OUT(19), 
                           SUM(18) => NPC_OUT(18), SUM(17) => NPC_OUT(17), 
                           SUM(16) => NPC_OUT(16), SUM(15) => NPC_OUT(15), 
                           SUM(14) => NPC_OUT(14), SUM(13) => NPC_OUT(13), 
                           SUM(12) => NPC_OUT(12), SUM(11) => NPC_OUT(11), 
                           SUM(10) => NPC_OUT(10), SUM(9) => NPC_OUT(9), SUM(8)
                           => NPC_OUT(8), SUM(7) => NPC_OUT(7), SUM(6) => 
                           NPC_OUT(6), SUM(5) => NPC_OUT(5), SUM(4) => 
                           NPC_OUT(4), SUM(3) => NPC_OUT(3), SUM(2) => 
                           NPC_OUT(2), SUM(1) => NPC_OUT(1), SUM(0) => 
                           NPC_OUT(0), CO => n_1598);
   U6 : NOR2_X1 port map( A1 => ZERO_FLAG, A2 => n4, ZN => sig_RST);
   U7 : INV_X1 port map( A => RST, ZN => n4);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity hardwired_cu_NBIT32 is

   port( MUX_A_SEL : out std_logic;  MUX_B_SEL : out std_logic_vector (1 downto
         0);  ALU_OPC : out std_logic_vector (0 to 4);  ALU_OUTREG_EN, 
         DRAM_R_IN : out std_logic;  JUMP_TYPE : out std_logic_vector (1 downto
         0);  MEM_EN_IN, DRAM_W_IN, RF_WE : out std_logic;  LOAD_TYPE_IN : out 
         std_logic_vector (1 downto 0);  STORE_TYPE_IN, WB_MUX_SEL : out 
         std_logic;  INS_IN : in std_logic_vector (31 downto 0);  Bubble, Clk, 
         Rst : in std_logic);

end hardwired_cu_NBIT32;

architecture SYN_bhv of hardwired_cu_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal AluOP_E_4_port, AluOP_E_3_port, AluOP_E_2_port, AluOP_E_1_port, 
      AluOP_E_0_port, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, 
      n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n_1599, n_1600, n_1601, n_1602, n_1603 : std_logic;

begin
   
   ALU_OPC_reg_4_inst : DFFR_X1 port map( D => AluOP_E_4_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(0), QN => n_1599);
   ALU_OPC_reg_3_inst : DFFR_X1 port map( D => AluOP_E_3_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(1), QN => n_1600);
   ALU_OPC_reg_2_inst : DFFR_X1 port map( D => AluOP_E_2_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(2), QN => n_1601);
   ALU_OPC_reg_1_inst : DFFR_X1 port map( D => AluOP_E_1_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(3), QN => n_1602);
   WB_MUX_SEL <= '0';
   STORE_TYPE_IN <= '0';
   LOAD_TYPE_IN(0) <= '0';
   LOAD_TYPE_IN(1) <= '0';
   RF_WE <= '0';
   DRAM_W_IN <= '0';
   MEM_EN_IN <= '0';
   JUMP_TYPE(0) <= '0';
   JUMP_TYPE(1) <= '0';
   DRAM_R_IN <= '0';
   ALU_OUTREG_EN <= '0';
   MUX_B_SEL(0) <= '0';
   MUX_B_SEL(1) <= '0';
   MUX_A_SEL <= '0';
   U126 : NAND3_X1 port map( A1 => INS_IN(1), A2 => n25, A3 => INS_IN(0), ZN =>
                           n65);
   U127 : NAND3_X1 port map( A1 => n87, A2 => n64, A3 => n88, ZN => n51);
   U128 : XOR2_X1 port map( A => n28, B => INS_IN(1), Z => n91);
   U129 : NAND3_X1 port map( A1 => n92, A2 => n27, A3 => INS_IN(0), ZN => n37);
   U130 : NAND3_X1 port map( A1 => n10, A2 => n7, A3 => n33, ZN => n103);
   U131 : NAND3_X1 port map( A1 => n28, A2 => n27, A3 => n92, ZN => n39);
   U132 : NAND3_X1 port map( A1 => n110, A2 => n25, A3 => INS_IN(1), ZN => n38)
                           ;
   U133 : NAND3_X1 port map( A1 => n26, A2 => n27, A3 => n53, ZN => n106);
   U134 : NAND3_X1 port map( A1 => INS_IN(1), A2 => n28, A3 => n92, ZN => n43);
   U135 : NAND3_X1 port map( A1 => n23, A2 => n21, A3 => n113, ZN => n112);
   ALU_OPC_reg_0_inst : DFFR_X2 port map( D => AluOP_E_0_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(4), QN => n_1603);
   U17 : INV_X1 port map( A => n77, ZN => n11);
   U18 : INV_X1 port map( A => n79, ZN => n4);
   U19 : INV_X1 port map( A => n59, ZN => n14);
   U20 : NAND2_X1 port map( A1 => n82, A2 => n66, ZN => n73);
   U21 : INV_X1 port map( A => n82, ZN => n5);
   U22 : INV_X1 port map( A => n66, ZN => n2);
   U23 : INV_X1 port map( A => n51, ZN => n17);
   U24 : INV_X1 port map( A => n34, ZN => n13);
   U25 : AOI21_X1 port map( B1 => n44, B2 => n45, A => Bubble, ZN => 
                           AluOP_E_3_port);
   U26 : AOI211_X1 port map( C1 => n14, C2 => n4, A => n54, B => n1, ZN => n44)
                           ;
   U27 : AOI221_X1 port map( B1 => n46, B2 => n34, C1 => n35, C2 => n47, A => 
                           n48, ZN => n45);
   U28 : OAI21_X1 port map( B1 => n49, B2 => n50, A => n17, ZN => n47);
   U29 : AOI21_X1 port map( B1 => n71, B2 => n72, A => Bubble, ZN => 
                           AluOP_E_1_port);
   U30 : AOI221_X1 port map( B1 => n46, B2 => n34, C1 => n14, C2 => n73, A => 
                           n32, ZN => n72);
   U31 : AOI221_X1 port map( B1 => n35, B2 => n76, C1 => n5, C2 => n77, A => 
                           n67, ZN => n71);
   U32 : NAND4_X1 port map( A1 => n43, A2 => n37, A3 => n83, A4 => n84, ZN => 
                           n76);
   U33 : AOI21_X1 port map( B1 => n93, B2 => n94, A => Bubble, ZN => 
                           AluOP_E_0_port);
   U34 : NOR3_X1 port map( A1 => n95, A2 => n6, A3 => n96, ZN => n94);
   U35 : AOI221_X1 port map( B1 => n35, B2 => n104, C1 => n77, C2 => n4, A => 
                           n1, ZN => n93);
   U36 : INV_X1 port map( A => n68, ZN => n6);
   U37 : NOR3_X1 port map( A1 => n33, A2 => n99, A3 => n11, ZN => n81);
   U38 : NAND2_X1 port map( A1 => n52, A2 => n89, ZN => n83);
   U39 : NAND4_X1 port map( A1 => n37, A2 => n38, A3 => n39, A4 => n40, ZN => 
                           n36);
   U40 : AOI21_X1 port map( B1 => n41, B2 => n42, A => n20, ZN => n40);
   U41 : INV_X1 port map( A => n43, ZN => n20);
   U42 : OAI21_X1 port map( B1 => n52, B2 => n41, A => n27, ZN => n90);
   U43 : NAND2_X1 port map( A1 => n70, A2 => n8, ZN => n79);
   U44 : NAND2_X1 port map( A1 => n70, A2 => n9, ZN => n82);
   U45 : OAI21_X1 port map( B1 => n100, B2 => n75, A => n101, ZN => n95);
   U46 : NOR3_X1 port map( A1 => n102, A2 => n4, A3 => n46, ZN => n100);
   U47 : OAI21_X1 port map( B1 => n14, B2 => n57, A => n73, ZN => n101);
   U48 : OAI21_X1 port map( B1 => n3, B2 => n60, A => n103, ZN => n102);
   U49 : AND4_X1 port map( A1 => n70, A2 => n57, A3 => n10, A4 => n7, ZN => n35
                           );
   U50 : NAND2_X1 port map( A1 => n75, A2 => n59, ZN => n34);
   U51 : AOI21_X1 port map( B1 => n55, B2 => n56, A => Bubble, ZN => 
                           AluOP_E_2_port);
   U52 : AOI211_X1 port map( C1 => n5, C2 => n12, A => n67, B => n54, ZN => n55
                           );
   U53 : AOI221_X1 port map( B1 => n2, B2 => n57, C1 => n35, C2 => n16, A => 
                           n58, ZN => n56);
   U54 : NOR3_X1 port map( A1 => n59, A2 => n33, A3 => n60, ZN => n58);
   U55 : INV_X1 port map( A => n60, ZN => n9);
   U56 : NAND2_X1 port map( A1 => n9, A2 => n74, ZN => n66);
   U57 : NAND2_X1 port map( A1 => n89, A2 => n110, ZN => n87);
   U58 : NAND2_X1 port map( A1 => n89, A2 => n41, ZN => n64);
   U59 : INV_X1 port map( A => n75, ZN => n12);
   U60 : AOI21_X1 port map( B1 => n29, B2 => n30, A => Bubble, ZN => 
                           AluOP_E_4_port);
   U61 : AOI211_X1 port map( C1 => n31, C2 => n9, A => n2, B => n32, ZN => n30)
                           ;
   U62 : AOI22_X1 port map( A1 => n35, A2 => n36, B1 => n12, B2 => n4, ZN => 
                           n29);
   U63 : NOR2_X1 port map( A1 => n13, A2 => n33, ZN => n31);
   U64 : OAI221_X1 port map( B1 => n78, B2 => n79, C1 => n66, C2 => n11, A => 
                           n80, ZN => n67);
   U65 : NOR3_X1 port map( A1 => n77, A2 => n57, A3 => n12, ZN => n78);
   U66 : NOR2_X1 port map( A1 => n48, A2 => n81, ZN => n80);
   U67 : AND3_X1 port map( A1 => n8, A2 => n74, A3 => n57, ZN => n32);
   U68 : AND3_X1 port map( A1 => n8, A2 => n74, A3 => n77, ZN => n48);
   U69 : INV_X1 port map( A => n99, ZN => n8);
   U70 : INV_X1 port map( A => n105, ZN => n1);
   U71 : AOI21_X1 port map( B1 => n57, B2 => n46, A => n81, ZN => n105);
   U72 : INV_X1 port map( A => n53, ZN => n19);
   U73 : INV_X1 port map( A => n38, ZN => n18);
   U74 : AND2_X1 port map( A1 => n41, A2 => n25, ZN => n92);
   U75 : INV_X1 port map( A => n50, ZN => n26);
   U76 : NOR3_X1 port map( A1 => n22, A2 => INS_IN(3), A3 => n112, ZN => n52);
   U77 : NOR3_X1 port map( A1 => n22, A2 => n24, A3 => n112, ZN => n41);
   U78 : INV_X1 port map( A => INS_IN(3), ZN => n24);
   U79 : NOR3_X1 port map( A1 => INS_IN(3), A2 => INS_IN(5), A3 => n112, ZN => 
                           n53);
   U80 : NOR3_X1 port map( A1 => n28, A2 => INS_IN(1), A3 => n25, ZN => n89);
   U81 : NOR4_X1 port map( A1 => INS_IN(7), A2 => INS_IN(10), A3 => INS_IN(9), 
                           A4 => INS_IN(8), ZN => n113);
   U82 : AOI221_X1 port map( B1 => n85, B2 => n52, C1 => n26, C2 => n86, A => 
                           n51, ZN => n84);
   U83 : NOR2_X1 port map( A1 => INS_IN(2), A2 => n91, ZN => n85);
   U84 : OAI21_X1 port map( B1 => n27, B2 => n19, A => n90, ZN => n86);
   U85 : NAND4_X1 port map( A1 => n88, A2 => n43, A3 => n106, A4 => n107, ZN =>
                           n104);
   U86 : AOI221_X1 port map( B1 => n108, B2 => n52, C1 => n18, C2 => INS_IN(0),
                           A => n62, ZN => n107);
   U87 : NOR2_X1 port map( A1 => INS_IN(2), A2 => INS_IN(0), ZN => n108);
   U88 : AOI22_X1 port map( A1 => n98, A2 => n77, B1 => n57, B2 => n99, ZN => 
                           n97);
   U89 : OAI21_X1 port map( B1 => INS_IN(1), B2 => n50, A => n65, ZN => n42);
   U90 : NAND4_X1 port map( A1 => n53, A2 => INS_IN(2), A3 => INS_IN(0), A4 => 
                           INS_IN(1), ZN => n88);
   U91 : NAND2_X1 port map( A1 => INS_IN(2), A2 => n28, ZN => n50);
   U92 : INV_X1 port map( A => INS_IN(1), ZN => n27);
   U93 : AOI21_X1 port map( B1 => n52, B2 => INS_IN(1), A => n53, ZN => n49);
   U94 : NAND4_X1 port map( A1 => n109, A2 => n83, A3 => n87, A4 => n39, ZN => 
                           n62);
   U95 : NAND4_X1 port map( A1 => INS_IN(3), A2 => n22, A3 => INS_IN(1), A4 => 
                           n111, ZN => n109);
   U96 : NOR2_X1 port map( A1 => n112, A2 => n50, ZN => n111);
   U97 : INV_X1 port map( A => INS_IN(0), ZN => n28);
   U98 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => n54);
   U99 : INV_X1 port map( A => INS_IN(5), ZN => n22);
   U100 : AND4_X1 port map( A1 => n113, A2 => n21, A3 => INS_IN(3), A4 => n114,
                           ZN => n110);
   U101 : NOR2_X1 port map( A1 => n23, A2 => n22, ZN => n114);
   U102 : INV_X1 port map( A => INS_IN(2), ZN => n25);
   U103 : INV_X1 port map( A => INS_IN(4), ZN => n23);
   U104 : INV_X1 port map( A => INS_IN(6), ZN => n21);
   U105 : INV_X1 port map( A => n61, ZN => n16);
   U106 : AOI211_X1 port map( C1 => n42, C2 => n52, A => n62, B => n63, ZN => 
                           n61);
   U107 : OAI211_X1 port map( C1 => n38, C2 => INS_IN(0), A => n37, B => n64, 
                           ZN => n63);
   U108 : NOR2_X1 port map( A1 => INS_IN(29), A2 => n10, ZN => n98);
   U109 : INV_X1 port map( A => INS_IN(29), ZN => n7);
   U110 : NAND2_X1 port map( A1 => INS_IN(29), A2 => n10, ZN => n60);
   U111 : NOR3_X1 port map( A1 => n3, A2 => INS_IN(30), A3 => n97, ZN => n96);
   U112 : AND2_X1 port map( A1 => INS_IN(30), A2 => n3, ZN => n74);
   U113 : NAND2_X1 port map( A1 => INS_IN(27), A2 => n15, ZN => n59);
   U114 : NOR2_X1 port map( A1 => n15, A2 => INS_IN(27), ZN => n77);
   U115 : NAND4_X1 port map( A1 => n70, A2 => n57, A3 => INS_IN(28), A4 => n7, 
                           ZN => n69);
   U116 : NAND4_X1 port map( A1 => n77, A2 => n70, A3 => INS_IN(28), A4 => n7, 
                           ZN => n68);
   U117 : AND3_X1 port map( A1 => INS_IN(28), A2 => n7, A3 => n74, ZN => n46);
   U118 : NAND2_X1 port map( A1 => INS_IN(29), A2 => INS_IN(28), ZN => n99);
   U119 : INV_X1 port map( A => INS_IN(28), ZN => n10);
   U120 : NOR2_X1 port map( A1 => INS_IN(27), A2 => INS_IN(26), ZN => n57);
   U121 : NAND2_X1 port map( A1 => INS_IN(26), A2 => INS_IN(27), ZN => n75);
   U122 : INV_X1 port map( A => INS_IN(26), ZN => n15);
   U123 : NAND2_X1 port map( A1 => INS_IN(31), A2 => INS_IN(30), ZN => n33);
   U124 : NOR2_X1 port map( A1 => INS_IN(31), A2 => INS_IN(30), ZN => n70);
   U125 : INV_X1 port map( A => INS_IN(31), ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Datapath is

   port( CLK, RST : in std_logic;  INS_IN, DATA_IN : in std_logic_vector (31 
         downto 0);  MUX_A_SEL : in std_logic;  MUX_B_SEL : in std_logic_vector
         (1 downto 0);  ALU_OPC : in std_logic_vector (0 to 4);  ALU_OUTREG_EN 
         : in std_logic;  JUMP_TYPE : in std_logic_vector (1 downto 0);  
         DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, RF_WE : in std_logic;  LOAD_TYPE_IN :
         in std_logic_vector (1 downto 0);  STORE_TYPE_IN, WB_MUX_SEL : in 
         std_logic;  INS_OUT, IRAM_ADDR_OUT, DRAM_ADDR_OUT, DATA_OUT : out 
         std_logic_vector (31 downto 0);  DRAM_R_OUT, DRAM_W_OUT, Bubble_out : 
         out std_logic;  LOAD_TYPE_OUT : out std_logic_vector (1 downto 0);  
         STORE_TYPE_OUT : out std_logic);

end Datapath;

architecture SYN_struct of Datapath is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HazardDetection
      port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : in std_logic_vector
            (4 downto 0);  DRAM_R : in std_logic;  INS_IN, PC_IN : in 
            std_logic_vector (31 downto 0);  Bubble : out std_logic;  
            HDU_INS_OUT, HDU_PC_OUT, HDU_NPC_OUT : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Writeback
      port( WB_MUX_SEL : in std_logic;  DATA_IN, ALU_RES_IN : in 
            std_logic_vector (31 downto 0);  ADD_WR_IN : in std_logic_vector (4
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0);  
            ADD_WR_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component ff_2
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Memory
      port( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN : in std_logic;  PC_SEL :
            in std_logic_vector (1 downto 0);  NPC_IN, NPC_ABS, NPC_REL, 
            ALU_RES_IN, B_IN : in std_logic_vector (31 downto 0);  ADD_WR_IN : 
            in std_logic_vector (4 downto 0);  DRAM_DATA_IN : in 
            std_logic_vector (31 downto 0);  LOAD_TYPE_IN : in std_logic_vector
            (1 downto 0);  STORE_TYPE_IN : in std_logic;  PC_OUT : out 
            std_logic_vector (31 downto 0);  DRAM_R_OUT, DRAM_W_OUT : out 
            std_logic;  DRAM_ADDR_OUT, DRAM_DATA_OUT, DATA_OUT, ALU_RES_OUT, 
            OP_MEM : out std_logic_vector (31 downto 0);  ADD_WR_MEM, 
            ADD_WR_OUT : out std_logic_vector (4 downto 0);  LOAD_TYPE_OUT : 
            out std_logic_vector (1 downto 0);  STORE_TYPE_OUT : out std_logic
            );
   end component;
   
   component ff_0
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Execute
      port( CLK, RST, MUX_A_SEL : in std_logic;  MUX_B_SEL : in 
            std_logic_vector (1 downto 0);  ALU_OPC : in std_logic_vector (0 to
            4);  ALU_OUTREG_EN : in std_logic;  JUMP_TYPE : in std_logic_vector
            (1 downto 0);  PC_IN, A_IN, B_IN, IMM_IN : in std_logic_vector (31 
            downto 0);  ADD_WR_IN, ADD_RS1_IN, ADD_RS2_IN, ADD_WR_MEM, 
            ADD_WR_WB : in std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB 
            : in std_logic;  OP_MEM, OP_WB : in std_logic_vector (31 downto 0);
            PC_SEL : out std_logic_vector (1 downto 0);  ZERO_FLAG : out 
            std_logic;  NPC_ABS, NPC_REL, ALU_RES, B_OUT : out std_logic_vector
            (31 downto 0);  ADD_WR_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component Decode
      port( CLK, RST, Bubble, RF_WE, ZERO_FLAG : in std_logic;  PC_IN, INS_IN :
            in std_logic_vector (31 downto 0);  ADD_WR : in std_logic_vector (4
            downto 0);  DATA_WR_IN : in std_logic_vector (31 downto 0);  PC_OUT
            , A_OUT, B_OUT, IMM_OUT : out std_logic_vector (31 downto 0);  
            ADD_RS1_HDU, ADD_RS2_HDU, ADD_WR_OUT, ADD_RS1_OUT, ADD_RS2_OUT : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component Fetch
      port( CLK, RST, ZERO_FLAG : in std_logic;  PC_EXT, INS_IN : in 
            std_logic_vector (31 downto 0);  Bubble_in : in std_logic;  
            HDU_INS_IN, HDU_PC_IN, HDU_NPC_IN : in std_logic_vector (31 downto 
            0);  PC_OUT, ADDR_OUT, NPC_OUT, INS_OUT : out std_logic_vector (31 
            downto 0));
   end component;
   
   signal X_Logic1_port, n6, INS_OUT_30_port, n7, n8, n9, n10, INS_OUT_25_port,
      INS_OUT_24_port, INS_OUT_23_port, INS_OUT_22_port, INS_OUT_21_port, 
      INS_OUT_20_port, INS_OUT_19_port, INS_OUT_18_port, INS_OUT_17_port, 
      INS_OUT_16_port, INS_OUT_15_port, INS_OUT_14_port, INS_OUT_13_port, 
      INS_OUT_12_port, INS_OUT_11_port, INS_OUT_10_port, INS_OUT_9_port, 
      INS_OUT_8_port, INS_OUT_7_port, INS_OUT_6_port, INS_OUT_5_port, 
      INS_OUT_4_port, INS_OUT_3_port, INS_OUT_2_port, INS_OUT_1_port, 
      INS_OUT_0_port, Bubble_out_port, ZERO_FLAG_EX, PC_MEM_OUT_31_port, 
      PC_MEM_OUT_30_port, PC_MEM_OUT_29_port, PC_MEM_OUT_28_port, 
      PC_MEM_OUT_27_port, PC_MEM_OUT_26_port, PC_MEM_OUT_25_port, 
      PC_MEM_OUT_24_port, PC_MEM_OUT_23_port, PC_MEM_OUT_22_port, 
      PC_MEM_OUT_21_port, PC_MEM_OUT_20_port, PC_MEM_OUT_19_port, 
      PC_MEM_OUT_18_port, PC_MEM_OUT_17_port, PC_MEM_OUT_16_port, 
      PC_MEM_OUT_15_port, PC_MEM_OUT_14_port, PC_MEM_OUT_13_port, 
      PC_MEM_OUT_12_port, PC_MEM_OUT_11_port, PC_MEM_OUT_10_port, 
      PC_MEM_OUT_9_port, PC_MEM_OUT_8_port, PC_MEM_OUT_7_port, 
      PC_MEM_OUT_6_port, PC_MEM_OUT_5_port, PC_MEM_OUT_4_port, 
      PC_MEM_OUT_3_port, PC_MEM_OUT_2_port, PC_MEM_OUT_1_port, 
      PC_MEM_OUT_0_port, sig_HDU_INS_OUT_31_port, sig_HDU_INS_OUT_30_port, 
      sig_HDU_INS_OUT_29_port, sig_HDU_INS_OUT_28_port, sig_HDU_INS_OUT_27_port
      , sig_HDU_INS_OUT_26_port, sig_HDU_INS_OUT_25_port, 
      sig_HDU_INS_OUT_24_port, sig_HDU_INS_OUT_23_port, sig_HDU_INS_OUT_22_port
      , sig_HDU_INS_OUT_21_port, sig_HDU_INS_OUT_20_port, 
      sig_HDU_INS_OUT_19_port, sig_HDU_INS_OUT_18_port, sig_HDU_INS_OUT_17_port
      , sig_HDU_INS_OUT_16_port, sig_HDU_INS_OUT_15_port, 
      sig_HDU_INS_OUT_14_port, sig_HDU_INS_OUT_13_port, sig_HDU_INS_OUT_12_port
      , sig_HDU_INS_OUT_11_port, sig_HDU_INS_OUT_10_port, 
      sig_HDU_INS_OUT_9_port, sig_HDU_INS_OUT_8_port, sig_HDU_INS_OUT_7_port, 
      sig_HDU_INS_OUT_6_port, sig_HDU_INS_OUT_5_port, sig_HDU_INS_OUT_4_port, 
      sig_HDU_INS_OUT_3_port, sig_HDU_INS_OUT_2_port, sig_HDU_INS_OUT_1_port, 
      sig_HDU_INS_OUT_0_port, sig_HDU_PC_OUT_31_port, sig_HDU_PC_OUT_30_port, 
      sig_HDU_PC_OUT_29_port, sig_HDU_PC_OUT_28_port, sig_HDU_PC_OUT_27_port, 
      sig_HDU_PC_OUT_26_port, sig_HDU_PC_OUT_25_port, sig_HDU_PC_OUT_24_port, 
      sig_HDU_PC_OUT_23_port, sig_HDU_PC_OUT_22_port, sig_HDU_PC_OUT_21_port, 
      sig_HDU_PC_OUT_20_port, sig_HDU_PC_OUT_19_port, sig_HDU_PC_OUT_18_port, 
      sig_HDU_PC_OUT_17_port, sig_HDU_PC_OUT_16_port, sig_HDU_PC_OUT_15_port, 
      sig_HDU_PC_OUT_14_port, sig_HDU_PC_OUT_13_port, sig_HDU_PC_OUT_12_port, 
      sig_HDU_PC_OUT_11_port, sig_HDU_PC_OUT_10_port, sig_HDU_PC_OUT_9_port, 
      sig_HDU_PC_OUT_8_port, sig_HDU_PC_OUT_7_port, sig_HDU_PC_OUT_6_port, 
      sig_HDU_PC_OUT_5_port, sig_HDU_PC_OUT_4_port, sig_HDU_PC_OUT_3_port, 
      sig_HDU_PC_OUT_2_port, sig_HDU_PC_OUT_1_port, sig_HDU_PC_OUT_0_port, 
      sig_HDU_NPC_OUT_31_port, sig_HDU_NPC_OUT_30_port, sig_HDU_NPC_OUT_29_port
      , sig_HDU_NPC_OUT_28_port, sig_HDU_NPC_OUT_27_port, 
      sig_HDU_NPC_OUT_26_port, sig_HDU_NPC_OUT_25_port, sig_HDU_NPC_OUT_24_port
      , sig_HDU_NPC_OUT_23_port, sig_HDU_NPC_OUT_22_port, 
      sig_HDU_NPC_OUT_21_port, sig_HDU_NPC_OUT_20_port, sig_HDU_NPC_OUT_19_port
      , sig_HDU_NPC_OUT_18_port, sig_HDU_NPC_OUT_17_port, 
      sig_HDU_NPC_OUT_16_port, sig_HDU_NPC_OUT_15_port, sig_HDU_NPC_OUT_14_port
      , sig_HDU_NPC_OUT_13_port, sig_HDU_NPC_OUT_12_port, 
      sig_HDU_NPC_OUT_11_port, sig_HDU_NPC_OUT_10_port, sig_HDU_NPC_OUT_9_port,
      sig_HDU_NPC_OUT_8_port, sig_HDU_NPC_OUT_7_port, sig_HDU_NPC_OUT_6_port, 
      sig_HDU_NPC_OUT_5_port, sig_HDU_NPC_OUT_4_port, sig_HDU_NPC_OUT_3_port, 
      sig_HDU_NPC_OUT_2_port, sig_HDU_NPC_OUT_1_port, sig_HDU_NPC_OUT_0_port, 
      PC_FETCH_OUT_31_port, PC_FETCH_OUT_30_port, PC_FETCH_OUT_29_port, 
      PC_FETCH_OUT_28_port, PC_FETCH_OUT_27_port, PC_FETCH_OUT_26_port, 
      PC_FETCH_OUT_25_port, PC_FETCH_OUT_24_port, PC_FETCH_OUT_23_port, 
      PC_FETCH_OUT_22_port, PC_FETCH_OUT_21_port, PC_FETCH_OUT_20_port, 
      PC_FETCH_OUT_19_port, PC_FETCH_OUT_18_port, PC_FETCH_OUT_17_port, 
      PC_FETCH_OUT_16_port, PC_FETCH_OUT_15_port, PC_FETCH_OUT_14_port, 
      PC_FETCH_OUT_13_port, PC_FETCH_OUT_12_port, PC_FETCH_OUT_11_port, 
      PC_FETCH_OUT_10_port, PC_FETCH_OUT_9_port, PC_FETCH_OUT_8_port, 
      PC_FETCH_OUT_7_port, PC_FETCH_OUT_6_port, PC_FETCH_OUT_5_port, 
      PC_FETCH_OUT_4_port, PC_FETCH_OUT_3_port, PC_FETCH_OUT_2_port, 
      PC_FETCH_OUT_1_port, PC_FETCH_OUT_0_port, NPC_FETCH_OUT_31_port, 
      NPC_FETCH_OUT_30_port, NPC_FETCH_OUT_29_port, NPC_FETCH_OUT_28_port, 
      NPC_FETCH_OUT_27_port, NPC_FETCH_OUT_26_port, NPC_FETCH_OUT_25_port, 
      NPC_FETCH_OUT_24_port, NPC_FETCH_OUT_23_port, NPC_FETCH_OUT_22_port, 
      NPC_FETCH_OUT_21_port, NPC_FETCH_OUT_20_port, NPC_FETCH_OUT_19_port, 
      NPC_FETCH_OUT_18_port, NPC_FETCH_OUT_17_port, NPC_FETCH_OUT_16_port, 
      NPC_FETCH_OUT_15_port, NPC_FETCH_OUT_14_port, NPC_FETCH_OUT_13_port, 
      NPC_FETCH_OUT_12_port, NPC_FETCH_OUT_11_port, NPC_FETCH_OUT_10_port, 
      NPC_FETCH_OUT_9_port, NPC_FETCH_OUT_8_port, NPC_FETCH_OUT_7_port, 
      NPC_FETCH_OUT_6_port, NPC_FETCH_OUT_5_port, NPC_FETCH_OUT_4_port, 
      NPC_FETCH_OUT_3_port, NPC_FETCH_OUT_2_port, NPC_FETCH_OUT_1_port, 
      NPC_FETCH_OUT_0_port, RF_WE_WB, ADD_WR_WB_4_port, ADD_WR_WB_3_port, 
      ADD_WR_WB_2_port, ADD_WR_WB_1_port, ADD_WR_WB_0_port, OP_WB_31_port, 
      OP_WB_30_port, OP_WB_29_port, OP_WB_28_port, OP_WB_27_port, OP_WB_26_port
      , OP_WB_25_port, OP_WB_24_port, OP_WB_23_port, OP_WB_22_port, 
      OP_WB_21_port, OP_WB_20_port, OP_WB_19_port, OP_WB_18_port, OP_WB_17_port
      , OP_WB_16_port, OP_WB_15_port, OP_WB_14_port, OP_WB_13_port, 
      OP_WB_12_port, OP_WB_11_port, OP_WB_10_port, OP_WB_9_port, OP_WB_8_port, 
      OP_WB_7_port, OP_WB_6_port, OP_WB_5_port, OP_WB_4_port, OP_WB_3_port, 
      OP_WB_2_port, OP_WB_1_port, OP_WB_0_port, PC_DECODE_OUT_31_port, 
      PC_DECODE_OUT_30_port, PC_DECODE_OUT_29_port, PC_DECODE_OUT_28_port, 
      PC_DECODE_OUT_27_port, PC_DECODE_OUT_26_port, PC_DECODE_OUT_25_port, 
      PC_DECODE_OUT_24_port, PC_DECODE_OUT_23_port, PC_DECODE_OUT_22_port, 
      PC_DECODE_OUT_21_port, PC_DECODE_OUT_20_port, PC_DECODE_OUT_19_port, 
      PC_DECODE_OUT_18_port, PC_DECODE_OUT_17_port, PC_DECODE_OUT_16_port, 
      PC_DECODE_OUT_15_port, PC_DECODE_OUT_14_port, PC_DECODE_OUT_13_port, 
      PC_DECODE_OUT_12_port, PC_DECODE_OUT_11_port, PC_DECODE_OUT_10_port, 
      PC_DECODE_OUT_9_port, PC_DECODE_OUT_8_port, PC_DECODE_OUT_7_port, 
      PC_DECODE_OUT_6_port, PC_DECODE_OUT_5_port, PC_DECODE_OUT_4_port, 
      PC_DECODE_OUT_3_port, PC_DECODE_OUT_2_port, PC_DECODE_OUT_1_port, 
      PC_DECODE_OUT_0_port, A_DECODE_OUT_31_port, A_DECODE_OUT_30_port, 
      A_DECODE_OUT_29_port, A_DECODE_OUT_28_port, A_DECODE_OUT_27_port, 
      A_DECODE_OUT_26_port, A_DECODE_OUT_25_port, A_DECODE_OUT_24_port, 
      A_DECODE_OUT_23_port, A_DECODE_OUT_22_port, A_DECODE_OUT_21_port, 
      A_DECODE_OUT_20_port, A_DECODE_OUT_19_port, A_DECODE_OUT_18_port, 
      A_DECODE_OUT_17_port, A_DECODE_OUT_16_port, A_DECODE_OUT_15_port, 
      A_DECODE_OUT_14_port, A_DECODE_OUT_13_port, A_DECODE_OUT_12_port, 
      A_DECODE_OUT_11_port, A_DECODE_OUT_10_port, A_DECODE_OUT_9_port, 
      A_DECODE_OUT_8_port, A_DECODE_OUT_7_port, A_DECODE_OUT_6_port, 
      A_DECODE_OUT_5_port, A_DECODE_OUT_4_port, A_DECODE_OUT_3_port, 
      A_DECODE_OUT_2_port, A_DECODE_OUT_1_port, A_DECODE_OUT_0_port, 
      B_DECODE_OUT_31_port, B_DECODE_OUT_30_port, B_DECODE_OUT_29_port, 
      B_DECODE_OUT_28_port, B_DECODE_OUT_27_port, B_DECODE_OUT_26_port, 
      B_DECODE_OUT_25_port, B_DECODE_OUT_24_port, B_DECODE_OUT_23_port, 
      B_DECODE_OUT_22_port, B_DECODE_OUT_21_port, B_DECODE_OUT_20_port, 
      B_DECODE_OUT_19_port, B_DECODE_OUT_18_port, B_DECODE_OUT_17_port, 
      B_DECODE_OUT_16_port, B_DECODE_OUT_15_port, B_DECODE_OUT_14_port, 
      B_DECODE_OUT_13_port, B_DECODE_OUT_12_port, B_DECODE_OUT_11_port, 
      B_DECODE_OUT_10_port, B_DECODE_OUT_9_port, B_DECODE_OUT_8_port, 
      B_DECODE_OUT_7_port, B_DECODE_OUT_6_port, B_DECODE_OUT_5_port, 
      B_DECODE_OUT_4_port, B_DECODE_OUT_3_port, B_DECODE_OUT_2_port, 
      B_DECODE_OUT_1_port, B_DECODE_OUT_0_port, IMM_DECODE_OUT_31_port, 
      IMM_DECODE_OUT_30_port, IMM_DECODE_OUT_29_port, IMM_DECODE_OUT_28_port, 
      IMM_DECODE_OUT_27_port, IMM_DECODE_OUT_26_port, IMM_DECODE_OUT_25_port, 
      IMM_DECODE_OUT_24_port, IMM_DECODE_OUT_23_port, IMM_DECODE_OUT_22_port, 
      IMM_DECODE_OUT_21_port, IMM_DECODE_OUT_20_port, IMM_DECODE_OUT_19_port, 
      IMM_DECODE_OUT_18_port, IMM_DECODE_OUT_17_port, IMM_DECODE_OUT_16_port, 
      IMM_DECODE_OUT_15_port, IMM_DECODE_OUT_14_port, IMM_DECODE_OUT_13_port, 
      IMM_DECODE_OUT_12_port, IMM_DECODE_OUT_11_port, IMM_DECODE_OUT_10_port, 
      IMM_DECODE_OUT_9_port, IMM_DECODE_OUT_8_port, IMM_DECODE_OUT_7_port, 
      IMM_DECODE_OUT_6_port, IMM_DECODE_OUT_5_port, IMM_DECODE_OUT_4_port, 
      IMM_DECODE_OUT_3_port, IMM_DECODE_OUT_2_port, IMM_DECODE_OUT_1_port, 
      IMM_DECODE_OUT_0_port, ADD_RS1_HDU_4_port, ADD_RS1_HDU_3_port, 
      ADD_RS1_HDU_2_port, ADD_RS1_HDU_1_port, ADD_RS1_HDU_0_port, 
      ADD_RS2_HDU_4_port, ADD_RS2_HDU_3_port, ADD_RS2_HDU_2_port, 
      ADD_RS2_HDU_1_port, ADD_RS2_HDU_0_port, ADD_WR_DECODE_OUT_4_port, 
      ADD_WR_DECODE_OUT_3_port, ADD_WR_DECODE_OUT_2_port, 
      ADD_WR_DECODE_OUT_1_port, ADD_WR_DECODE_OUT_0_port, 
      ADD_RS1_DECODE_OUT_4_port, ADD_RS1_DECODE_OUT_3_port, 
      ADD_RS1_DECODE_OUT_2_port, ADD_RS1_DECODE_OUT_1_port, 
      ADD_RS1_DECODE_OUT_0_port, ADD_RS2_DECODE_OUT_4_port, 
      ADD_RS2_DECODE_OUT_3_port, ADD_RS2_DECODE_OUT_2_port, 
      ADD_RS2_DECODE_OUT_1_port, ADD_RS2_DECODE_OUT_0_port, ADD_WR_MEM_4_port, 
      ADD_WR_MEM_3_port, ADD_WR_MEM_2_port, ADD_WR_MEM_1_port, 
      ADD_WR_MEM_0_port, OP_MEM_31_port, OP_MEM_30_port, OP_MEM_29_port, 
      OP_MEM_28_port, OP_MEM_27_port, OP_MEM_26_port, OP_MEM_25_port, 
      OP_MEM_24_port, OP_MEM_23_port, OP_MEM_22_port, OP_MEM_21_port, 
      OP_MEM_20_port, OP_MEM_19_port, OP_MEM_18_port, OP_MEM_17_port, 
      OP_MEM_16_port, OP_MEM_15_port, OP_MEM_14_port, OP_MEM_13_port, 
      OP_MEM_12_port, OP_MEM_11_port, OP_MEM_10_port, OP_MEM_9_port, 
      OP_MEM_8_port, OP_MEM_7_port, OP_MEM_6_port, OP_MEM_5_port, OP_MEM_4_port
      , OP_MEM_3_port, OP_MEM_2_port, OP_MEM_1_port, OP_MEM_0_port, 
      PC_SEL_EX_1_port, PC_SEL_EX_0_port, NPC_ABS_EX_31_port, 
      NPC_ABS_EX_30_port, NPC_ABS_EX_29_port, NPC_ABS_EX_28_port, 
      NPC_ABS_EX_27_port, NPC_ABS_EX_26_port, NPC_ABS_EX_25_port, 
      NPC_ABS_EX_24_port, NPC_ABS_EX_23_port, NPC_ABS_EX_22_port, 
      NPC_ABS_EX_21_port, NPC_ABS_EX_20_port, NPC_ABS_EX_19_port, 
      NPC_ABS_EX_18_port, NPC_ABS_EX_17_port, NPC_ABS_EX_16_port, 
      NPC_ABS_EX_15_port, NPC_ABS_EX_14_port, NPC_ABS_EX_13_port, 
      NPC_ABS_EX_12_port, NPC_ABS_EX_11_port, NPC_ABS_EX_10_port, 
      NPC_ABS_EX_9_port, NPC_ABS_EX_8_port, NPC_ABS_EX_7_port, 
      NPC_ABS_EX_6_port, NPC_ABS_EX_5_port, NPC_ABS_EX_4_port, 
      NPC_ABS_EX_3_port, NPC_ABS_EX_2_port, NPC_ABS_EX_1_port, 
      NPC_ABS_EX_0_port, NPC_REL_EX_31_port, NPC_REL_EX_30_port, 
      NPC_REL_EX_29_port, NPC_REL_EX_28_port, NPC_REL_EX_27_port, 
      NPC_REL_EX_26_port, NPC_REL_EX_25_port, NPC_REL_EX_24_port, 
      NPC_REL_EX_23_port, NPC_REL_EX_22_port, NPC_REL_EX_21_port, 
      NPC_REL_EX_20_port, NPC_REL_EX_19_port, NPC_REL_EX_18_port, 
      NPC_REL_EX_17_port, NPC_REL_EX_16_port, NPC_REL_EX_15_port, 
      NPC_REL_EX_14_port, NPC_REL_EX_13_port, NPC_REL_EX_12_port, 
      NPC_REL_EX_11_port, NPC_REL_EX_10_port, NPC_REL_EX_9_port, 
      NPC_REL_EX_8_port, NPC_REL_EX_7_port, NPC_REL_EX_6_port, 
      NPC_REL_EX_5_port, NPC_REL_EX_4_port, NPC_REL_EX_3_port, 
      NPC_REL_EX_2_port, NPC_REL_EX_1_port, NPC_REL_EX_0_port, 
      ALU_RES_EX_31_port, ALU_RES_EX_30_port, ALU_RES_EX_29_port, 
      ALU_RES_EX_28_port, ALU_RES_EX_27_port, ALU_RES_EX_26_port, 
      ALU_RES_EX_25_port, ALU_RES_EX_24_port, ALU_RES_EX_23_port, 
      ALU_RES_EX_22_port, ALU_RES_EX_21_port, ALU_RES_EX_20_port, 
      ALU_RES_EX_19_port, ALU_RES_EX_18_port, ALU_RES_EX_17_port, 
      ALU_RES_EX_16_port, ALU_RES_EX_15_port, ALU_RES_EX_14_port, 
      ALU_RES_EX_13_port, ALU_RES_EX_12_port, ALU_RES_EX_11_port, 
      ALU_RES_EX_10_port, ALU_RES_EX_9_port, ALU_RES_EX_8_port, 
      ALU_RES_EX_7_port, ALU_RES_EX_6_port, ALU_RES_EX_5_port, 
      ALU_RES_EX_4_port, ALU_RES_EX_3_port, ALU_RES_EX_2_port, 
      ALU_RES_EX_1_port, ALU_RES_EX_0_port, B_EX_OUT_31_port, B_EX_OUT_30_port,
      B_EX_OUT_29_port, B_EX_OUT_28_port, B_EX_OUT_27_port, B_EX_OUT_26_port, 
      B_EX_OUT_25_port, B_EX_OUT_24_port, B_EX_OUT_23_port, B_EX_OUT_22_port, 
      B_EX_OUT_21_port, B_EX_OUT_20_port, B_EX_OUT_19_port, B_EX_OUT_18_port, 
      B_EX_OUT_17_port, B_EX_OUT_16_port, B_EX_OUT_15_port, B_EX_OUT_14_port, 
      B_EX_OUT_13_port, B_EX_OUT_12_port, B_EX_OUT_11_port, B_EX_OUT_10_port, 
      B_EX_OUT_9_port, B_EX_OUT_8_port, B_EX_OUT_7_port, B_EX_OUT_6_port, 
      B_EX_OUT_5_port, B_EX_OUT_4_port, B_EX_OUT_3_port, B_EX_OUT_2_port, 
      B_EX_OUT_1_port, B_EX_OUT_0_port, ADD_WR_EX_OUT_4_port, 
      ADD_WR_EX_OUT_3_port, ADD_WR_EX_OUT_2_port, ADD_WR_EX_OUT_1_port, 
      ADD_WR_EX_OUT_0_port, DRAM_R_MEM, DATA_MEM_OUT_31_port, 
      DATA_MEM_OUT_30_port, DATA_MEM_OUT_29_port, DATA_MEM_OUT_28_port, 
      DATA_MEM_OUT_27_port, DATA_MEM_OUT_26_port, DATA_MEM_OUT_25_port, 
      DATA_MEM_OUT_24_port, DATA_MEM_OUT_23_port, DATA_MEM_OUT_22_port, 
      DATA_MEM_OUT_21_port, DATA_MEM_OUT_20_port, DATA_MEM_OUT_19_port, 
      DATA_MEM_OUT_18_port, DATA_MEM_OUT_17_port, DATA_MEM_OUT_16_port, 
      DATA_MEM_OUT_15_port, DATA_MEM_OUT_14_port, DATA_MEM_OUT_13_port, 
      DATA_MEM_OUT_12_port, DATA_MEM_OUT_11_port, DATA_MEM_OUT_10_port, 
      DATA_MEM_OUT_9_port, DATA_MEM_OUT_8_port, DATA_MEM_OUT_7_port, 
      DATA_MEM_OUT_6_port, DATA_MEM_OUT_5_port, DATA_MEM_OUT_4_port, 
      DATA_MEM_OUT_3_port, DATA_MEM_OUT_2_port, DATA_MEM_OUT_1_port, 
      DATA_MEM_OUT_0_port, ALU_RES_MEM_31_port, ALU_RES_MEM_30_port, 
      ALU_RES_MEM_29_port, ALU_RES_MEM_28_port, ALU_RES_MEM_27_port, 
      ALU_RES_MEM_26_port, ALU_RES_MEM_25_port, ALU_RES_MEM_24_port, 
      ALU_RES_MEM_23_port, ALU_RES_MEM_22_port, ALU_RES_MEM_21_port, 
      ALU_RES_MEM_20_port, ALU_RES_MEM_19_port, ALU_RES_MEM_18_port, 
      ALU_RES_MEM_17_port, ALU_RES_MEM_16_port, ALU_RES_MEM_15_port, 
      ALU_RES_MEM_14_port, ALU_RES_MEM_13_port, ALU_RES_MEM_12_port, 
      ALU_RES_MEM_11_port, ALU_RES_MEM_10_port, ALU_RES_MEM_9_port, 
      ALU_RES_MEM_8_port, ALU_RES_MEM_7_port, ALU_RES_MEM_6_port, 
      ALU_RES_MEM_5_port, ALU_RES_MEM_4_port, ALU_RES_MEM_3_port, 
      ALU_RES_MEM_2_port, ALU_RES_MEM_1_port, ALU_RES_MEM_0_port, 
      ADD_WR_MEM_OUT_4_port, ADD_WR_MEM_OUT_3_port, ADD_WR_MEM_OUT_2_port, 
      ADD_WR_MEM_OUT_1_port, ADD_WR_MEM_OUT_0_port, INS_OUT_29_port, 
      INS_OUT_28_port, INS_OUT_26_port, INS_OUT_31_port, INS_OUT_27_port : 
      std_logic;

begin
   INS_OUT <= ( INS_OUT_31_port, INS_OUT_30_port, INS_OUT_29_port, 
      INS_OUT_28_port, INS_OUT_27_port, INS_OUT_26_port, INS_OUT_25_port, 
      INS_OUT_24_port, INS_OUT_23_port, INS_OUT_22_port, INS_OUT_21_port, 
      INS_OUT_20_port, INS_OUT_19_port, INS_OUT_18_port, INS_OUT_17_port, 
      INS_OUT_16_port, INS_OUT_15_port, INS_OUT_14_port, INS_OUT_13_port, 
      INS_OUT_12_port, INS_OUT_11_port, INS_OUT_10_port, INS_OUT_9_port, 
      INS_OUT_8_port, INS_OUT_7_port, INS_OUT_6_port, INS_OUT_5_port, 
      INS_OUT_4_port, INS_OUT_3_port, INS_OUT_2_port, INS_OUT_1_port, 
      INS_OUT_0_port );
   Bubble_out <= Bubble_out_port;
   
   X_Logic1_port <= '1';
   FetchStage : Fetch port map( CLK => CLK, RST => RST, ZERO_FLAG => 
                           ZERO_FLAG_EX, PC_EXT(31) => PC_MEM_OUT_31_port, 
                           PC_EXT(30) => PC_MEM_OUT_30_port, PC_EXT(29) => 
                           PC_MEM_OUT_29_port, PC_EXT(28) => PC_MEM_OUT_28_port
                           , PC_EXT(27) => PC_MEM_OUT_27_port, PC_EXT(26) => 
                           PC_MEM_OUT_26_port, PC_EXT(25) => PC_MEM_OUT_25_port
                           , PC_EXT(24) => PC_MEM_OUT_24_port, PC_EXT(23) => 
                           PC_MEM_OUT_23_port, PC_EXT(22) => PC_MEM_OUT_22_port
                           , PC_EXT(21) => PC_MEM_OUT_21_port, PC_EXT(20) => 
                           PC_MEM_OUT_20_port, PC_EXT(19) => PC_MEM_OUT_19_port
                           , PC_EXT(18) => PC_MEM_OUT_18_port, PC_EXT(17) => 
                           PC_MEM_OUT_17_port, PC_EXT(16) => PC_MEM_OUT_16_port
                           , PC_EXT(15) => PC_MEM_OUT_15_port, PC_EXT(14) => 
                           PC_MEM_OUT_14_port, PC_EXT(13) => PC_MEM_OUT_13_port
                           , PC_EXT(12) => PC_MEM_OUT_12_port, PC_EXT(11) => 
                           PC_MEM_OUT_11_port, PC_EXT(10) => PC_MEM_OUT_10_port
                           , PC_EXT(9) => PC_MEM_OUT_9_port, PC_EXT(8) => 
                           PC_MEM_OUT_8_port, PC_EXT(7) => PC_MEM_OUT_7_port, 
                           PC_EXT(6) => PC_MEM_OUT_6_port, PC_EXT(5) => 
                           PC_MEM_OUT_5_port, PC_EXT(4) => PC_MEM_OUT_4_port, 
                           PC_EXT(3) => PC_MEM_OUT_3_port, PC_EXT(2) => 
                           PC_MEM_OUT_2_port, PC_EXT(1) => PC_MEM_OUT_1_port, 
                           PC_EXT(0) => PC_MEM_OUT_0_port, INS_IN(31) => 
                           INS_IN(31), INS_IN(30) => INS_IN(30), INS_IN(29) => 
                           INS_IN(29), INS_IN(28) => INS_IN(28), INS_IN(27) => 
                           INS_IN(27), INS_IN(26) => INS_IN(26), INS_IN(25) => 
                           INS_IN(25), INS_IN(24) => INS_IN(24), INS_IN(23) => 
                           INS_IN(23), INS_IN(22) => INS_IN(22), INS_IN(21) => 
                           INS_IN(21), INS_IN(20) => INS_IN(20), INS_IN(19) => 
                           INS_IN(19), INS_IN(18) => INS_IN(18), INS_IN(17) => 
                           INS_IN(17), INS_IN(16) => INS_IN(16), INS_IN(15) => 
                           INS_IN(15), INS_IN(14) => INS_IN(14), INS_IN(13) => 
                           INS_IN(13), INS_IN(12) => INS_IN(12), INS_IN(11) => 
                           INS_IN(11), INS_IN(10) => INS_IN(10), INS_IN(9) => 
                           INS_IN(9), INS_IN(8) => INS_IN(8), INS_IN(7) => 
                           INS_IN(7), INS_IN(6) => INS_IN(6), INS_IN(5) => 
                           INS_IN(5), INS_IN(4) => INS_IN(4), INS_IN(3) => 
                           INS_IN(3), INS_IN(2) => INS_IN(2), INS_IN(1) => 
                           INS_IN(1), INS_IN(0) => INS_IN(0), Bubble_in => 
                           Bubble_out_port, HDU_INS_IN(31) => 
                           sig_HDU_INS_OUT_31_port, HDU_INS_IN(30) => 
                           sig_HDU_INS_OUT_30_port, HDU_INS_IN(29) => 
                           sig_HDU_INS_OUT_29_port, HDU_INS_IN(28) => 
                           sig_HDU_INS_OUT_28_port, HDU_INS_IN(27) => 
                           sig_HDU_INS_OUT_27_port, HDU_INS_IN(26) => 
                           sig_HDU_INS_OUT_26_port, HDU_INS_IN(25) => 
                           sig_HDU_INS_OUT_25_port, HDU_INS_IN(24) => 
                           sig_HDU_INS_OUT_24_port, HDU_INS_IN(23) => 
                           sig_HDU_INS_OUT_23_port, HDU_INS_IN(22) => 
                           sig_HDU_INS_OUT_22_port, HDU_INS_IN(21) => 
                           sig_HDU_INS_OUT_21_port, HDU_INS_IN(20) => 
                           sig_HDU_INS_OUT_20_port, HDU_INS_IN(19) => 
                           sig_HDU_INS_OUT_19_port, HDU_INS_IN(18) => 
                           sig_HDU_INS_OUT_18_port, HDU_INS_IN(17) => 
                           sig_HDU_INS_OUT_17_port, HDU_INS_IN(16) => 
                           sig_HDU_INS_OUT_16_port, HDU_INS_IN(15) => 
                           sig_HDU_INS_OUT_15_port, HDU_INS_IN(14) => 
                           sig_HDU_INS_OUT_14_port, HDU_INS_IN(13) => 
                           sig_HDU_INS_OUT_13_port, HDU_INS_IN(12) => 
                           sig_HDU_INS_OUT_12_port, HDU_INS_IN(11) => 
                           sig_HDU_INS_OUT_11_port, HDU_INS_IN(10) => 
                           sig_HDU_INS_OUT_10_port, HDU_INS_IN(9) => 
                           sig_HDU_INS_OUT_9_port, HDU_INS_IN(8) => 
                           sig_HDU_INS_OUT_8_port, HDU_INS_IN(7) => 
                           sig_HDU_INS_OUT_7_port, HDU_INS_IN(6) => 
                           sig_HDU_INS_OUT_6_port, HDU_INS_IN(5) => 
                           sig_HDU_INS_OUT_5_port, HDU_INS_IN(4) => 
                           sig_HDU_INS_OUT_4_port, HDU_INS_IN(3) => 
                           sig_HDU_INS_OUT_3_port, HDU_INS_IN(2) => 
                           sig_HDU_INS_OUT_2_port, HDU_INS_IN(1) => 
                           sig_HDU_INS_OUT_1_port, HDU_INS_IN(0) => 
                           sig_HDU_INS_OUT_0_port, HDU_PC_IN(31) => 
                           sig_HDU_PC_OUT_31_port, HDU_PC_IN(30) => 
                           sig_HDU_PC_OUT_30_port, HDU_PC_IN(29) => 
                           sig_HDU_PC_OUT_29_port, HDU_PC_IN(28) => 
                           sig_HDU_PC_OUT_28_port, HDU_PC_IN(27) => 
                           sig_HDU_PC_OUT_27_port, HDU_PC_IN(26) => 
                           sig_HDU_PC_OUT_26_port, HDU_PC_IN(25) => 
                           sig_HDU_PC_OUT_25_port, HDU_PC_IN(24) => 
                           sig_HDU_PC_OUT_24_port, HDU_PC_IN(23) => 
                           sig_HDU_PC_OUT_23_port, HDU_PC_IN(22) => 
                           sig_HDU_PC_OUT_22_port, HDU_PC_IN(21) => 
                           sig_HDU_PC_OUT_21_port, HDU_PC_IN(20) => 
                           sig_HDU_PC_OUT_20_port, HDU_PC_IN(19) => 
                           sig_HDU_PC_OUT_19_port, HDU_PC_IN(18) => 
                           sig_HDU_PC_OUT_18_port, HDU_PC_IN(17) => 
                           sig_HDU_PC_OUT_17_port, HDU_PC_IN(16) => 
                           sig_HDU_PC_OUT_16_port, HDU_PC_IN(15) => 
                           sig_HDU_PC_OUT_15_port, HDU_PC_IN(14) => 
                           sig_HDU_PC_OUT_14_port, HDU_PC_IN(13) => 
                           sig_HDU_PC_OUT_13_port, HDU_PC_IN(12) => 
                           sig_HDU_PC_OUT_12_port, HDU_PC_IN(11) => 
                           sig_HDU_PC_OUT_11_port, HDU_PC_IN(10) => 
                           sig_HDU_PC_OUT_10_port, HDU_PC_IN(9) => 
                           sig_HDU_PC_OUT_9_port, HDU_PC_IN(8) => 
                           sig_HDU_PC_OUT_8_port, HDU_PC_IN(7) => 
                           sig_HDU_PC_OUT_7_port, HDU_PC_IN(6) => 
                           sig_HDU_PC_OUT_6_port, HDU_PC_IN(5) => 
                           sig_HDU_PC_OUT_5_port, HDU_PC_IN(4) => 
                           sig_HDU_PC_OUT_4_port, HDU_PC_IN(3) => 
                           sig_HDU_PC_OUT_3_port, HDU_PC_IN(2) => 
                           sig_HDU_PC_OUT_2_port, HDU_PC_IN(1) => 
                           sig_HDU_PC_OUT_1_port, HDU_PC_IN(0) => 
                           sig_HDU_PC_OUT_0_port, HDU_NPC_IN(31) => 
                           sig_HDU_NPC_OUT_31_port, HDU_NPC_IN(30) => 
                           sig_HDU_NPC_OUT_30_port, HDU_NPC_IN(29) => 
                           sig_HDU_NPC_OUT_29_port, HDU_NPC_IN(28) => 
                           sig_HDU_NPC_OUT_28_port, HDU_NPC_IN(27) => 
                           sig_HDU_NPC_OUT_27_port, HDU_NPC_IN(26) => 
                           sig_HDU_NPC_OUT_26_port, HDU_NPC_IN(25) => 
                           sig_HDU_NPC_OUT_25_port, HDU_NPC_IN(24) => 
                           sig_HDU_NPC_OUT_24_port, HDU_NPC_IN(23) => 
                           sig_HDU_NPC_OUT_23_port, HDU_NPC_IN(22) => 
                           sig_HDU_NPC_OUT_22_port, HDU_NPC_IN(21) => 
                           sig_HDU_NPC_OUT_21_port, HDU_NPC_IN(20) => 
                           sig_HDU_NPC_OUT_20_port, HDU_NPC_IN(19) => 
                           sig_HDU_NPC_OUT_19_port, HDU_NPC_IN(18) => 
                           sig_HDU_NPC_OUT_18_port, HDU_NPC_IN(17) => 
                           sig_HDU_NPC_OUT_17_port, HDU_NPC_IN(16) => 
                           sig_HDU_NPC_OUT_16_port, HDU_NPC_IN(15) => 
                           sig_HDU_NPC_OUT_15_port, HDU_NPC_IN(14) => 
                           sig_HDU_NPC_OUT_14_port, HDU_NPC_IN(13) => 
                           sig_HDU_NPC_OUT_13_port, HDU_NPC_IN(12) => 
                           sig_HDU_NPC_OUT_12_port, HDU_NPC_IN(11) => 
                           sig_HDU_NPC_OUT_11_port, HDU_NPC_IN(10) => 
                           sig_HDU_NPC_OUT_10_port, HDU_NPC_IN(9) => 
                           sig_HDU_NPC_OUT_9_port, HDU_NPC_IN(8) => 
                           sig_HDU_NPC_OUT_8_port, HDU_NPC_IN(7) => 
                           sig_HDU_NPC_OUT_7_port, HDU_NPC_IN(6) => 
                           sig_HDU_NPC_OUT_6_port, HDU_NPC_IN(5) => 
                           sig_HDU_NPC_OUT_5_port, HDU_NPC_IN(4) => 
                           sig_HDU_NPC_OUT_4_port, HDU_NPC_IN(3) => 
                           sig_HDU_NPC_OUT_3_port, HDU_NPC_IN(2) => 
                           sig_HDU_NPC_OUT_2_port, HDU_NPC_IN(1) => 
                           sig_HDU_NPC_OUT_1_port, HDU_NPC_IN(0) => 
                           sig_HDU_NPC_OUT_0_port, PC_OUT(31) => 
                           PC_FETCH_OUT_31_port, PC_OUT(30) => 
                           PC_FETCH_OUT_30_port, PC_OUT(29) => 
                           PC_FETCH_OUT_29_port, PC_OUT(28) => 
                           PC_FETCH_OUT_28_port, PC_OUT(27) => 
                           PC_FETCH_OUT_27_port, PC_OUT(26) => 
                           PC_FETCH_OUT_26_port, PC_OUT(25) => 
                           PC_FETCH_OUT_25_port, PC_OUT(24) => 
                           PC_FETCH_OUT_24_port, PC_OUT(23) => 
                           PC_FETCH_OUT_23_port, PC_OUT(22) => 
                           PC_FETCH_OUT_22_port, PC_OUT(21) => 
                           PC_FETCH_OUT_21_port, PC_OUT(20) => 
                           PC_FETCH_OUT_20_port, PC_OUT(19) => 
                           PC_FETCH_OUT_19_port, PC_OUT(18) => 
                           PC_FETCH_OUT_18_port, PC_OUT(17) => 
                           PC_FETCH_OUT_17_port, PC_OUT(16) => 
                           PC_FETCH_OUT_16_port, PC_OUT(15) => 
                           PC_FETCH_OUT_15_port, PC_OUT(14) => 
                           PC_FETCH_OUT_14_port, PC_OUT(13) => 
                           PC_FETCH_OUT_13_port, PC_OUT(12) => 
                           PC_FETCH_OUT_12_port, PC_OUT(11) => 
                           PC_FETCH_OUT_11_port, PC_OUT(10) => 
                           PC_FETCH_OUT_10_port, PC_OUT(9) => 
                           PC_FETCH_OUT_9_port, PC_OUT(8) => 
                           PC_FETCH_OUT_8_port, PC_OUT(7) => 
                           PC_FETCH_OUT_7_port, PC_OUT(6) => 
                           PC_FETCH_OUT_6_port, PC_OUT(5) => 
                           PC_FETCH_OUT_5_port, PC_OUT(4) => 
                           PC_FETCH_OUT_4_port, PC_OUT(3) => 
                           PC_FETCH_OUT_3_port, PC_OUT(2) => 
                           PC_FETCH_OUT_2_port, PC_OUT(1) => 
                           PC_FETCH_OUT_1_port, PC_OUT(0) => 
                           PC_FETCH_OUT_0_port, ADDR_OUT(31) => 
                           IRAM_ADDR_OUT(31), ADDR_OUT(30) => IRAM_ADDR_OUT(30)
                           , ADDR_OUT(29) => IRAM_ADDR_OUT(29), ADDR_OUT(28) =>
                           IRAM_ADDR_OUT(28), ADDR_OUT(27) => IRAM_ADDR_OUT(27)
                           , ADDR_OUT(26) => IRAM_ADDR_OUT(26), ADDR_OUT(25) =>
                           IRAM_ADDR_OUT(25), ADDR_OUT(24) => IRAM_ADDR_OUT(24)
                           , ADDR_OUT(23) => IRAM_ADDR_OUT(23), ADDR_OUT(22) =>
                           IRAM_ADDR_OUT(22), ADDR_OUT(21) => IRAM_ADDR_OUT(21)
                           , ADDR_OUT(20) => IRAM_ADDR_OUT(20), ADDR_OUT(19) =>
                           IRAM_ADDR_OUT(19), ADDR_OUT(18) => IRAM_ADDR_OUT(18)
                           , ADDR_OUT(17) => IRAM_ADDR_OUT(17), ADDR_OUT(16) =>
                           IRAM_ADDR_OUT(16), ADDR_OUT(15) => IRAM_ADDR_OUT(15)
                           , ADDR_OUT(14) => IRAM_ADDR_OUT(14), ADDR_OUT(13) =>
                           IRAM_ADDR_OUT(13), ADDR_OUT(12) => IRAM_ADDR_OUT(12)
                           , ADDR_OUT(11) => IRAM_ADDR_OUT(11), ADDR_OUT(10) =>
                           IRAM_ADDR_OUT(10), ADDR_OUT(9) => IRAM_ADDR_OUT(9), 
                           ADDR_OUT(8) => IRAM_ADDR_OUT(8), ADDR_OUT(7) => 
                           IRAM_ADDR_OUT(7), ADDR_OUT(6) => IRAM_ADDR_OUT(6), 
                           ADDR_OUT(5) => IRAM_ADDR_OUT(5), ADDR_OUT(4) => 
                           IRAM_ADDR_OUT(4), ADDR_OUT(3) => IRAM_ADDR_OUT(3), 
                           ADDR_OUT(2) => IRAM_ADDR_OUT(2), ADDR_OUT(1) => 
                           IRAM_ADDR_OUT(1), ADDR_OUT(0) => IRAM_ADDR_OUT(0), 
                           NPC_OUT(31) => NPC_FETCH_OUT_31_port, NPC_OUT(30) =>
                           NPC_FETCH_OUT_30_port, NPC_OUT(29) => 
                           NPC_FETCH_OUT_29_port, NPC_OUT(28) => 
                           NPC_FETCH_OUT_28_port, NPC_OUT(27) => 
                           NPC_FETCH_OUT_27_port, NPC_OUT(26) => 
                           NPC_FETCH_OUT_26_port, NPC_OUT(25) => 
                           NPC_FETCH_OUT_25_port, NPC_OUT(24) => 
                           NPC_FETCH_OUT_24_port, NPC_OUT(23) => 
                           NPC_FETCH_OUT_23_port, NPC_OUT(22) => 
                           NPC_FETCH_OUT_22_port, NPC_OUT(21) => 
                           NPC_FETCH_OUT_21_port, NPC_OUT(20) => 
                           NPC_FETCH_OUT_20_port, NPC_OUT(19) => 
                           NPC_FETCH_OUT_19_port, NPC_OUT(18) => 
                           NPC_FETCH_OUT_18_port, NPC_OUT(17) => 
                           NPC_FETCH_OUT_17_port, NPC_OUT(16) => 
                           NPC_FETCH_OUT_16_port, NPC_OUT(15) => 
                           NPC_FETCH_OUT_15_port, NPC_OUT(14) => 
                           NPC_FETCH_OUT_14_port, NPC_OUT(13) => 
                           NPC_FETCH_OUT_13_port, NPC_OUT(12) => 
                           NPC_FETCH_OUT_12_port, NPC_OUT(11) => 
                           NPC_FETCH_OUT_11_port, NPC_OUT(10) => 
                           NPC_FETCH_OUT_10_port, NPC_OUT(9) => 
                           NPC_FETCH_OUT_9_port, NPC_OUT(8) => 
                           NPC_FETCH_OUT_8_port, NPC_OUT(7) => 
                           NPC_FETCH_OUT_7_port, NPC_OUT(6) => 
                           NPC_FETCH_OUT_6_port, NPC_OUT(5) => 
                           NPC_FETCH_OUT_5_port, NPC_OUT(4) => 
                           NPC_FETCH_OUT_4_port, NPC_OUT(3) => 
                           NPC_FETCH_OUT_3_port, NPC_OUT(2) => 
                           NPC_FETCH_OUT_2_port, NPC_OUT(1) => 
                           NPC_FETCH_OUT_1_port, NPC_OUT(0) => 
                           NPC_FETCH_OUT_0_port, INS_OUT(31) => n6, INS_OUT(30)
                           => INS_OUT_30_port, INS_OUT(29) => n7, INS_OUT(28) 
                           => n8, INS_OUT(27) => n9, INS_OUT(26) => n10, 
                           INS_OUT(25) => INS_OUT_25_port, INS_OUT(24) => 
                           INS_OUT_24_port, INS_OUT(23) => INS_OUT_23_port, 
                           INS_OUT(22) => INS_OUT_22_port, INS_OUT(21) => 
                           INS_OUT_21_port, INS_OUT(20) => INS_OUT_20_port, 
                           INS_OUT(19) => INS_OUT_19_port, INS_OUT(18) => 
                           INS_OUT_18_port, INS_OUT(17) => INS_OUT_17_port, 
                           INS_OUT(16) => INS_OUT_16_port, INS_OUT(15) => 
                           INS_OUT_15_port, INS_OUT(14) => INS_OUT_14_port, 
                           INS_OUT(13) => INS_OUT_13_port, INS_OUT(12) => 
                           INS_OUT_12_port, INS_OUT(11) => INS_OUT_11_port, 
                           INS_OUT(10) => INS_OUT_10_port, INS_OUT(9) => 
                           INS_OUT_9_port, INS_OUT(8) => INS_OUT_8_port, 
                           INS_OUT(7) => INS_OUT_7_port, INS_OUT(6) => 
                           INS_OUT_6_port, INS_OUT(5) => INS_OUT_5_port, 
                           INS_OUT(4) => INS_OUT_4_port, INS_OUT(3) => 
                           INS_OUT_3_port, INS_OUT(2) => INS_OUT_2_port, 
                           INS_OUT(1) => INS_OUT_1_port, INS_OUT(0) => 
                           INS_OUT_0_port);
   DecodeStage : Decode port map( CLK => CLK, RST => RST, Bubble => 
                           Bubble_out_port, RF_WE => RF_WE_WB, ZERO_FLAG => 
                           ZERO_FLAG_EX, PC_IN(31) => PC_FETCH_OUT_31_port, 
                           PC_IN(30) => PC_FETCH_OUT_30_port, PC_IN(29) => 
                           PC_FETCH_OUT_29_port, PC_IN(28) => 
                           PC_FETCH_OUT_28_port, PC_IN(27) => 
                           PC_FETCH_OUT_27_port, PC_IN(26) => 
                           PC_FETCH_OUT_26_port, PC_IN(25) => 
                           PC_FETCH_OUT_25_port, PC_IN(24) => 
                           PC_FETCH_OUT_24_port, PC_IN(23) => 
                           PC_FETCH_OUT_23_port, PC_IN(22) => 
                           PC_FETCH_OUT_22_port, PC_IN(21) => 
                           PC_FETCH_OUT_21_port, PC_IN(20) => 
                           PC_FETCH_OUT_20_port, PC_IN(19) => 
                           PC_FETCH_OUT_19_port, PC_IN(18) => 
                           PC_FETCH_OUT_18_port, PC_IN(17) => 
                           PC_FETCH_OUT_17_port, PC_IN(16) => 
                           PC_FETCH_OUT_16_port, PC_IN(15) => 
                           PC_FETCH_OUT_15_port, PC_IN(14) => 
                           PC_FETCH_OUT_14_port, PC_IN(13) => 
                           PC_FETCH_OUT_13_port, PC_IN(12) => 
                           PC_FETCH_OUT_12_port, PC_IN(11) => 
                           PC_FETCH_OUT_11_port, PC_IN(10) => 
                           PC_FETCH_OUT_10_port, PC_IN(9) => 
                           PC_FETCH_OUT_9_port, PC_IN(8) => PC_FETCH_OUT_8_port
                           , PC_IN(7) => PC_FETCH_OUT_7_port, PC_IN(6) => 
                           PC_FETCH_OUT_6_port, PC_IN(5) => PC_FETCH_OUT_5_port
                           , PC_IN(4) => PC_FETCH_OUT_4_port, PC_IN(3) => 
                           PC_FETCH_OUT_3_port, PC_IN(2) => PC_FETCH_OUT_2_port
                           , PC_IN(1) => PC_FETCH_OUT_1_port, PC_IN(0) => 
                           PC_FETCH_OUT_0_port, INS_IN(31) => n6, INS_IN(30) =>
                           INS_OUT_30_port, INS_IN(29) => n7, INS_IN(28) => n8,
                           INS_IN(27) => n9, INS_IN(26) => n10, INS_IN(25) => 
                           INS_OUT_25_port, INS_IN(24) => INS_OUT_24_port, 
                           INS_IN(23) => INS_OUT_23_port, INS_IN(22) => 
                           INS_OUT_22_port, INS_IN(21) => INS_OUT_21_port, 
                           INS_IN(20) => INS_OUT_20_port, INS_IN(19) => 
                           INS_OUT_19_port, INS_IN(18) => INS_OUT_18_port, 
                           INS_IN(17) => INS_OUT_17_port, INS_IN(16) => 
                           INS_OUT_16_port, INS_IN(15) => INS_OUT_15_port, 
                           INS_IN(14) => INS_OUT_14_port, INS_IN(13) => 
                           INS_OUT_13_port, INS_IN(12) => INS_OUT_12_port, 
                           INS_IN(11) => INS_OUT_11_port, INS_IN(10) => 
                           INS_OUT_10_port, INS_IN(9) => INS_OUT_9_port, 
                           INS_IN(8) => INS_OUT_8_port, INS_IN(7) => 
                           INS_OUT_7_port, INS_IN(6) => INS_OUT_6_port, 
                           INS_IN(5) => INS_OUT_5_port, INS_IN(4) => 
                           INS_OUT_4_port, INS_IN(3) => INS_OUT_3_port, 
                           INS_IN(2) => INS_OUT_2_port, INS_IN(1) => 
                           INS_OUT_1_port, INS_IN(0) => INS_OUT_0_port, 
                           ADD_WR(4) => ADD_WR_WB_4_port, ADD_WR(3) => 
                           ADD_WR_WB_3_port, ADD_WR(2) => ADD_WR_WB_2_port, 
                           ADD_WR(1) => ADD_WR_WB_1_port, ADD_WR(0) => 
                           ADD_WR_WB_0_port, DATA_WR_IN(31) => OP_WB_31_port, 
                           DATA_WR_IN(30) => OP_WB_30_port, DATA_WR_IN(29) => 
                           OP_WB_29_port, DATA_WR_IN(28) => OP_WB_28_port, 
                           DATA_WR_IN(27) => OP_WB_27_port, DATA_WR_IN(26) => 
                           OP_WB_26_port, DATA_WR_IN(25) => OP_WB_25_port, 
                           DATA_WR_IN(24) => OP_WB_24_port, DATA_WR_IN(23) => 
                           OP_WB_23_port, DATA_WR_IN(22) => OP_WB_22_port, 
                           DATA_WR_IN(21) => OP_WB_21_port, DATA_WR_IN(20) => 
                           OP_WB_20_port, DATA_WR_IN(19) => OP_WB_19_port, 
                           DATA_WR_IN(18) => OP_WB_18_port, DATA_WR_IN(17) => 
                           OP_WB_17_port, DATA_WR_IN(16) => OP_WB_16_port, 
                           DATA_WR_IN(15) => OP_WB_15_port, DATA_WR_IN(14) => 
                           OP_WB_14_port, DATA_WR_IN(13) => OP_WB_13_port, 
                           DATA_WR_IN(12) => OP_WB_12_port, DATA_WR_IN(11) => 
                           OP_WB_11_port, DATA_WR_IN(10) => OP_WB_10_port, 
                           DATA_WR_IN(9) => OP_WB_9_port, DATA_WR_IN(8) => 
                           OP_WB_8_port, DATA_WR_IN(7) => OP_WB_7_port, 
                           DATA_WR_IN(6) => OP_WB_6_port, DATA_WR_IN(5) => 
                           OP_WB_5_port, DATA_WR_IN(4) => OP_WB_4_port, 
                           DATA_WR_IN(3) => OP_WB_3_port, DATA_WR_IN(2) => 
                           OP_WB_2_port, DATA_WR_IN(1) => OP_WB_1_port, 
                           DATA_WR_IN(0) => OP_WB_0_port, PC_OUT(31) => 
                           PC_DECODE_OUT_31_port, PC_OUT(30) => 
                           PC_DECODE_OUT_30_port, PC_OUT(29) => 
                           PC_DECODE_OUT_29_port, PC_OUT(28) => 
                           PC_DECODE_OUT_28_port, PC_OUT(27) => 
                           PC_DECODE_OUT_27_port, PC_OUT(26) => 
                           PC_DECODE_OUT_26_port, PC_OUT(25) => 
                           PC_DECODE_OUT_25_port, PC_OUT(24) => 
                           PC_DECODE_OUT_24_port, PC_OUT(23) => 
                           PC_DECODE_OUT_23_port, PC_OUT(22) => 
                           PC_DECODE_OUT_22_port, PC_OUT(21) => 
                           PC_DECODE_OUT_21_port, PC_OUT(20) => 
                           PC_DECODE_OUT_20_port, PC_OUT(19) => 
                           PC_DECODE_OUT_19_port, PC_OUT(18) => 
                           PC_DECODE_OUT_18_port, PC_OUT(17) => 
                           PC_DECODE_OUT_17_port, PC_OUT(16) => 
                           PC_DECODE_OUT_16_port, PC_OUT(15) => 
                           PC_DECODE_OUT_15_port, PC_OUT(14) => 
                           PC_DECODE_OUT_14_port, PC_OUT(13) => 
                           PC_DECODE_OUT_13_port, PC_OUT(12) => 
                           PC_DECODE_OUT_12_port, PC_OUT(11) => 
                           PC_DECODE_OUT_11_port, PC_OUT(10) => 
                           PC_DECODE_OUT_10_port, PC_OUT(9) => 
                           PC_DECODE_OUT_9_port, PC_OUT(8) => 
                           PC_DECODE_OUT_8_port, PC_OUT(7) => 
                           PC_DECODE_OUT_7_port, PC_OUT(6) => 
                           PC_DECODE_OUT_6_port, PC_OUT(5) => 
                           PC_DECODE_OUT_5_port, PC_OUT(4) => 
                           PC_DECODE_OUT_4_port, PC_OUT(3) => 
                           PC_DECODE_OUT_3_port, PC_OUT(2) => 
                           PC_DECODE_OUT_2_port, PC_OUT(1) => 
                           PC_DECODE_OUT_1_port, PC_OUT(0) => 
                           PC_DECODE_OUT_0_port, A_OUT(31) => 
                           A_DECODE_OUT_31_port, A_OUT(30) => 
                           A_DECODE_OUT_30_port, A_OUT(29) => 
                           A_DECODE_OUT_29_port, A_OUT(28) => 
                           A_DECODE_OUT_28_port, A_OUT(27) => 
                           A_DECODE_OUT_27_port, A_OUT(26) => 
                           A_DECODE_OUT_26_port, A_OUT(25) => 
                           A_DECODE_OUT_25_port, A_OUT(24) => 
                           A_DECODE_OUT_24_port, A_OUT(23) => 
                           A_DECODE_OUT_23_port, A_OUT(22) => 
                           A_DECODE_OUT_22_port, A_OUT(21) => 
                           A_DECODE_OUT_21_port, A_OUT(20) => 
                           A_DECODE_OUT_20_port, A_OUT(19) => 
                           A_DECODE_OUT_19_port, A_OUT(18) => 
                           A_DECODE_OUT_18_port, A_OUT(17) => 
                           A_DECODE_OUT_17_port, A_OUT(16) => 
                           A_DECODE_OUT_16_port, A_OUT(15) => 
                           A_DECODE_OUT_15_port, A_OUT(14) => 
                           A_DECODE_OUT_14_port, A_OUT(13) => 
                           A_DECODE_OUT_13_port, A_OUT(12) => 
                           A_DECODE_OUT_12_port, A_OUT(11) => 
                           A_DECODE_OUT_11_port, A_OUT(10) => 
                           A_DECODE_OUT_10_port, A_OUT(9) => 
                           A_DECODE_OUT_9_port, A_OUT(8) => A_DECODE_OUT_8_port
                           , A_OUT(7) => A_DECODE_OUT_7_port, A_OUT(6) => 
                           A_DECODE_OUT_6_port, A_OUT(5) => A_DECODE_OUT_5_port
                           , A_OUT(4) => A_DECODE_OUT_4_port, A_OUT(3) => 
                           A_DECODE_OUT_3_port, A_OUT(2) => A_DECODE_OUT_2_port
                           , A_OUT(1) => A_DECODE_OUT_1_port, A_OUT(0) => 
                           A_DECODE_OUT_0_port, B_OUT(31) => 
                           B_DECODE_OUT_31_port, B_OUT(30) => 
                           B_DECODE_OUT_30_port, B_OUT(29) => 
                           B_DECODE_OUT_29_port, B_OUT(28) => 
                           B_DECODE_OUT_28_port, B_OUT(27) => 
                           B_DECODE_OUT_27_port, B_OUT(26) => 
                           B_DECODE_OUT_26_port, B_OUT(25) => 
                           B_DECODE_OUT_25_port, B_OUT(24) => 
                           B_DECODE_OUT_24_port, B_OUT(23) => 
                           B_DECODE_OUT_23_port, B_OUT(22) => 
                           B_DECODE_OUT_22_port, B_OUT(21) => 
                           B_DECODE_OUT_21_port, B_OUT(20) => 
                           B_DECODE_OUT_20_port, B_OUT(19) => 
                           B_DECODE_OUT_19_port, B_OUT(18) => 
                           B_DECODE_OUT_18_port, B_OUT(17) => 
                           B_DECODE_OUT_17_port, B_OUT(16) => 
                           B_DECODE_OUT_16_port, B_OUT(15) => 
                           B_DECODE_OUT_15_port, B_OUT(14) => 
                           B_DECODE_OUT_14_port, B_OUT(13) => 
                           B_DECODE_OUT_13_port, B_OUT(12) => 
                           B_DECODE_OUT_12_port, B_OUT(11) => 
                           B_DECODE_OUT_11_port, B_OUT(10) => 
                           B_DECODE_OUT_10_port, B_OUT(9) => 
                           B_DECODE_OUT_9_port, B_OUT(8) => B_DECODE_OUT_8_port
                           , B_OUT(7) => B_DECODE_OUT_7_port, B_OUT(6) => 
                           B_DECODE_OUT_6_port, B_OUT(5) => B_DECODE_OUT_5_port
                           , B_OUT(4) => B_DECODE_OUT_4_port, B_OUT(3) => 
                           B_DECODE_OUT_3_port, B_OUT(2) => B_DECODE_OUT_2_port
                           , B_OUT(1) => B_DECODE_OUT_1_port, B_OUT(0) => 
                           B_DECODE_OUT_0_port, IMM_OUT(31) => 
                           IMM_DECODE_OUT_31_port, IMM_OUT(30) => 
                           IMM_DECODE_OUT_30_port, IMM_OUT(29) => 
                           IMM_DECODE_OUT_29_port, IMM_OUT(28) => 
                           IMM_DECODE_OUT_28_port, IMM_OUT(27) => 
                           IMM_DECODE_OUT_27_port, IMM_OUT(26) => 
                           IMM_DECODE_OUT_26_port, IMM_OUT(25) => 
                           IMM_DECODE_OUT_25_port, IMM_OUT(24) => 
                           IMM_DECODE_OUT_24_port, IMM_OUT(23) => 
                           IMM_DECODE_OUT_23_port, IMM_OUT(22) => 
                           IMM_DECODE_OUT_22_port, IMM_OUT(21) => 
                           IMM_DECODE_OUT_21_port, IMM_OUT(20) => 
                           IMM_DECODE_OUT_20_port, IMM_OUT(19) => 
                           IMM_DECODE_OUT_19_port, IMM_OUT(18) => 
                           IMM_DECODE_OUT_18_port, IMM_OUT(17) => 
                           IMM_DECODE_OUT_17_port, IMM_OUT(16) => 
                           IMM_DECODE_OUT_16_port, IMM_OUT(15) => 
                           IMM_DECODE_OUT_15_port, IMM_OUT(14) => 
                           IMM_DECODE_OUT_14_port, IMM_OUT(13) => 
                           IMM_DECODE_OUT_13_port, IMM_OUT(12) => 
                           IMM_DECODE_OUT_12_port, IMM_OUT(11) => 
                           IMM_DECODE_OUT_11_port, IMM_OUT(10) => 
                           IMM_DECODE_OUT_10_port, IMM_OUT(9) => 
                           IMM_DECODE_OUT_9_port, IMM_OUT(8) => 
                           IMM_DECODE_OUT_8_port, IMM_OUT(7) => 
                           IMM_DECODE_OUT_7_port, IMM_OUT(6) => 
                           IMM_DECODE_OUT_6_port, IMM_OUT(5) => 
                           IMM_DECODE_OUT_5_port, IMM_OUT(4) => 
                           IMM_DECODE_OUT_4_port, IMM_OUT(3) => 
                           IMM_DECODE_OUT_3_port, IMM_OUT(2) => 
                           IMM_DECODE_OUT_2_port, IMM_OUT(1) => 
                           IMM_DECODE_OUT_1_port, IMM_OUT(0) => 
                           IMM_DECODE_OUT_0_port, ADD_RS1_HDU(4) => 
                           ADD_RS1_HDU_4_port, ADD_RS1_HDU(3) => 
                           ADD_RS1_HDU_3_port, ADD_RS1_HDU(2) => 
                           ADD_RS1_HDU_2_port, ADD_RS1_HDU(1) => 
                           ADD_RS1_HDU_1_port, ADD_RS1_HDU(0) => 
                           ADD_RS1_HDU_0_port, ADD_RS2_HDU(4) => 
                           ADD_RS2_HDU_4_port, ADD_RS2_HDU(3) => 
                           ADD_RS2_HDU_3_port, ADD_RS2_HDU(2) => 
                           ADD_RS2_HDU_2_port, ADD_RS2_HDU(1) => 
                           ADD_RS2_HDU_1_port, ADD_RS2_HDU(0) => 
                           ADD_RS2_HDU_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_DECODE_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_DECODE_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_DECODE_OUT_0_port, ADD_RS1_OUT(4) => 
                           ADD_RS1_DECODE_OUT_4_port, ADD_RS1_OUT(3) => 
                           ADD_RS1_DECODE_OUT_3_port, ADD_RS1_OUT(2) => 
                           ADD_RS1_DECODE_OUT_2_port, ADD_RS1_OUT(1) => 
                           ADD_RS1_DECODE_OUT_1_port, ADD_RS1_OUT(0) => 
                           ADD_RS1_DECODE_OUT_0_port, ADD_RS2_OUT(4) => 
                           ADD_RS2_DECODE_OUT_4_port, ADD_RS2_OUT(3) => 
                           ADD_RS2_DECODE_OUT_3_port, ADD_RS2_OUT(2) => 
                           ADD_RS2_DECODE_OUT_2_port, ADD_RS2_OUT(1) => 
                           ADD_RS2_DECODE_OUT_1_port, ADD_RS2_OUT(0) => 
                           ADD_RS2_DECODE_OUT_0_port);
   ExecuteStage : Execute port map( CLK => CLK, RST => RST, MUX_A_SEL => 
                           MUX_A_SEL, MUX_B_SEL(1) => MUX_B_SEL(1), 
                           MUX_B_SEL(0) => MUX_B_SEL(0), ALU_OPC(0) => 
                           ALU_OPC(0), ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => 
                           ALU_OPC(2), ALU_OPC(3) => ALU_OPC(3), ALU_OPC(4) => 
                           ALU_OPC(4), ALU_OUTREG_EN => ALU_OUTREG_EN, 
                           JUMP_TYPE(1) => JUMP_TYPE(1), JUMP_TYPE(0) => 
                           JUMP_TYPE(0), PC_IN(31) => PC_DECODE_OUT_31_port, 
                           PC_IN(30) => PC_DECODE_OUT_30_port, PC_IN(29) => 
                           PC_DECODE_OUT_29_port, PC_IN(28) => 
                           PC_DECODE_OUT_28_port, PC_IN(27) => 
                           PC_DECODE_OUT_27_port, PC_IN(26) => 
                           PC_DECODE_OUT_26_port, PC_IN(25) => 
                           PC_DECODE_OUT_25_port, PC_IN(24) => 
                           PC_DECODE_OUT_24_port, PC_IN(23) => 
                           PC_DECODE_OUT_23_port, PC_IN(22) => 
                           PC_DECODE_OUT_22_port, PC_IN(21) => 
                           PC_DECODE_OUT_21_port, PC_IN(20) => 
                           PC_DECODE_OUT_20_port, PC_IN(19) => 
                           PC_DECODE_OUT_19_port, PC_IN(18) => 
                           PC_DECODE_OUT_18_port, PC_IN(17) => 
                           PC_DECODE_OUT_17_port, PC_IN(16) => 
                           PC_DECODE_OUT_16_port, PC_IN(15) => 
                           PC_DECODE_OUT_15_port, PC_IN(14) => 
                           PC_DECODE_OUT_14_port, PC_IN(13) => 
                           PC_DECODE_OUT_13_port, PC_IN(12) => 
                           PC_DECODE_OUT_12_port, PC_IN(11) => 
                           PC_DECODE_OUT_11_port, PC_IN(10) => 
                           PC_DECODE_OUT_10_port, PC_IN(9) => 
                           PC_DECODE_OUT_9_port, PC_IN(8) => 
                           PC_DECODE_OUT_8_port, PC_IN(7) => 
                           PC_DECODE_OUT_7_port, PC_IN(6) => 
                           PC_DECODE_OUT_6_port, PC_IN(5) => 
                           PC_DECODE_OUT_5_port, PC_IN(4) => 
                           PC_DECODE_OUT_4_port, PC_IN(3) => 
                           PC_DECODE_OUT_3_port, PC_IN(2) => 
                           PC_DECODE_OUT_2_port, PC_IN(1) => 
                           PC_DECODE_OUT_1_port, PC_IN(0) => 
                           PC_DECODE_OUT_0_port, A_IN(31) => 
                           A_DECODE_OUT_31_port, A_IN(30) => 
                           A_DECODE_OUT_30_port, A_IN(29) => 
                           A_DECODE_OUT_29_port, A_IN(28) => 
                           A_DECODE_OUT_28_port, A_IN(27) => 
                           A_DECODE_OUT_27_port, A_IN(26) => 
                           A_DECODE_OUT_26_port, A_IN(25) => 
                           A_DECODE_OUT_25_port, A_IN(24) => 
                           A_DECODE_OUT_24_port, A_IN(23) => 
                           A_DECODE_OUT_23_port, A_IN(22) => 
                           A_DECODE_OUT_22_port, A_IN(21) => 
                           A_DECODE_OUT_21_port, A_IN(20) => 
                           A_DECODE_OUT_20_port, A_IN(19) => 
                           A_DECODE_OUT_19_port, A_IN(18) => 
                           A_DECODE_OUT_18_port, A_IN(17) => 
                           A_DECODE_OUT_17_port, A_IN(16) => 
                           A_DECODE_OUT_16_port, A_IN(15) => 
                           A_DECODE_OUT_15_port, A_IN(14) => 
                           A_DECODE_OUT_14_port, A_IN(13) => 
                           A_DECODE_OUT_13_port, A_IN(12) => 
                           A_DECODE_OUT_12_port, A_IN(11) => 
                           A_DECODE_OUT_11_port, A_IN(10) => 
                           A_DECODE_OUT_10_port, A_IN(9) => A_DECODE_OUT_9_port
                           , A_IN(8) => A_DECODE_OUT_8_port, A_IN(7) => 
                           A_DECODE_OUT_7_port, A_IN(6) => A_DECODE_OUT_6_port,
                           A_IN(5) => A_DECODE_OUT_5_port, A_IN(4) => 
                           A_DECODE_OUT_4_port, A_IN(3) => A_DECODE_OUT_3_port,
                           A_IN(2) => A_DECODE_OUT_2_port, A_IN(1) => 
                           A_DECODE_OUT_1_port, A_IN(0) => A_DECODE_OUT_0_port,
                           B_IN(31) => B_DECODE_OUT_31_port, B_IN(30) => 
                           B_DECODE_OUT_30_port, B_IN(29) => 
                           B_DECODE_OUT_29_port, B_IN(28) => 
                           B_DECODE_OUT_28_port, B_IN(27) => 
                           B_DECODE_OUT_27_port, B_IN(26) => 
                           B_DECODE_OUT_26_port, B_IN(25) => 
                           B_DECODE_OUT_25_port, B_IN(24) => 
                           B_DECODE_OUT_24_port, B_IN(23) => 
                           B_DECODE_OUT_23_port, B_IN(22) => 
                           B_DECODE_OUT_22_port, B_IN(21) => 
                           B_DECODE_OUT_21_port, B_IN(20) => 
                           B_DECODE_OUT_20_port, B_IN(19) => 
                           B_DECODE_OUT_19_port, B_IN(18) => 
                           B_DECODE_OUT_18_port, B_IN(17) => 
                           B_DECODE_OUT_17_port, B_IN(16) => 
                           B_DECODE_OUT_16_port, B_IN(15) => 
                           B_DECODE_OUT_15_port, B_IN(14) => 
                           B_DECODE_OUT_14_port, B_IN(13) => 
                           B_DECODE_OUT_13_port, B_IN(12) => 
                           B_DECODE_OUT_12_port, B_IN(11) => 
                           B_DECODE_OUT_11_port, B_IN(10) => 
                           B_DECODE_OUT_10_port, B_IN(9) => B_DECODE_OUT_9_port
                           , B_IN(8) => B_DECODE_OUT_8_port, B_IN(7) => 
                           B_DECODE_OUT_7_port, B_IN(6) => B_DECODE_OUT_6_port,
                           B_IN(5) => B_DECODE_OUT_5_port, B_IN(4) => 
                           B_DECODE_OUT_4_port, B_IN(3) => B_DECODE_OUT_3_port,
                           B_IN(2) => B_DECODE_OUT_2_port, B_IN(1) => 
                           B_DECODE_OUT_1_port, B_IN(0) => B_DECODE_OUT_0_port,
                           IMM_IN(31) => IMM_DECODE_OUT_31_port, IMM_IN(30) => 
                           IMM_DECODE_OUT_30_port, IMM_IN(29) => 
                           IMM_DECODE_OUT_29_port, IMM_IN(28) => 
                           IMM_DECODE_OUT_28_port, IMM_IN(27) => 
                           IMM_DECODE_OUT_27_port, IMM_IN(26) => 
                           IMM_DECODE_OUT_26_port, IMM_IN(25) => 
                           IMM_DECODE_OUT_25_port, IMM_IN(24) => 
                           IMM_DECODE_OUT_24_port, IMM_IN(23) => 
                           IMM_DECODE_OUT_23_port, IMM_IN(22) => 
                           IMM_DECODE_OUT_22_port, IMM_IN(21) => 
                           IMM_DECODE_OUT_21_port, IMM_IN(20) => 
                           IMM_DECODE_OUT_20_port, IMM_IN(19) => 
                           IMM_DECODE_OUT_19_port, IMM_IN(18) => 
                           IMM_DECODE_OUT_18_port, IMM_IN(17) => 
                           IMM_DECODE_OUT_17_port, IMM_IN(16) => 
                           IMM_DECODE_OUT_16_port, IMM_IN(15) => 
                           IMM_DECODE_OUT_15_port, IMM_IN(14) => 
                           IMM_DECODE_OUT_14_port, IMM_IN(13) => 
                           IMM_DECODE_OUT_13_port, IMM_IN(12) => 
                           IMM_DECODE_OUT_12_port, IMM_IN(11) => 
                           IMM_DECODE_OUT_11_port, IMM_IN(10) => 
                           IMM_DECODE_OUT_10_port, IMM_IN(9) => 
                           IMM_DECODE_OUT_9_port, IMM_IN(8) => 
                           IMM_DECODE_OUT_8_port, IMM_IN(7) => 
                           IMM_DECODE_OUT_7_port, IMM_IN(6) => 
                           IMM_DECODE_OUT_6_port, IMM_IN(5) => 
                           IMM_DECODE_OUT_5_port, IMM_IN(4) => 
                           IMM_DECODE_OUT_4_port, IMM_IN(3) => 
                           IMM_DECODE_OUT_3_port, IMM_IN(2) => 
                           IMM_DECODE_OUT_2_port, IMM_IN(1) => 
                           IMM_DECODE_OUT_1_port, IMM_IN(0) => 
                           IMM_DECODE_OUT_0_port, ADD_WR_IN(4) => 
                           ADD_WR_DECODE_OUT_4_port, ADD_WR_IN(3) => 
                           ADD_WR_DECODE_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_DECODE_OUT_0_port, ADD_RS1_IN(4) => 
                           ADD_RS1_DECODE_OUT_4_port, ADD_RS1_IN(3) => 
                           ADD_RS1_DECODE_OUT_3_port, ADD_RS1_IN(2) => 
                           ADD_RS1_DECODE_OUT_2_port, ADD_RS1_IN(1) => 
                           ADD_RS1_DECODE_OUT_1_port, ADD_RS1_IN(0) => 
                           ADD_RS1_DECODE_OUT_0_port, ADD_RS2_IN(4) => 
                           ADD_RS2_DECODE_OUT_4_port, ADD_RS2_IN(3) => 
                           ADD_RS2_DECODE_OUT_3_port, ADD_RS2_IN(2) => 
                           ADD_RS2_DECODE_OUT_2_port, ADD_RS2_IN(1) => 
                           ADD_RS2_DECODE_OUT_1_port, ADD_RS2_IN(0) => 
                           ADD_RS2_DECODE_OUT_0_port, ADD_WR_MEM(4) => 
                           ADD_WR_MEM_4_port, ADD_WR_MEM(3) => 
                           ADD_WR_MEM_3_port, ADD_WR_MEM(2) => 
                           ADD_WR_MEM_2_port, ADD_WR_MEM(1) => 
                           ADD_WR_MEM_1_port, ADD_WR_MEM(0) => 
                           ADD_WR_MEM_0_port, ADD_WR_WB(4) => ADD_WR_WB_4_port,
                           ADD_WR_WB(3) => ADD_WR_WB_3_port, ADD_WR_WB(2) => 
                           ADD_WR_WB_2_port, ADD_WR_WB(1) => ADD_WR_WB_1_port, 
                           ADD_WR_WB(0) => ADD_WR_WB_0_port, RF_WE_MEM => RF_WE
                           , RF_WE_WB => RF_WE_WB, OP_MEM(31) => OP_MEM_31_port
                           , OP_MEM(30) => OP_MEM_30_port, OP_MEM(29) => 
                           OP_MEM_29_port, OP_MEM(28) => OP_MEM_28_port, 
                           OP_MEM(27) => OP_MEM_27_port, OP_MEM(26) => 
                           OP_MEM_26_port, OP_MEM(25) => OP_MEM_25_port, 
                           OP_MEM(24) => OP_MEM_24_port, OP_MEM(23) => 
                           OP_MEM_23_port, OP_MEM(22) => OP_MEM_22_port, 
                           OP_MEM(21) => OP_MEM_21_port, OP_MEM(20) => 
                           OP_MEM_20_port, OP_MEM(19) => OP_MEM_19_port, 
                           OP_MEM(18) => OP_MEM_18_port, OP_MEM(17) => 
                           OP_MEM_17_port, OP_MEM(16) => OP_MEM_16_port, 
                           OP_MEM(15) => OP_MEM_15_port, OP_MEM(14) => 
                           OP_MEM_14_port, OP_MEM(13) => OP_MEM_13_port, 
                           OP_MEM(12) => OP_MEM_12_port, OP_MEM(11) => 
                           OP_MEM_11_port, OP_MEM(10) => OP_MEM_10_port, 
                           OP_MEM(9) => OP_MEM_9_port, OP_MEM(8) => 
                           OP_MEM_8_port, OP_MEM(7) => OP_MEM_7_port, OP_MEM(6)
                           => OP_MEM_6_port, OP_MEM(5) => OP_MEM_5_port, 
                           OP_MEM(4) => OP_MEM_4_port, OP_MEM(3) => 
                           OP_MEM_3_port, OP_MEM(2) => OP_MEM_2_port, OP_MEM(1)
                           => OP_MEM_1_port, OP_MEM(0) => OP_MEM_0_port, 
                           OP_WB(31) => OP_WB_31_port, OP_WB(30) => 
                           OP_WB_30_port, OP_WB(29) => OP_WB_29_port, OP_WB(28)
                           => OP_WB_28_port, OP_WB(27) => OP_WB_27_port, 
                           OP_WB(26) => OP_WB_26_port, OP_WB(25) => 
                           OP_WB_25_port, OP_WB(24) => OP_WB_24_port, OP_WB(23)
                           => OP_WB_23_port, OP_WB(22) => OP_WB_22_port, 
                           OP_WB(21) => OP_WB_21_port, OP_WB(20) => 
                           OP_WB_20_port, OP_WB(19) => OP_WB_19_port, OP_WB(18)
                           => OP_WB_18_port, OP_WB(17) => OP_WB_17_port, 
                           OP_WB(16) => OP_WB_16_port, OP_WB(15) => 
                           OP_WB_15_port, OP_WB(14) => OP_WB_14_port, OP_WB(13)
                           => OP_WB_13_port, OP_WB(12) => OP_WB_12_port, 
                           OP_WB(11) => OP_WB_11_port, OP_WB(10) => 
                           OP_WB_10_port, OP_WB(9) => OP_WB_9_port, OP_WB(8) =>
                           OP_WB_8_port, OP_WB(7) => OP_WB_7_port, OP_WB(6) => 
                           OP_WB_6_port, OP_WB(5) => OP_WB_5_port, OP_WB(4) => 
                           OP_WB_4_port, OP_WB(3) => OP_WB_3_port, OP_WB(2) => 
                           OP_WB_2_port, OP_WB(1) => OP_WB_1_port, OP_WB(0) => 
                           OP_WB_0_port, PC_SEL(1) => PC_SEL_EX_1_port, 
                           PC_SEL(0) => PC_SEL_EX_0_port, ZERO_FLAG => 
                           ZERO_FLAG_EX, NPC_ABS(31) => NPC_ABS_EX_31_port, 
                           NPC_ABS(30) => NPC_ABS_EX_30_port, NPC_ABS(29) => 
                           NPC_ABS_EX_29_port, NPC_ABS(28) => 
                           NPC_ABS_EX_28_port, NPC_ABS(27) => 
                           NPC_ABS_EX_27_port, NPC_ABS(26) => 
                           NPC_ABS_EX_26_port, NPC_ABS(25) => 
                           NPC_ABS_EX_25_port, NPC_ABS(24) => 
                           NPC_ABS_EX_24_port, NPC_ABS(23) => 
                           NPC_ABS_EX_23_port, NPC_ABS(22) => 
                           NPC_ABS_EX_22_port, NPC_ABS(21) => 
                           NPC_ABS_EX_21_port, NPC_ABS(20) => 
                           NPC_ABS_EX_20_port, NPC_ABS(19) => 
                           NPC_ABS_EX_19_port, NPC_ABS(18) => 
                           NPC_ABS_EX_18_port, NPC_ABS(17) => 
                           NPC_ABS_EX_17_port, NPC_ABS(16) => 
                           NPC_ABS_EX_16_port, NPC_ABS(15) => 
                           NPC_ABS_EX_15_port, NPC_ABS(14) => 
                           NPC_ABS_EX_14_port, NPC_ABS(13) => 
                           NPC_ABS_EX_13_port, NPC_ABS(12) => 
                           NPC_ABS_EX_12_port, NPC_ABS(11) => 
                           NPC_ABS_EX_11_port, NPC_ABS(10) => 
                           NPC_ABS_EX_10_port, NPC_ABS(9) => NPC_ABS_EX_9_port,
                           NPC_ABS(8) => NPC_ABS_EX_8_port, NPC_ABS(7) => 
                           NPC_ABS_EX_7_port, NPC_ABS(6) => NPC_ABS_EX_6_port, 
                           NPC_ABS(5) => NPC_ABS_EX_5_port, NPC_ABS(4) => 
                           NPC_ABS_EX_4_port, NPC_ABS(3) => NPC_ABS_EX_3_port, 
                           NPC_ABS(2) => NPC_ABS_EX_2_port, NPC_ABS(1) => 
                           NPC_ABS_EX_1_port, NPC_ABS(0) => NPC_ABS_EX_0_port, 
                           NPC_REL(31) => NPC_REL_EX_31_port, NPC_REL(30) => 
                           NPC_REL_EX_30_port, NPC_REL(29) => 
                           NPC_REL_EX_29_port, NPC_REL(28) => 
                           NPC_REL_EX_28_port, NPC_REL(27) => 
                           NPC_REL_EX_27_port, NPC_REL(26) => 
                           NPC_REL_EX_26_port, NPC_REL(25) => 
                           NPC_REL_EX_25_port, NPC_REL(24) => 
                           NPC_REL_EX_24_port, NPC_REL(23) => 
                           NPC_REL_EX_23_port, NPC_REL(22) => 
                           NPC_REL_EX_22_port, NPC_REL(21) => 
                           NPC_REL_EX_21_port, NPC_REL(20) => 
                           NPC_REL_EX_20_port, NPC_REL(19) => 
                           NPC_REL_EX_19_port, NPC_REL(18) => 
                           NPC_REL_EX_18_port, NPC_REL(17) => 
                           NPC_REL_EX_17_port, NPC_REL(16) => 
                           NPC_REL_EX_16_port, NPC_REL(15) => 
                           NPC_REL_EX_15_port, NPC_REL(14) => 
                           NPC_REL_EX_14_port, NPC_REL(13) => 
                           NPC_REL_EX_13_port, NPC_REL(12) => 
                           NPC_REL_EX_12_port, NPC_REL(11) => 
                           NPC_REL_EX_11_port, NPC_REL(10) => 
                           NPC_REL_EX_10_port, NPC_REL(9) => NPC_REL_EX_9_port,
                           NPC_REL(8) => NPC_REL_EX_8_port, NPC_REL(7) => 
                           NPC_REL_EX_7_port, NPC_REL(6) => NPC_REL_EX_6_port, 
                           NPC_REL(5) => NPC_REL_EX_5_port, NPC_REL(4) => 
                           NPC_REL_EX_4_port, NPC_REL(3) => NPC_REL_EX_3_port, 
                           NPC_REL(2) => NPC_REL_EX_2_port, NPC_REL(1) => 
                           NPC_REL_EX_1_port, NPC_REL(0) => NPC_REL_EX_0_port, 
                           ALU_RES(31) => ALU_RES_EX_31_port, ALU_RES(30) => 
                           ALU_RES_EX_30_port, ALU_RES(29) => 
                           ALU_RES_EX_29_port, ALU_RES(28) => 
                           ALU_RES_EX_28_port, ALU_RES(27) => 
                           ALU_RES_EX_27_port, ALU_RES(26) => 
                           ALU_RES_EX_26_port, ALU_RES(25) => 
                           ALU_RES_EX_25_port, ALU_RES(24) => 
                           ALU_RES_EX_24_port, ALU_RES(23) => 
                           ALU_RES_EX_23_port, ALU_RES(22) => 
                           ALU_RES_EX_22_port, ALU_RES(21) => 
                           ALU_RES_EX_21_port, ALU_RES(20) => 
                           ALU_RES_EX_20_port, ALU_RES(19) => 
                           ALU_RES_EX_19_port, ALU_RES(18) => 
                           ALU_RES_EX_18_port, ALU_RES(17) => 
                           ALU_RES_EX_17_port, ALU_RES(16) => 
                           ALU_RES_EX_16_port, ALU_RES(15) => 
                           ALU_RES_EX_15_port, ALU_RES(14) => 
                           ALU_RES_EX_14_port, ALU_RES(13) => 
                           ALU_RES_EX_13_port, ALU_RES(12) => 
                           ALU_RES_EX_12_port, ALU_RES(11) => 
                           ALU_RES_EX_11_port, ALU_RES(10) => 
                           ALU_RES_EX_10_port, ALU_RES(9) => ALU_RES_EX_9_port,
                           ALU_RES(8) => ALU_RES_EX_8_port, ALU_RES(7) => 
                           ALU_RES_EX_7_port, ALU_RES(6) => ALU_RES_EX_6_port, 
                           ALU_RES(5) => ALU_RES_EX_5_port, ALU_RES(4) => 
                           ALU_RES_EX_4_port, ALU_RES(3) => ALU_RES_EX_3_port, 
                           ALU_RES(2) => ALU_RES_EX_2_port, ALU_RES(1) => 
                           ALU_RES_EX_1_port, ALU_RES(0) => ALU_RES_EX_0_port, 
                           B_OUT(31) => B_EX_OUT_31_port, B_OUT(30) => 
                           B_EX_OUT_30_port, B_OUT(29) => B_EX_OUT_29_port, 
                           B_OUT(28) => B_EX_OUT_28_port, B_OUT(27) => 
                           B_EX_OUT_27_port, B_OUT(26) => B_EX_OUT_26_port, 
                           B_OUT(25) => B_EX_OUT_25_port, B_OUT(24) => 
                           B_EX_OUT_24_port, B_OUT(23) => B_EX_OUT_23_port, 
                           B_OUT(22) => B_EX_OUT_22_port, B_OUT(21) => 
                           B_EX_OUT_21_port, B_OUT(20) => B_EX_OUT_20_port, 
                           B_OUT(19) => B_EX_OUT_19_port, B_OUT(18) => 
                           B_EX_OUT_18_port, B_OUT(17) => B_EX_OUT_17_port, 
                           B_OUT(16) => B_EX_OUT_16_port, B_OUT(15) => 
                           B_EX_OUT_15_port, B_OUT(14) => B_EX_OUT_14_port, 
                           B_OUT(13) => B_EX_OUT_13_port, B_OUT(12) => 
                           B_EX_OUT_12_port, B_OUT(11) => B_EX_OUT_11_port, 
                           B_OUT(10) => B_EX_OUT_10_port, B_OUT(9) => 
                           B_EX_OUT_9_port, B_OUT(8) => B_EX_OUT_8_port, 
                           B_OUT(7) => B_EX_OUT_7_port, B_OUT(6) => 
                           B_EX_OUT_6_port, B_OUT(5) => B_EX_OUT_5_port, 
                           B_OUT(4) => B_EX_OUT_4_port, B_OUT(3) => 
                           B_EX_OUT_3_port, B_OUT(2) => B_EX_OUT_2_port, 
                           B_OUT(1) => B_EX_OUT_1_port, B_OUT(0) => 
                           B_EX_OUT_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_EX_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_EX_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_EX_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_EX_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_EX_OUT_0_port);
   DRAM_R_ff : ff_0 port map( D => DRAM_R_IN, CLK => CLK, EN => X_Logic1_port, 
                           RST => RST, Q => DRAM_R_MEM);
   MemoryStage : Memory port map( CLK => CLK, RST => RST, MEM_EN_IN => 
                           MEM_EN_IN, DRAM_R_IN => DRAM_R_MEM, DRAM_W_IN => 
                           DRAM_W_IN, PC_SEL(1) => PC_SEL_EX_1_port, PC_SEL(0) 
                           => PC_SEL_EX_0_port, NPC_IN(31) => 
                           NPC_FETCH_OUT_31_port, NPC_IN(30) => 
                           NPC_FETCH_OUT_30_port, NPC_IN(29) => 
                           NPC_FETCH_OUT_29_port, NPC_IN(28) => 
                           NPC_FETCH_OUT_28_port, NPC_IN(27) => 
                           NPC_FETCH_OUT_27_port, NPC_IN(26) => 
                           NPC_FETCH_OUT_26_port, NPC_IN(25) => 
                           NPC_FETCH_OUT_25_port, NPC_IN(24) => 
                           NPC_FETCH_OUT_24_port, NPC_IN(23) => 
                           NPC_FETCH_OUT_23_port, NPC_IN(22) => 
                           NPC_FETCH_OUT_22_port, NPC_IN(21) => 
                           NPC_FETCH_OUT_21_port, NPC_IN(20) => 
                           NPC_FETCH_OUT_20_port, NPC_IN(19) => 
                           NPC_FETCH_OUT_19_port, NPC_IN(18) => 
                           NPC_FETCH_OUT_18_port, NPC_IN(17) => 
                           NPC_FETCH_OUT_17_port, NPC_IN(16) => 
                           NPC_FETCH_OUT_16_port, NPC_IN(15) => 
                           NPC_FETCH_OUT_15_port, NPC_IN(14) => 
                           NPC_FETCH_OUT_14_port, NPC_IN(13) => 
                           NPC_FETCH_OUT_13_port, NPC_IN(12) => 
                           NPC_FETCH_OUT_12_port, NPC_IN(11) => 
                           NPC_FETCH_OUT_11_port, NPC_IN(10) => 
                           NPC_FETCH_OUT_10_port, NPC_IN(9) => 
                           NPC_FETCH_OUT_9_port, NPC_IN(8) => 
                           NPC_FETCH_OUT_8_port, NPC_IN(7) => 
                           NPC_FETCH_OUT_7_port, NPC_IN(6) => 
                           NPC_FETCH_OUT_6_port, NPC_IN(5) => 
                           NPC_FETCH_OUT_5_port, NPC_IN(4) => 
                           NPC_FETCH_OUT_4_port, NPC_IN(3) => 
                           NPC_FETCH_OUT_3_port, NPC_IN(2) => 
                           NPC_FETCH_OUT_2_port, NPC_IN(1) => 
                           NPC_FETCH_OUT_1_port, NPC_IN(0) => 
                           NPC_FETCH_OUT_0_port, NPC_ABS(31) => 
                           NPC_ABS_EX_31_port, NPC_ABS(30) => 
                           NPC_ABS_EX_30_port, NPC_ABS(29) => 
                           NPC_ABS_EX_29_port, NPC_ABS(28) => 
                           NPC_ABS_EX_28_port, NPC_ABS(27) => 
                           NPC_ABS_EX_27_port, NPC_ABS(26) => 
                           NPC_ABS_EX_26_port, NPC_ABS(25) => 
                           NPC_ABS_EX_25_port, NPC_ABS(24) => 
                           NPC_ABS_EX_24_port, NPC_ABS(23) => 
                           NPC_ABS_EX_23_port, NPC_ABS(22) => 
                           NPC_ABS_EX_22_port, NPC_ABS(21) => 
                           NPC_ABS_EX_21_port, NPC_ABS(20) => 
                           NPC_ABS_EX_20_port, NPC_ABS(19) => 
                           NPC_ABS_EX_19_port, NPC_ABS(18) => 
                           NPC_ABS_EX_18_port, NPC_ABS(17) => 
                           NPC_ABS_EX_17_port, NPC_ABS(16) => 
                           NPC_ABS_EX_16_port, NPC_ABS(15) => 
                           NPC_ABS_EX_15_port, NPC_ABS(14) => 
                           NPC_ABS_EX_14_port, NPC_ABS(13) => 
                           NPC_ABS_EX_13_port, NPC_ABS(12) => 
                           NPC_ABS_EX_12_port, NPC_ABS(11) => 
                           NPC_ABS_EX_11_port, NPC_ABS(10) => 
                           NPC_ABS_EX_10_port, NPC_ABS(9) => NPC_ABS_EX_9_port,
                           NPC_ABS(8) => NPC_ABS_EX_8_port, NPC_ABS(7) => 
                           NPC_ABS_EX_7_port, NPC_ABS(6) => NPC_ABS_EX_6_port, 
                           NPC_ABS(5) => NPC_ABS_EX_5_port, NPC_ABS(4) => 
                           NPC_ABS_EX_4_port, NPC_ABS(3) => NPC_ABS_EX_3_port, 
                           NPC_ABS(2) => NPC_ABS_EX_2_port, NPC_ABS(1) => 
                           NPC_ABS_EX_1_port, NPC_ABS(0) => NPC_ABS_EX_0_port, 
                           NPC_REL(31) => NPC_REL_EX_31_port, NPC_REL(30) => 
                           NPC_REL_EX_30_port, NPC_REL(29) => 
                           NPC_REL_EX_29_port, NPC_REL(28) => 
                           NPC_REL_EX_28_port, NPC_REL(27) => 
                           NPC_REL_EX_27_port, NPC_REL(26) => 
                           NPC_REL_EX_26_port, NPC_REL(25) => 
                           NPC_REL_EX_25_port, NPC_REL(24) => 
                           NPC_REL_EX_24_port, NPC_REL(23) => 
                           NPC_REL_EX_23_port, NPC_REL(22) => 
                           NPC_REL_EX_22_port, NPC_REL(21) => 
                           NPC_REL_EX_21_port, NPC_REL(20) => 
                           NPC_REL_EX_20_port, NPC_REL(19) => 
                           NPC_REL_EX_19_port, NPC_REL(18) => 
                           NPC_REL_EX_18_port, NPC_REL(17) => 
                           NPC_REL_EX_17_port, NPC_REL(16) => 
                           NPC_REL_EX_16_port, NPC_REL(15) => 
                           NPC_REL_EX_15_port, NPC_REL(14) => 
                           NPC_REL_EX_14_port, NPC_REL(13) => 
                           NPC_REL_EX_13_port, NPC_REL(12) => 
                           NPC_REL_EX_12_port, NPC_REL(11) => 
                           NPC_REL_EX_11_port, NPC_REL(10) => 
                           NPC_REL_EX_10_port, NPC_REL(9) => NPC_REL_EX_9_port,
                           NPC_REL(8) => NPC_REL_EX_8_port, NPC_REL(7) => 
                           NPC_REL_EX_7_port, NPC_REL(6) => NPC_REL_EX_6_port, 
                           NPC_REL(5) => NPC_REL_EX_5_port, NPC_REL(4) => 
                           NPC_REL_EX_4_port, NPC_REL(3) => NPC_REL_EX_3_port, 
                           NPC_REL(2) => NPC_REL_EX_2_port, NPC_REL(1) => 
                           NPC_REL_EX_1_port, NPC_REL(0) => NPC_REL_EX_0_port, 
                           ALU_RES_IN(31) => ALU_RES_EX_31_port, ALU_RES_IN(30)
                           => ALU_RES_EX_30_port, ALU_RES_IN(29) => 
                           ALU_RES_EX_29_port, ALU_RES_IN(28) => 
                           ALU_RES_EX_28_port, ALU_RES_IN(27) => 
                           ALU_RES_EX_27_port, ALU_RES_IN(26) => 
                           ALU_RES_EX_26_port, ALU_RES_IN(25) => 
                           ALU_RES_EX_25_port, ALU_RES_IN(24) => 
                           ALU_RES_EX_24_port, ALU_RES_IN(23) => 
                           ALU_RES_EX_23_port, ALU_RES_IN(22) => 
                           ALU_RES_EX_22_port, ALU_RES_IN(21) => 
                           ALU_RES_EX_21_port, ALU_RES_IN(20) => 
                           ALU_RES_EX_20_port, ALU_RES_IN(19) => 
                           ALU_RES_EX_19_port, ALU_RES_IN(18) => 
                           ALU_RES_EX_18_port, ALU_RES_IN(17) => 
                           ALU_RES_EX_17_port, ALU_RES_IN(16) => 
                           ALU_RES_EX_16_port, ALU_RES_IN(15) => 
                           ALU_RES_EX_15_port, ALU_RES_IN(14) => 
                           ALU_RES_EX_14_port, ALU_RES_IN(13) => 
                           ALU_RES_EX_13_port, ALU_RES_IN(12) => 
                           ALU_RES_EX_12_port, ALU_RES_IN(11) => 
                           ALU_RES_EX_11_port, ALU_RES_IN(10) => 
                           ALU_RES_EX_10_port, ALU_RES_IN(9) => 
                           ALU_RES_EX_9_port, ALU_RES_IN(8) => 
                           ALU_RES_EX_8_port, ALU_RES_IN(7) => 
                           ALU_RES_EX_7_port, ALU_RES_IN(6) => 
                           ALU_RES_EX_6_port, ALU_RES_IN(5) => 
                           ALU_RES_EX_5_port, ALU_RES_IN(4) => 
                           ALU_RES_EX_4_port, ALU_RES_IN(3) => 
                           ALU_RES_EX_3_port, ALU_RES_IN(2) => 
                           ALU_RES_EX_2_port, ALU_RES_IN(1) => 
                           ALU_RES_EX_1_port, ALU_RES_IN(0) => 
                           ALU_RES_EX_0_port, B_IN(31) => B_EX_OUT_31_port, 
                           B_IN(30) => B_EX_OUT_30_port, B_IN(29) => 
                           B_EX_OUT_29_port, B_IN(28) => B_EX_OUT_28_port, 
                           B_IN(27) => B_EX_OUT_27_port, B_IN(26) => 
                           B_EX_OUT_26_port, B_IN(25) => B_EX_OUT_25_port, 
                           B_IN(24) => B_EX_OUT_24_port, B_IN(23) => 
                           B_EX_OUT_23_port, B_IN(22) => B_EX_OUT_22_port, 
                           B_IN(21) => B_EX_OUT_21_port, B_IN(20) => 
                           B_EX_OUT_20_port, B_IN(19) => B_EX_OUT_19_port, 
                           B_IN(18) => B_EX_OUT_18_port, B_IN(17) => 
                           B_EX_OUT_17_port, B_IN(16) => B_EX_OUT_16_port, 
                           B_IN(15) => B_EX_OUT_15_port, B_IN(14) => 
                           B_EX_OUT_14_port, B_IN(13) => B_EX_OUT_13_port, 
                           B_IN(12) => B_EX_OUT_12_port, B_IN(11) => 
                           B_EX_OUT_11_port, B_IN(10) => B_EX_OUT_10_port, 
                           B_IN(9) => B_EX_OUT_9_port, B_IN(8) => 
                           B_EX_OUT_8_port, B_IN(7) => B_EX_OUT_7_port, B_IN(6)
                           => B_EX_OUT_6_port, B_IN(5) => B_EX_OUT_5_port, 
                           B_IN(4) => B_EX_OUT_4_port, B_IN(3) => 
                           B_EX_OUT_3_port, B_IN(2) => B_EX_OUT_2_port, B_IN(1)
                           => B_EX_OUT_1_port, B_IN(0) => B_EX_OUT_0_port, 
                           ADD_WR_IN(4) => ADD_WR_EX_OUT_4_port, ADD_WR_IN(3) 
                           => ADD_WR_EX_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_EX_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_EX_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_EX_OUT_0_port, DRAM_DATA_IN(31) => 
                           DATA_IN(31), DRAM_DATA_IN(30) => DATA_IN(30), 
                           DRAM_DATA_IN(29) => DATA_IN(29), DRAM_DATA_IN(28) =>
                           DATA_IN(28), DRAM_DATA_IN(27) => DATA_IN(27), 
                           DRAM_DATA_IN(26) => DATA_IN(26), DRAM_DATA_IN(25) =>
                           DATA_IN(25), DRAM_DATA_IN(24) => DATA_IN(24), 
                           DRAM_DATA_IN(23) => DATA_IN(23), DRAM_DATA_IN(22) =>
                           DATA_IN(22), DRAM_DATA_IN(21) => DATA_IN(21), 
                           DRAM_DATA_IN(20) => DATA_IN(20), DRAM_DATA_IN(19) =>
                           DATA_IN(19), DRAM_DATA_IN(18) => DATA_IN(18), 
                           DRAM_DATA_IN(17) => DATA_IN(17), DRAM_DATA_IN(16) =>
                           DATA_IN(16), DRAM_DATA_IN(15) => DATA_IN(15), 
                           DRAM_DATA_IN(14) => DATA_IN(14), DRAM_DATA_IN(13) =>
                           DATA_IN(13), DRAM_DATA_IN(12) => DATA_IN(12), 
                           DRAM_DATA_IN(11) => DATA_IN(11), DRAM_DATA_IN(10) =>
                           DATA_IN(10), DRAM_DATA_IN(9) => DATA_IN(9), 
                           DRAM_DATA_IN(8) => DATA_IN(8), DRAM_DATA_IN(7) => 
                           DATA_IN(7), DRAM_DATA_IN(6) => DATA_IN(6), 
                           DRAM_DATA_IN(5) => DATA_IN(5), DRAM_DATA_IN(4) => 
                           DATA_IN(4), DRAM_DATA_IN(3) => DATA_IN(3), 
                           DRAM_DATA_IN(2) => DATA_IN(2), DRAM_DATA_IN(1) => 
                           DATA_IN(1), DRAM_DATA_IN(0) => DATA_IN(0), 
                           LOAD_TYPE_IN(1) => LOAD_TYPE_IN(1), LOAD_TYPE_IN(0) 
                           => LOAD_TYPE_IN(0), STORE_TYPE_IN => STORE_TYPE_IN, 
                           PC_OUT(31) => PC_MEM_OUT_31_port, PC_OUT(30) => 
                           PC_MEM_OUT_30_port, PC_OUT(29) => PC_MEM_OUT_29_port
                           , PC_OUT(28) => PC_MEM_OUT_28_port, PC_OUT(27) => 
                           PC_MEM_OUT_27_port, PC_OUT(26) => PC_MEM_OUT_26_port
                           , PC_OUT(25) => PC_MEM_OUT_25_port, PC_OUT(24) => 
                           PC_MEM_OUT_24_port, PC_OUT(23) => PC_MEM_OUT_23_port
                           , PC_OUT(22) => PC_MEM_OUT_22_port, PC_OUT(21) => 
                           PC_MEM_OUT_21_port, PC_OUT(20) => PC_MEM_OUT_20_port
                           , PC_OUT(19) => PC_MEM_OUT_19_port, PC_OUT(18) => 
                           PC_MEM_OUT_18_port, PC_OUT(17) => PC_MEM_OUT_17_port
                           , PC_OUT(16) => PC_MEM_OUT_16_port, PC_OUT(15) => 
                           PC_MEM_OUT_15_port, PC_OUT(14) => PC_MEM_OUT_14_port
                           , PC_OUT(13) => PC_MEM_OUT_13_port, PC_OUT(12) => 
                           PC_MEM_OUT_12_port, PC_OUT(11) => PC_MEM_OUT_11_port
                           , PC_OUT(10) => PC_MEM_OUT_10_port, PC_OUT(9) => 
                           PC_MEM_OUT_9_port, PC_OUT(8) => PC_MEM_OUT_8_port, 
                           PC_OUT(7) => PC_MEM_OUT_7_port, PC_OUT(6) => 
                           PC_MEM_OUT_6_port, PC_OUT(5) => PC_MEM_OUT_5_port, 
                           PC_OUT(4) => PC_MEM_OUT_4_port, PC_OUT(3) => 
                           PC_MEM_OUT_3_port, PC_OUT(2) => PC_MEM_OUT_2_port, 
                           PC_OUT(1) => PC_MEM_OUT_1_port, PC_OUT(0) => 
                           PC_MEM_OUT_0_port, DRAM_R_OUT => DRAM_R_OUT, 
                           DRAM_W_OUT => DRAM_W_OUT, DRAM_ADDR_OUT(31) => 
                           DRAM_ADDR_OUT(31), DRAM_ADDR_OUT(30) => 
                           DRAM_ADDR_OUT(30), DRAM_ADDR_OUT(29) => 
                           DRAM_ADDR_OUT(29), DRAM_ADDR_OUT(28) => 
                           DRAM_ADDR_OUT(28), DRAM_ADDR_OUT(27) => 
                           DRAM_ADDR_OUT(27), DRAM_ADDR_OUT(26) => 
                           DRAM_ADDR_OUT(26), DRAM_ADDR_OUT(25) => 
                           DRAM_ADDR_OUT(25), DRAM_ADDR_OUT(24) => 
                           DRAM_ADDR_OUT(24), DRAM_ADDR_OUT(23) => 
                           DRAM_ADDR_OUT(23), DRAM_ADDR_OUT(22) => 
                           DRAM_ADDR_OUT(22), DRAM_ADDR_OUT(21) => 
                           DRAM_ADDR_OUT(21), DRAM_ADDR_OUT(20) => 
                           DRAM_ADDR_OUT(20), DRAM_ADDR_OUT(19) => 
                           DRAM_ADDR_OUT(19), DRAM_ADDR_OUT(18) => 
                           DRAM_ADDR_OUT(18), DRAM_ADDR_OUT(17) => 
                           DRAM_ADDR_OUT(17), DRAM_ADDR_OUT(16) => 
                           DRAM_ADDR_OUT(16), DRAM_ADDR_OUT(15) => 
                           DRAM_ADDR_OUT(15), DRAM_ADDR_OUT(14) => 
                           DRAM_ADDR_OUT(14), DRAM_ADDR_OUT(13) => 
                           DRAM_ADDR_OUT(13), DRAM_ADDR_OUT(12) => 
                           DRAM_ADDR_OUT(12), DRAM_ADDR_OUT(11) => 
                           DRAM_ADDR_OUT(11), DRAM_ADDR_OUT(10) => 
                           DRAM_ADDR_OUT(10), DRAM_ADDR_OUT(9) => 
                           DRAM_ADDR_OUT(9), DRAM_ADDR_OUT(8) => 
                           DRAM_ADDR_OUT(8), DRAM_ADDR_OUT(7) => 
                           DRAM_ADDR_OUT(7), DRAM_ADDR_OUT(6) => 
                           DRAM_ADDR_OUT(6), DRAM_ADDR_OUT(5) => 
                           DRAM_ADDR_OUT(5), DRAM_ADDR_OUT(4) => 
                           DRAM_ADDR_OUT(4), DRAM_ADDR_OUT(3) => 
                           DRAM_ADDR_OUT(3), DRAM_ADDR_OUT(2) => 
                           DRAM_ADDR_OUT(2), DRAM_ADDR_OUT(1) => 
                           DRAM_ADDR_OUT(1), DRAM_ADDR_OUT(0) => 
                           DRAM_ADDR_OUT(0), DRAM_DATA_OUT(31) => DATA_OUT(31),
                           DRAM_DATA_OUT(30) => DATA_OUT(30), DRAM_DATA_OUT(29)
                           => DATA_OUT(29), DRAM_DATA_OUT(28) => DATA_OUT(28), 
                           DRAM_DATA_OUT(27) => DATA_OUT(27), DRAM_DATA_OUT(26)
                           => DATA_OUT(26), DRAM_DATA_OUT(25) => DATA_OUT(25), 
                           DRAM_DATA_OUT(24) => DATA_OUT(24), DRAM_DATA_OUT(23)
                           => DATA_OUT(23), DRAM_DATA_OUT(22) => DATA_OUT(22), 
                           DRAM_DATA_OUT(21) => DATA_OUT(21), DRAM_DATA_OUT(20)
                           => DATA_OUT(20), DRAM_DATA_OUT(19) => DATA_OUT(19), 
                           DRAM_DATA_OUT(18) => DATA_OUT(18), DRAM_DATA_OUT(17)
                           => DATA_OUT(17), DRAM_DATA_OUT(16) => DATA_OUT(16), 
                           DRAM_DATA_OUT(15) => DATA_OUT(15), DRAM_DATA_OUT(14)
                           => DATA_OUT(14), DRAM_DATA_OUT(13) => DATA_OUT(13), 
                           DRAM_DATA_OUT(12) => DATA_OUT(12), DRAM_DATA_OUT(11)
                           => DATA_OUT(11), DRAM_DATA_OUT(10) => DATA_OUT(10), 
                           DRAM_DATA_OUT(9) => DATA_OUT(9), DRAM_DATA_OUT(8) =>
                           DATA_OUT(8), DRAM_DATA_OUT(7) => DATA_OUT(7), 
                           DRAM_DATA_OUT(6) => DATA_OUT(6), DRAM_DATA_OUT(5) =>
                           DATA_OUT(5), DRAM_DATA_OUT(4) => DATA_OUT(4), 
                           DRAM_DATA_OUT(3) => DATA_OUT(3), DRAM_DATA_OUT(2) =>
                           DATA_OUT(2), DRAM_DATA_OUT(1) => DATA_OUT(1), 
                           DRAM_DATA_OUT(0) => DATA_OUT(0), DATA_OUT(31) => 
                           DATA_MEM_OUT_31_port, DATA_OUT(30) => 
                           DATA_MEM_OUT_30_port, DATA_OUT(29) => 
                           DATA_MEM_OUT_29_port, DATA_OUT(28) => 
                           DATA_MEM_OUT_28_port, DATA_OUT(27) => 
                           DATA_MEM_OUT_27_port, DATA_OUT(26) => 
                           DATA_MEM_OUT_26_port, DATA_OUT(25) => 
                           DATA_MEM_OUT_25_port, DATA_OUT(24) => 
                           DATA_MEM_OUT_24_port, DATA_OUT(23) => 
                           DATA_MEM_OUT_23_port, DATA_OUT(22) => 
                           DATA_MEM_OUT_22_port, DATA_OUT(21) => 
                           DATA_MEM_OUT_21_port, DATA_OUT(20) => 
                           DATA_MEM_OUT_20_port, DATA_OUT(19) => 
                           DATA_MEM_OUT_19_port, DATA_OUT(18) => 
                           DATA_MEM_OUT_18_port, DATA_OUT(17) => 
                           DATA_MEM_OUT_17_port, DATA_OUT(16) => 
                           DATA_MEM_OUT_16_port, DATA_OUT(15) => 
                           DATA_MEM_OUT_15_port, DATA_OUT(14) => 
                           DATA_MEM_OUT_14_port, DATA_OUT(13) => 
                           DATA_MEM_OUT_13_port, DATA_OUT(12) => 
                           DATA_MEM_OUT_12_port, DATA_OUT(11) => 
                           DATA_MEM_OUT_11_port, DATA_OUT(10) => 
                           DATA_MEM_OUT_10_port, DATA_OUT(9) => 
                           DATA_MEM_OUT_9_port, DATA_OUT(8) => 
                           DATA_MEM_OUT_8_port, DATA_OUT(7) => 
                           DATA_MEM_OUT_7_port, DATA_OUT(6) => 
                           DATA_MEM_OUT_6_port, DATA_OUT(5) => 
                           DATA_MEM_OUT_5_port, DATA_OUT(4) => 
                           DATA_MEM_OUT_4_port, DATA_OUT(3) => 
                           DATA_MEM_OUT_3_port, DATA_OUT(2) => 
                           DATA_MEM_OUT_2_port, DATA_OUT(1) => 
                           DATA_MEM_OUT_1_port, DATA_OUT(0) => 
                           DATA_MEM_OUT_0_port, ALU_RES_OUT(31) => 
                           ALU_RES_MEM_31_port, ALU_RES_OUT(30) => 
                           ALU_RES_MEM_30_port, ALU_RES_OUT(29) => 
                           ALU_RES_MEM_29_port, ALU_RES_OUT(28) => 
                           ALU_RES_MEM_28_port, ALU_RES_OUT(27) => 
                           ALU_RES_MEM_27_port, ALU_RES_OUT(26) => 
                           ALU_RES_MEM_26_port, ALU_RES_OUT(25) => 
                           ALU_RES_MEM_25_port, ALU_RES_OUT(24) => 
                           ALU_RES_MEM_24_port, ALU_RES_OUT(23) => 
                           ALU_RES_MEM_23_port, ALU_RES_OUT(22) => 
                           ALU_RES_MEM_22_port, ALU_RES_OUT(21) => 
                           ALU_RES_MEM_21_port, ALU_RES_OUT(20) => 
                           ALU_RES_MEM_20_port, ALU_RES_OUT(19) => 
                           ALU_RES_MEM_19_port, ALU_RES_OUT(18) => 
                           ALU_RES_MEM_18_port, ALU_RES_OUT(17) => 
                           ALU_RES_MEM_17_port, ALU_RES_OUT(16) => 
                           ALU_RES_MEM_16_port, ALU_RES_OUT(15) => 
                           ALU_RES_MEM_15_port, ALU_RES_OUT(14) => 
                           ALU_RES_MEM_14_port, ALU_RES_OUT(13) => 
                           ALU_RES_MEM_13_port, ALU_RES_OUT(12) => 
                           ALU_RES_MEM_12_port, ALU_RES_OUT(11) => 
                           ALU_RES_MEM_11_port, ALU_RES_OUT(10) => 
                           ALU_RES_MEM_10_port, ALU_RES_OUT(9) => 
                           ALU_RES_MEM_9_port, ALU_RES_OUT(8) => 
                           ALU_RES_MEM_8_port, ALU_RES_OUT(7) => 
                           ALU_RES_MEM_7_port, ALU_RES_OUT(6) => 
                           ALU_RES_MEM_6_port, ALU_RES_OUT(5) => 
                           ALU_RES_MEM_5_port, ALU_RES_OUT(4) => 
                           ALU_RES_MEM_4_port, ALU_RES_OUT(3) => 
                           ALU_RES_MEM_3_port, ALU_RES_OUT(2) => 
                           ALU_RES_MEM_2_port, ALU_RES_OUT(1) => 
                           ALU_RES_MEM_1_port, ALU_RES_OUT(0) => 
                           ALU_RES_MEM_0_port, OP_MEM(31) => OP_MEM_31_port, 
                           OP_MEM(30) => OP_MEM_30_port, OP_MEM(29) => 
                           OP_MEM_29_port, OP_MEM(28) => OP_MEM_28_port, 
                           OP_MEM(27) => OP_MEM_27_port, OP_MEM(26) => 
                           OP_MEM_26_port, OP_MEM(25) => OP_MEM_25_port, 
                           OP_MEM(24) => OP_MEM_24_port, OP_MEM(23) => 
                           OP_MEM_23_port, OP_MEM(22) => OP_MEM_22_port, 
                           OP_MEM(21) => OP_MEM_21_port, OP_MEM(20) => 
                           OP_MEM_20_port, OP_MEM(19) => OP_MEM_19_port, 
                           OP_MEM(18) => OP_MEM_18_port, OP_MEM(17) => 
                           OP_MEM_17_port, OP_MEM(16) => OP_MEM_16_port, 
                           OP_MEM(15) => OP_MEM_15_port, OP_MEM(14) => 
                           OP_MEM_14_port, OP_MEM(13) => OP_MEM_13_port, 
                           OP_MEM(12) => OP_MEM_12_port, OP_MEM(11) => 
                           OP_MEM_11_port, OP_MEM(10) => OP_MEM_10_port, 
                           OP_MEM(9) => OP_MEM_9_port, OP_MEM(8) => 
                           OP_MEM_8_port, OP_MEM(7) => OP_MEM_7_port, OP_MEM(6)
                           => OP_MEM_6_port, OP_MEM(5) => OP_MEM_5_port, 
                           OP_MEM(4) => OP_MEM_4_port, OP_MEM(3) => 
                           OP_MEM_3_port, OP_MEM(2) => OP_MEM_2_port, OP_MEM(1)
                           => OP_MEM_1_port, OP_MEM(0) => OP_MEM_0_port, 
                           ADD_WR_MEM(4) => ADD_WR_MEM_4_port, ADD_WR_MEM(3) =>
                           ADD_WR_MEM_3_port, ADD_WR_MEM(2) => 
                           ADD_WR_MEM_2_port, ADD_WR_MEM(1) => 
                           ADD_WR_MEM_1_port, ADD_WR_MEM(0) => 
                           ADD_WR_MEM_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_MEM_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_MEM_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_MEM_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_MEM_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_MEM_OUT_0_port, LOAD_TYPE_OUT(1) => 
                           LOAD_TYPE_OUT(1), LOAD_TYPE_OUT(0) => 
                           LOAD_TYPE_OUT(0), STORE_TYPE_OUT => STORE_TYPE_OUT);
   RF_WE_ff : ff_2 port map( D => RF_WE, CLK => CLK, EN => X_Logic1_port, RST 
                           => RST, Q => RF_WE_WB);
   WritebackStage : Writeback port map( WB_MUX_SEL => WB_MUX_SEL, DATA_IN(31) 
                           => DATA_MEM_OUT_31_port, DATA_IN(30) => 
                           DATA_MEM_OUT_30_port, DATA_IN(29) => 
                           DATA_MEM_OUT_29_port, DATA_IN(28) => 
                           DATA_MEM_OUT_28_port, DATA_IN(27) => 
                           DATA_MEM_OUT_27_port, DATA_IN(26) => 
                           DATA_MEM_OUT_26_port, DATA_IN(25) => 
                           DATA_MEM_OUT_25_port, DATA_IN(24) => 
                           DATA_MEM_OUT_24_port, DATA_IN(23) => 
                           DATA_MEM_OUT_23_port, DATA_IN(22) => 
                           DATA_MEM_OUT_22_port, DATA_IN(21) => 
                           DATA_MEM_OUT_21_port, DATA_IN(20) => 
                           DATA_MEM_OUT_20_port, DATA_IN(19) => 
                           DATA_MEM_OUT_19_port, DATA_IN(18) => 
                           DATA_MEM_OUT_18_port, DATA_IN(17) => 
                           DATA_MEM_OUT_17_port, DATA_IN(16) => 
                           DATA_MEM_OUT_16_port, DATA_IN(15) => 
                           DATA_MEM_OUT_15_port, DATA_IN(14) => 
                           DATA_MEM_OUT_14_port, DATA_IN(13) => 
                           DATA_MEM_OUT_13_port, DATA_IN(12) => 
                           DATA_MEM_OUT_12_port, DATA_IN(11) => 
                           DATA_MEM_OUT_11_port, DATA_IN(10) => 
                           DATA_MEM_OUT_10_port, DATA_IN(9) => 
                           DATA_MEM_OUT_9_port, DATA_IN(8) => 
                           DATA_MEM_OUT_8_port, DATA_IN(7) => 
                           DATA_MEM_OUT_7_port, DATA_IN(6) => 
                           DATA_MEM_OUT_6_port, DATA_IN(5) => 
                           DATA_MEM_OUT_5_port, DATA_IN(4) => 
                           DATA_MEM_OUT_4_port, DATA_IN(3) => 
                           DATA_MEM_OUT_3_port, DATA_IN(2) => 
                           DATA_MEM_OUT_2_port, DATA_IN(1) => 
                           DATA_MEM_OUT_1_port, DATA_IN(0) => 
                           DATA_MEM_OUT_0_port, ALU_RES_IN(31) => 
                           ALU_RES_MEM_31_port, ALU_RES_IN(30) => 
                           ALU_RES_MEM_30_port, ALU_RES_IN(29) => 
                           ALU_RES_MEM_29_port, ALU_RES_IN(28) => 
                           ALU_RES_MEM_28_port, ALU_RES_IN(27) => 
                           ALU_RES_MEM_27_port, ALU_RES_IN(26) => 
                           ALU_RES_MEM_26_port, ALU_RES_IN(25) => 
                           ALU_RES_MEM_25_port, ALU_RES_IN(24) => 
                           ALU_RES_MEM_24_port, ALU_RES_IN(23) => 
                           ALU_RES_MEM_23_port, ALU_RES_IN(22) => 
                           ALU_RES_MEM_22_port, ALU_RES_IN(21) => 
                           ALU_RES_MEM_21_port, ALU_RES_IN(20) => 
                           ALU_RES_MEM_20_port, ALU_RES_IN(19) => 
                           ALU_RES_MEM_19_port, ALU_RES_IN(18) => 
                           ALU_RES_MEM_18_port, ALU_RES_IN(17) => 
                           ALU_RES_MEM_17_port, ALU_RES_IN(16) => 
                           ALU_RES_MEM_16_port, ALU_RES_IN(15) => 
                           ALU_RES_MEM_15_port, ALU_RES_IN(14) => 
                           ALU_RES_MEM_14_port, ALU_RES_IN(13) => 
                           ALU_RES_MEM_13_port, ALU_RES_IN(12) => 
                           ALU_RES_MEM_12_port, ALU_RES_IN(11) => 
                           ALU_RES_MEM_11_port, ALU_RES_IN(10) => 
                           ALU_RES_MEM_10_port, ALU_RES_IN(9) => 
                           ALU_RES_MEM_9_port, ALU_RES_IN(8) => 
                           ALU_RES_MEM_8_port, ALU_RES_IN(7) => 
                           ALU_RES_MEM_7_port, ALU_RES_IN(6) => 
                           ALU_RES_MEM_6_port, ALU_RES_IN(5) => 
                           ALU_RES_MEM_5_port, ALU_RES_IN(4) => 
                           ALU_RES_MEM_4_port, ALU_RES_IN(3) => 
                           ALU_RES_MEM_3_port, ALU_RES_IN(2) => 
                           ALU_RES_MEM_2_port, ALU_RES_IN(1) => 
                           ALU_RES_MEM_1_port, ALU_RES_IN(0) => 
                           ALU_RES_MEM_0_port, ADD_WR_IN(4) => 
                           ADD_WR_MEM_OUT_4_port, ADD_WR_IN(3) => 
                           ADD_WR_MEM_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_MEM_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_MEM_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_MEM_OUT_0_port, DATA_OUT(31) => OP_WB_31_port
                           , DATA_OUT(30) => OP_WB_30_port, DATA_OUT(29) => 
                           OP_WB_29_port, DATA_OUT(28) => OP_WB_28_port, 
                           DATA_OUT(27) => OP_WB_27_port, DATA_OUT(26) => 
                           OP_WB_26_port, DATA_OUT(25) => OP_WB_25_port, 
                           DATA_OUT(24) => OP_WB_24_port, DATA_OUT(23) => 
                           OP_WB_23_port, DATA_OUT(22) => OP_WB_22_port, 
                           DATA_OUT(21) => OP_WB_21_port, DATA_OUT(20) => 
                           OP_WB_20_port, DATA_OUT(19) => OP_WB_19_port, 
                           DATA_OUT(18) => OP_WB_18_port, DATA_OUT(17) => 
                           OP_WB_17_port, DATA_OUT(16) => OP_WB_16_port, 
                           DATA_OUT(15) => OP_WB_15_port, DATA_OUT(14) => 
                           OP_WB_14_port, DATA_OUT(13) => OP_WB_13_port, 
                           DATA_OUT(12) => OP_WB_12_port, DATA_OUT(11) => 
                           OP_WB_11_port, DATA_OUT(10) => OP_WB_10_port, 
                           DATA_OUT(9) => OP_WB_9_port, DATA_OUT(8) => 
                           OP_WB_8_port, DATA_OUT(7) => OP_WB_7_port, 
                           DATA_OUT(6) => OP_WB_6_port, DATA_OUT(5) => 
                           OP_WB_5_port, DATA_OUT(4) => OP_WB_4_port, 
                           DATA_OUT(3) => OP_WB_3_port, DATA_OUT(2) => 
                           OP_WB_2_port, DATA_OUT(1) => OP_WB_1_port, 
                           DATA_OUT(0) => OP_WB_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_WB_4_port, ADD_WR_OUT(3) => ADD_WR_WB_3_port,
                           ADD_WR_OUT(2) => ADD_WR_WB_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_WB_1_port, ADD_WR_OUT(0) => ADD_WR_WB_0_port)
                           ;
   HDU : HazardDetection port map( RST => RST, ADD_RS1(4) => ADD_RS1_HDU_4_port
                           , ADD_RS1(3) => ADD_RS1_HDU_3_port, ADD_RS1(2) => 
                           ADD_RS1_HDU_2_port, ADD_RS1(1) => ADD_RS1_HDU_1_port
                           , ADD_RS1(0) => ADD_RS1_HDU_0_port, ADD_RS2(4) => 
                           ADD_RS2_HDU_4_port, ADD_RS2(3) => ADD_RS2_HDU_3_port
                           , ADD_RS2(2) => ADD_RS2_HDU_2_port, ADD_RS2(1) => 
                           ADD_RS2_HDU_1_port, ADD_RS2(0) => ADD_RS2_HDU_0_port
                           , ADD_WR(4) => ADD_WR_DECODE_OUT_4_port, ADD_WR(3) 
                           => ADD_WR_DECODE_OUT_3_port, ADD_WR(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR(0) => 
                           ADD_WR_DECODE_OUT_0_port, DRAM_R => DRAM_R_IN, 
                           INS_IN(31) => INS_OUT_31_port, INS_IN(30) => 
                           INS_OUT_30_port, INS_IN(29) => INS_OUT_29_port, 
                           INS_IN(28) => INS_OUT_28_port, INS_IN(27) => 
                           INS_OUT_27_port, INS_IN(26) => INS_OUT_26_port, 
                           INS_IN(25) => INS_OUT_25_port, INS_IN(24) => 
                           INS_OUT_24_port, INS_IN(23) => INS_OUT_23_port, 
                           INS_IN(22) => INS_OUT_22_port, INS_IN(21) => 
                           INS_OUT_21_port, INS_IN(20) => INS_OUT_20_port, 
                           INS_IN(19) => INS_OUT_19_port, INS_IN(18) => 
                           INS_OUT_18_port, INS_IN(17) => INS_OUT_17_port, 
                           INS_IN(16) => INS_OUT_16_port, INS_IN(15) => 
                           INS_OUT_15_port, INS_IN(14) => INS_OUT_14_port, 
                           INS_IN(13) => INS_OUT_13_port, INS_IN(12) => 
                           INS_OUT_12_port, INS_IN(11) => INS_OUT_11_port, 
                           INS_IN(10) => INS_OUT_10_port, INS_IN(9) => 
                           INS_OUT_9_port, INS_IN(8) => INS_OUT_8_port, 
                           INS_IN(7) => INS_OUT_7_port, INS_IN(6) => 
                           INS_OUT_6_port, INS_IN(5) => INS_OUT_5_port, 
                           INS_IN(4) => INS_OUT_4_port, INS_IN(3) => 
                           INS_OUT_3_port, INS_IN(2) => INS_OUT_2_port, 
                           INS_IN(1) => INS_OUT_1_port, INS_IN(0) => 
                           INS_OUT_0_port, PC_IN(31) => PC_FETCH_OUT_31_port, 
                           PC_IN(30) => PC_FETCH_OUT_30_port, PC_IN(29) => 
                           PC_FETCH_OUT_29_port, PC_IN(28) => 
                           PC_FETCH_OUT_28_port, PC_IN(27) => 
                           PC_FETCH_OUT_27_port, PC_IN(26) => 
                           PC_FETCH_OUT_26_port, PC_IN(25) => 
                           PC_FETCH_OUT_25_port, PC_IN(24) => 
                           PC_FETCH_OUT_24_port, PC_IN(23) => 
                           PC_FETCH_OUT_23_port, PC_IN(22) => 
                           PC_FETCH_OUT_22_port, PC_IN(21) => 
                           PC_FETCH_OUT_21_port, PC_IN(20) => 
                           PC_FETCH_OUT_20_port, PC_IN(19) => 
                           PC_FETCH_OUT_19_port, PC_IN(18) => 
                           PC_FETCH_OUT_18_port, PC_IN(17) => 
                           PC_FETCH_OUT_17_port, PC_IN(16) => 
                           PC_FETCH_OUT_16_port, PC_IN(15) => 
                           PC_FETCH_OUT_15_port, PC_IN(14) => 
                           PC_FETCH_OUT_14_port, PC_IN(13) => 
                           PC_FETCH_OUT_13_port, PC_IN(12) => 
                           PC_FETCH_OUT_12_port, PC_IN(11) => 
                           PC_FETCH_OUT_11_port, PC_IN(10) => 
                           PC_FETCH_OUT_10_port, PC_IN(9) => 
                           PC_FETCH_OUT_9_port, PC_IN(8) => PC_FETCH_OUT_8_port
                           , PC_IN(7) => PC_FETCH_OUT_7_port, PC_IN(6) => 
                           PC_FETCH_OUT_6_port, PC_IN(5) => PC_FETCH_OUT_5_port
                           , PC_IN(4) => PC_FETCH_OUT_4_port, PC_IN(3) => 
                           PC_FETCH_OUT_3_port, PC_IN(2) => PC_FETCH_OUT_2_port
                           , PC_IN(1) => PC_FETCH_OUT_1_port, PC_IN(0) => 
                           PC_FETCH_OUT_0_port, Bubble => Bubble_out_port, 
                           HDU_INS_OUT(31) => sig_HDU_INS_OUT_31_port, 
                           HDU_INS_OUT(30) => sig_HDU_INS_OUT_30_port, 
                           HDU_INS_OUT(29) => sig_HDU_INS_OUT_29_port, 
                           HDU_INS_OUT(28) => sig_HDU_INS_OUT_28_port, 
                           HDU_INS_OUT(27) => sig_HDU_INS_OUT_27_port, 
                           HDU_INS_OUT(26) => sig_HDU_INS_OUT_26_port, 
                           HDU_INS_OUT(25) => sig_HDU_INS_OUT_25_port, 
                           HDU_INS_OUT(24) => sig_HDU_INS_OUT_24_port, 
                           HDU_INS_OUT(23) => sig_HDU_INS_OUT_23_port, 
                           HDU_INS_OUT(22) => sig_HDU_INS_OUT_22_port, 
                           HDU_INS_OUT(21) => sig_HDU_INS_OUT_21_port, 
                           HDU_INS_OUT(20) => sig_HDU_INS_OUT_20_port, 
                           HDU_INS_OUT(19) => sig_HDU_INS_OUT_19_port, 
                           HDU_INS_OUT(18) => sig_HDU_INS_OUT_18_port, 
                           HDU_INS_OUT(17) => sig_HDU_INS_OUT_17_port, 
                           HDU_INS_OUT(16) => sig_HDU_INS_OUT_16_port, 
                           HDU_INS_OUT(15) => sig_HDU_INS_OUT_15_port, 
                           HDU_INS_OUT(14) => sig_HDU_INS_OUT_14_port, 
                           HDU_INS_OUT(13) => sig_HDU_INS_OUT_13_port, 
                           HDU_INS_OUT(12) => sig_HDU_INS_OUT_12_port, 
                           HDU_INS_OUT(11) => sig_HDU_INS_OUT_11_port, 
                           HDU_INS_OUT(10) => sig_HDU_INS_OUT_10_port, 
                           HDU_INS_OUT(9) => sig_HDU_INS_OUT_9_port, 
                           HDU_INS_OUT(8) => sig_HDU_INS_OUT_8_port, 
                           HDU_INS_OUT(7) => sig_HDU_INS_OUT_7_port, 
                           HDU_INS_OUT(6) => sig_HDU_INS_OUT_6_port, 
                           HDU_INS_OUT(5) => sig_HDU_INS_OUT_5_port, 
                           HDU_INS_OUT(4) => sig_HDU_INS_OUT_4_port, 
                           HDU_INS_OUT(3) => sig_HDU_INS_OUT_3_port, 
                           HDU_INS_OUT(2) => sig_HDU_INS_OUT_2_port, 
                           HDU_INS_OUT(1) => sig_HDU_INS_OUT_1_port, 
                           HDU_INS_OUT(0) => sig_HDU_INS_OUT_0_port, 
                           HDU_PC_OUT(31) => sig_HDU_PC_OUT_31_port, 
                           HDU_PC_OUT(30) => sig_HDU_PC_OUT_30_port, 
                           HDU_PC_OUT(29) => sig_HDU_PC_OUT_29_port, 
                           HDU_PC_OUT(28) => sig_HDU_PC_OUT_28_port, 
                           HDU_PC_OUT(27) => sig_HDU_PC_OUT_27_port, 
                           HDU_PC_OUT(26) => sig_HDU_PC_OUT_26_port, 
                           HDU_PC_OUT(25) => sig_HDU_PC_OUT_25_port, 
                           HDU_PC_OUT(24) => sig_HDU_PC_OUT_24_port, 
                           HDU_PC_OUT(23) => sig_HDU_PC_OUT_23_port, 
                           HDU_PC_OUT(22) => sig_HDU_PC_OUT_22_port, 
                           HDU_PC_OUT(21) => sig_HDU_PC_OUT_21_port, 
                           HDU_PC_OUT(20) => sig_HDU_PC_OUT_20_port, 
                           HDU_PC_OUT(19) => sig_HDU_PC_OUT_19_port, 
                           HDU_PC_OUT(18) => sig_HDU_PC_OUT_18_port, 
                           HDU_PC_OUT(17) => sig_HDU_PC_OUT_17_port, 
                           HDU_PC_OUT(16) => sig_HDU_PC_OUT_16_port, 
                           HDU_PC_OUT(15) => sig_HDU_PC_OUT_15_port, 
                           HDU_PC_OUT(14) => sig_HDU_PC_OUT_14_port, 
                           HDU_PC_OUT(13) => sig_HDU_PC_OUT_13_port, 
                           HDU_PC_OUT(12) => sig_HDU_PC_OUT_12_port, 
                           HDU_PC_OUT(11) => sig_HDU_PC_OUT_11_port, 
                           HDU_PC_OUT(10) => sig_HDU_PC_OUT_10_port, 
                           HDU_PC_OUT(9) => sig_HDU_PC_OUT_9_port, 
                           HDU_PC_OUT(8) => sig_HDU_PC_OUT_8_port, 
                           HDU_PC_OUT(7) => sig_HDU_PC_OUT_7_port, 
                           HDU_PC_OUT(6) => sig_HDU_PC_OUT_6_port, 
                           HDU_PC_OUT(5) => sig_HDU_PC_OUT_5_port, 
                           HDU_PC_OUT(4) => sig_HDU_PC_OUT_4_port, 
                           HDU_PC_OUT(3) => sig_HDU_PC_OUT_3_port, 
                           HDU_PC_OUT(2) => sig_HDU_PC_OUT_2_port, 
                           HDU_PC_OUT(1) => sig_HDU_PC_OUT_1_port, 
                           HDU_PC_OUT(0) => sig_HDU_PC_OUT_0_port, 
                           HDU_NPC_OUT(31) => sig_HDU_NPC_OUT_31_port, 
                           HDU_NPC_OUT(30) => sig_HDU_NPC_OUT_30_port, 
                           HDU_NPC_OUT(29) => sig_HDU_NPC_OUT_29_port, 
                           HDU_NPC_OUT(28) => sig_HDU_NPC_OUT_28_port, 
                           HDU_NPC_OUT(27) => sig_HDU_NPC_OUT_27_port, 
                           HDU_NPC_OUT(26) => sig_HDU_NPC_OUT_26_port, 
                           HDU_NPC_OUT(25) => sig_HDU_NPC_OUT_25_port, 
                           HDU_NPC_OUT(24) => sig_HDU_NPC_OUT_24_port, 
                           HDU_NPC_OUT(23) => sig_HDU_NPC_OUT_23_port, 
                           HDU_NPC_OUT(22) => sig_HDU_NPC_OUT_22_port, 
                           HDU_NPC_OUT(21) => sig_HDU_NPC_OUT_21_port, 
                           HDU_NPC_OUT(20) => sig_HDU_NPC_OUT_20_port, 
                           HDU_NPC_OUT(19) => sig_HDU_NPC_OUT_19_port, 
                           HDU_NPC_OUT(18) => sig_HDU_NPC_OUT_18_port, 
                           HDU_NPC_OUT(17) => sig_HDU_NPC_OUT_17_port, 
                           HDU_NPC_OUT(16) => sig_HDU_NPC_OUT_16_port, 
                           HDU_NPC_OUT(15) => sig_HDU_NPC_OUT_15_port, 
                           HDU_NPC_OUT(14) => sig_HDU_NPC_OUT_14_port, 
                           HDU_NPC_OUT(13) => sig_HDU_NPC_OUT_13_port, 
                           HDU_NPC_OUT(12) => sig_HDU_NPC_OUT_12_port, 
                           HDU_NPC_OUT(11) => sig_HDU_NPC_OUT_11_port, 
                           HDU_NPC_OUT(10) => sig_HDU_NPC_OUT_10_port, 
                           HDU_NPC_OUT(9) => sig_HDU_NPC_OUT_9_port, 
                           HDU_NPC_OUT(8) => sig_HDU_NPC_OUT_8_port, 
                           HDU_NPC_OUT(7) => sig_HDU_NPC_OUT_7_port, 
                           HDU_NPC_OUT(6) => sig_HDU_NPC_OUT_6_port, 
                           HDU_NPC_OUT(5) => sig_HDU_NPC_OUT_5_port, 
                           HDU_NPC_OUT(4) => sig_HDU_NPC_OUT_4_port, 
                           HDU_NPC_OUT(3) => sig_HDU_NPC_OUT_3_port, 
                           HDU_NPC_OUT(2) => sig_HDU_NPC_OUT_2_port, 
                           HDU_NPC_OUT(1) => sig_HDU_NPC_OUT_1_port, 
                           HDU_NPC_OUT(0) => sig_HDU_NPC_OUT_0_port);
   U2 : CLKBUF_X1 port map( A => n7, Z => INS_OUT_29_port);
   U3 : CLKBUF_X1 port map( A => n8, Z => INS_OUT_28_port);
   U4 : CLKBUF_X1 port map( A => n10, Z => INS_OUT_26_port);
   U5 : CLKBUF_X1 port map( A => n6, Z => INS_OUT_31_port);
   U6 : CLKBUF_X1 port map( A => n9, Z => INS_OUT_27_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( Clk, Rst : in std_logic);

end DLX;

architecture SYN_dlx_rtl of DLX is

   component DRAM
      port( Clk, Rst : in std_logic;  ADDR_IN, DATA_IN : in std_logic_vector 
            (31 downto 0);  LOAD_TYPE : in std_logic_vector (1 downto 0);  
            STORE_TYPE, DRAM_W, DRAM_R : in std_logic;  DATA_OUT : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component IRAM
      port( Rst : in std_logic;  Addr : in std_logic_vector (31 downto 0);  
            Iout : out std_logic_vector (31 downto 0));
   end component;
   
   component hardwired_cu_NBIT32
      port( MUX_A_SEL : out std_logic;  MUX_B_SEL : out std_logic_vector (1 
            downto 0);  ALU_OPC : out std_logic_vector (0 to 4);  ALU_OUTREG_EN
            , DRAM_R_IN : out std_logic;  JUMP_TYPE : out std_logic_vector (1 
            downto 0);  MEM_EN_IN, DRAM_W_IN, RF_WE : out std_logic;  
            LOAD_TYPE_IN : out std_logic_vector (1 downto 0);  STORE_TYPE_IN, 
            WB_MUX_SEL : out std_logic;  INS_IN : in std_logic_vector (31 
            downto 0);  Bubble, Clk, Rst : in std_logic);
   end component;
   
   component Datapath
      port( CLK, RST : in std_logic;  INS_IN, DATA_IN : in std_logic_vector (31
            downto 0);  MUX_A_SEL : in std_logic;  MUX_B_SEL : in 
            std_logic_vector (1 downto 0);  ALU_OPC : in std_logic_vector (0 to
            4);  ALU_OUTREG_EN : in std_logic;  JUMP_TYPE : in std_logic_vector
            (1 downto 0);  DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, RF_WE : in 
            std_logic;  LOAD_TYPE_IN : in std_logic_vector (1 downto 0);  
            STORE_TYPE_IN, WB_MUX_SEL : in std_logic;  INS_OUT, IRAM_ADDR_OUT, 
            DRAM_ADDR_OUT, DATA_OUT : out std_logic_vector (31 downto 0);  
            DRAM_R_OUT, DRAM_W_OUT, Bubble_out : out std_logic;  LOAD_TYPE_OUT 
            : out std_logic_vector (1 downto 0);  STORE_TYPE_OUT : out 
            std_logic);
   end component;
   
   signal INS_IN_31_port, INS_IN_30_port, INS_IN_29_port, INS_IN_28_port, 
      INS_IN_27_port, INS_IN_26_port, INS_IN_25_port, INS_IN_24_port, 
      INS_IN_23_port, INS_IN_22_port, INS_IN_21_port, INS_IN_20_port, 
      INS_IN_19_port, INS_IN_18_port, INS_IN_17_port, INS_IN_16_port, 
      INS_IN_15_port, INS_IN_14_port, INS_IN_13_port, INS_IN_12_port, 
      INS_IN_11_port, INS_IN_10_port, INS_IN_9_port, INS_IN_8_port, 
      INS_IN_7_port, INS_IN_6_port, INS_IN_5_port, INS_IN_4_port, INS_IN_3_port
      , INS_IN_2_port, INS_IN_1_port, INS_IN_0_port, DATA_IN_31_port, 
      DATA_IN_30_port, DATA_IN_29_port, DATA_IN_28_port, DATA_IN_27_port, 
      DATA_IN_26_port, DATA_IN_25_port, DATA_IN_24_port, DATA_IN_23_port, 
      DATA_IN_22_port, DATA_IN_21_port, DATA_IN_20_port, DATA_IN_19_port, 
      DATA_IN_18_port, DATA_IN_17_port, DATA_IN_16_port, DATA_IN_15_port, 
      DATA_IN_14_port, DATA_IN_13_port, DATA_IN_12_port, DATA_IN_11_port, 
      DATA_IN_10_port, DATA_IN_9_port, DATA_IN_8_port, DATA_IN_7_port, 
      DATA_IN_6_port, DATA_IN_5_port, DATA_IN_4_port, DATA_IN_3_port, 
      DATA_IN_2_port, DATA_IN_1_port, DATA_IN_0_port, MUX_A_SEL, 
      MUX_B_SEL_1_port, MUX_B_SEL_0_port, ALU_OPC_4_port, ALU_OPC_3_port, 
      ALU_OPC_2_port, ALU_OPC_1_port, ALU_OPC_0_port, ALU_OUTREG_EN, 
      JUMP_TYPE_1_port, JUMP_TYPE_0_port, DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, 
      RF_WE, LOAD_TYPE_IN_1_port, LOAD_TYPE_IN_0_port, STORE_TYPE_IN, 
      WB_MUX_SEL, INST_31_port, INST_30_port, INST_29_port, INST_28_port, 
      INST_27_port, INST_26_port, INST_25_port, INST_24_port, INST_23_port, 
      INST_22_port, INST_21_port, INST_20_port, INST_19_port, INST_18_port, 
      INST_17_port, INST_16_port, INST_15_port, INST_14_port, INST_13_port, 
      INST_12_port, INST_11_port, INST_10_port, INST_9_port, INST_8_port, 
      INST_7_port, INST_6_port, INST_5_port, INST_4_port, INST_3_port, 
      INST_2_port, INST_1_port, INST_0_port, IRAM_ADDR_OUT_31_port, 
      IRAM_ADDR_OUT_30_port, IRAM_ADDR_OUT_29_port, IRAM_ADDR_OUT_28_port, 
      IRAM_ADDR_OUT_27_port, IRAM_ADDR_OUT_26_port, IRAM_ADDR_OUT_25_port, 
      IRAM_ADDR_OUT_24_port, IRAM_ADDR_OUT_23_port, IRAM_ADDR_OUT_22_port, 
      IRAM_ADDR_OUT_21_port, IRAM_ADDR_OUT_20_port, IRAM_ADDR_OUT_19_port, 
      IRAM_ADDR_OUT_18_port, IRAM_ADDR_OUT_17_port, IRAM_ADDR_OUT_16_port, 
      IRAM_ADDR_OUT_15_port, IRAM_ADDR_OUT_14_port, IRAM_ADDR_OUT_13_port, 
      IRAM_ADDR_OUT_12_port, IRAM_ADDR_OUT_11_port, IRAM_ADDR_OUT_10_port, 
      IRAM_ADDR_OUT_9_port, IRAM_ADDR_OUT_8_port, IRAM_ADDR_OUT_7_port, 
      IRAM_ADDR_OUT_6_port, IRAM_ADDR_OUT_5_port, IRAM_ADDR_OUT_4_port, 
      IRAM_ADDR_OUT_3_port, IRAM_ADDR_OUT_2_port, IRAM_ADDR_OUT_1_port, 
      IRAM_ADDR_OUT_0_port, DRAM_ADDR_OUT_31_port, DRAM_ADDR_OUT_30_port, 
      DRAM_ADDR_OUT_29_port, DRAM_ADDR_OUT_28_port, DRAM_ADDR_OUT_27_port, 
      DRAM_ADDR_OUT_26_port, DRAM_ADDR_OUT_25_port, DRAM_ADDR_OUT_24_port, 
      DRAM_ADDR_OUT_23_port, DRAM_ADDR_OUT_22_port, DRAM_ADDR_OUT_21_port, 
      DRAM_ADDR_OUT_20_port, DRAM_ADDR_OUT_19_port, DRAM_ADDR_OUT_18_port, 
      DRAM_ADDR_OUT_17_port, DRAM_ADDR_OUT_16_port, DRAM_ADDR_OUT_15_port, 
      DRAM_ADDR_OUT_14_port, DRAM_ADDR_OUT_13_port, DRAM_ADDR_OUT_12_port, 
      DRAM_ADDR_OUT_11_port, DRAM_ADDR_OUT_10_port, DRAM_ADDR_OUT_9_port, 
      DRAM_ADDR_OUT_8_port, DRAM_ADDR_OUT_7_port, DRAM_ADDR_OUT_6_port, 
      DRAM_ADDR_OUT_5_port, DRAM_ADDR_OUT_4_port, DRAM_ADDR_OUT_3_port, 
      DRAM_ADDR_OUT_2_port, DRAM_ADDR_OUT_1_port, DRAM_ADDR_OUT_0_port, 
      DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, DATA_OUT_28_port, 
      DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, DATA_OUT_24_port, 
      DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, DATA_OUT_20_port, 
      DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, DATA_OUT_16_port, 
      DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, DATA_OUT_12_port, 
      DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, DATA_OUT_8_port, 
      DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, DATA_OUT_4_port, 
      DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, DATA_OUT_0_port, 
      DRAM_R_OUT, DRAM_W_OUT, Bubble, LOAD_TYPE_OUT_1_port, 
      LOAD_TYPE_OUT_0_port, STORE_TYPE_OUT, n_1604, n_1605, n_1606, n_1607, 
      n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, 
      n_1617 : std_logic;

begin
   
   DP : Datapath port map( CLK => Clk, RST => Rst, INS_IN(31) => INS_IN_31_port
                           , INS_IN(30) => INS_IN_30_port, INS_IN(29) => 
                           INS_IN_29_port, INS_IN(28) => INS_IN_28_port, 
                           INS_IN(27) => INS_IN_27_port, INS_IN(26) => 
                           INS_IN_26_port, INS_IN(25) => INS_IN_25_port, 
                           INS_IN(24) => INS_IN_24_port, INS_IN(23) => 
                           INS_IN_23_port, INS_IN(22) => INS_IN_22_port, 
                           INS_IN(21) => INS_IN_21_port, INS_IN(20) => 
                           INS_IN_20_port, INS_IN(19) => INS_IN_19_port, 
                           INS_IN(18) => INS_IN_18_port, INS_IN(17) => 
                           INS_IN_17_port, INS_IN(16) => INS_IN_16_port, 
                           INS_IN(15) => INS_IN_15_port, INS_IN(14) => 
                           INS_IN_14_port, INS_IN(13) => INS_IN_13_port, 
                           INS_IN(12) => INS_IN_12_port, INS_IN(11) => 
                           INS_IN_11_port, INS_IN(10) => INS_IN_10_port, 
                           INS_IN(9) => INS_IN_9_port, INS_IN(8) => 
                           INS_IN_8_port, INS_IN(7) => INS_IN_7_port, INS_IN(6)
                           => INS_IN_6_port, INS_IN(5) => INS_IN_5_port, 
                           INS_IN(4) => INS_IN_4_port, INS_IN(3) => 
                           INS_IN_3_port, INS_IN(2) => INS_IN_2_port, INS_IN(1)
                           => INS_IN_1_port, INS_IN(0) => INS_IN_0_port, 
                           DATA_IN(31) => DATA_IN_31_port, DATA_IN(30) => 
                           DATA_IN_30_port, DATA_IN(29) => DATA_IN_29_port, 
                           DATA_IN(28) => DATA_IN_28_port, DATA_IN(27) => 
                           DATA_IN_27_port, DATA_IN(26) => DATA_IN_26_port, 
                           DATA_IN(25) => DATA_IN_25_port, DATA_IN(24) => 
                           DATA_IN_24_port, DATA_IN(23) => DATA_IN_23_port, 
                           DATA_IN(22) => DATA_IN_22_port, DATA_IN(21) => 
                           DATA_IN_21_port, DATA_IN(20) => DATA_IN_20_port, 
                           DATA_IN(19) => DATA_IN_19_port, DATA_IN(18) => 
                           DATA_IN_18_port, DATA_IN(17) => DATA_IN_17_port, 
                           DATA_IN(16) => DATA_IN_16_port, DATA_IN(15) => 
                           DATA_IN_15_port, DATA_IN(14) => DATA_IN_14_port, 
                           DATA_IN(13) => DATA_IN_13_port, DATA_IN(12) => 
                           DATA_IN_12_port, DATA_IN(11) => DATA_IN_11_port, 
                           DATA_IN(10) => DATA_IN_10_port, DATA_IN(9) => 
                           DATA_IN_9_port, DATA_IN(8) => DATA_IN_8_port, 
                           DATA_IN(7) => DATA_IN_7_port, DATA_IN(6) => 
                           DATA_IN_6_port, DATA_IN(5) => DATA_IN_5_port, 
                           DATA_IN(4) => DATA_IN_4_port, DATA_IN(3) => 
                           DATA_IN_3_port, DATA_IN(2) => DATA_IN_2_port, 
                           DATA_IN(1) => DATA_IN_1_port, DATA_IN(0) => 
                           DATA_IN_0_port, MUX_A_SEL => MUX_A_SEL, MUX_B_SEL(1)
                           => MUX_B_SEL_1_port, MUX_B_SEL(0) => 
                           MUX_B_SEL_0_port, ALU_OPC(0) => ALU_OPC_4_port, 
                           ALU_OPC(1) => ALU_OPC_3_port, ALU_OPC(2) => 
                           ALU_OPC_2_port, ALU_OPC(3) => ALU_OPC_1_port, 
                           ALU_OPC(4) => ALU_OPC_0_port, ALU_OUTREG_EN => 
                           ALU_OUTREG_EN, JUMP_TYPE(1) => JUMP_TYPE_1_port, 
                           JUMP_TYPE(0) => JUMP_TYPE_0_port, DRAM_R_IN => 
                           DRAM_R_IN, MEM_EN_IN => MEM_EN_IN, DRAM_W_IN => 
                           DRAM_W_IN, RF_WE => RF_WE, LOAD_TYPE_IN(1) => 
                           LOAD_TYPE_IN_1_port, LOAD_TYPE_IN(0) => 
                           LOAD_TYPE_IN_0_port, STORE_TYPE_IN => STORE_TYPE_IN,
                           WB_MUX_SEL => WB_MUX_SEL, INS_OUT(31) => 
                           INST_31_port, INS_OUT(30) => INST_30_port, 
                           INS_OUT(29) => INST_29_port, INS_OUT(28) => 
                           INST_28_port, INS_OUT(27) => INST_27_port, 
                           INS_OUT(26) => INST_26_port, INS_OUT(25) => 
                           INST_25_port, INS_OUT(24) => INST_24_port, 
                           INS_OUT(23) => INST_23_port, INS_OUT(22) => 
                           INST_22_port, INS_OUT(21) => INST_21_port, 
                           INS_OUT(20) => INST_20_port, INS_OUT(19) => 
                           INST_19_port, INS_OUT(18) => INST_18_port, 
                           INS_OUT(17) => INST_17_port, INS_OUT(16) => 
                           INST_16_port, INS_OUT(15) => INST_15_port, 
                           INS_OUT(14) => INST_14_port, INS_OUT(13) => 
                           INST_13_port, INS_OUT(12) => INST_12_port, 
                           INS_OUT(11) => INST_11_port, INS_OUT(10) => 
                           INST_10_port, INS_OUT(9) => INST_9_port, INS_OUT(8) 
                           => INST_8_port, INS_OUT(7) => INST_7_port, 
                           INS_OUT(6) => INST_6_port, INS_OUT(5) => INST_5_port
                           , INS_OUT(4) => INST_4_port, INS_OUT(3) => 
                           INST_3_port, INS_OUT(2) => INST_2_port, INS_OUT(1) 
                           => INST_1_port, INS_OUT(0) => INST_0_port, 
                           IRAM_ADDR_OUT(31) => IRAM_ADDR_OUT_31_port, 
                           IRAM_ADDR_OUT(30) => IRAM_ADDR_OUT_30_port, 
                           IRAM_ADDR_OUT(29) => IRAM_ADDR_OUT_29_port, 
                           IRAM_ADDR_OUT(28) => IRAM_ADDR_OUT_28_port, 
                           IRAM_ADDR_OUT(27) => IRAM_ADDR_OUT_27_port, 
                           IRAM_ADDR_OUT(26) => IRAM_ADDR_OUT_26_port, 
                           IRAM_ADDR_OUT(25) => IRAM_ADDR_OUT_25_port, 
                           IRAM_ADDR_OUT(24) => IRAM_ADDR_OUT_24_port, 
                           IRAM_ADDR_OUT(23) => IRAM_ADDR_OUT_23_port, 
                           IRAM_ADDR_OUT(22) => IRAM_ADDR_OUT_22_port, 
                           IRAM_ADDR_OUT(21) => IRAM_ADDR_OUT_21_port, 
                           IRAM_ADDR_OUT(20) => IRAM_ADDR_OUT_20_port, 
                           IRAM_ADDR_OUT(19) => IRAM_ADDR_OUT_19_port, 
                           IRAM_ADDR_OUT(18) => IRAM_ADDR_OUT_18_port, 
                           IRAM_ADDR_OUT(17) => IRAM_ADDR_OUT_17_port, 
                           IRAM_ADDR_OUT(16) => IRAM_ADDR_OUT_16_port, 
                           IRAM_ADDR_OUT(15) => IRAM_ADDR_OUT_15_port, 
                           IRAM_ADDR_OUT(14) => IRAM_ADDR_OUT_14_port, 
                           IRAM_ADDR_OUT(13) => IRAM_ADDR_OUT_13_port, 
                           IRAM_ADDR_OUT(12) => IRAM_ADDR_OUT_12_port, 
                           IRAM_ADDR_OUT(11) => IRAM_ADDR_OUT_11_port, 
                           IRAM_ADDR_OUT(10) => IRAM_ADDR_OUT_10_port, 
                           IRAM_ADDR_OUT(9) => IRAM_ADDR_OUT_9_port, 
                           IRAM_ADDR_OUT(8) => IRAM_ADDR_OUT_8_port, 
                           IRAM_ADDR_OUT(7) => IRAM_ADDR_OUT_7_port, 
                           IRAM_ADDR_OUT(6) => IRAM_ADDR_OUT_6_port, 
                           IRAM_ADDR_OUT(5) => IRAM_ADDR_OUT_5_port, 
                           IRAM_ADDR_OUT(4) => IRAM_ADDR_OUT_4_port, 
                           IRAM_ADDR_OUT(3) => IRAM_ADDR_OUT_3_port, 
                           IRAM_ADDR_OUT(2) => IRAM_ADDR_OUT_2_port, 
                           IRAM_ADDR_OUT(1) => IRAM_ADDR_OUT_1_port, 
                           IRAM_ADDR_OUT(0) => IRAM_ADDR_OUT_0_port, 
                           DRAM_ADDR_OUT(31) => DRAM_ADDR_OUT_31_port, 
                           DRAM_ADDR_OUT(30) => DRAM_ADDR_OUT_30_port, 
                           DRAM_ADDR_OUT(29) => DRAM_ADDR_OUT_29_port, 
                           DRAM_ADDR_OUT(28) => DRAM_ADDR_OUT_28_port, 
                           DRAM_ADDR_OUT(27) => DRAM_ADDR_OUT_27_port, 
                           DRAM_ADDR_OUT(26) => DRAM_ADDR_OUT_26_port, 
                           DRAM_ADDR_OUT(25) => DRAM_ADDR_OUT_25_port, 
                           DRAM_ADDR_OUT(24) => DRAM_ADDR_OUT_24_port, 
                           DRAM_ADDR_OUT(23) => DRAM_ADDR_OUT_23_port, 
                           DRAM_ADDR_OUT(22) => DRAM_ADDR_OUT_22_port, 
                           DRAM_ADDR_OUT(21) => DRAM_ADDR_OUT_21_port, 
                           DRAM_ADDR_OUT(20) => DRAM_ADDR_OUT_20_port, 
                           DRAM_ADDR_OUT(19) => DRAM_ADDR_OUT_19_port, 
                           DRAM_ADDR_OUT(18) => DRAM_ADDR_OUT_18_port, 
                           DRAM_ADDR_OUT(17) => DRAM_ADDR_OUT_17_port, 
                           DRAM_ADDR_OUT(16) => DRAM_ADDR_OUT_16_port, 
                           DRAM_ADDR_OUT(15) => DRAM_ADDR_OUT_15_port, 
                           DRAM_ADDR_OUT(14) => DRAM_ADDR_OUT_14_port, 
                           DRAM_ADDR_OUT(13) => DRAM_ADDR_OUT_13_port, 
                           DRAM_ADDR_OUT(12) => DRAM_ADDR_OUT_12_port, 
                           DRAM_ADDR_OUT(11) => DRAM_ADDR_OUT_11_port, 
                           DRAM_ADDR_OUT(10) => DRAM_ADDR_OUT_10_port, 
                           DRAM_ADDR_OUT(9) => DRAM_ADDR_OUT_9_port, 
                           DRAM_ADDR_OUT(8) => DRAM_ADDR_OUT_8_port, 
                           DRAM_ADDR_OUT(7) => DRAM_ADDR_OUT_7_port, 
                           DRAM_ADDR_OUT(6) => DRAM_ADDR_OUT_6_port, 
                           DRAM_ADDR_OUT(5) => DRAM_ADDR_OUT_5_port, 
                           DRAM_ADDR_OUT(4) => DRAM_ADDR_OUT_4_port, 
                           DRAM_ADDR_OUT(3) => DRAM_ADDR_OUT_3_port, 
                           DRAM_ADDR_OUT(2) => DRAM_ADDR_OUT_2_port, 
                           DRAM_ADDR_OUT(1) => DRAM_ADDR_OUT_1_port, 
                           DRAM_ADDR_OUT(0) => DRAM_ADDR_OUT_0_port, 
                           DATA_OUT(31) => DATA_OUT_31_port, DATA_OUT(30) => 
                           DATA_OUT_30_port, DATA_OUT(29) => DATA_OUT_29_port, 
                           DATA_OUT(28) => DATA_OUT_28_port, DATA_OUT(27) => 
                           DATA_OUT_27_port, DATA_OUT(26) => DATA_OUT_26_port, 
                           DATA_OUT(25) => DATA_OUT_25_port, DATA_OUT(24) => 
                           DATA_OUT_24_port, DATA_OUT(23) => DATA_OUT_23_port, 
                           DATA_OUT(22) => DATA_OUT_22_port, DATA_OUT(21) => 
                           DATA_OUT_21_port, DATA_OUT(20) => DATA_OUT_20_port, 
                           DATA_OUT(19) => DATA_OUT_19_port, DATA_OUT(18) => 
                           DATA_OUT_18_port, DATA_OUT(17) => DATA_OUT_17_port, 
                           DATA_OUT(16) => DATA_OUT_16_port, DATA_OUT(15) => 
                           DATA_OUT_15_port, DATA_OUT(14) => DATA_OUT_14_port, 
                           DATA_OUT(13) => DATA_OUT_13_port, DATA_OUT(12) => 
                           DATA_OUT_12_port, DATA_OUT(11) => DATA_OUT_11_port, 
                           DATA_OUT(10) => DATA_OUT_10_port, DATA_OUT(9) => 
                           DATA_OUT_9_port, DATA_OUT(8) => DATA_OUT_8_port, 
                           DATA_OUT(7) => DATA_OUT_7_port, DATA_OUT(6) => 
                           DATA_OUT_6_port, DATA_OUT(5) => DATA_OUT_5_port, 
                           DATA_OUT(4) => DATA_OUT_4_port, DATA_OUT(3) => 
                           DATA_OUT_3_port, DATA_OUT(2) => DATA_OUT_2_port, 
                           DATA_OUT(1) => DATA_OUT_1_port, DATA_OUT(0) => 
                           DATA_OUT_0_port, DRAM_R_OUT => DRAM_R_OUT, 
                           DRAM_W_OUT => DRAM_W_OUT, Bubble_out => Bubble, 
                           LOAD_TYPE_OUT(1) => LOAD_TYPE_OUT_1_port, 
                           LOAD_TYPE_OUT(0) => LOAD_TYPE_OUT_0_port, 
                           STORE_TYPE_OUT => STORE_TYPE_OUT);
   CU : hardwired_cu_NBIT32 port map( MUX_A_SEL => n_1604, MUX_B_SEL(1) => 
                           n_1605, MUX_B_SEL(0) => n_1606, ALU_OPC(0) => 
                           ALU_OPC_4_port, ALU_OPC(1) => ALU_OPC_3_port, 
                           ALU_OPC(2) => ALU_OPC_2_port, ALU_OPC(3) => 
                           ALU_OPC_1_port, ALU_OPC(4) => ALU_OPC_0_port, 
                           ALU_OUTREG_EN => n_1607, DRAM_R_IN => n_1608, 
                           JUMP_TYPE(1) => n_1609, JUMP_TYPE(0) => n_1610, 
                           MEM_EN_IN => n_1611, DRAM_W_IN => n_1612, RF_WE => 
                           n_1613, LOAD_TYPE_IN(1) => n_1614, LOAD_TYPE_IN(0) 
                           => n_1615, STORE_TYPE_IN => n_1616, WB_MUX_SEL => 
                           n_1617, INS_IN(31) => INST_31_port, INS_IN(30) => 
                           INST_30_port, INS_IN(29) => INST_29_port, INS_IN(28)
                           => INST_28_port, INS_IN(27) => INST_27_port, 
                           INS_IN(26) => INST_26_port, INS_IN(25) => 
                           INST_25_port, INS_IN(24) => INST_24_port, INS_IN(23)
                           => INST_23_port, INS_IN(22) => INST_22_port, 
                           INS_IN(21) => INST_21_port, INS_IN(20) => 
                           INST_20_port, INS_IN(19) => INST_19_port, INS_IN(18)
                           => INST_18_port, INS_IN(17) => INST_17_port, 
                           INS_IN(16) => INST_16_port, INS_IN(15) => 
                           INST_15_port, INS_IN(14) => INST_14_port, INS_IN(13)
                           => INST_13_port, INS_IN(12) => INST_12_port, 
                           INS_IN(11) => INST_11_port, INS_IN(10) => 
                           INST_10_port, INS_IN(9) => INST_9_port, INS_IN(8) =>
                           INST_8_port, INS_IN(7) => INST_7_port, INS_IN(6) => 
                           INST_6_port, INS_IN(5) => INST_5_port, INS_IN(4) => 
                           INST_4_port, INS_IN(3) => INST_3_port, INS_IN(2) => 
                           INST_2_port, INS_IN(1) => INST_1_port, INS_IN(0) => 
                           INST_0_port, Bubble => Bubble, Clk => Clk, Rst => 
                           Rst);
   IRAM_I : IRAM port map( Rst => Rst, Addr(31) => IRAM_ADDR_OUT_31_port, 
                           Addr(30) => IRAM_ADDR_OUT_30_port, Addr(29) => 
                           IRAM_ADDR_OUT_29_port, Addr(28) => 
                           IRAM_ADDR_OUT_28_port, Addr(27) => 
                           IRAM_ADDR_OUT_27_port, Addr(26) => 
                           IRAM_ADDR_OUT_26_port, Addr(25) => 
                           IRAM_ADDR_OUT_25_port, Addr(24) => 
                           IRAM_ADDR_OUT_24_port, Addr(23) => 
                           IRAM_ADDR_OUT_23_port, Addr(22) => 
                           IRAM_ADDR_OUT_22_port, Addr(21) => 
                           IRAM_ADDR_OUT_21_port, Addr(20) => 
                           IRAM_ADDR_OUT_20_port, Addr(19) => 
                           IRAM_ADDR_OUT_19_port, Addr(18) => 
                           IRAM_ADDR_OUT_18_port, Addr(17) => 
                           IRAM_ADDR_OUT_17_port, Addr(16) => 
                           IRAM_ADDR_OUT_16_port, Addr(15) => 
                           IRAM_ADDR_OUT_15_port, Addr(14) => 
                           IRAM_ADDR_OUT_14_port, Addr(13) => 
                           IRAM_ADDR_OUT_13_port, Addr(12) => 
                           IRAM_ADDR_OUT_12_port, Addr(11) => 
                           IRAM_ADDR_OUT_11_port, Addr(10) => 
                           IRAM_ADDR_OUT_10_port, Addr(9) => 
                           IRAM_ADDR_OUT_9_port, Addr(8) => 
                           IRAM_ADDR_OUT_8_port, Addr(7) => 
                           IRAM_ADDR_OUT_7_port, Addr(6) => 
                           IRAM_ADDR_OUT_6_port, Addr(5) => 
                           IRAM_ADDR_OUT_5_port, Addr(4) => 
                           IRAM_ADDR_OUT_4_port, Addr(3) => 
                           IRAM_ADDR_OUT_3_port, Addr(2) => 
                           IRAM_ADDR_OUT_2_port, Addr(1) => 
                           IRAM_ADDR_OUT_1_port, Addr(0) => 
                           IRAM_ADDR_OUT_0_port, Iout(31) => INS_IN_31_port, 
                           Iout(30) => INS_IN_30_port, Iout(29) => 
                           INS_IN_29_port, Iout(28) => INS_IN_28_port, Iout(27)
                           => INS_IN_27_port, Iout(26) => INS_IN_26_port, 
                           Iout(25) => INS_IN_25_port, Iout(24) => 
                           INS_IN_24_port, Iout(23) => INS_IN_23_port, Iout(22)
                           => INS_IN_22_port, Iout(21) => INS_IN_21_port, 
                           Iout(20) => INS_IN_20_port, Iout(19) => 
                           INS_IN_19_port, Iout(18) => INS_IN_18_port, Iout(17)
                           => INS_IN_17_port, Iout(16) => INS_IN_16_port, 
                           Iout(15) => INS_IN_15_port, Iout(14) => 
                           INS_IN_14_port, Iout(13) => INS_IN_13_port, Iout(12)
                           => INS_IN_12_port, Iout(11) => INS_IN_11_port, 
                           Iout(10) => INS_IN_10_port, Iout(9) => INS_IN_9_port
                           , Iout(8) => INS_IN_8_port, Iout(7) => INS_IN_7_port
                           , Iout(6) => INS_IN_6_port, Iout(5) => INS_IN_5_port
                           , Iout(4) => INS_IN_4_port, Iout(3) => INS_IN_3_port
                           , Iout(2) => INS_IN_2_port, Iout(1) => INS_IN_1_port
                           , Iout(0) => INS_IN_0_port);
   DRAM_I : DRAM port map( Clk => Clk, Rst => Rst, ADDR_IN(31) => 
                           DRAM_ADDR_OUT_31_port, ADDR_IN(30) => 
                           DRAM_ADDR_OUT_30_port, ADDR_IN(29) => 
                           DRAM_ADDR_OUT_29_port, ADDR_IN(28) => 
                           DRAM_ADDR_OUT_28_port, ADDR_IN(27) => 
                           DRAM_ADDR_OUT_27_port, ADDR_IN(26) => 
                           DRAM_ADDR_OUT_26_port, ADDR_IN(25) => 
                           DRAM_ADDR_OUT_25_port, ADDR_IN(24) => 
                           DRAM_ADDR_OUT_24_port, ADDR_IN(23) => 
                           DRAM_ADDR_OUT_23_port, ADDR_IN(22) => 
                           DRAM_ADDR_OUT_22_port, ADDR_IN(21) => 
                           DRAM_ADDR_OUT_21_port, ADDR_IN(20) => 
                           DRAM_ADDR_OUT_20_port, ADDR_IN(19) => 
                           DRAM_ADDR_OUT_19_port, ADDR_IN(18) => 
                           DRAM_ADDR_OUT_18_port, ADDR_IN(17) => 
                           DRAM_ADDR_OUT_17_port, ADDR_IN(16) => 
                           DRAM_ADDR_OUT_16_port, ADDR_IN(15) => 
                           DRAM_ADDR_OUT_15_port, ADDR_IN(14) => 
                           DRAM_ADDR_OUT_14_port, ADDR_IN(13) => 
                           DRAM_ADDR_OUT_13_port, ADDR_IN(12) => 
                           DRAM_ADDR_OUT_12_port, ADDR_IN(11) => 
                           DRAM_ADDR_OUT_11_port, ADDR_IN(10) => 
                           DRAM_ADDR_OUT_10_port, ADDR_IN(9) => 
                           DRAM_ADDR_OUT_9_port, ADDR_IN(8) => 
                           DRAM_ADDR_OUT_8_port, ADDR_IN(7) => 
                           DRAM_ADDR_OUT_7_port, ADDR_IN(6) => 
                           DRAM_ADDR_OUT_6_port, ADDR_IN(5) => 
                           DRAM_ADDR_OUT_5_port, ADDR_IN(4) => 
                           DRAM_ADDR_OUT_4_port, ADDR_IN(3) => 
                           DRAM_ADDR_OUT_3_port, ADDR_IN(2) => 
                           DRAM_ADDR_OUT_2_port, ADDR_IN(1) => 
                           DRAM_ADDR_OUT_1_port, ADDR_IN(0) => 
                           DRAM_ADDR_OUT_0_port, DATA_IN(31) => 
                           DATA_OUT_31_port, DATA_IN(30) => DATA_OUT_30_port, 
                           DATA_IN(29) => DATA_OUT_29_port, DATA_IN(28) => 
                           DATA_OUT_28_port, DATA_IN(27) => DATA_OUT_27_port, 
                           DATA_IN(26) => DATA_OUT_26_port, DATA_IN(25) => 
                           DATA_OUT_25_port, DATA_IN(24) => DATA_OUT_24_port, 
                           DATA_IN(23) => DATA_OUT_23_port, DATA_IN(22) => 
                           DATA_OUT_22_port, DATA_IN(21) => DATA_OUT_21_port, 
                           DATA_IN(20) => DATA_OUT_20_port, DATA_IN(19) => 
                           DATA_OUT_19_port, DATA_IN(18) => DATA_OUT_18_port, 
                           DATA_IN(17) => DATA_OUT_17_port, DATA_IN(16) => 
                           DATA_OUT_16_port, DATA_IN(15) => DATA_OUT_15_port, 
                           DATA_IN(14) => DATA_OUT_14_port, DATA_IN(13) => 
                           DATA_OUT_13_port, DATA_IN(12) => DATA_OUT_12_port, 
                           DATA_IN(11) => DATA_OUT_11_port, DATA_IN(10) => 
                           DATA_OUT_10_port, DATA_IN(9) => DATA_OUT_9_port, 
                           DATA_IN(8) => DATA_OUT_8_port, DATA_IN(7) => 
                           DATA_OUT_7_port, DATA_IN(6) => DATA_OUT_6_port, 
                           DATA_IN(5) => DATA_OUT_5_port, DATA_IN(4) => 
                           DATA_OUT_4_port, DATA_IN(3) => DATA_OUT_3_port, 
                           DATA_IN(2) => DATA_OUT_2_port, DATA_IN(1) => 
                           DATA_OUT_1_port, DATA_IN(0) => DATA_OUT_0_port, 
                           LOAD_TYPE(1) => LOAD_TYPE_OUT_1_port, LOAD_TYPE(0) 
                           => LOAD_TYPE_OUT_0_port, STORE_TYPE => 
                           STORE_TYPE_OUT, DRAM_W => DRAM_W_OUT, DRAM_R => 
                           DRAM_R_OUT, DATA_OUT(31) => DATA_IN_31_port, 
                           DATA_OUT(30) => DATA_IN_30_port, DATA_OUT(29) => 
                           DATA_IN_29_port, DATA_OUT(28) => DATA_IN_28_port, 
                           DATA_OUT(27) => DATA_IN_27_port, DATA_OUT(26) => 
                           DATA_IN_26_port, DATA_OUT(25) => DATA_IN_25_port, 
                           DATA_OUT(24) => DATA_IN_24_port, DATA_OUT(23) => 
                           DATA_IN_23_port, DATA_OUT(22) => DATA_IN_22_port, 
                           DATA_OUT(21) => DATA_IN_21_port, DATA_OUT(20) => 
                           DATA_IN_20_port, DATA_OUT(19) => DATA_IN_19_port, 
                           DATA_OUT(18) => DATA_IN_18_port, DATA_OUT(17) => 
                           DATA_IN_17_port, DATA_OUT(16) => DATA_IN_16_port, 
                           DATA_OUT(15) => DATA_IN_15_port, DATA_OUT(14) => 
                           DATA_IN_14_port, DATA_OUT(13) => DATA_IN_13_port, 
                           DATA_OUT(12) => DATA_IN_12_port, DATA_OUT(11) => 
                           DATA_IN_11_port, DATA_OUT(10) => DATA_IN_10_port, 
                           DATA_OUT(9) => DATA_IN_9_port, DATA_OUT(8) => 
                           DATA_IN_8_port, DATA_OUT(7) => DATA_IN_7_port, 
                           DATA_OUT(6) => DATA_IN_6_port, DATA_OUT(5) => 
                           DATA_IN_5_port, DATA_OUT(4) => DATA_IN_4_port, 
                           DATA_OUT(3) => DATA_IN_3_port, DATA_OUT(2) => 
                           DATA_IN_2_port, DATA_OUT(1) => DATA_IN_1_port, 
                           DATA_OUT(0) => DATA_IN_0_port);
   WB_MUX_SEL <= '0';
   STORE_TYPE_IN <= '0';
   LOAD_TYPE_IN_0_port <= '0';
   LOAD_TYPE_IN_1_port <= '0';
   RF_WE <= '0';
   DRAM_W_IN <= '0';
   MEM_EN_IN <= '0';
   JUMP_TYPE_0_port <= '0';
   JUMP_TYPE_1_port <= '0';
   DRAM_R_IN <= '0';
   ALU_OUTREG_EN <= '0';
   MUX_B_SEL_0_port <= '0';
   MUX_B_SEL_1_port <= '0';
   MUX_A_SEL <= '0';

end SYN_dlx_rtl;
