
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type VHDLOUT_TYPE is range 0 to 5;
type aluOp is (NOP, ADDS, ADDUS, SUBS, SUBUS, MULTS, ANDS, ORS, XORS, SLLS, 
   SRLS, SRAS, BEQZS, BNEZS, SGES, SGEUS, SGTS, SGTUS, SLES, SLTS, SLTUS, SEQS,
   NEQS, LHIS);
attribute ENUM_ENCODING of aluOp : type is 
   "00000 00001 00010 00011 00100 00101 00110 00111 01000 01001 01010 01011 01100 01101 01110 01111 10000 10001 10010 10011 10100 10101 10110 10111";
   
   -- Declarations for conversion functions.
   function integer_to_unsigned(arg, size : in INTEGER) return std_logic_vector
               ;
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
               return aluOp;
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX;

package body CONV_PACK_DLX is
   
   -- integer type to std_logic_vector function
   function integer_to_unsigned(arg, size : in INTEGER) return std_logic_vector
   is 
      variable result: std_logic_vector(size-1 downto 0);
      variable temp: INTEGER;
      -- synopsys built_in SYN_INTEGER_TO_UNSIGNED
   begin
      temp := arg;
      for i in 0 to size-1 loop
         if (temp mod 2) = 1 then
            result(i) := '1';
         else
            result(i) := '0';
         end if;
         temp := temp / 2;
      end loop;
      return result;
   end;
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
   return aluOp is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "00000" => return NOP;
         when "00001" => return ADDS;
         when "00010" => return ADDUS;
         when "00011" => return SUBS;
         when "00100" => return SUBUS;
         when "00101" => return MULTS;
         when "00110" => return ANDS;
         when "00111" => return ORS;
         when "01000" => return XORS;
         when "01001" => return SLLS;
         when "01010" => return SRLS;
         when "01011" => return SRAS;
         when "01100" => return BEQZS;
         when "01101" => return BNEZS;
         when "01110" => return SGES;
         when "01111" => return SGEUS;
         when "10000" => return SGTS;
         when "10001" => return SGTUS;
         when "10010" => return SLES;
         when "10011" => return SLTS;
         when "10100" => return SLTUS;
         when "10101" => return SEQS;
         when "10110" => return NEQS;
         when "10111" => return LHIS;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "00000";
         when ADDS => return "00001";
         when ADDUS => return "00010";
         when SUBS => return "00011";
         when SUBUS => return "00100";
         when MULTS => return "00101";
         when ANDS => return "00110";
         when ORS => return "00111";
         when XORS => return "01000";
         when SLLS => return "01001";
         when SRLS => return "01010";
         when SRAS => return "01011";
         when BEQZS => return "01100";
         when BNEZS => return "01101";
         when SGES => return "01110";
         when SGEUS => return "01111";
         when SGTS => return "10000";
         when SGTUS => return "10001";
         when SLES => return "10010";
         when SLTS => return "10011";
         when SLTUS => return "10100";
         when SEQS => return "10101";
         when NEQS => return "10110";
         when LHIS => return "10111";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "00000";
      end case;
   end;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Fetch_DW01_add_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Fetch_DW01_add_1;

architecture SYN_cla of Fetch_DW01_add_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, SUM_2_port, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, 
      n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71 : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U2 : XOR2_X1 port map( A => n1, B => n18, Z => SUM_31_port);
   U3 : NAND2_X1 port map( A1 => n19, A2 => A(30), ZN => n1);
   U4 : NOR2_X1 port map( A1 => n69, A2 => n52, ZN => n13);
   U5 : AND2_X1 port map( A1 => n13, A2 => n11, ZN => n58);
   U6 : NOR2_X1 port map( A1 => n70, A2 => n12, ZN => n62);
   U7 : INV_X1 port map( A => n32, ZN => n36);
   U8 : INV_X1 port map( A => n25, ZN => n29);
   U9 : INV_X1 port map( A => n40, ZN => n44);
   U10 : OR2_X1 port map( A1 => n32, A2 => n33, ZN => n2);
   U11 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => n3);
   U12 : NAND3_X1 port map( A1 => n50, A2 => n51, A3 => n11, ZN => n4);
   U13 : OR2_X1 port map( A1 => n48, A2 => n49, ZN => n5);
   U14 : AND2_X1 port map( A1 => n57, A2 => A(13), ZN => n54);
   U15 : AND2_X1 port map( A1 => n15, A2 => A(5), ZN => n14);
   U16 : NOR2_X1 port map( A1 => n32, A2 => n33, ZN => n30);
   U17 : NOR2_X1 port map( A1 => n9, A2 => n21, ZN => n19);
   U18 : AND2_X1 port map( A1 => A(12), A2 => n58, ZN => n57);
   U19 : NOR2_X1 port map( A1 => n68, A2 => n69, ZN => n15);
   U20 : NOR2_X1 port map( A1 => n40, A2 => n41, ZN => n37);
   U21 : AND4_X1 port map( A1 => A(11), A2 => A(10), A3 => A(9), A4 => A(8), ZN
                           => n11);
   U22 : NOR2_X1 port map( A1 => n25, A2 => n26, ZN => n23);
   U23 : NOR2_X1 port map( A1 => SUM_2_port, A2 => n16, ZN => n51);
   U24 : AND2_X1 port map( A1 => n54, A2 => A(14), ZN => n53);
   U25 : AND2_X1 port map( A1 => n62, A2 => A(10), ZN => n61);
   U26 : AND2_X1 port map( A1 => n8, A2 => A(18), ZN => n42);
   U27 : NAND2_X1 port map( A1 => n13, A2 => A(8), ZN => n12);
   U28 : AND2_X1 port map( A1 => A(21), A2 => n36, ZN => n6);
   U29 : AND2_X1 port map( A1 => A(25), A2 => n29, ZN => n7);
   U30 : AND2_X1 port map( A1 => A(17), A2 => n44, ZN => n8);
   U31 : NAND2_X1 port map( A1 => A(22), A2 => n6, ZN => n34);
   U32 : NAND2_X1 port map( A1 => A(26), A2 => n7, ZN => n27);
   U33 : NAND2_X1 port map( A1 => A(12), A2 => A(13), ZN => n49);
   U34 : NAND2_X1 port map( A1 => A(14), A2 => A(15), ZN => n48);
   U35 : NAND2_X1 port map( A1 => n23, A2 => A(28), ZN => n9);
   U36 : AND2_X1 port map( A1 => A(6), A2 => n14, ZN => n10);
   U37 : INV_X1 port map( A => A(14), ZN => n56);
   U38 : INV_X1 port map( A => A(3), ZN => n16);
   U39 : INV_X1 port map( A => A(29), ZN => n21);
   U40 : XNOR2_X1 port map( A => n65, B => n10, ZN => SUM_7_port);
   U41 : XNOR2_X1 port map( A => n68, B => n51, ZN => SUM_4_port);
   U42 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U43 : INV_X1 port map( A => A(13), ZN => n59);
   U44 : INV_X1 port map( A => A(12), ZN => n60);
   U45 : INV_X1 port map( A => A(17), ZN => n46);
   U46 : INV_X1 port map( A => A(25), ZN => n31);
   U47 : INV_X1 port map( A => A(26), ZN => n28);
   U48 : INV_X1 port map( A => A(18), ZN => n45);
   U49 : INV_X1 port map( A => A(15), ZN => n55);
   U50 : XNOR2_X1 port map( A => n66, B => n14, ZN => SUM_6_port);
   U51 : XNOR2_X1 port map( A => n56, B => n54, ZN => SUM_14_port);
   U52 : XNOR2_X1 port map( A => n16, B => A(2), ZN => SUM_3_port);
   U53 : XNOR2_X1 port map( A => n60, B => n58, ZN => SUM_12_port);
   U54 : XNOR2_X1 port map( A => n6, B => n35, ZN => SUM_22_port);
   U55 : XNOR2_X1 port map( A => n34, B => A(23), ZN => SUM_23_port);
   U56 : XNOR2_X1 port map( A => n2, B => A(24), ZN => SUM_24_port);
   U57 : XNOR2_X1 port map( A => n31, B => n29, ZN => SUM_25_port);
   U58 : XNOR2_X1 port map( A => n7, B => n28, ZN => SUM_26_port);
   U59 : XNOR2_X1 port map( A => n24, B => A(28), ZN => SUM_28_port);
   U60 : XNOR2_X1 port map( A => n21, B => n22, ZN => SUM_29_port);
   U61 : XNOR2_X1 port map( A => n27, B => A(27), ZN => SUM_27_port);
   U62 : XNOR2_X1 port map( A => n38, B => n36, ZN => SUM_21_port);
   U63 : XNOR2_X1 port map( A => n45, B => n8, ZN => SUM_18_port);
   U64 : XNOR2_X1 port map( A => n46, B => n44, ZN => SUM_17_port);
   U65 : INV_X1 port map( A => A(19), ZN => n43);
   U66 : INV_X1 port map( A => A(11), ZN => n63);
   U67 : INV_X1 port map( A => A(21), ZN => n38);
   U68 : INV_X1 port map( A => A(22), ZN => n35);
   U69 : INV_X1 port map( A => A(31), ZN => n18);
   U70 : INV_X1 port map( A => A(6), ZN => n66);
   U71 : INV_X1 port map( A => A(4), ZN => n68);
   U72 : INV_X1 port map( A => n9, ZN => n22);
   U73 : INV_X1 port map( A => A(7), ZN => n65);
   U74 : INV_X1 port map( A => A(5), ZN => n67);
   U75 : INV_X1 port map( A => A(9), ZN => n70);
   U76 : INV_X1 port map( A => A(10), ZN => n71);
   U77 : NAND4_X1 port map( A1 => A(4), A2 => A(5), A3 => A(6), A4 => A(7), ZN 
                           => n52);
   U78 : NAND2_X1 port map( A1 => n37, A2 => A(20), ZN => n32);
   U79 : NAND2_X1 port map( A1 => n30, A2 => A(24), ZN => n25);
   U80 : NAND2_X1 port map( A1 => n3, A2 => A(16), ZN => n40);
   U81 : XNOR2_X1 port map( A => n20, B => A(30), ZN => SUM_30_port);
   U82 : INV_X1 port map( A => A(8), ZN => n64);
   U83 : XNOR2_X1 port map( A => n12, B => A(9), ZN => SUM_9_port);
   U84 : XNOR2_X1 port map( A => n64, B => n13, ZN => SUM_8_port);
   U85 : XNOR2_X1 port map( A => n67, B => n15, ZN => SUM_5_port);
   U86 : INV_X1 port map( A => n19, ZN => n20);
   U87 : INV_X1 port map( A => n23, ZN => n24);
   U88 : NAND3_X1 port map( A1 => A(26), A2 => A(27), A3 => A(25), ZN => n26);
   U89 : NAND3_X1 port map( A1 => A(22), A2 => A(23), A3 => A(21), ZN => n33);
   U90 : XNOR2_X1 port map( A => n39, B => A(20), ZN => SUM_20_port);
   U91 : INV_X1 port map( A => n37, ZN => n39);
   U92 : NAND3_X1 port map( A1 => A(18), A2 => A(19), A3 => A(17), ZN => n41);
   U93 : XNOR2_X1 port map( A => n43, B => n42, ZN => SUM_19_port);
   U94 : XNOR2_X1 port map( A => n47, B => A(16), ZN => SUM_16_port);
   U95 : INV_X1 port map( A => n3, ZN => n47);
   U96 : INV_X1 port map( A => n52, ZN => n50);
   U97 : XNOR2_X1 port map( A => n55, B => n53, ZN => SUM_15_port);
   U98 : XNOR2_X1 port map( A => n59, B => n57, ZN => SUM_13_port);
   U99 : XNOR2_X1 port map( A => n63, B => n61, ZN => SUM_11_port);
   U100 : XNOR2_X1 port map( A => n71, B => n62, ZN => SUM_10_port);
   U101 : INV_X1 port map( A => n51, ZN => n69);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute_DW01_add_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Execute_DW01_add_1;

architecture SYN_rpl of Execute_DW01_add_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_3_port, SUM_4_port, SUM_5_port, SUM_6_port, 
      SUM_7_port, SUM_8_port, SUM_9_port, SUM_10_port, SUM_11_port, SUM_12_port
      , SUM_13_port, SUM_14_port, SUM_15_port, SUM_16_port, SUM_17_port, 
      SUM_18_port, SUM_19_port, SUM_20_port, SUM_21_port, SUM_22_port, 
      SUM_23_port, SUM_24_port, SUM_25_port, SUM_26_port, SUM_27_port, 
      SUM_28_port, SUM_29_port, SUM_30_port, n30, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n54, n55, n56, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, B(1), B(0) );
   
   U1 : XNOR2_X1 port map( A => B(31), B => n57, ZN => SUM_31_port);
   U2 : NAND2_X1 port map( A1 => B(30), A2 => n56, ZN => n57);
   U3 : INV_X1 port map( A => B(2), ZN => SUM_2_port);
   U4 : XOR2_X1 port map( A => B(3), B => B(2), Z => SUM_3_port);
   U5 : XOR2_X1 port map( A => B(4), B => n30, Z => SUM_4_port);
   U6 : XOR2_X1 port map( A => B(5), B => n31, Z => SUM_5_port);
   U7 : XOR2_X1 port map( A => B(6), B => n32, Z => SUM_6_port);
   U8 : XOR2_X1 port map( A => B(7), B => n33, Z => SUM_7_port);
   U9 : XOR2_X1 port map( A => B(8), B => n34, Z => SUM_8_port);
   U10 : XOR2_X1 port map( A => B(9), B => n35, Z => SUM_9_port);
   U11 : XOR2_X1 port map( A => B(10), B => n36, Z => SUM_10_port);
   U12 : XOR2_X1 port map( A => B(11), B => n37, Z => SUM_11_port);
   U13 : XOR2_X1 port map( A => B(12), B => n38, Z => SUM_12_port);
   U14 : XOR2_X1 port map( A => B(13), B => n39, Z => SUM_13_port);
   U15 : XOR2_X1 port map( A => B(14), B => n40, Z => SUM_14_port);
   U16 : XOR2_X1 port map( A => B(15), B => n41, Z => SUM_15_port);
   U17 : XOR2_X1 port map( A => B(16), B => n42, Z => SUM_16_port);
   U18 : XOR2_X1 port map( A => B(17), B => n43, Z => SUM_17_port);
   U19 : XOR2_X1 port map( A => B(18), B => n44, Z => SUM_18_port);
   U20 : XOR2_X1 port map( A => B(19), B => n45, Z => SUM_19_port);
   U21 : XOR2_X1 port map( A => B(20), B => n46, Z => SUM_20_port);
   U22 : XOR2_X1 port map( A => B(21), B => n47, Z => SUM_21_port);
   U23 : XOR2_X1 port map( A => B(22), B => n48, Z => SUM_22_port);
   U24 : XOR2_X1 port map( A => B(23), B => n49, Z => SUM_23_port);
   U25 : XOR2_X1 port map( A => B(24), B => n50, Z => SUM_24_port);
   U26 : XOR2_X1 port map( A => B(25), B => n51, Z => SUM_25_port);
   U27 : XOR2_X1 port map( A => B(26), B => n52, Z => SUM_26_port);
   U28 : XOR2_X1 port map( A => B(27), B => n53, Z => SUM_27_port);
   U29 : XOR2_X1 port map( A => B(28), B => n54, Z => SUM_28_port);
   U30 : XOR2_X1 port map( A => B(29), B => n55, Z => SUM_29_port);
   U31 : XOR2_X1 port map( A => B(30), B => n56, Z => SUM_30_port);
   U32 : AND2_X1 port map( A1 => B(3), A2 => B(2), ZN => n30);
   U33 : AND2_X1 port map( A1 => B(4), A2 => n30, ZN => n31);
   U34 : AND2_X1 port map( A1 => B(5), A2 => n31, ZN => n32);
   U35 : AND2_X1 port map( A1 => B(6), A2 => n32, ZN => n33);
   U36 : AND2_X1 port map( A1 => B(7), A2 => n33, ZN => n34);
   U37 : AND2_X1 port map( A1 => B(8), A2 => n34, ZN => n35);
   U38 : AND2_X1 port map( A1 => B(9), A2 => n35, ZN => n36);
   U39 : AND2_X1 port map( A1 => B(10), A2 => n36, ZN => n37);
   U40 : AND2_X1 port map( A1 => B(11), A2 => n37, ZN => n38);
   U41 : AND2_X1 port map( A1 => B(12), A2 => n38, ZN => n39);
   U42 : AND2_X1 port map( A1 => B(13), A2 => n39, ZN => n40);
   U43 : AND2_X1 port map( A1 => B(14), A2 => n40, ZN => n41);
   U44 : AND2_X1 port map( A1 => B(15), A2 => n41, ZN => n42);
   U45 : AND2_X1 port map( A1 => B(16), A2 => n42, ZN => n43);
   U46 : AND2_X1 port map( A1 => B(17), A2 => n43, ZN => n44);
   U47 : AND2_X1 port map( A1 => B(18), A2 => n44, ZN => n45);
   U48 : AND2_X1 port map( A1 => B(19), A2 => n45, ZN => n46);
   U49 : AND2_X1 port map( A1 => B(20), A2 => n46, ZN => n47);
   U50 : AND2_X1 port map( A1 => B(21), A2 => n47, ZN => n48);
   U51 : AND2_X1 port map( A1 => B(22), A2 => n48, ZN => n49);
   U52 : AND2_X1 port map( A1 => B(23), A2 => n49, ZN => n50);
   U53 : AND2_X1 port map( A1 => B(24), A2 => n50, ZN => n51);
   U54 : AND2_X1 port map( A1 => B(25), A2 => n51, ZN => n52);
   U55 : AND2_X1 port map( A1 => B(26), A2 => n52, ZN => n53);
   U56 : AND2_X1 port map( A1 => B(27), A2 => n53, ZN => n54);
   U57 : AND2_X1 port map( A1 => B(28), A2 => n54, ZN => n55);
   U58 : AND2_X1 port map( A1 => B(29), A2 => n55, ZN => n56);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Execute_DW01_add_0;

architecture SYN_rpl of Execute_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n2, n_1070 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1070, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n2, CO => carry_2_port, S
                           => SUM(1));
   U1 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U2 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n2);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity comparator_NBIT32_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end comparator_NBIT32_DW01_cmp6_0;

architecture SYN_rpl of comparator_NBIT32_DW01_cmp6_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal GT_port, GE_port, NE_port, LE_port, n3, n5, n6, n7, n8, n9, n10, n11,
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55
      , n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, 
      n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84
      , n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, 
      n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202 : std_logic;

begin
   GT <= GT_port;
   LE <= LE_port;
   GE <= GE_port;
   NE <= NE_port;
   
   U1 : INV_X1 port map( A => NE_port, ZN => EQ);
   U2 : INV_X1 port map( A => n142, ZN => n55);
   U3 : INV_X1 port map( A => n130, ZN => n7);
   U4 : INV_X1 port map( A => n118, ZN => n15);
   U5 : INV_X1 port map( A => n106, ZN => n23);
   U6 : INV_X1 port map( A => n94, ZN => n31);
   U7 : INV_X1 port map( A => n82, ZN => n39);
   U8 : INV_X1 port map( A => n139, ZN => n58);
   U9 : INV_X1 port map( A => n127, ZN => n10);
   U10 : INV_X1 port map( A => n115, ZN => n18);
   U11 : INV_X1 port map( A => n103, ZN => n26);
   U12 : INV_X1 port map( A => n91, ZN => n34);
   U13 : INV_X1 port map( A => n79, ZN => n42);
   U14 : INV_X1 port map( A => GT_port, ZN => LE_port);
   U15 : INV_X1 port map( A => n132, ZN => n61);
   U16 : INV_X1 port map( A => n141, ZN => n56);
   U17 : INV_X1 port map( A => n144, ZN => n53);
   U18 : INV_X1 port map( A => n120, ZN => n13);
   U19 : INV_X1 port map( A => n108, ZN => n21);
   U20 : INV_X1 port map( A => n96, ZN => n29);
   U21 : INV_X1 port map( A => n84, ZN => n37);
   U22 : INV_X1 port map( A => n129, ZN => n8);
   U23 : INV_X1 port map( A => n117, ZN => n16);
   U24 : INV_X1 port map( A => n105, ZN => n24);
   U25 : INV_X1 port map( A => n93, ZN => n32);
   U26 : INV_X1 port map( A => n81, ZN => n40);
   U27 : INV_X1 port map( A => n154, ZN => n47);
   U28 : INV_X1 port map( A => n68, ZN => n5);
   U29 : INV_X1 port map( A => A(30), ZN => n49);
   U30 : INV_X1 port map( A => n72, ZN => n45);
   U31 : INV_X1 port map( A => n151, ZN => n50);
   U32 : INV_X1 port map( A => B(30), ZN => n64);
   U33 : INV_X1 port map( A => n202, ZN => n3);
   U34 : INV_X1 port map( A => B(1), ZN => n63);
   U35 : INV_X1 port map( A => A(0), ZN => n6);
   U36 : INV_X1 port map( A => A(3), ZN => n51);
   U37 : INV_X1 port map( A => A(5), ZN => n54);
   U38 : INV_X1 port map( A => A(7), ZN => n59);
   U39 : INV_X1 port map( A => A(9), ZN => n62);
   U40 : INV_X1 port map( A => A(11), ZN => n11);
   U41 : INV_X1 port map( A => A(13), ZN => n14);
   U42 : INV_X1 port map( A => A(15), ZN => n19);
   U43 : INV_X1 port map( A => B(31), ZN => n65);
   U44 : INV_X1 port map( A => A(17), ZN => n22);
   U45 : INV_X1 port map( A => A(19), ZN => n27);
   U46 : INV_X1 port map( A => A(21), ZN => n30);
   U47 : INV_X1 port map( A => A(23), ZN => n35);
   U48 : INV_X1 port map( A => A(25), ZN => n38);
   U49 : INV_X1 port map( A => A(27), ZN => n43);
   U50 : INV_X1 port map( A => A(29), ZN => n46);
   U51 : INV_X1 port map( A => A(4), ZN => n52);
   U52 : INV_X1 port map( A => A(8), ZN => n60);
   U53 : INV_X1 port map( A => A(12), ZN => n12);
   U54 : INV_X1 port map( A => A(2), ZN => n48);
   U55 : INV_X1 port map( A => A(6), ZN => n57);
   U56 : INV_X1 port map( A => A(10), ZN => n9);
   U57 : INV_X1 port map( A => A(14), ZN => n17);
   U58 : INV_X1 port map( A => A(16), ZN => n20);
   U59 : INV_X1 port map( A => A(20), ZN => n28);
   U60 : INV_X1 port map( A => A(24), ZN => n36);
   U61 : INV_X1 port map( A => A(28), ZN => n44);
   U62 : INV_X1 port map( A => A(18), ZN => n25);
   U63 : INV_X1 port map( A => A(22), ZN => n33);
   U64 : INV_X1 port map( A => A(26), ZN => n41);
   U65 : INV_X1 port map( A => GE_port, ZN => LT);
   U66 : NAND2_X1 port map( A1 => LE_port, A2 => GE_port, ZN => NE_port);
   U67 : AOI21_X1 port map( B1 => n66, B2 => n5, A => n67, ZN => GE_port);
   U68 : AOI22_X1 port map( A1 => B(30), A2 => n49, B1 => n69, B2 => n70, ZN =>
                           n68);
   U69 : AOI21_X1 port map( B1 => n71, B2 => n72, A => n73, ZN => n69);
   U70 : AOI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => n71);
   U71 : AOI21_X1 port map( B1 => n77, B2 => n78, A => n79, ZN => n74);
   U72 : AOI21_X1 port map( B1 => n80, B2 => n39, A => n40, ZN => n77);
   U73 : AOI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n80);
   U74 : AOI21_X1 port map( B1 => n86, B2 => n87, A => n88, ZN => n83);
   U75 : AOI21_X1 port map( B1 => n89, B2 => n90, A => n91, ZN => n86);
   U76 : AOI21_X1 port map( B1 => n92, B2 => n31, A => n32, ZN => n89);
   U77 : AOI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n92);
   U78 : AOI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => n95);
   U79 : AOI21_X1 port map( B1 => n101, B2 => n102, A => n103, ZN => n98);
   U80 : AOI21_X1 port map( B1 => n104, B2 => n23, A => n24, ZN => n101);
   U81 : AOI21_X1 port map( B1 => n107, B2 => n108, A => n109, ZN => n104);
   U82 : AOI21_X1 port map( B1 => n110, B2 => n111, A => n112, ZN => n107);
   U83 : AOI21_X1 port map( B1 => n113, B2 => n114, A => n115, ZN => n110);
   U84 : AOI21_X1 port map( B1 => n116, B2 => n15, A => n16, ZN => n113);
   U85 : AOI21_X1 port map( B1 => n119, B2 => n120, A => n121, ZN => n116);
   U86 : AOI21_X1 port map( B1 => n122, B2 => n123, A => n124, ZN => n119);
   U87 : AOI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n122);
   U88 : AOI21_X1 port map( B1 => n128, B2 => n7, A => n8, ZN => n125);
   U89 : AOI21_X1 port map( B1 => n131, B2 => n132, A => n133, ZN => n128);
   U90 : AOI21_X1 port map( B1 => n134, B2 => n135, A => n136, ZN => n131);
   U91 : AOI21_X1 port map( B1 => n137, B2 => n138, A => n139, ZN => n134);
   U92 : AOI21_X1 port map( B1 => n140, B2 => n55, A => n56, ZN => n137);
   U93 : AOI21_X1 port map( B1 => n143, B2 => n144, A => n145, ZN => n140);
   U94 : AOI21_X1 port map( B1 => n146, B2 => n147, A => n148, ZN => n143);
   U95 : AOI21_X1 port map( B1 => n149, B2 => n150, A => n151, ZN => n146);
   U96 : AOI21_X1 port map( B1 => n152, B2 => n153, A => n47, ZN => n149);
   U97 : AOI22_X1 port map( A1 => n155, A2 => n63, B1 => A(1), B2 => n156, ZN 
                           => n152);
   U98 : OR2_X1 port map( A1 => n156, A2 => A(1), ZN => n155);
   U99 : NAND2_X1 port map( A1 => B(0), A2 => n6, ZN => n156);
   U100 : OAI21_X1 port map( B1 => n67, B2 => n157, A => n66, ZN => GT_port);
   U101 : NAND2_X1 port map( A1 => A(31), A2 => n65, ZN => n66);
   U102 : AOI22_X1 port map( A1 => A(30), A2 => n64, B1 => n158, B2 => n70, ZN 
                           => n157);
   U103 : XOR2_X1 port map( A => A(30), B => n64, Z => n70);
   U104 : AOI21_X1 port map( B1 => n159, B2 => n160, A => n45, ZN => n158);
   U105 : NAND2_X1 port map( A1 => B(29), A2 => n46, ZN => n72);
   U106 : OAI211_X1 port map( C1 => n161, C2 => n162, A => n78, B => n75, ZN =>
                           n160);
   U107 : NOR2_X1 port map( A1 => n163, A2 => n76, ZN => n75);
   U108 : AND2_X1 port map( A1 => B(28), A2 => n44, ZN => n76);
   U109 : NAND2_X1 port map( A1 => B(27), A2 => n43, ZN => n78);
   U110 : NAND2_X1 port map( A1 => n42, A2 => n164, ZN => n162);
   U111 : NOR2_X1 port map( A1 => n43, A2 => B(27), ZN => n79);
   U112 : AOI211_X1 port map( C1 => n165, C2 => n166, A => n82, B => n37, ZN =>
                           n161);
   U113 : NAND2_X1 port map( A1 => B(25), A2 => n38, ZN => n84);
   U114 : NAND2_X1 port map( A1 => n164, A2 => n81, ZN => n82);
   U115 : NAND2_X1 port map( A1 => B(26), A2 => n41, ZN => n81);
   U116 : OR2_X1 port map( A1 => n41, A2 => B(26), ZN => n164);
   U117 : OAI211_X1 port map( C1 => n167, C2 => n168, A => n90, B => n87, ZN =>
                           n166);
   U118 : NOR2_X1 port map( A1 => n169, A2 => n88, ZN => n87);
   U119 : AND2_X1 port map( A1 => B(24), A2 => n36, ZN => n88);
   U120 : NAND2_X1 port map( A1 => B(23), A2 => n35, ZN => n90);
   U121 : NAND2_X1 port map( A1 => n34, A2 => n170, ZN => n168);
   U122 : NOR2_X1 port map( A1 => n35, A2 => B(23), ZN => n91);
   U123 : AOI211_X1 port map( C1 => n171, C2 => n172, A => n94, B => n29, ZN =>
                           n167);
   U124 : NAND2_X1 port map( A1 => B(21), A2 => n30, ZN => n96);
   U125 : NAND2_X1 port map( A1 => n170, A2 => n93, ZN => n94);
   U126 : NAND2_X1 port map( A1 => B(22), A2 => n33, ZN => n93);
   U127 : OR2_X1 port map( A1 => n33, A2 => B(22), ZN => n170);
   U128 : OAI211_X1 port map( C1 => n173, C2 => n174, A => n102, B => n99, ZN 
                           => n172);
   U129 : NOR2_X1 port map( A1 => n175, A2 => n100, ZN => n99);
   U130 : AND2_X1 port map( A1 => B(20), A2 => n28, ZN => n100);
   U131 : NAND2_X1 port map( A1 => B(19), A2 => n27, ZN => n102);
   U132 : NAND2_X1 port map( A1 => n26, A2 => n176, ZN => n174);
   U133 : NOR2_X1 port map( A1 => n27, A2 => B(19), ZN => n103);
   U134 : AOI211_X1 port map( C1 => n177, C2 => n178, A => n106, B => n21, ZN 
                           => n173);
   U135 : NAND2_X1 port map( A1 => B(17), A2 => n22, ZN => n108);
   U136 : NAND2_X1 port map( A1 => n176, A2 => n105, ZN => n106);
   U137 : NAND2_X1 port map( A1 => B(18), A2 => n25, ZN => n105);
   U138 : OR2_X1 port map( A1 => n25, A2 => B(18), ZN => n176);
   U139 : OAI211_X1 port map( C1 => n179, C2 => n180, A => n114, B => n111, ZN 
                           => n178);
   U140 : NOR2_X1 port map( A1 => n181, A2 => n112, ZN => n111);
   U141 : AND2_X1 port map( A1 => B(16), A2 => n20, ZN => n112);
   U142 : NAND2_X1 port map( A1 => B(15), A2 => n19, ZN => n114);
   U143 : NAND2_X1 port map( A1 => n18, A2 => n182, ZN => n180);
   U144 : NOR2_X1 port map( A1 => n19, A2 => B(15), ZN => n115);
   U145 : AOI211_X1 port map( C1 => n183, C2 => n184, A => n118, B => n13, ZN 
                           => n179);
   U146 : NAND2_X1 port map( A1 => B(13), A2 => n14, ZN => n120);
   U147 : NAND2_X1 port map( A1 => n182, A2 => n117, ZN => n118);
   U148 : NAND2_X1 port map( A1 => B(14), A2 => n17, ZN => n117);
   U149 : OR2_X1 port map( A1 => n17, A2 => B(14), ZN => n182);
   U150 : OAI211_X1 port map( C1 => n185, C2 => n186, A => n126, B => n123, ZN 
                           => n184);
   U151 : NOR2_X1 port map( A1 => n187, A2 => n124, ZN => n123);
   U152 : AND2_X1 port map( A1 => B(12), A2 => n12, ZN => n124);
   U153 : NAND2_X1 port map( A1 => B(11), A2 => n11, ZN => n126);
   U154 : NAND2_X1 port map( A1 => n10, A2 => n188, ZN => n186);
   U155 : NOR2_X1 port map( A1 => n11, A2 => B(11), ZN => n127);
   U156 : AOI211_X1 port map( C1 => n189, C2 => n190, A => n130, B => n61, ZN 
                           => n185);
   U157 : NAND2_X1 port map( A1 => B(9), A2 => n62, ZN => n132);
   U158 : NAND2_X1 port map( A1 => n188, A2 => n129, ZN => n130);
   U159 : NAND2_X1 port map( A1 => B(10), A2 => n9, ZN => n129);
   U160 : OR2_X1 port map( A1 => n9, A2 => B(10), ZN => n188);
   U161 : OAI211_X1 port map( C1 => n191, C2 => n192, A => n138, B => n135, ZN 
                           => n190);
   U162 : NOR2_X1 port map( A1 => n193, A2 => n136, ZN => n135);
   U163 : AND2_X1 port map( A1 => B(8), A2 => n60, ZN => n136);
   U164 : NAND2_X1 port map( A1 => B(7), A2 => n59, ZN => n138);
   U165 : NAND2_X1 port map( A1 => n58, A2 => n194, ZN => n192);
   U166 : NOR2_X1 port map( A1 => n59, A2 => B(7), ZN => n139);
   U167 : AOI211_X1 port map( C1 => n195, C2 => n196, A => n142, B => n53, ZN 
                           => n191);
   U168 : NAND2_X1 port map( A1 => B(5), A2 => n54, ZN => n144);
   U169 : NAND2_X1 port map( A1 => n194, A2 => n141, ZN => n142);
   U170 : NAND2_X1 port map( A1 => B(6), A2 => n57, ZN => n141);
   U171 : OR2_X1 port map( A1 => n57, A2 => B(6), ZN => n194);
   U172 : NAND3_X1 port map( A1 => n197, A2 => n150, A3 => n147, ZN => n196);
   U173 : NOR2_X1 port map( A1 => n198, A2 => n148, ZN => n147);
   U174 : AND2_X1 port map( A1 => B(4), A2 => n52, ZN => n148);
   U175 : NAND2_X1 port map( A1 => B(3), A2 => n51, ZN => n150);
   U176 : NAND3_X1 port map( A1 => n50, A2 => n199, A3 => n200, ZN => n197);
   U177 : OAI211_X1 port map( C1 => A(1), C2 => n201, A => n3, B => n153, ZN =>
                           n200);
   U178 : AND2_X1 port map( A1 => n199, A2 => n154, ZN => n153);
   U179 : NAND2_X1 port map( A1 => B(2), A2 => n48, ZN => n154);
   U180 : AOI21_X1 port map( B1 => A(1), B2 => n201, A => n63, ZN => n202);
   U181 : NOR2_X1 port map( A1 => n6, A2 => B(0), ZN => n201);
   U182 : OR2_X1 port map( A1 => n48, A2 => B(2), ZN => n199);
   U183 : NOR2_X1 port map( A1 => n51, A2 => B(3), ZN => n151);
   U184 : NOR2_X1 port map( A1 => n198, A2 => n145, ZN => n195);
   U185 : NOR2_X1 port map( A1 => n54, A2 => B(5), ZN => n145);
   U186 : NOR2_X1 port map( A1 => n52, A2 => B(4), ZN => n198);
   U187 : NOR2_X1 port map( A1 => n193, A2 => n133, ZN => n189);
   U188 : NOR2_X1 port map( A1 => n62, A2 => B(9), ZN => n133);
   U189 : NOR2_X1 port map( A1 => n60, A2 => B(8), ZN => n193);
   U190 : NOR2_X1 port map( A1 => n187, A2 => n121, ZN => n183);
   U191 : NOR2_X1 port map( A1 => n14, A2 => B(13), ZN => n121);
   U192 : NOR2_X1 port map( A1 => n12, A2 => B(12), ZN => n187);
   U193 : NOR2_X1 port map( A1 => n181, A2 => n109, ZN => n177);
   U194 : NOR2_X1 port map( A1 => n22, A2 => B(17), ZN => n109);
   U195 : NOR2_X1 port map( A1 => n20, A2 => B(16), ZN => n181);
   U196 : NOR2_X1 port map( A1 => n175, A2 => n97, ZN => n171);
   U197 : NOR2_X1 port map( A1 => n30, A2 => B(21), ZN => n97);
   U198 : NOR2_X1 port map( A1 => n28, A2 => B(20), ZN => n175);
   U199 : NOR2_X1 port map( A1 => n169, A2 => n85, ZN => n165);
   U200 : NOR2_X1 port map( A1 => n38, A2 => B(25), ZN => n85);
   U201 : NOR2_X1 port map( A1 => n36, A2 => B(24), ZN => n169);
   U202 : NOR2_X1 port map( A1 => n163, A2 => n73, ZN => n159);
   U203 : NOR2_X1 port map( A1 => n46, A2 => B(29), ZN => n73);
   U204 : NOR2_X1 port map( A1 => n44, A2 => B(28), ZN => n163);
   U205 : NOR2_X1 port map( A1 => n65, A2 => A(31), ZN => n67);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_0_DW01_add_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end rca_bhv_numBit32_0_DW01_add_0;

architecture SYN_rpl of rca_bhv_numBit32_0_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1075 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1075, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_6_DW01_add_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end rca_bhv_numBit32_6_DW01_add_0;

architecture SYN_rpl of rca_bhv_numBit32_6_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1079 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1079, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_5_DW01_add_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end rca_bhv_numBit32_5_DW01_add_0;

architecture SYN_rpl of rca_bhv_numBit32_5_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1083 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1083, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_4_DW01_add_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end rca_bhv_numBit32_4_DW01_add_0;

architecture SYN_rpl of rca_bhv_numBit32_4_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1087 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1087, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_3_DW01_add_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end rca_bhv_numBit32_3_DW01_add_0;

architecture SYN_rpl of rca_bhv_numBit32_3_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1091 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1091, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_2_DW01_add_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end rca_bhv_numBit32_2_DW01_add_0;

architecture SYN_rpl of rca_bhv_numBit32_2_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1095 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1095, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_1_DW01_add_0 is

   port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (32 downto 0);  CO : out std_logic);

end rca_bhv_numBit32_1_DW01_add_0;

architecture SYN_rpl of rca_bhv_numBit32_1_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1099 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1099, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HazardDetection_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end HazardDetection_DW01_add_0;

architecture SYN_rpl of HazardDetection_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_30_port, SUM_16_port, SUM_17_port, SUM_18_port, 
      SUM_19_port, SUM_20_port, SUM_21_port, SUM_22_port, SUM_23_port, 
      SUM_24_port, SUM_25_port, SUM_26_port, SUM_27_port, SUM_28_port, 
      SUM_29_port, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , SUM_3_port, SUM_9_port, SUM_11_port, SUM_12_port, SUM_13_port, 
      SUM_14_port, SUM_15_port, SUM_4_port, SUM_5_port, SUM_6_port, SUM_7_port,
      SUM_8_port, SUM_10_port, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U1 : XNOR2_X1 port map( A => A(31), B => n57, ZN => SUM_31_port);
   U2 : XOR2_X1 port map( A => A(30), B => n35, Z => SUM_30_port);
   U3 : XOR2_X1 port map( A => A(16), B => n21, Z => SUM_16_port);
   U4 : XOR2_X1 port map( A => A(17), B => n22, Z => SUM_17_port);
   U5 : XOR2_X1 port map( A => A(18), B => n23, Z => SUM_18_port);
   U6 : XOR2_X1 port map( A => A(19), B => n24, Z => SUM_19_port);
   U7 : XOR2_X1 port map( A => A(20), B => n25, Z => SUM_20_port);
   U8 : XOR2_X1 port map( A => A(21), B => n26, Z => SUM_21_port);
   U9 : XOR2_X1 port map( A => A(22), B => n27, Z => SUM_22_port);
   U10 : XOR2_X1 port map( A => A(23), B => n28, Z => SUM_23_port);
   U11 : XOR2_X1 port map( A => A(24), B => n29, Z => SUM_24_port);
   U12 : XOR2_X1 port map( A => A(25), B => n30, Z => SUM_25_port);
   U13 : XOR2_X1 port map( A => A(26), B => n31, Z => SUM_26_port);
   U14 : XOR2_X1 port map( A => A(27), B => n32, Z => SUM_27_port);
   U15 : XOR2_X1 port map( A => A(28), B => n33, Z => SUM_28_port);
   U16 : XOR2_X1 port map( A => A(29), B => n34, Z => SUM_29_port);
   U17 : NAND2_X1 port map( A1 => A(30), A2 => n35, ZN => n57);
   U18 : AND2_X1 port map( A1 => A(11), A2 => n43, ZN => n17);
   U19 : AND2_X1 port map( A1 => A(12), A2 => n17, ZN => n18);
   U20 : AND2_X1 port map( A1 => A(13), A2 => n18, ZN => n19);
   U21 : AND2_X1 port map( A1 => A(14), A2 => n19, ZN => n20);
   U22 : AND2_X1 port map( A1 => A(15), A2 => n20, ZN => n21);
   U23 : AND2_X1 port map( A1 => A(16), A2 => n21, ZN => n22);
   U24 : AND2_X1 port map( A1 => A(17), A2 => n22, ZN => n23);
   U25 : AND2_X1 port map( A1 => A(18), A2 => n23, ZN => n24);
   U26 : AND2_X1 port map( A1 => A(19), A2 => n24, ZN => n25);
   U27 : AND2_X1 port map( A1 => A(20), A2 => n25, ZN => n26);
   U28 : AND2_X1 port map( A1 => A(21), A2 => n26, ZN => n27);
   U29 : AND2_X1 port map( A1 => A(22), A2 => n27, ZN => n28);
   U30 : AND2_X1 port map( A1 => A(23), A2 => n28, ZN => n29);
   U31 : AND2_X1 port map( A1 => A(24), A2 => n29, ZN => n30);
   U32 : AND2_X1 port map( A1 => A(25), A2 => n30, ZN => n31);
   U33 : AND2_X1 port map( A1 => A(26), A2 => n31, ZN => n32);
   U34 : AND2_X1 port map( A1 => A(27), A2 => n32, ZN => n33);
   U35 : AND2_X1 port map( A1 => A(28), A2 => n33, ZN => n34);
   U36 : AND2_X1 port map( A1 => A(29), A2 => n34, ZN => n35);
   U37 : AND2_X1 port map( A1 => A(9), A2 => n42, ZN => n36);
   U38 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n37);
   U39 : AND2_X1 port map( A1 => A(4), A2 => n37, ZN => n38);
   U40 : AND2_X1 port map( A1 => A(5), A2 => n38, ZN => n39);
   U41 : AND2_X1 port map( A1 => A(6), A2 => n39, ZN => n40);
   U42 : AND2_X1 port map( A1 => A(7), A2 => n40, ZN => n41);
   U43 : AND2_X1 port map( A1 => A(8), A2 => n41, ZN => n42);
   U44 : AND2_X1 port map( A1 => A(10), A2 => n36, ZN => n43);
   U45 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U46 : XOR2_X1 port map( A => A(3), B => A(2), Z => SUM_3_port);
   U47 : XOR2_X1 port map( A => A(9), B => n42, Z => SUM_9_port);
   U48 : XOR2_X1 port map( A => A(11), B => n43, Z => SUM_11_port);
   U49 : XOR2_X1 port map( A => A(12), B => n17, Z => SUM_12_port);
   U50 : XOR2_X1 port map( A => A(13), B => n18, Z => SUM_13_port);
   U51 : XOR2_X1 port map( A => A(14), B => n19, Z => SUM_14_port);
   U52 : XOR2_X1 port map( A => A(15), B => n20, Z => SUM_15_port);
   U53 : XOR2_X1 port map( A => A(4), B => n37, Z => SUM_4_port);
   U54 : XOR2_X1 port map( A => A(5), B => n38, Z => SUM_5_port);
   U55 : XOR2_X1 port map( A => A(6), B => n39, Z => SUM_6_port);
   U56 : XOR2_X1 port map( A => A(7), B => n40, Z => SUM_7_port);
   U57 : XOR2_X1 port map( A => A(8), B => n41, Z => SUM_8_port);
   U58 : XOR2_X1 port map( A => A(10), B => n36, Z => SUM_10_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_15;

architecture SYN_STRUCTURAL of RCA_N4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_14;

architecture SYN_STRUCTURAL of RCA_N4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_13;

architecture SYN_STRUCTURAL of RCA_N4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_12;

architecture SYN_STRUCTURAL of RCA_N4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_11;

architecture SYN_STRUCTURAL of RCA_N4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_10;

architecture SYN_STRUCTURAL of RCA_N4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_9;

architecture SYN_STRUCTURAL of RCA_N4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_8;

architecture SYN_STRUCTURAL of RCA_N4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_7;

architecture SYN_STRUCTURAL of RCA_N4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_6;

architecture SYN_STRUCTURAL of RCA_N4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_5;

architecture SYN_STRUCTURAL of RCA_N4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_4;

architecture SYN_STRUCTURAL of RCA_N4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_3;

architecture SYN_STRUCTURAL of RCA_N4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_2;

architecture SYN_STRUCTURAL of RCA_N4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_1;

architecture SYN_STRUCTURAL of RCA_N4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_7;

architecture SYN_struct of carry_select_basic_N4_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1134, n_1135 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1134);
   RCA1 : RCA_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1135);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n11, ZN => S(1));
   U5 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n13, ZN => S(3));
   U9 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_6;

architecture SYN_struct of carry_select_basic_N4_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1136, n_1137 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1136);
   RCA1 : RCA_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1137);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n11, ZN => S(1));
   U5 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n13, ZN => S(3));
   U9 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_5;

architecture SYN_struct of carry_select_basic_N4_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1138, n_1139 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1138);
   RCA1 : RCA_N4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1139);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n11, ZN => S(1));
   U5 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n13, ZN => S(3));
   U9 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_4;

architecture SYN_struct of carry_select_basic_N4_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1140, n_1141 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1140);
   RCA1 : RCA_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1141);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n11, ZN => S(1));
   U5 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n13, ZN => S(3));
   U9 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_3;

architecture SYN_struct of carry_select_basic_N4_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1142, n_1143 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1142);
   RCA1 : RCA_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1143);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n11, ZN => S(1));
   U5 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n13, ZN => S(3));
   U9 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_2;

architecture SYN_struct of carry_select_basic_N4_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1144, n_1145 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1144);
   RCA1 : RCA_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1145);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n11, ZN => S(1));
   U5 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U6 : INV_X1 port map( A => n12, ZN => S(2));
   U7 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U8 : INV_X1 port map( A => n13, ZN => S(3));
   U9 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_1;

architecture SYN_struct of carry_select_basic_N4_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n5, n10, n11, n12,
      n13, n_1146, n_1147 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1146);
   RCA1 : RCA_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1147);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n13, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n13);
   U6 : INV_X1 port map( A => n11, ZN => S(1));
   U7 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n11);
   U8 : INV_X1 port map( A => n12, ZN => S(2));
   U9 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n12);
   U10 : INV_X1 port map( A => n10, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_26 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_26;

architecture SYN_bhv of PGblock_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_25 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_25;

architecture SYN_bhv of PGblock_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_24 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_24;

architecture SYN_bhv of PGblock_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_23 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_23;

architecture SYN_bhv of PGblock_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_22 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_22;

architecture SYN_bhv of PGblock_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_21 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_21;

architecture SYN_bhv of PGblock_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_20 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_20;

architecture SYN_bhv of PGblock_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_19 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_19;

architecture SYN_bhv of PGblock_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_18 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_18;

architecture SYN_bhv of PGblock_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_17 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_17;

architecture SYN_bhv of PGblock_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_16 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_16;

architecture SYN_bhv of PGblock_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_15 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_15;

architecture SYN_bhv of PGblock_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_14 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_14;

architecture SYN_bhv of PGblock_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_13 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_13;

architecture SYN_bhv of PGblock_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_12 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_12;

architecture SYN_bhv of PGblock_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_11 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_11;

architecture SYN_bhv of PGblock_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_10 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_10;

architecture SYN_bhv of PGblock_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_9 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_9;

architecture SYN_bhv of PGblock_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_8 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_8;

architecture SYN_bhv of PGblock_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_7 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_7;

architecture SYN_bhv of PGblock_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_6 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_6;

architecture SYN_bhv of PGblock_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_5 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_5;

architecture SYN_bhv of PGblock_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_4 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_4;

architecture SYN_bhv of PGblock_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_3 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_3;

architecture SYN_bhv of PGblock_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U2 : INV_X1 port map( A => n3, ZN => Gij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_2 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_2;

architecture SYN_bhv of PGblock_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_1 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_1;

architecture SYN_bhv of PGblock_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);
   U3 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_8 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_8;

architecture SYN_bhv of Gblock_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_7 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_7;

architecture SYN_bhv of Gblock_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_6 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_6;

architecture SYN_bhv of Gblock_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_5 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_5;

architecture SYN_bhv of Gblock_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_4 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_4;

architecture SYN_bhv of Gblock_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_3 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_3;

architecture SYN_bhv of Gblock_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_2 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_2;

architecture SYN_bhv of Gblock_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_1 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_1;

architecture SYN_bhv of Gblock_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_30 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_30;

architecture SYN_bhv of PG_net_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_29 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_29;

architecture SYN_bhv of PG_net_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_28 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_28;

architecture SYN_bhv of PG_net_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_27 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_27;

architecture SYN_bhv of PG_net_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_26 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_26;

architecture SYN_bhv of PG_net_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_25 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_25;

architecture SYN_bhv of PG_net_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_24 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_24;

architecture SYN_bhv of PG_net_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_23 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_23;

architecture SYN_bhv of PG_net_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_22 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_22;

architecture SYN_bhv of PG_net_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_21 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_21;

architecture SYN_bhv of PG_net_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_20 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_20;

architecture SYN_bhv of PG_net_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_19 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_19;

architecture SYN_bhv of PG_net_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_18 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_18;

architecture SYN_bhv of PG_net_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_17 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_17;

architecture SYN_bhv of PG_net_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_16 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_16;

architecture SYN_bhv of PG_net_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_15 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_15;

architecture SYN_bhv of PG_net_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_14 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_14;

architecture SYN_bhv of PG_net_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_13 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_13;

architecture SYN_bhv of PG_net_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_12 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_12;

architecture SYN_bhv of PG_net_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_11 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_11;

architecture SYN_bhv of PG_net_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_10 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_10;

architecture SYN_bhv of PG_net_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_9 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_9;

architecture SYN_bhv of PG_net_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_8 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_8;

architecture SYN_bhv of PG_net_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_7 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_7;

architecture SYN_bhv of PG_net_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_6 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_6;

architecture SYN_bhv of PG_net_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_5 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_5;

architecture SYN_bhv of PG_net_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_4 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_4;

architecture SYN_bhv of PG_net_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_3 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_3;

architecture SYN_bhv of PG_net_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_2 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_2;

architecture SYN_bhv of PG_net_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_1 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_1;

architecture SYN_bhv of PG_net_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_6 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end rca_bhv_numBit32_6;

architecture SYN_BEHAVIORAL of rca_bhv_numBit32_6 is

   component rca_bhv_numBit32_6_DW01_add_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   signal n_1148 : std_logic;

begin
   
   add_1_root_add_35_2 : rca_bhv_numBit32_6_DW01_add_0 port map( A(32) => A(31)
                           , A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(32) => Co, SUM(31)
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1148);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end rca_bhv_numBit32_5;

architecture SYN_BEHAVIORAL of rca_bhv_numBit32_5 is

   component rca_bhv_numBit32_5_DW01_add_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   signal n_1149 : std_logic;

begin
   
   add_1_root_add_35_2 : rca_bhv_numBit32_5_DW01_add_0 port map( A(32) => A(31)
                           , A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(32) => Co, SUM(31)
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1149);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end rca_bhv_numBit32_4;

architecture SYN_BEHAVIORAL of rca_bhv_numBit32_4 is

   component rca_bhv_numBit32_4_DW01_add_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   signal n_1150 : std_logic;

begin
   
   add_1_root_add_35_2 : rca_bhv_numBit32_4_DW01_add_0 port map( A(32) => A(31)
                           , A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(32) => Co, SUM(31)
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1150);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end rca_bhv_numBit32_3;

architecture SYN_BEHAVIORAL of rca_bhv_numBit32_3 is

   component rca_bhv_numBit32_3_DW01_add_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   signal n_1151 : std_logic;

begin
   
   add_1_root_add_35_2 : rca_bhv_numBit32_3_DW01_add_0 port map( A(32) => A(31)
                           , A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(32) => Co, SUM(31)
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1151);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end rca_bhv_numBit32_2;

architecture SYN_BEHAVIORAL of rca_bhv_numBit32_2 is

   component rca_bhv_numBit32_2_DW01_add_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   signal n_1152 : std_logic;

begin
   
   add_1_root_add_35_2 : rca_bhv_numBit32_2_DW01_add_0 port map( A(32) => A(31)
                           , A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(32) => Co, SUM(31)
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1152);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end rca_bhv_numBit32_1;

architecture SYN_BEHAVIORAL of rca_bhv_numBit32_1 is

   component rca_bhv_numBit32_1_DW01_add_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   signal n_1153 : std_logic;

begin
   
   add_1_root_add_35_2 : rca_bhv_numBit32_1_DW01_add_0 port map( A(32) => A(31)
                           , A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(32) => Co, SUM(31)
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1153);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_7 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_7;

architecture SYN_bhv of mux5to1_numBit32_7 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n91, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n160);
   U2 : BUF_X1 port map( A => n158, Z => n4);
   U3 : BUF_X1 port map( A => n158, Z => n77);
   U4 : BUF_X1 port map( A => n158, Z => n78);
   U5 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84,
                           C1 => IN5(25), C2 => n81, ZN => n146);
   U6 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84,
                           C1 => IN5(26), C2 => n81, ZN => n148);
   U7 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84,
                           C1 => IN5(27), C2 => n81, ZN => n150);
   U8 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => n84,
                           C1 => IN5(28), C2 => n81, ZN => n152);
   U9 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => n84,
                           C1 => IN5(29), C2 => n81, ZN => n154);
   U10 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => n84
                           , C1 => IN5(30), C2 => n81, ZN => n156);
   U11 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n132);
   U12 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n134);
   U13 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n136);
   U14 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n138);
   U15 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n140);
   U16 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n142);
   U17 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n144);
   U18 : BUF_X1 port map( A => n89, Z => n1);
   U19 : BUF_X1 port map( A => n89, Z => n2);
   U20 : NOR2_X1 port map( A1 => n88, A2 => n93, ZN => n158);
   U21 : INV_X1 port map( A => n94, ZN => n88);
   U22 : BUF_X1 port map( A => n89, Z => n3);
   U23 : NOR4_X1 port map( A1 => n92, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n94);
   U24 : BUF_X1 port map( A => n160, Z => n82);
   U25 : BUF_X1 port map( A => n160, Z => n83);
   U26 : BUF_X1 port map( A => n159, Z => n79);
   U27 : BUF_X1 port map( A => n159, Z => n80);
   U28 : BUF_X1 port map( A => n161, Z => n85);
   U29 : BUF_X1 port map( A => n161, Z => n86);
   U30 : BUF_X1 port map( A => n160, Z => n84);
   U31 : NOR2_X1 port map( A1 => n91, A2 => n90, ZN => n93);
   U32 : BUF_X1 port map( A => n159, Z => n81);
   U33 : BUF_X1 port map( A => n161, Z => n87);
   U34 : INV_X1 port map( A => n95, ZN => n89);
   U35 : AOI21_X1 port map( B1 => n94, B2 => n93, A => n92, ZN => n95);
   U36 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82, 
                           C1 => IN5(4), C2 => n79, ZN => n104);
   U37 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82, 
                           C1 => IN5(5), C2 => n79, ZN => n106);
   U38 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82, 
                           C1 => IN5(6), C2 => n79, ZN => n108);
   U39 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82, 
                           C1 => IN5(7), C2 => n79, ZN => n110);
   U40 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82, 
                           C1 => IN5(8), C2 => n79, ZN => n112);
   U41 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82, 
                           C1 => IN5(9), C2 => n79, ZN => n114);
   U42 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => n82
                           , C1 => IN5(10), C2 => n79, ZN => n116);
   U43 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => n82
                           , C1 => IN5(11), C2 => n79, ZN => n118);
   U44 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => n83
                           , C1 => IN5(12), C2 => n80, ZN => n120);
   U45 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => n83
                           , C1 => IN5(13), C2 => n80, ZN => n122);
   U46 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n124);
   U47 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n126);
   U48 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n128);
   U49 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n130);
   U50 : NOR3_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => n90, ZN => n161);
   U51 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n92);
   U52 : INV_X1 port map( A => SEL_in(0), ZN => n90);
   U53 : AND3_X1 port map( A1 => n90, A2 => n91, A3 => SEL_in(2), ZN => n159);
   U54 : INV_X1 port map( A => SEL_in(1), ZN => n91);
   U55 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(3));
   U56 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82, 
                           C1 => IN5(3), C2 => n79, ZN => n102);
   U57 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN 
                           => n103);
   U58 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2, 
                           ZN => n129);
   U59 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82, 
                           C1 => IN5(2), C2 => n79, ZN => n100);
   U60 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2, 
                           ZN => n131);
   U61 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2, 
                           ZN => n133);
   U62 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(4));
   U63 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN 
                           => n105);
   U64 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(5));
   U65 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN 
                           => n107);
   U66 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(6));
   U67 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN 
                           => n109);
   U68 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(7));
   U69 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN 
                           => n111);
   U70 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(8));
   U71 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN 
                           => n113);
   U72 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(9));
   U73 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN 
                           => n115);
   U74 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(10));
   U75 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n117);
   U76 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(11));
   U77 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n119);
   U78 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(12));
   U79 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2, 
                           ZN => n121);
   U80 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(13));
   U81 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2, 
                           ZN => n123);
   U82 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(14));
   U83 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n125);
   U84 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(15));
   U85 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n127);
   U86 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(16));
   U87 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(17));
   U88 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(18));
   U89 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(19));
   U90 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n135);
   U91 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(20));
   U92 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n137);
   U93 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(21));
   U94 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n139);
   U95 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(22));
   U96 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n141);
   U97 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(23));
   U98 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n143);
   U99 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Z(24));
   U100 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3,
                           ZN => n145);
   U101 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Z(25));
   U102 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3,
                           ZN => n147);
   U103 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(26));
   U104 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3,
                           ZN => n149);
   U105 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Z(27));
   U106 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3,
                           ZN => n151);
   U107 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Z(28));
   U108 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3,
                           ZN => n153);
   U110 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Z(29));
   U111 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3,
                           ZN => n155);
   U112 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => Z(30));
   U113 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3,
                           ZN => n157);
   U114 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(2));
   U115 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN
                           => n101);
   U116 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(0));
   U117 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN
                           => n97);
   U118 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(1));
   U119 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN
                           => n99);
   U120 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => Z(31));
   U121 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n163);
   U122 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => 
                           n84, C1 => IN5(31), C2 => n81, ZN => n162);
   U123 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82,
                           C1 => IN5(0), C2 => n79, ZN => n96);
   U124 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82,
                           C1 => IN5(1), C2 => n79, ZN => n98);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_6 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_6;

architecture SYN_bhv of mux5to1_numBit32_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n91, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n160);
   U2 : BUF_X1 port map( A => n158, Z => n4);
   U3 : BUF_X1 port map( A => n158, Z => n77);
   U4 : BUF_X1 port map( A => n158, Z => n78);
   U5 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => n84,
                           C1 => IN5(31), C2 => n81, ZN => n162);
   U6 : BUF_X1 port map( A => n89, Z => n1);
   U7 : BUF_X1 port map( A => n89, Z => n2);
   U8 : NOR2_X1 port map( A1 => n88, A2 => n93, ZN => n158);
   U9 : INV_X1 port map( A => n94, ZN => n88);
   U10 : BUF_X1 port map( A => n89, Z => n3);
   U11 : NOR4_X1 port map( A1 => n92, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n94);
   U12 : BUF_X1 port map( A => n160, Z => n82);
   U13 : BUF_X1 port map( A => n160, Z => n83);
   U14 : BUF_X1 port map( A => n159, Z => n79);
   U15 : BUF_X1 port map( A => n159, Z => n80);
   U16 : BUF_X1 port map( A => n161, Z => n85);
   U17 : BUF_X1 port map( A => n161, Z => n86);
   U18 : BUF_X1 port map( A => n160, Z => n84);
   U19 : NOR2_X1 port map( A1 => n91, A2 => n90, ZN => n93);
   U20 : BUF_X1 port map( A => n159, Z => n81);
   U21 : BUF_X1 port map( A => n161, Z => n87);
   U22 : INV_X1 port map( A => n95, ZN => n89);
   U23 : AOI21_X1 port map( B1 => n94, B2 => n93, A => n92, ZN => n95);
   U24 : NOR3_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => n90, ZN => n161);
   U25 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n92);
   U26 : INV_X1 port map( A => SEL_in(0), ZN => n90);
   U27 : AND3_X1 port map( A1 => n90, A2 => n91, A3 => SEL_in(2), ZN => n159);
   U28 : INV_X1 port map( A => SEL_in(1), ZN => n91);
   U29 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(5));
   U30 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82, 
                           C1 => IN5(5), C2 => n79, ZN => n106);
   U31 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN 
                           => n107);
   U32 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(6));
   U33 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN 
                           => n109);
   U34 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82, 
                           C1 => IN5(6), C2 => n79, ZN => n108);
   U35 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(7));
   U36 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN 
                           => n111);
   U37 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82, 
                           C1 => IN5(7), C2 => n79, ZN => n110);
   U38 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(8));
   U39 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN 
                           => n113);
   U40 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82, 
                           C1 => IN5(8), C2 => n79, ZN => n112);
   U41 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(9));
   U42 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN 
                           => n115);
   U43 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82, 
                           C1 => IN5(9), C2 => n79, ZN => n114);
   U44 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(10));
   U45 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n117);
   U46 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => n82
                           , C1 => IN5(10), C2 => n79, ZN => n116);
   U47 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(11));
   U48 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n119);
   U49 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => n82
                           , C1 => IN5(11), C2 => n79, ZN => n118);
   U50 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(12));
   U51 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2, 
                           ZN => n121);
   U52 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => n83
                           , C1 => IN5(12), C2 => n80, ZN => n120);
   U53 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(13));
   U54 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2, 
                           ZN => n123);
   U55 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => n83
                           , C1 => IN5(13), C2 => n80, ZN => n122);
   U56 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(14));
   U57 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n125);
   U58 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n124);
   U59 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(15));
   U60 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n127);
   U61 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n126);
   U62 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(16));
   U63 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2, 
                           ZN => n129);
   U64 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n128);
   U65 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(17));
   U66 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2, 
                           ZN => n131);
   U67 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n130);
   U68 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(18));
   U69 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2, 
                           ZN => n133);
   U70 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n132);
   U71 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(19));
   U72 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n135);
   U73 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n134);
   U74 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(20));
   U75 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n137);
   U76 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n136);
   U77 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(21));
   U78 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n139);
   U79 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n138);
   U80 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(22));
   U81 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n141);
   U82 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n140);
   U83 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(23));
   U84 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n143);
   U85 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n142);
   U86 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Z(24));
   U87 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3, 
                           ZN => n145);
   U88 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n144);
   U89 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Z(25));
   U90 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3, 
                           ZN => n147);
   U91 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84
                           , C1 => IN5(25), C2 => n81, ZN => n146);
   U92 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(26));
   U93 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3, 
                           ZN => n149);
   U94 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84
                           , C1 => IN5(26), C2 => n81, ZN => n148);
   U95 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Z(27));
   U96 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3, 
                           ZN => n151);
   U97 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84
                           , C1 => IN5(27), C2 => n81, ZN => n150);
   U98 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Z(28));
   U99 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3, 
                           ZN => n153);
   U100 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => 
                           n84, C1 => IN5(28), C2 => n81, ZN => n152);
   U101 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Z(29));
   U102 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3,
                           ZN => n155);
   U103 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => 
                           n84, C1 => IN5(29), C2 => n81, ZN => n154);
   U104 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => Z(30));
   U105 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3,
                           ZN => n157);
   U106 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => 
                           n84, C1 => IN5(30), C2 => n81, ZN => n156);
   U107 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(4));
   U108 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN
                           => n105);
   U110 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82,
                           C1 => IN5(4), C2 => n79, ZN => n104);
   U111 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(0));
   U112 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN
                           => n97);
   U113 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82,
                           C1 => IN5(0), C2 => n79, ZN => n96);
   U114 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(1));
   U115 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN
                           => n99);
   U116 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82,
                           C1 => IN5(1), C2 => n79, ZN => n98);
   U117 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(2));
   U118 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN
                           => n101);
   U119 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82,
                           C1 => IN5(2), C2 => n79, ZN => n100);
   U120 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(3));
   U121 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN
                           => n103);
   U122 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82,
                           C1 => IN5(3), C2 => n79, ZN => n102);
   U123 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => Z(31));
   U124 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n163);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_5 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_5;

architecture SYN_bhv of mux5to1_numBit32_5 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n91, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n160);
   U2 : BUF_X1 port map( A => n158, Z => n4);
   U3 : BUF_X1 port map( A => n158, Z => n77);
   U4 : BUF_X1 port map( A => n158, Z => n78);
   U5 : BUF_X1 port map( A => n89, Z => n1);
   U6 : BUF_X1 port map( A => n89, Z => n2);
   U7 : NOR2_X1 port map( A1 => n88, A2 => n93, ZN => n158);
   U8 : INV_X1 port map( A => n94, ZN => n88);
   U9 : BUF_X1 port map( A => n89, Z => n3);
   U10 : NOR4_X1 port map( A1 => n92, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n94);
   U11 : BUF_X1 port map( A => n160, Z => n82);
   U12 : BUF_X1 port map( A => n160, Z => n83);
   U13 : BUF_X1 port map( A => n159, Z => n79);
   U14 : BUF_X1 port map( A => n159, Z => n80);
   U15 : BUF_X1 port map( A => n161, Z => n85);
   U16 : BUF_X1 port map( A => n161, Z => n86);
   U17 : BUF_X1 port map( A => n160, Z => n84);
   U18 : NOR2_X1 port map( A1 => n91, A2 => n90, ZN => n93);
   U19 : BUF_X1 port map( A => n159, Z => n81);
   U20 : BUF_X1 port map( A => n161, Z => n87);
   U21 : INV_X1 port map( A => n95, ZN => n89);
   U22 : AOI21_X1 port map( B1 => n94, B2 => n93, A => n92, ZN => n95);
   U23 : NOR3_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => n90, ZN => n161);
   U24 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n92);
   U25 : INV_X1 port map( A => SEL_in(0), ZN => n90);
   U26 : AND3_X1 port map( A1 => n90, A2 => n91, A3 => SEL_in(2), ZN => n159);
   U27 : INV_X1 port map( A => SEL_in(1), ZN => n91);
   U28 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(7));
   U29 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82, 
                           C1 => IN5(7), C2 => n79, ZN => n110);
   U30 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN 
                           => n111);
   U31 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(8));
   U32 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN 
                           => n113);
   U33 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82, 
                           C1 => IN5(8), C2 => n79, ZN => n112);
   U34 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(9));
   U35 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN 
                           => n115);
   U36 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82, 
                           C1 => IN5(9), C2 => n79, ZN => n114);
   U37 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(10));
   U38 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n117);
   U39 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => n82
                           , C1 => IN5(10), C2 => n79, ZN => n116);
   U40 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(11));
   U41 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n119);
   U42 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => n82
                           , C1 => IN5(11), C2 => n79, ZN => n118);
   U43 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(12));
   U44 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2, 
                           ZN => n121);
   U45 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => n83
                           , C1 => IN5(12), C2 => n80, ZN => n120);
   U46 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(13));
   U47 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2, 
                           ZN => n123);
   U48 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => n83
                           , C1 => IN5(13), C2 => n80, ZN => n122);
   U49 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(14));
   U50 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n125);
   U51 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n124);
   U52 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(15));
   U53 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n127);
   U54 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n126);
   U55 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(16));
   U56 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2, 
                           ZN => n129);
   U57 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n128);
   U58 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(17));
   U59 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2, 
                           ZN => n131);
   U60 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n130);
   U61 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(18));
   U62 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2, 
                           ZN => n133);
   U63 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n132);
   U64 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(19));
   U65 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n135);
   U66 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n134);
   U67 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(20));
   U68 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n137);
   U69 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n136);
   U70 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(21));
   U71 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n139);
   U72 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n138);
   U73 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(22));
   U74 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n141);
   U75 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n140);
   U76 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(23));
   U77 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n143);
   U78 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n142);
   U79 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Z(24));
   U80 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3, 
                           ZN => n145);
   U81 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n144);
   U82 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Z(25));
   U83 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3, 
                           ZN => n147);
   U84 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84
                           , C1 => IN5(25), C2 => n81, ZN => n146);
   U85 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(26));
   U86 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3, 
                           ZN => n149);
   U87 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84
                           , C1 => IN5(26), C2 => n81, ZN => n148);
   U88 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Z(27));
   U89 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3, 
                           ZN => n151);
   U90 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84
                           , C1 => IN5(27), C2 => n81, ZN => n150);
   U91 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Z(28));
   U92 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3, 
                           ZN => n153);
   U93 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => n84
                           , C1 => IN5(28), C2 => n81, ZN => n152);
   U94 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Z(29));
   U95 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3, 
                           ZN => n155);
   U96 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => n84
                           , C1 => IN5(29), C2 => n81, ZN => n154);
   U97 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => Z(30));
   U98 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3, 
                           ZN => n157);
   U99 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => n84
                           , C1 => IN5(30), C2 => n81, ZN => n156);
   U100 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(6));
   U101 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN
                           => n109);
   U102 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82,
                           C1 => IN5(6), C2 => n79, ZN => n108);
   U103 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(0));
   U104 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN
                           => n97);
   U105 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82,
                           C1 => IN5(0), C2 => n79, ZN => n96);
   U106 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(1));
   U107 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN
                           => n99);
   U108 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82,
                           C1 => IN5(1), C2 => n79, ZN => n98);
   U110 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(2));
   U111 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN
                           => n101);
   U112 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82,
                           C1 => IN5(2), C2 => n79, ZN => n100);
   U113 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(3));
   U114 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN
                           => n103);
   U115 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82,
                           C1 => IN5(3), C2 => n79, ZN => n102);
   U116 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(4));
   U117 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN
                           => n105);
   U118 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82,
                           C1 => IN5(4), C2 => n79, ZN => n104);
   U119 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(5));
   U120 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN
                           => n107);
   U121 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82,
                           C1 => IN5(5), C2 => n79, ZN => n106);
   U122 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => Z(31));
   U123 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n163);
   U124 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => 
                           n84, C1 => IN5(31), C2 => n81, ZN => n162);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_4 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_4;

architecture SYN_bhv of mux5to1_numBit32_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n91, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n160);
   U2 : BUF_X1 port map( A => n158, Z => n4);
   U3 : BUF_X1 port map( A => n158, Z => n77);
   U4 : BUF_X1 port map( A => n158, Z => n78);
   U5 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => n84,
                           C1 => IN5(31), C2 => n81, ZN => n162);
   U6 : BUF_X1 port map( A => n89, Z => n1);
   U7 : BUF_X1 port map( A => n89, Z => n2);
   U8 : NOR2_X1 port map( A1 => n88, A2 => n93, ZN => n158);
   U9 : INV_X1 port map( A => n94, ZN => n88);
   U10 : BUF_X1 port map( A => n89, Z => n3);
   U11 : NOR4_X1 port map( A1 => n92, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n94);
   U12 : BUF_X1 port map( A => n160, Z => n82);
   U13 : BUF_X1 port map( A => n160, Z => n83);
   U14 : BUF_X1 port map( A => n159, Z => n79);
   U15 : BUF_X1 port map( A => n159, Z => n80);
   U16 : BUF_X1 port map( A => n161, Z => n85);
   U17 : BUF_X1 port map( A => n161, Z => n86);
   U18 : BUF_X1 port map( A => n160, Z => n84);
   U19 : NOR2_X1 port map( A1 => n91, A2 => n90, ZN => n93);
   U20 : BUF_X1 port map( A => n159, Z => n81);
   U21 : BUF_X1 port map( A => n161, Z => n87);
   U22 : INV_X1 port map( A => n95, ZN => n89);
   U23 : AOI21_X1 port map( B1 => n94, B2 => n93, A => n92, ZN => n95);
   U24 : NOR3_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => n90, ZN => n161);
   U25 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n92);
   U26 : INV_X1 port map( A => SEL_in(0), ZN => n90);
   U27 : AND3_X1 port map( A1 => n90, A2 => n91, A3 => SEL_in(2), ZN => n159);
   U28 : INV_X1 port map( A => SEL_in(1), ZN => n91);
   U29 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(9));
   U30 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82, 
                           C1 => IN5(9), C2 => n79, ZN => n114);
   U31 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN 
                           => n115);
   U32 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(10));
   U33 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n117);
   U34 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => n82
                           , C1 => IN5(10), C2 => n79, ZN => n116);
   U35 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(11));
   U36 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n119);
   U37 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => n82
                           , C1 => IN5(11), C2 => n79, ZN => n118);
   U38 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(12));
   U39 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2, 
                           ZN => n121);
   U40 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => n83
                           , C1 => IN5(12), C2 => n80, ZN => n120);
   U41 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(13));
   U42 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2, 
                           ZN => n123);
   U43 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => n83
                           , C1 => IN5(13), C2 => n80, ZN => n122);
   U44 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(14));
   U45 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n125);
   U46 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n124);
   U47 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(15));
   U48 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n127);
   U49 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n126);
   U50 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(16));
   U51 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2, 
                           ZN => n129);
   U52 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n128);
   U53 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(17));
   U54 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2, 
                           ZN => n131);
   U55 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n130);
   U56 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(18));
   U57 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2, 
                           ZN => n133);
   U58 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n132);
   U59 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(19));
   U60 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n135);
   U61 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n134);
   U62 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(20));
   U63 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n137);
   U64 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n136);
   U65 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(21));
   U66 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n139);
   U67 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n138);
   U68 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(22));
   U69 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n141);
   U70 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n140);
   U71 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(23));
   U72 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n143);
   U73 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n142);
   U74 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Z(24));
   U75 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3, 
                           ZN => n145);
   U76 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n144);
   U77 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Z(25));
   U78 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3, 
                           ZN => n147);
   U79 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84
                           , C1 => IN5(25), C2 => n81, ZN => n146);
   U80 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(26));
   U81 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3, 
                           ZN => n149);
   U82 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84
                           , C1 => IN5(26), C2 => n81, ZN => n148);
   U83 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Z(27));
   U84 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3, 
                           ZN => n151);
   U85 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84
                           , C1 => IN5(27), C2 => n81, ZN => n150);
   U86 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Z(28));
   U87 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3, 
                           ZN => n153);
   U88 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => n84
                           , C1 => IN5(28), C2 => n81, ZN => n152);
   U89 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Z(29));
   U90 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3, 
                           ZN => n155);
   U91 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => n84
                           , C1 => IN5(29), C2 => n81, ZN => n154);
   U92 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => Z(30));
   U93 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3, 
                           ZN => n157);
   U94 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => n84
                           , C1 => IN5(30), C2 => n81, ZN => n156);
   U95 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(8));
   U96 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN 
                           => n113);
   U97 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82, 
                           C1 => IN5(8), C2 => n79, ZN => n112);
   U98 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(0));
   U99 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN 
                           => n97);
   U100 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82,
                           C1 => IN5(0), C2 => n79, ZN => n96);
   U101 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(1));
   U102 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN
                           => n99);
   U103 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82,
                           C1 => IN5(1), C2 => n79, ZN => n98);
   U104 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(2));
   U105 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN
                           => n101);
   U106 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82,
                           C1 => IN5(2), C2 => n79, ZN => n100);
   U107 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(3));
   U108 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN
                           => n103);
   U110 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82,
                           C1 => IN5(3), C2 => n79, ZN => n102);
   U111 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(4));
   U112 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN
                           => n105);
   U113 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82,
                           C1 => IN5(4), C2 => n79, ZN => n104);
   U114 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(5));
   U115 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN
                           => n107);
   U116 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82,
                           C1 => IN5(5), C2 => n79, ZN => n106);
   U117 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(6));
   U118 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN
                           => n109);
   U119 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82,
                           C1 => IN5(6), C2 => n79, ZN => n108);
   U120 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(7));
   U121 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN
                           => n111);
   U122 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82,
                           C1 => IN5(7), C2 => n79, ZN => n110);
   U123 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => Z(31));
   U124 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n163);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_3 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_3;

architecture SYN_bhv of mux5to1_numBit32_3 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n90, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n160);
   U2 : BUF_X1 port map( A => n158, Z => n4);
   U3 : BUF_X1 port map( A => n158, Z => n77);
   U4 : BUF_X1 port map( A => n158, Z => n78);
   U5 : BUF_X1 port map( A => n89, Z => n1);
   U6 : BUF_X1 port map( A => n89, Z => n2);
   U7 : NOR2_X1 port map( A1 => n88, A2 => n93, ZN => n158);
   U8 : INV_X1 port map( A => n94, ZN => n88);
   U9 : BUF_X1 port map( A => n89, Z => n3);
   U10 : NOR4_X1 port map( A1 => n92, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n94);
   U11 : BUF_X1 port map( A => n160, Z => n82);
   U12 : BUF_X1 port map( A => n160, Z => n83);
   U13 : BUF_X1 port map( A => n159, Z => n79);
   U14 : BUF_X1 port map( A => n159, Z => n80);
   U15 : BUF_X1 port map( A => n161, Z => n85);
   U16 : BUF_X1 port map( A => n161, Z => n86);
   U17 : BUF_X1 port map( A => n160, Z => n84);
   U18 : NOR2_X1 port map( A1 => n90, A2 => n91, ZN => n93);
   U19 : BUF_X1 port map( A => n159, Z => n81);
   U20 : BUF_X1 port map( A => n161, Z => n87);
   U21 : INV_X1 port map( A => n95, ZN => n89);
   U22 : AOI21_X1 port map( B1 => n94, B2 => n93, A => n92, ZN => n95);
   U23 : NOR3_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => n91, ZN => n161);
   U24 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n92);
   U25 : INV_X1 port map( A => SEL_in(0), ZN => n91);
   U26 : AND3_X1 port map( A1 => n91, A2 => n90, A3 => SEL_in(2), ZN => n159);
   U27 : INV_X1 port map( A => SEL_in(1), ZN => n90);
   U28 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(11));
   U29 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => n82
                           , C1 => IN5(11), C2 => n79, ZN => n118);
   U30 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n119);
   U31 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(12));
   U32 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2, 
                           ZN => n121);
   U33 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => n83
                           , C1 => IN5(12), C2 => n80, ZN => n120);
   U34 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(13));
   U35 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2, 
                           ZN => n123);
   U36 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => n83
                           , C1 => IN5(13), C2 => n80, ZN => n122);
   U37 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(14));
   U38 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n125);
   U39 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n124);
   U40 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(15));
   U41 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n127);
   U42 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n126);
   U43 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(16));
   U44 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2, 
                           ZN => n129);
   U45 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n128);
   U46 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(17));
   U47 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2, 
                           ZN => n131);
   U48 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n130);
   U49 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(18));
   U50 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2, 
                           ZN => n133);
   U51 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n132);
   U52 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(19));
   U53 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n135);
   U54 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n134);
   U55 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(20));
   U56 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n137);
   U57 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n136);
   U58 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(21));
   U59 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n139);
   U60 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n138);
   U61 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(22));
   U62 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n141);
   U63 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n140);
   U64 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(23));
   U65 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n143);
   U66 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n142);
   U67 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Z(24));
   U68 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3, 
                           ZN => n145);
   U69 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n144);
   U70 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Z(25));
   U71 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3, 
                           ZN => n147);
   U72 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84
                           , C1 => IN5(25), C2 => n81, ZN => n146);
   U73 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(26));
   U74 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3, 
                           ZN => n149);
   U75 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84
                           , C1 => IN5(26), C2 => n81, ZN => n148);
   U76 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Z(27));
   U77 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3, 
                           ZN => n151);
   U78 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84
                           , C1 => IN5(27), C2 => n81, ZN => n150);
   U79 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Z(28));
   U80 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3, 
                           ZN => n153);
   U81 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => n84
                           , C1 => IN5(28), C2 => n81, ZN => n152);
   U82 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Z(29));
   U83 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3, 
                           ZN => n155);
   U84 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => n84
                           , C1 => IN5(29), C2 => n81, ZN => n154);
   U85 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => Z(30));
   U86 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3, 
                           ZN => n157);
   U87 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => n84
                           , C1 => IN5(30), C2 => n81, ZN => n156);
   U88 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(10));
   U89 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n117);
   U90 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => n82
                           , C1 => IN5(10), C2 => n79, ZN => n116);
   U91 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(0));
   U92 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN 
                           => n97);
   U93 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82, 
                           C1 => IN5(0), C2 => n79, ZN => n96);
   U94 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(1));
   U95 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN 
                           => n99);
   U96 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82, 
                           C1 => IN5(1), C2 => n79, ZN => n98);
   U97 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(2));
   U98 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN 
                           => n101);
   U99 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82, 
                           C1 => IN5(2), C2 => n79, ZN => n100);
   U100 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(3));
   U101 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN
                           => n103);
   U102 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82,
                           C1 => IN5(3), C2 => n79, ZN => n102);
   U103 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(4));
   U104 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN
                           => n105);
   U105 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82,
                           C1 => IN5(4), C2 => n79, ZN => n104);
   U106 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(5));
   U107 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN
                           => n107);
   U108 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82,
                           C1 => IN5(5), C2 => n79, ZN => n106);
   U110 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(6));
   U111 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN
                           => n109);
   U112 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82,
                           C1 => IN5(6), C2 => n79, ZN => n108);
   U113 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(7));
   U114 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN
                           => n111);
   U115 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82,
                           C1 => IN5(7), C2 => n79, ZN => n110);
   U116 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(8));
   U117 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN
                           => n113);
   U118 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82,
                           C1 => IN5(8), C2 => n79, ZN => n112);
   U119 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(9));
   U120 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN
                           => n115);
   U121 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82,
                           C1 => IN5(9), C2 => n79, ZN => n114);
   U122 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => Z(31));
   U123 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n163);
   U124 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => 
                           n84, C1 => IN5(31), C2 => n81, ZN => n162);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_2 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_2;

architecture SYN_bhv of mux5to1_numBit32_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n91, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n160);
   U2 : BUF_X1 port map( A => n158, Z => n4);
   U3 : BUF_X1 port map( A => n158, Z => n77);
   U4 : BUF_X1 port map( A => n158, Z => n78);
   U5 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => n84,
                           C1 => IN5(31), C2 => n81, ZN => n162);
   U6 : BUF_X1 port map( A => n89, Z => n1);
   U7 : BUF_X1 port map( A => n89, Z => n2);
   U8 : NOR2_X1 port map( A1 => n88, A2 => n93, ZN => n158);
   U9 : INV_X1 port map( A => n94, ZN => n88);
   U10 : BUF_X1 port map( A => n89, Z => n3);
   U11 : NOR4_X1 port map( A1 => n92, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n94);
   U12 : BUF_X1 port map( A => n160, Z => n82);
   U13 : BUF_X1 port map( A => n160, Z => n83);
   U14 : BUF_X1 port map( A => n159, Z => n79);
   U15 : BUF_X1 port map( A => n159, Z => n80);
   U16 : BUF_X1 port map( A => n161, Z => n85);
   U17 : BUF_X1 port map( A => n161, Z => n86);
   U18 : BUF_X1 port map( A => n160, Z => n84);
   U19 : NOR2_X1 port map( A1 => n91, A2 => n90, ZN => n93);
   U20 : BUF_X1 port map( A => n159, Z => n81);
   U21 : BUF_X1 port map( A => n161, Z => n87);
   U22 : INV_X1 port map( A => n95, ZN => n89);
   U23 : AOI21_X1 port map( B1 => n94, B2 => n93, A => n92, ZN => n95);
   U24 : NOR3_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => n90, ZN => n161);
   U25 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n92);
   U26 : INV_X1 port map( A => SEL_in(0), ZN => n90);
   U27 : AND3_X1 port map( A1 => n90, A2 => n91, A3 => SEL_in(2), ZN => n159);
   U28 : INV_X1 port map( A => SEL_in(1), ZN => n91);
   U29 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(13));
   U30 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => n83
                           , C1 => IN5(13), C2 => n80, ZN => n122);
   U31 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2, 
                           ZN => n123);
   U32 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(14));
   U33 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n125);
   U34 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n124);
   U35 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(15));
   U36 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n127);
   U37 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n126);
   U38 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(16));
   U39 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2, 
                           ZN => n129);
   U40 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n128);
   U41 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(17));
   U42 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2, 
                           ZN => n131);
   U43 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n130);
   U44 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(18));
   U45 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2, 
                           ZN => n133);
   U46 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n132);
   U47 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(19));
   U48 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n135);
   U49 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n134);
   U50 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(20));
   U51 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n137);
   U52 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n136);
   U53 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(21));
   U54 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n139);
   U55 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n138);
   U56 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(22));
   U57 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n141);
   U58 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n140);
   U59 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(23));
   U60 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n143);
   U61 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n142);
   U62 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Z(24));
   U63 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3, 
                           ZN => n145);
   U64 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n144);
   U65 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Z(25));
   U66 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3, 
                           ZN => n147);
   U67 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84
                           , C1 => IN5(25), C2 => n81, ZN => n146);
   U68 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(26));
   U69 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3, 
                           ZN => n149);
   U70 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84
                           , C1 => IN5(26), C2 => n81, ZN => n148);
   U71 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Z(27));
   U72 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3, 
                           ZN => n151);
   U73 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84
                           , C1 => IN5(27), C2 => n81, ZN => n150);
   U74 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Z(28));
   U75 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3, 
                           ZN => n153);
   U76 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => n84
                           , C1 => IN5(28), C2 => n81, ZN => n152);
   U77 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Z(29));
   U78 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3, 
                           ZN => n155);
   U79 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => n84
                           , C1 => IN5(29), C2 => n81, ZN => n154);
   U80 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => Z(30));
   U81 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3, 
                           ZN => n157);
   U82 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => n84
                           , C1 => IN5(30), C2 => n81, ZN => n156);
   U83 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(12));
   U84 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2, 
                           ZN => n121);
   U85 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => n83
                           , C1 => IN5(12), C2 => n80, ZN => n120);
   U86 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(0));
   U87 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN 
                           => n97);
   U88 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82, 
                           C1 => IN5(0), C2 => n79, ZN => n96);
   U89 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(1));
   U90 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN 
                           => n99);
   U91 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82, 
                           C1 => IN5(1), C2 => n79, ZN => n98);
   U92 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(2));
   U93 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN 
                           => n101);
   U94 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82, 
                           C1 => IN5(2), C2 => n79, ZN => n100);
   U95 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(3));
   U96 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN 
                           => n103);
   U97 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82, 
                           C1 => IN5(3), C2 => n79, ZN => n102);
   U98 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(4));
   U99 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN 
                           => n105);
   U100 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82,
                           C1 => IN5(4), C2 => n79, ZN => n104);
   U101 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(5));
   U102 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN
                           => n107);
   U103 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82,
                           C1 => IN5(5), C2 => n79, ZN => n106);
   U104 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(6));
   U105 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN
                           => n109);
   U106 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82,
                           C1 => IN5(6), C2 => n79, ZN => n108);
   U107 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(7));
   U108 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN
                           => n111);
   U110 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82,
                           C1 => IN5(7), C2 => n79, ZN => n110);
   U111 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(8));
   U112 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN
                           => n113);
   U113 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82,
                           C1 => IN5(8), C2 => n79, ZN => n112);
   U114 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(9));
   U115 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN
                           => n115);
   U116 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82,
                           C1 => IN5(9), C2 => n79, ZN => n114);
   U117 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(10));
   U118 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n117);
   U119 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => 
                           n82, C1 => IN5(10), C2 => n79, ZN => n116);
   U120 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(11));
   U121 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n119);
   U122 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => 
                           n82, C1 => IN5(11), C2 => n79, ZN => n118);
   U123 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => Z(31));
   U124 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n163);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_1 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_1;

architecture SYN_bhv of mux5to1_numBit32_1 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n91, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n160);
   U2 : BUF_X1 port map( A => n158, Z => n4);
   U3 : BUF_X1 port map( A => n158, Z => n77);
   U4 : BUF_X1 port map( A => n158, Z => n78);
   U5 : BUF_X1 port map( A => n89, Z => n1);
   U6 : BUF_X1 port map( A => n89, Z => n2);
   U7 : NOR2_X1 port map( A1 => n88, A2 => n93, ZN => n158);
   U8 : INV_X1 port map( A => n94, ZN => n88);
   U9 : BUF_X1 port map( A => n89, Z => n3);
   U10 : NOR4_X1 port map( A1 => n92, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n94);
   U11 : BUF_X1 port map( A => n160, Z => n82);
   U12 : BUF_X1 port map( A => n160, Z => n83);
   U13 : BUF_X1 port map( A => n159, Z => n79);
   U14 : BUF_X1 port map( A => n159, Z => n80);
   U15 : BUF_X1 port map( A => n161, Z => n85);
   U16 : BUF_X1 port map( A => n161, Z => n86);
   U17 : BUF_X1 port map( A => n160, Z => n84);
   U18 : NOR2_X1 port map( A1 => n91, A2 => n90, ZN => n93);
   U19 : BUF_X1 port map( A => n159, Z => n81);
   U20 : BUF_X1 port map( A => n161, Z => n87);
   U21 : INV_X1 port map( A => n95, ZN => n89);
   U22 : AOI21_X1 port map( B1 => n94, B2 => n93, A => n92, ZN => n95);
   U23 : NOR3_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => n90, ZN => n161);
   U24 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n92);
   U25 : INV_X1 port map( A => SEL_in(0), ZN => n90);
   U26 : AND3_X1 port map( A1 => n90, A2 => n91, A3 => SEL_in(2), ZN => n159);
   U27 : INV_X1 port map( A => SEL_in(1), ZN => n91);
   U28 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(15));
   U29 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n126);
   U30 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n127);
   U31 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(16));
   U32 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2, 
                           ZN => n129);
   U33 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n128);
   U34 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(17));
   U35 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2, 
                           ZN => n131);
   U36 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n130);
   U37 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(18));
   U38 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2, 
                           ZN => n133);
   U39 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n132);
   U40 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(19));
   U41 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n135);
   U42 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n134);
   U43 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(20));
   U44 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n137);
   U45 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n136);
   U46 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(21));
   U47 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n139);
   U48 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n138);
   U49 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(22));
   U50 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n141);
   U51 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n140);
   U52 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(23));
   U53 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n143);
   U54 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n142);
   U55 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => Z(24));
   U56 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3, 
                           ZN => n145);
   U57 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n144);
   U58 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => Z(25));
   U59 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3, 
                           ZN => n147);
   U60 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84
                           , C1 => IN5(25), C2 => n81, ZN => n146);
   U61 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(26));
   U62 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3, 
                           ZN => n149);
   U63 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84
                           , C1 => IN5(26), C2 => n81, ZN => n148);
   U64 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => Z(27));
   U65 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3, 
                           ZN => n151);
   U66 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84
                           , C1 => IN5(27), C2 => n81, ZN => n150);
   U67 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => Z(28));
   U68 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3, 
                           ZN => n153);
   U69 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => n84
                           , C1 => IN5(28), C2 => n81, ZN => n152);
   U70 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Z(29));
   U71 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3, 
                           ZN => n155);
   U72 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => n84
                           , C1 => IN5(29), C2 => n81, ZN => n154);
   U73 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => Z(30));
   U74 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3, 
                           ZN => n157);
   U75 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => n84
                           , C1 => IN5(30), C2 => n81, ZN => n156);
   U76 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(14));
   U77 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n125);
   U78 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n124);
   U79 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(0));
   U80 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN 
                           => n97);
   U81 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82, 
                           C1 => IN5(0), C2 => n79, ZN => n96);
   U82 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(1));
   U83 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN 
                           => n99);
   U84 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82, 
                           C1 => IN5(1), C2 => n79, ZN => n98);
   U85 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(2));
   U86 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN 
                           => n101);
   U87 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82, 
                           C1 => IN5(2), C2 => n79, ZN => n100);
   U88 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(3));
   U89 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN 
                           => n103);
   U90 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82, 
                           C1 => IN5(3), C2 => n79, ZN => n102);
   U91 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(4));
   U92 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN 
                           => n105);
   U93 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82, 
                           C1 => IN5(4), C2 => n79, ZN => n104);
   U94 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(5));
   U95 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN 
                           => n107);
   U96 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82, 
                           C1 => IN5(5), C2 => n79, ZN => n106);
   U97 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(6));
   U98 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN 
                           => n109);
   U99 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82, 
                           C1 => IN5(6), C2 => n79, ZN => n108);
   U100 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(7));
   U101 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN
                           => n111);
   U102 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82,
                           C1 => IN5(7), C2 => n79, ZN => n110);
   U103 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(8));
   U104 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN
                           => n113);
   U105 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82,
                           C1 => IN5(8), C2 => n79, ZN => n112);
   U106 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(9));
   U107 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN
                           => n115);
   U108 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82,
                           C1 => IN5(9), C2 => n79, ZN => n114);
   U110 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(10));
   U111 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n117);
   U112 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => 
                           n82, C1 => IN5(10), C2 => n79, ZN => n116);
   U113 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(11));
   U114 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n119);
   U115 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => 
                           n82, C1 => IN5(11), C2 => n79, ZN => n118);
   U116 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(12));
   U117 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2,
                           ZN => n121);
   U118 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => 
                           n83, C1 => IN5(12), C2 => n80, ZN => n120);
   U119 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(13));
   U120 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2,
                           ZN => n123);
   U121 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => 
                           n83, C1 => IN5(13), C2 => n80, ZN => n122);
   U122 : NAND2_X1 port map( A1 => n163, A2 => n162, ZN => Z(31));
   U123 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n163);
   U124 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => 
                           n84, C1 => IN5(31), C2 => n81, ZN => n162);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_4 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_4;

architecture SYN_bhv of mux41_NBIT32_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n145, Z => n73);
   U2 : BUF_X1 port map( A => n147, Z => n79);
   U3 : BUF_X1 port map( A => n144, Z => n70);
   U4 : BUF_X1 port map( A => n146, Z => n76);
   U5 : BUF_X1 port map( A => n145, Z => n72);
   U6 : BUF_X1 port map( A => n147, Z => n78);
   U7 : BUF_X1 port map( A => n144, Z => n1);
   U8 : BUF_X1 port map( A => n146, Z => n75);
   U9 : BUF_X1 port map( A => n145, Z => n74);
   U10 : BUF_X1 port map( A => n147, Z => n80);
   U11 : BUF_X1 port map( A => n144, Z => n71);
   U12 : BUF_X1 port map( A => n146, Z => n77);
   U13 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n145);
   U14 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n144);
   U15 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n147);
   U16 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n146);
   U17 : INV_X1 port map( A => S(0), ZN => n81);
   U18 : NAND2_X1 port map( A1 => n83, A2 => n82, ZN => Z(0));
   U19 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(3));
   U20 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(1));
   U21 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(4));
   U22 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN =>
                           n135);
   U23 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN =>
                           n134);
   U24 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(8));
   U25 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n143);
   U26 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n142);
   U27 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => Z(12));
   U28 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n89);
   U29 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN 
                           => n88);
   U30 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(16));
   U31 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n97);
   U32 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n96);
   U33 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(24));
   U34 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN 
                           => n115);
   U35 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN 
                           => n114);
   U36 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(5));
   U37 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN =>
                           n137);
   U38 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN =>
                           n136);
   U39 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(9));
   U40 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN =>
                           n149);
   U41 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN =>
                           n148);
   U42 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => Z(13));
   U43 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n91);
   U44 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN 
                           => n90);
   U45 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(17));
   U46 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n99);
   U47 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n98);
   U48 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(25));
   U49 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n117);
   U50 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n116);
   U51 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(2));
   U52 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN =>
                           n127);
   U53 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN =>
                           n126);
   U54 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(6));
   U55 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n139);
   U56 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n138);
   U57 : NAND2_X1 port map( A1 => n85, A2 => n84, ZN => Z(10));
   U58 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n85);
   U59 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN 
                           => n84);
   U60 : NAND2_X1 port map( A1 => n93, A2 => n92, ZN => Z(14));
   U61 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n93);
   U62 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN 
                           => n92);
   U63 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(18));
   U64 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n101);
   U65 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n100);
   U66 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(26));
   U67 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n119);
   U68 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n118);
   U69 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(22));
   U70 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n111);
   U71 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n110);
   U72 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(21));
   U73 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n109);
   U74 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n108);
   U75 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(20));
   U76 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN 
                           => n107);
   U77 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN 
                           => n106);
   U78 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(30));
   U79 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN 
                           => n129);
   U80 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN 
                           => n128);
   U81 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(29));
   U82 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n125);
   U83 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n124);
   U84 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(28));
   U85 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n123);
   U86 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n122);
   U87 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(7));
   U88 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n141);
   U89 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n140);
   U90 : NAND2_X1 port map( A1 => n87, A2 => n86, ZN => Z(11));
   U91 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n87);
   U92 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN 
                           => n86);
   U93 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => Z(15));
   U94 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n95);
   U95 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN 
                           => n94);
   U96 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(19));
   U97 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n103);
   U98 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN 
                           => n102);
   U99 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(23));
   U100 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN
                           => n113);
   U101 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN
                           => n112);
   U102 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(27));
   U103 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN
                           => n121);
   U104 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN
                           => n120);
   U105 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(31));
   U106 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN
                           => n131);
   U107 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN
                           => n130);
   U108 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN 
                           => n133);
   U109 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN 
                           => n132);
   U110 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN =>
                           n105);
   U111 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN 
                           => n104);
   U112 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN =>
                           n83);
   U113 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN 
                           => n82);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_3 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_3;

architecture SYN_bhv of mux41_NBIT32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n145, Z => n72);
   U2 : BUF_X1 port map( A => n147, Z => n78);
   U3 : BUF_X1 port map( A => n145, Z => n73);
   U4 : BUF_X1 port map( A => n147, Z => n79);
   U5 : BUF_X1 port map( A => n144, Z => n1);
   U6 : BUF_X1 port map( A => n146, Z => n75);
   U7 : BUF_X1 port map( A => n144, Z => n70);
   U8 : BUF_X1 port map( A => n146, Z => n76);
   U9 : BUF_X1 port map( A => n145, Z => n74);
   U10 : BUF_X1 port map( A => n147, Z => n80);
   U11 : BUF_X1 port map( A => n144, Z => n71);
   U12 : BUF_X1 port map( A => n146, Z => n77);
   U13 : NAND2_X1 port map( A1 => n83, A2 => n82, ZN => Z(0));
   U14 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n82);
   U15 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n83);
   U16 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(1));
   U17 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN =>
                           n104);
   U18 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN => 
                           n105);
   U19 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(3));
   U20 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN =>
                           n132);
   U21 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN =>
                           n133);
   U22 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(4));
   U23 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN =>
                           n134);
   U24 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN =>
                           n135);
   U25 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(8));
   U26 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n142);
   U27 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n143);
   U28 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => Z(12));
   U29 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN 
                           => n88);
   U30 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n89);
   U31 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(16));
   U32 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n96);
   U33 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n97);
   U34 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(24));
   U35 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN 
                           => n114);
   U36 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN 
                           => n115);
   U37 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(5));
   U38 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN =>
                           n136);
   U39 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN =>
                           n137);
   U40 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(9));
   U41 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN =>
                           n148);
   U42 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN =>
                           n149);
   U43 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => Z(13));
   U44 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN 
                           => n90);
   U45 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n91);
   U46 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(17));
   U47 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n98);
   U48 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n99);
   U49 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(25));
   U50 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n116);
   U51 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n117);
   U52 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(2));
   U53 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN =>
                           n126);
   U54 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN =>
                           n127);
   U55 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(6));
   U56 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n138);
   U57 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n139);
   U58 : NAND2_X1 port map( A1 => n85, A2 => n84, ZN => Z(10));
   U59 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN 
                           => n84);
   U60 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n85);
   U61 : NAND2_X1 port map( A1 => n93, A2 => n92, ZN => Z(14));
   U62 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN 
                           => n92);
   U63 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n93);
   U64 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(18));
   U65 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n100);
   U66 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n101);
   U67 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(26));
   U68 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n118);
   U69 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n119);
   U70 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(22));
   U71 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n110);
   U72 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n111);
   U73 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(21));
   U74 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n108);
   U75 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n109);
   U76 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(20));
   U77 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN 
                           => n106);
   U78 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN 
                           => n107);
   U79 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(30));
   U80 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN 
                           => n128);
   U81 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN 
                           => n129);
   U82 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(29));
   U83 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n124);
   U84 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n125);
   U85 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(28));
   U86 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n122);
   U87 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n123);
   U88 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(7));
   U89 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n140);
   U90 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n141);
   U91 : NAND2_X1 port map( A1 => n87, A2 => n86, ZN => Z(11));
   U92 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN 
                           => n86);
   U93 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n87);
   U94 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => Z(15));
   U95 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN 
                           => n94);
   U96 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n95);
   U97 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(19));
   U98 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN 
                           => n102);
   U99 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n103);
   U100 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(23));
   U101 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN
                           => n112);
   U102 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN
                           => n113);
   U103 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(27));
   U104 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN
                           => n120);
   U105 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN
                           => n121);
   U106 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(31));
   U107 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN
                           => n130);
   U108 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN
                           => n131);
   U109 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n145);
   U110 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n144);
   U111 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n147);
   U112 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n146);
   U113 : INV_X1 port map( A => S(0), ZN => n81);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_2 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_2;

architecture SYN_bhv of mux41_NBIT32_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n5, n6, n7, n20, n21, n22, n23, n26, n27, n28, n29, n30, n31,
      n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n48
      , n49, n50, n51, n52, n53, n54, n55, n70, n71, n72, n73, n74, n75, n76, 
      n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91
      , n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => S(1), A2 => n34, ZN => n1);
   U2 : AND2_X1 port map( A1 => S(0), A2 => n33, ZN => n4);
   U3 : AND2_X1 port map( A1 => n33, A2 => n34, ZN => n5);
   U4 : AND2_X1 port map( A1 => S(0), A2 => S(1), ZN => n6);
   U5 : BUF_X1 port map( A => n5, Z => n27);
   U6 : BUF_X1 port map( A => n5, Z => n28);
   U7 : BUF_X1 port map( A => n5, Z => n29);
   U8 : BUF_X1 port map( A => n1, Z => n7);
   U9 : BUF_X1 port map( A => n4, Z => n31);
   U10 : BUF_X1 port map( A => n4, Z => n30);
   U11 : BUF_X1 port map( A => n1, Z => n20);
   U12 : BUF_X1 port map( A => n4, Z => n32);
   U13 : BUF_X1 port map( A => n1, Z => n21);
   U14 : BUF_X1 port map( A => n6, Z => n22);
   U15 : BUF_X1 port map( A => n6, Z => n23);
   U16 : BUF_X1 port map( A => n6, Z => n26);
   U17 : NAND2_X1 port map( A1 => n88, A2 => n87, ZN => Z(11));
   U18 : AOI22_X1 port map( A1 => D(11), A2 => n22, B1 => C(11), B2 => n7, ZN 
                           => n87);
   U19 : AOI22_X1 port map( A1 => B(11), A2 => n30, B1 => A(11), B2 => n27, ZN 
                           => n88);
   U20 : NAND2_X1 port map( A1 => n106, A2 => n105, ZN => Z(5));
   U21 : AOI22_X1 port map( A1 => D(5), A2 => n22, B1 => C(5), B2 => n7, ZN => 
                           n105);
   U22 : AOI22_X1 port map( A1 => B(5), A2 => n30, B1 => A(5), B2 => n27, ZN =>
                           n106);
   U23 : NAND2_X1 port map( A1 => n112, A2 => n111, ZN => Z(8));
   U24 : AOI22_X1 port map( A1 => D(8), A2 => n23, B1 => C(8), B2 => n20, ZN =>
                           n111);
   U25 : AOI22_X1 port map( A1 => B(8), A2 => n31, B1 => A(8), B2 => n28, ZN =>
                           n112);
   U26 : NAND2_X1 port map( A1 => n110, A2 => n109, ZN => Z(7));
   U27 : AOI22_X1 port map( A1 => D(7), A2 => n23, B1 => C(7), B2 => n20, ZN =>
                           n109);
   U28 : AOI22_X1 port map( A1 => B(7), A2 => n31, B1 => A(7), B2 => n28, ZN =>
                           n110);
   U29 : NAND2_X1 port map( A1 => n104, A2 => n103, ZN => Z(4));
   U30 : AOI22_X1 port map( A1 => D(4), A2 => n22, B1 => C(4), B2 => n7, ZN => 
                           n103);
   U31 : AOI22_X1 port map( A1 => B(4), A2 => n30, B1 => A(4), B2 => n27, ZN =>
                           n104);
   U32 : AOI22_X1 port map( A1 => D(15), A2 => n22, B1 => C(15), B2 => n7, ZN 
                           => n95);
   U33 : NAND2_X1 port map( A1 => n108, A2 => n107, ZN => Z(6));
   U34 : AOI22_X1 port map( A1 => D(6), A2 => n23, B1 => C(6), B2 => n20, ZN =>
                           n107);
   U35 : AOI22_X1 port map( A1 => B(6), A2 => n31, B1 => A(6), B2 => n28, ZN =>
                           n108);
   U36 : NAND2_X1 port map( A1 => n114, A2 => n113, ZN => Z(9));
   U37 : AOI22_X1 port map( A1 => D(9), A2 => n23, B1 => C(9), B2 => n20, ZN =>
                           n113);
   U38 : AOI22_X1 port map( A1 => B(9), A2 => n31, B1 => A(9), B2 => n28, ZN =>
                           n114);
   U39 : NAND2_X1 port map( A1 => n92, A2 => n91, ZN => Z(13));
   U40 : AOI22_X1 port map( A1 => D(13), A2 => n22, B1 => C(13), B2 => n7, ZN 
                           => n91);
   U41 : AOI22_X1 port map( A1 => B(13), A2 => n30, B1 => A(13), B2 => n27, ZN 
                           => n92);
   U42 : NAND2_X1 port map( A1 => n94, A2 => n93, ZN => Z(14));
   U43 : AOI22_X1 port map( A1 => D(14), A2 => n22, B1 => C(14), B2 => n7, ZN 
                           => n93);
   U44 : AOI22_X1 port map( A1 => B(14), A2 => n30, B1 => A(14), B2 => n27, ZN 
                           => n94);
   U45 : NAND2_X1 port map( A1 => n84, A2 => n83, ZN => Z(0));
   U46 : AOI22_X1 port map( A1 => B(0), A2 => n30, B1 => A(0), B2 => n27, ZN =>
                           n84);
   U47 : AOI22_X1 port map( A1 => D(0), A2 => n22, B1 => C(0), B2 => n7, ZN => 
                           n83);
   U48 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => Z(1));
   U49 : AOI22_X1 port map( A1 => B(1), A2 => n30, B1 => A(1), B2 => n27, ZN =>
                           n98);
   U50 : AOI22_X1 port map( A1 => D(1), A2 => n22, B1 => C(1), B2 => n7, ZN => 
                           n97);
   U51 : NAND2_X1 port map( A1 => n100, A2 => n99, ZN => Z(2));
   U52 : AOI22_X1 port map( A1 => B(2), A2 => n30, B1 => A(2), B2 => n27, ZN =>
                           n100);
   U53 : AOI22_X1 port map( A1 => D(2), A2 => n22, B1 => C(2), B2 => n7, ZN => 
                           n99);
   U54 : NAND2_X1 port map( A1 => n102, A2 => n101, ZN => Z(3));
   U55 : AOI22_X1 port map( A1 => B(3), A2 => n30, B1 => A(3), B2 => n27, ZN =>
                           n102);
   U56 : AOI22_X1 port map( A1 => D(3), A2 => n22, B1 => C(3), B2 => n7, ZN => 
                           n101);
   U57 : NAND2_X1 port map( A1 => n86, A2 => n85, ZN => Z(10));
   U58 : AOI22_X1 port map( A1 => D(10), A2 => n22, B1 => C(10), B2 => n7, ZN 
                           => n85);
   U59 : AOI22_X1 port map( A1 => B(10), A2 => n30, B1 => A(10), B2 => n27, ZN 
                           => n86);
   U60 : NAND2_X1 port map( A1 => n90, A2 => n89, ZN => Z(12));
   U61 : AOI22_X1 port map( A1 => D(12), A2 => n22, B1 => C(12), B2 => n7, ZN 
                           => n89);
   U62 : AOI22_X1 port map( A1 => B(12), A2 => n30, B1 => A(12), B2 => n27, ZN 
                           => n90);
   U63 : NAND2_X1 port map( A1 => n96, A2 => n95, ZN => Z(15));
   U64 : AOI22_X1 port map( A1 => B(15), A2 => n30, B1 => A(15), B2 => n27, ZN 
                           => n96);
   U65 : INV_X1 port map( A => S(1), ZN => n33);
   U66 : INV_X1 port map( A => S(0), ZN => n34);
   U67 : AOI22_X1 port map( A1 => B(16), A2 => n32, B1 => A(16), B2 => n29, ZN 
                           => n36);
   U68 : AOI22_X1 port map( A1 => D(16), A2 => n26, B1 => C(16), B2 => n21, ZN 
                           => n35);
   U69 : NAND2_X1 port map( A1 => n36, A2 => n35, ZN => Z(16));
   U70 : AOI22_X1 port map( A1 => B(17), A2 => n32, B1 => A(17), B2 => n29, ZN 
                           => n38);
   U71 : AOI22_X1 port map( A1 => D(17), A2 => n26, B1 => C(17), B2 => n21, ZN 
                           => n37);
   U72 : NAND2_X1 port map( A1 => n38, A2 => n37, ZN => Z(17));
   U73 : AOI22_X1 port map( A1 => B(18), A2 => n32, B1 => A(18), B2 => n29, ZN 
                           => n40);
   U74 : AOI22_X1 port map( A1 => D(18), A2 => n26, B1 => C(18), B2 => n21, ZN 
                           => n39);
   U75 : NAND2_X1 port map( A1 => n40, A2 => n39, ZN => Z(18));
   U76 : AOI22_X1 port map( A1 => B(19), A2 => n31, B1 => A(19), B2 => n28, ZN 
                           => n42);
   U77 : AOI22_X1 port map( A1 => D(19), A2 => n23, B1 => C(19), B2 => n20, ZN 
                           => n41);
   U78 : NAND2_X1 port map( A1 => n42, A2 => n41, ZN => Z(19));
   U79 : AOI22_X1 port map( A1 => B(20), A2 => n31, B1 => A(20), B2 => n28, ZN 
                           => n44);
   U80 : AOI22_X1 port map( A1 => D(20), A2 => n23, B1 => C(20), B2 => n20, ZN 
                           => n43);
   U81 : NAND2_X1 port map( A1 => n44, A2 => n43, ZN => Z(20));
   U82 : AOI22_X1 port map( A1 => B(21), A2 => n31, B1 => A(21), B2 => n28, ZN 
                           => n48);
   U83 : AOI22_X1 port map( A1 => D(21), A2 => n23, B1 => C(21), B2 => n20, ZN 
                           => n45);
   U84 : NAND2_X1 port map( A1 => n48, A2 => n45, ZN => Z(21));
   U85 : AOI22_X1 port map( A1 => B(22), A2 => n31, B1 => A(22), B2 => n28, ZN 
                           => n50);
   U86 : AOI22_X1 port map( A1 => D(22), A2 => n23, B1 => C(22), B2 => n20, ZN 
                           => n49);
   U87 : NAND2_X1 port map( A1 => n50, A2 => n49, ZN => Z(22));
   U88 : AOI22_X1 port map( A1 => B(23), A2 => n31, B1 => A(23), B2 => n28, ZN 
                           => n52);
   U89 : AOI22_X1 port map( A1 => D(23), A2 => n23, B1 => C(23), B2 => n20, ZN 
                           => n51);
   U90 : NAND2_X1 port map( A1 => n52, A2 => n51, ZN => Z(23));
   U91 : AOI22_X1 port map( A1 => B(24), A2 => n31, B1 => A(24), B2 => n28, ZN 
                           => n54);
   U92 : AOI22_X1 port map( A1 => D(24), A2 => n23, B1 => C(24), B2 => n20, ZN 
                           => n53);
   U93 : NAND2_X1 port map( A1 => n54, A2 => n53, ZN => Z(24));
   U94 : AOI22_X1 port map( A1 => B(25), A2 => n31, B1 => A(25), B2 => n28, ZN 
                           => n70);
   U95 : AOI22_X1 port map( A1 => D(25), A2 => n23, B1 => C(25), B2 => n20, ZN 
                           => n55);
   U96 : NAND2_X1 port map( A1 => n70, A2 => n55, ZN => Z(25));
   U97 : AOI22_X1 port map( A1 => B(26), A2 => n31, B1 => A(26), B2 => n28, ZN 
                           => n72);
   U98 : AOI22_X1 port map( A1 => D(26), A2 => n23, B1 => C(26), B2 => n20, ZN 
                           => n71);
   U99 : NAND2_X1 port map( A1 => n72, A2 => n71, ZN => Z(26));
   U100 : AOI22_X1 port map( A1 => B(27), A2 => n31, B1 => A(27), B2 => n28, ZN
                           => n74);
   U101 : AOI22_X1 port map( A1 => D(27), A2 => n23, B1 => C(27), B2 => n20, ZN
                           => n73);
   U102 : NAND2_X1 port map( A1 => n74, A2 => n73, ZN => Z(27));
   U103 : AOI22_X1 port map( A1 => B(28), A2 => n31, B1 => A(28), B2 => n28, ZN
                           => n76);
   U104 : AOI22_X1 port map( A1 => D(28), A2 => n23, B1 => C(28), B2 => n20, ZN
                           => n75);
   U105 : NAND2_X1 port map( A1 => n76, A2 => n75, ZN => Z(28));
   U106 : AOI22_X1 port map( A1 => B(29), A2 => n31, B1 => A(29), B2 => n28, ZN
                           => n78);
   U107 : AOI22_X1 port map( A1 => D(29), A2 => n23, B1 => C(29), B2 => n20, ZN
                           => n77);
   U108 : NAND2_X1 port map( A1 => n78, A2 => n77, ZN => Z(29));
   U109 : AOI22_X1 port map( A1 => B(30), A2 => n31, B1 => A(30), B2 => n28, ZN
                           => n80);
   U110 : AOI22_X1 port map( A1 => D(30), A2 => n23, B1 => C(30), B2 => n20, ZN
                           => n79);
   U111 : NAND2_X1 port map( A1 => n80, A2 => n79, ZN => Z(30));
   U112 : AOI22_X1 port map( A1 => B(31), A2 => n31, B1 => A(31), B2 => n28, ZN
                           => n82);
   U113 : AOI22_X1 port map( A1 => D(31), A2 => n23, B1 => C(31), B2 => n20, ZN
                           => n81);
   U114 : NAND2_X1 port map( A1 => n82, A2 => n81, ZN => Z(31));

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_1 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_1;

architecture SYN_bhv of mux41_NBIT32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n145, Z => n72);
   U2 : BUF_X1 port map( A => n145, Z => n73);
   U3 : BUF_X1 port map( A => n146, Z => n75);
   U4 : BUF_X1 port map( A => n146, Z => n76);
   U5 : BUF_X1 port map( A => n145, Z => n74);
   U6 : BUF_X1 port map( A => n146, Z => n77);
   U7 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n145);
   U8 : BUF_X1 port map( A => n147, Z => n78);
   U9 : BUF_X1 port map( A => n147, Z => n79);
   U10 : BUF_X1 port map( A => n144, Z => n1);
   U11 : BUF_X1 port map( A => n144, Z => n70);
   U12 : BUF_X1 port map( A => n147, Z => n80);
   U13 : BUF_X1 port map( A => n144, Z => n71);
   U14 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n146);
   U15 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n144);
   U16 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n82);
   U17 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN =>
                           n137);
   U18 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n139);
   U19 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n141);
   U20 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN =>
                           n149);
   U21 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN 
                           => n131);
   U22 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n85);
   U23 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n87);
   U24 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n91);
   U25 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n93);
   U26 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n95);
   U27 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n99);
   U28 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n101);
   U29 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n103);
   U30 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n109);
   U31 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n111);
   U32 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN 
                           => n113);
   U33 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n117);
   U34 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n119);
   U35 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN 
                           => n121);
   U36 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n125);
   U37 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN 
                           => n129);
   U38 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n147);
   U39 : INV_X1 port map( A => S(0), ZN => n81);
   U40 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN =>
                           n133);
   U41 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN =>
                           n135);
   U42 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n143);
   U43 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN => 
                           n105);
   U44 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN =>
                           n127);
   U45 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n89);
   U46 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n97);
   U47 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN 
                           => n107);
   U48 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN 
                           => n115);
   U49 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n123);
   U50 : NAND2_X1 port map( A1 => n131, A2 => n130, ZN => Z(31));
   U51 : NAND2_X1 port map( A1 => n83, A2 => n82, ZN => Z(0));
   U52 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n83);
   U53 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN 
                           => n130);
   U54 : NAND2_X1 port map( A1 => n133, A2 => n132, ZN => Z(3));
   U55 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN =>
                           n132);
   U56 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => Z(4));
   U57 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN =>
                           n134);
   U58 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => Z(5));
   U59 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN =>
                           n136);
   U60 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => Z(6));
   U61 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n138);
   U62 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => Z(7));
   U63 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n140);
   U64 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => Z(8));
   U65 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n142);
   U66 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => Z(9));
   U67 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN =>
                           n148);
   U68 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => Z(15));
   U69 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN 
                           => n94);
   U70 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => Z(16));
   U71 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n96);
   U72 : NAND2_X1 port map( A1 => n99, A2 => n98, ZN => Z(17));
   U73 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n98);
   U74 : NAND2_X1 port map( A1 => n101, A2 => n100, ZN => Z(18));
   U75 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n100);
   U76 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => Z(19));
   U77 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN 
                           => n102);
   U78 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => Z(20));
   U79 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN 
                           => n106);
   U80 : NAND2_X1 port map( A1 => n109, A2 => n108, ZN => Z(21));
   U81 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n108);
   U82 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => Z(22));
   U83 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n110);
   U84 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => Z(23));
   U85 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN 
                           => n112);
   U86 : NAND2_X1 port map( A1 => n115, A2 => n114, ZN => Z(24));
   U87 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN 
                           => n114);
   U88 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => Z(25));
   U89 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n116);
   U90 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => Z(26));
   U91 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n118);
   U92 : NAND2_X1 port map( A1 => n121, A2 => n120, ZN => Z(27));
   U93 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN 
                           => n120);
   U94 : NAND2_X1 port map( A1 => n123, A2 => n122, ZN => Z(28));
   U95 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n122);
   U96 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => Z(29));
   U97 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n124);
   U98 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => Z(30));
   U99 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN 
                           => n128);
   U100 : NAND2_X1 port map( A1 => n93, A2 => n92, ZN => Z(14));
   U101 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN
                           => n92);
   U102 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => Z(1));
   U103 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN 
                           => n104);
   U104 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => Z(2));
   U105 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN 
                           => n126);
   U106 : NAND2_X1 port map( A1 => n85, A2 => n84, ZN => Z(10));
   U107 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN
                           => n84);
   U108 : NAND2_X1 port map( A1 => n87, A2 => n86, ZN => Z(11));
   U109 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN
                           => n86);
   U110 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => Z(12));
   U111 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN
                           => n88);
   U112 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => Z(13));
   U113 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN
                           => n90);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT5_2 is

   port( A, B : in std_logic_vector (4 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (4 downto 0));

end mux21_NBIT5_2;

architecture SYN_bhv of mux21_NBIT5_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n14, n15, n16, n17, n18 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => S, Z => n1);
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : INV_X1 port map( A => n18, ZN => Z(4));
   U4 : INV_X1 port map( A => n15, ZN => Z(1));
   U5 : INV_X1 port map( A => n16, ZN => Z(2));
   U6 : INV_X1 port map( A => n17, ZN => Z(3));
   U7 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => n1, ZN => 
                           n17);
   U8 : INV_X1 port map( A => n14, ZN => Z(0));
   U9 : AOI22_X1 port map( A1 => A(1), A2 => n3, B1 => B(1), B2 => n1, ZN => 
                           n15);
   U10 : AOI22_X1 port map( A1 => A(2), A2 => n3, B1 => B(2), B2 => n1, ZN => 
                           n16);
   U11 : AOI22_X1 port map( A1 => A(0), A2 => n3, B1 => B(0), B2 => n1, ZN => 
                           n14);
   U12 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => n2, B2 => B(4), ZN => 
                           n18);
   U13 : INV_X1 port map( A => n2, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT5_1 is

   port( A, B : in std_logic_vector (4 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (4 downto 0));

end mux21_NBIT5_1;

architecture SYN_bhv of mux21_NBIT5_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n14, n15, n16, n17, n18 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => S, Z => n1);
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : INV_X1 port map( A => n15, ZN => Z(1));
   U4 : AOI22_X1 port map( A1 => A(1), A2 => n3, B1 => B(1), B2 => n1, ZN => 
                           n15);
   U5 : INV_X1 port map( A => n16, ZN => Z(2));
   U6 : AOI22_X1 port map( A1 => A(2), A2 => n3, B1 => B(2), B2 => n1, ZN => 
                           n16);
   U7 : INV_X1 port map( A => n17, ZN => Z(3));
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => n1, ZN => 
                           n17);
   U9 : INV_X1 port map( A => n18, ZN => Z(4));
   U10 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => n2, B2 => B(4), ZN => 
                           n18);
   U11 : INV_X1 port map( A => n14, ZN => Z(0));
   U12 : AOI22_X1 port map( A1 => A(0), A2 => n3, B1 => B(0), B2 => n1, ZN => 
                           n14);
   U13 : INV_X1 port map( A => n2, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_4 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_4;

architecture SYN_bhv of regn_N5_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n16, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n21);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n17, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n22);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n18, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n23);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n19, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n24);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n20, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n25);
   U2 : OAI21_X1 port map( B1 => n21, B2 => EN, A => n26, ZN => n16);
   U3 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n26);
   U4 : OAI21_X1 port map( B1 => n24, B2 => EN, A => n29, ZN => n19);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n29);
   U6 : OAI21_X1 port map( B1 => n23, B2 => EN, A => n28, ZN => n18);
   U7 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n28);
   U8 : OAI21_X1 port map( B1 => n22, B2 => EN, A => n27, ZN => n17);
   U9 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n27);
   U10 : OAI21_X1 port map( B1 => n25, B2 => EN, A => n30, ZN => n20);
   U11 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n30);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_3 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_3;

architecture SYN_bhv of regn_N5_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n16, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n21);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n17, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n22);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n18, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n23);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n19, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n24);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n20, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n25);
   U2 : OAI21_X1 port map( B1 => n21, B2 => EN, A => n26, ZN => n16);
   U3 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n26);
   U4 : OAI21_X1 port map( B1 => n24, B2 => EN, A => n29, ZN => n19);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n29);
   U6 : OAI21_X1 port map( B1 => n23, B2 => EN, A => n28, ZN => n18);
   U7 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n28);
   U8 : OAI21_X1 port map( B1 => n22, B2 => EN, A => n27, ZN => n17);
   U9 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n27);
   U10 : OAI21_X1 port map( B1 => n25, B2 => EN, A => n30, ZN => n20);
   U11 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n30);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_2 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_2;

architecture SYN_bhv of regn_N5_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n16, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n21);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n17, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n22);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n18, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n23);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n19, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n24);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n20, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n25);
   U2 : OAI21_X1 port map( B1 => n24, B2 => EN, A => n29, ZN => n19);
   U3 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n29);
   U4 : OAI21_X1 port map( B1 => n23, B2 => EN, A => n28, ZN => n18);
   U5 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n28);
   U6 : OAI21_X1 port map( B1 => n22, B2 => EN, A => n27, ZN => n17);
   U7 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n27);
   U8 : OAI21_X1 port map( B1 => n21, B2 => EN, A => n26, ZN => n16);
   U9 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n26);
   U10 : OAI21_X1 port map( B1 => n25, B2 => EN, A => n30, ZN => n20);
   U11 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n30);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_1 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_1;

architecture SYN_bhv of regn_N5_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n16, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n21);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n17, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n22);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n18, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n23);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n19, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n24);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n20, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n25);
   U2 : OAI21_X1 port map( B1 => n25, B2 => EN, A => n30, ZN => n20);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n30);
   U4 : OAI21_X1 port map( B1 => n24, B2 => EN, A => n29, ZN => n19);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n29);
   U6 : OAI21_X1 port map( B1 => n23, B2 => EN, A => n28, ZN => n18);
   U7 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n28);
   U8 : OAI21_X1 port map( B1 => n22, B2 => EN, A => n27, ZN => n17);
   U9 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n27);
   U10 : OAI21_X1 port map( B1 => n21, B2 => EN, A => n26, ZN => n16);
   U11 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n26);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_9 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_9;

architecture SYN_bhv of regn_N32_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U6 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);
   U7 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U8 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U9 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U10 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U11 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U12 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U13 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U14 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U15 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U16 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U17 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U18 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U22 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U23 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U24 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U25 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U26 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U27 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U28 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U29 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U30 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U31 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U32 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U33 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U34 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U35 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U36 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U37 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U38 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U39 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U40 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U41 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U42 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U43 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U44 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U45 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U46 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U47 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U48 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U49 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U50 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U51 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U52 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U53 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U54 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U55 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U56 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U57 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U58 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U59 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U60 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U61 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U62 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U63 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U64 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U65 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U66 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U67 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U68 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_8 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_8;

architecture SYN_bhv of regn_N32_8 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110
      , n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n_1154 : std_logic;

begin
   
   DOUT_reg_25_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n101, Q => 
                           DOUT(25), QN => n140);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n101, Q => 
                           DOUT(24), QN => n141);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n100, Q => 
                           DOUT(23), QN => n142);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n100, Q => 
                           DOUT(22), QN => n143);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n100, Q => 
                           DOUT(21), QN => n144);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n100, Q => 
                           DOUT(20), QN => n145);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n100, Q => 
                           DOUT(19), QN => n146);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n100, Q => 
                           DOUT(18), QN => n147);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n100, Q => 
                           DOUT(17), QN => n148);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n100, Q => 
                           DOUT(16), QN => n149);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n100, Q => 
                           DOUT(15), QN => n150);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n100, Q => 
                           DOUT(14), QN => n151);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n100, Q => 
                           DOUT(13), QN => n152);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n100, Q => 
                           DOUT(12), QN => n153);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n99, Q => 
                           DOUT(11), QN => n154);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n99, Q => 
                           DOUT(10), QN => n155);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n99, Q => 
                           DOUT(9), QN => n156);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n99, Q => 
                           DOUT(8), QN => n157);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n99, Q => 
                           DOUT(7), QN => n158);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n99, Q => 
                           DOUT(6), QN => n159);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n99, Q => 
                           DOUT(5), QN => n160);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n99, Q => 
                           DOUT(4), QN => n161);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n99, Q => 
                           DOUT(3), QN => n162);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n99, Q => 
                           DOUT(2), QN => n163);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n132, CK => CLK, RN => n99, Q => 
                           DOUT(1), QN => n164);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n133, CK => CLK, RN => n99, Q => 
                           DOUT(0), QN => n165);
   DOUT_reg_31_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n101, Q => 
                           DOUT(31), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n101, Q => 
                           n_1154, QN => n137);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n101, Q => 
                           DOUT(30), QN => n135);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n101, Q => 
                           DOUT(29), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n101, Q => 
                           DOUT(26), QN => n139);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n101, Q => 
                           DOUT(27), QN => n138);
   U2 : INV_X2 port map( A => n137, ZN => DOUT(28));
   U3 : BUF_X1 port map( A => RST, Z => n99);
   U4 : BUF_X1 port map( A => RST, Z => n100);
   U5 : BUF_X1 port map( A => RST, Z => n101);
   U6 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n170);
   U7 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n171);
   U8 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n168);
   U9 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n167);
   U10 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n166);
   U11 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n169);
   U12 : OAI21_X1 port map( B1 => n164, B2 => EN, A => n196, ZN => n132);
   U13 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n196);
   U14 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U15 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n195);
   U16 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U17 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n194);
   U18 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U19 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n193);
   U20 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U21 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n192);
   U22 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U23 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n191);
   U24 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U25 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n190);
   U26 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U27 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n189);
   U28 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U29 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n187);
   U30 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U31 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n186);
   U32 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U33 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n185);
   U34 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U35 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n184);
   U36 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U37 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n183);
   U38 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U39 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n182);
   U40 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U41 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n181);
   U42 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U43 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n180);
   U44 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U45 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n179);
   U46 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U47 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n178);
   U48 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U49 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n177);
   U50 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U51 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n176);
   U52 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U53 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n175);
   U54 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U55 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n174);
   U56 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U57 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n173);
   U58 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U59 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n172);
   U60 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U61 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n188);
   U62 : OAI21_X1 port map( B1 => n165, B2 => EN, A => n197, ZN => n133);
   U63 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n197);
   U64 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U65 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U66 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U67 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U68 : OAI21_X1 port map( B1 => EN, B2 => n137, A => n169, ZN => n105);
   U69 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_7 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_7;

architecture SYN_bhv of regn_N32_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U6 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U7 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U8 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U9 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U10 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U11 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U12 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U13 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U14 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U15 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U16 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U17 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U18 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U19 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U20 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U21 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U22 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U23 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U24 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U25 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U26 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U27 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U28 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U29 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U30 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U31 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U32 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U33 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U34 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U35 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U36 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U37 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U38 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U39 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U40 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U41 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U42 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U43 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U44 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U45 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U46 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U47 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U48 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U49 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U50 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U51 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U52 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U53 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U54 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U55 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U56 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U57 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U58 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U59 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U60 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U61 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U62 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U63 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U64 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U65 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U66 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);
   U67 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U68 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_6 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_6;

architecture SYN_bhv of regn_N32_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U6 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U7 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U8 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U9 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U10 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U11 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U12 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U13 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U14 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U15 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U16 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U17 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U18 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);
   U19 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U20 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U21 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U22 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U23 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U24 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U25 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U26 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U27 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U28 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U29 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U30 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U31 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U32 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U33 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U34 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U35 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U36 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U37 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U38 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U39 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U40 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U41 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U42 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U43 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U44 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U45 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U46 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U47 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U48 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U49 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U50 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U51 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U52 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U53 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U54 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U55 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U56 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U57 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U58 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U59 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U60 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U61 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U62 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U63 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U64 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U65 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U66 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U67 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U68 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_5 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_5;

architecture SYN_bhv of regn_N32_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_4 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_4;

architecture SYN_bhv of regn_N32_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_3 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_3;

architecture SYN_bhv of regn_N32_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_2 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_2;

architecture SYN_bhv of regn_N32_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : BUF_X1 port map( A => RST, Z => n97);
   U3 : BUF_X1 port map( A => RST, Z => n98);
   U4 : BUF_X1 port map( A => RST, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_1 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_1;

architecture SYN_bhv of regn_N32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n99, Q => 
                           DOUT(31), QN => n132);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n99, Q => 
                           DOUT(30), QN => n133);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n99, Q => 
                           DOUT(29), QN => n134);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n99, Q => 
                           DOUT(28), QN => n135);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n104, CK => CLK, RN => n99, Q => 
                           DOUT(27), QN => n136);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n105, CK => CLK, RN => n99, Q => 
                           DOUT(26), QN => n137);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n106, CK => CLK, RN => n99, Q => 
                           DOUT(25), QN => n138);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n107, CK => CLK, RN => n99, Q => 
                           DOUT(24), QN => n139);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n108, CK => CLK, RN => n98, Q => 
                           DOUT(23), QN => n140);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n109, CK => CLK, RN => n98, Q => 
                           DOUT(22), QN => n141);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n110, CK => CLK, RN => n98, Q => 
                           DOUT(21), QN => n142);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n111, CK => CLK, RN => n98, Q => 
                           DOUT(20), QN => n143);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n112, CK => CLK, RN => n98, Q => 
                           DOUT(19), QN => n144);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n113, CK => CLK, RN => n98, Q => 
                           DOUT(18), QN => n145);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n114, CK => CLK, RN => n98, Q => 
                           DOUT(17), QN => n146);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n115, CK => CLK, RN => n98, Q => 
                           DOUT(16), QN => n147);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n116, CK => CLK, RN => n98, Q => 
                           DOUT(15), QN => n148);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n117, CK => CLK, RN => n98, Q => 
                           DOUT(14), QN => n149);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n118, CK => CLK, RN => n98, Q => 
                           DOUT(13), QN => n150);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n119, CK => CLK, RN => n98, Q => 
                           DOUT(12), QN => n151);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n120, CK => CLK, RN => n97, Q => 
                           DOUT(11), QN => n152);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n121, CK => CLK, RN => n97, Q => 
                           DOUT(10), QN => n153);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n122, CK => CLK, RN => n97, Q => 
                           DOUT(9), QN => n154);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n123, CK => CLK, RN => n97, Q => 
                           DOUT(8), QN => n155);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n124, CK => CLK, RN => n97, Q => 
                           DOUT(7), QN => n156);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n125, CK => CLK, RN => n97, Q => 
                           DOUT(6), QN => n157);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n126, CK => CLK, RN => n97, Q => 
                           DOUT(5), QN => n158);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n127, CK => CLK, RN => n97, Q => 
                           DOUT(4), QN => n159);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n128, CK => CLK, RN => n97, Q => 
                           DOUT(3), QN => n160);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n129, CK => CLK, RN => n97, Q => 
                           DOUT(2), QN => n161);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n130, CK => CLK, RN => n97, Q => 
                           DOUT(1), QN => n162);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n131, CK => CLK, RN => n97, Q => 
                           DOUT(0), QN => n163);
   U2 : OAI21_X1 port map( B1 => n163, B2 => EN, A => n195, ZN => n131);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n195);
   U4 : OAI21_X1 port map( B1 => n162, B2 => EN, A => n194, ZN => n130);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n194);
   U6 : OAI21_X1 port map( B1 => n161, B2 => EN, A => n193, ZN => n129);
   U7 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n193);
   U8 : OAI21_X1 port map( B1 => n160, B2 => EN, A => n192, ZN => n128);
   U9 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n192);
   U10 : OAI21_X1 port map( B1 => n159, B2 => EN, A => n191, ZN => n127);
   U11 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n191);
   U12 : OAI21_X1 port map( B1 => n158, B2 => EN, A => n190, ZN => n126);
   U13 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n190);
   U14 : OAI21_X1 port map( B1 => n157, B2 => EN, A => n189, ZN => n125);
   U15 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n189);
   U16 : OAI21_X1 port map( B1 => n156, B2 => EN, A => n188, ZN => n124);
   U17 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n188);
   U18 : OAI21_X1 port map( B1 => n155, B2 => EN, A => n187, ZN => n123);
   U19 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n187);
   U20 : OAI21_X1 port map( B1 => n154, B2 => EN, A => n186, ZN => n122);
   U21 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n186);
   U22 : OAI21_X1 port map( B1 => n153, B2 => EN, A => n185, ZN => n121);
   U23 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n185);
   U24 : OAI21_X1 port map( B1 => n152, B2 => EN, A => n184, ZN => n120);
   U25 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n184);
   U26 : OAI21_X1 port map( B1 => n151, B2 => EN, A => n183, ZN => n119);
   U27 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n183);
   U28 : OAI21_X1 port map( B1 => n150, B2 => EN, A => n182, ZN => n118);
   U29 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n182);
   U30 : OAI21_X1 port map( B1 => n149, B2 => EN, A => n181, ZN => n117);
   U31 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n181);
   U32 : OAI21_X1 port map( B1 => n148, B2 => EN, A => n180, ZN => n116);
   U33 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n180);
   U34 : OAI21_X1 port map( B1 => n147, B2 => EN, A => n179, ZN => n115);
   U35 : NAND2_X1 port map( A1 => DIN(16), A2 => EN, ZN => n179);
   U36 : OAI21_X1 port map( B1 => n146, B2 => EN, A => n178, ZN => n114);
   U37 : NAND2_X1 port map( A1 => DIN(17), A2 => EN, ZN => n178);
   U38 : OAI21_X1 port map( B1 => n145, B2 => EN, A => n177, ZN => n113);
   U39 : NAND2_X1 port map( A1 => DIN(18), A2 => EN, ZN => n177);
   U40 : OAI21_X1 port map( B1 => n144, B2 => EN, A => n176, ZN => n112);
   U41 : NAND2_X1 port map( A1 => DIN(19), A2 => EN, ZN => n176);
   U42 : OAI21_X1 port map( B1 => n143, B2 => EN, A => n175, ZN => n111);
   U43 : NAND2_X1 port map( A1 => DIN(20), A2 => EN, ZN => n175);
   U44 : OAI21_X1 port map( B1 => n142, B2 => EN, A => n174, ZN => n110);
   U45 : NAND2_X1 port map( A1 => DIN(21), A2 => EN, ZN => n174);
   U46 : OAI21_X1 port map( B1 => n141, B2 => EN, A => n173, ZN => n109);
   U47 : NAND2_X1 port map( A1 => DIN(22), A2 => EN, ZN => n173);
   U48 : OAI21_X1 port map( B1 => n140, B2 => EN, A => n172, ZN => n108);
   U49 : NAND2_X1 port map( A1 => DIN(23), A2 => EN, ZN => n172);
   U50 : OAI21_X1 port map( B1 => n139, B2 => EN, A => n171, ZN => n107);
   U51 : NAND2_X1 port map( A1 => DIN(24), A2 => EN, ZN => n171);
   U52 : OAI21_X1 port map( B1 => n138, B2 => EN, A => n170, ZN => n106);
   U53 : NAND2_X1 port map( A1 => DIN(25), A2 => EN, ZN => n170);
   U54 : OAI21_X1 port map( B1 => n137, B2 => EN, A => n169, ZN => n105);
   U55 : NAND2_X1 port map( A1 => DIN(26), A2 => EN, ZN => n169);
   U56 : OAI21_X1 port map( B1 => n136, B2 => EN, A => n168, ZN => n104);
   U57 : NAND2_X1 port map( A1 => DIN(27), A2 => EN, ZN => n168);
   U58 : OAI21_X1 port map( B1 => n135, B2 => EN, A => n167, ZN => n103);
   U59 : NAND2_X1 port map( A1 => DIN(28), A2 => EN, ZN => n167);
   U60 : OAI21_X1 port map( B1 => n134, B2 => EN, A => n166, ZN => n102);
   U61 : NAND2_X1 port map( A1 => DIN(29), A2 => EN, ZN => n166);
   U62 : OAI21_X1 port map( B1 => n133, B2 => EN, A => n165, ZN => n101);
   U63 : NAND2_X1 port map( A1 => DIN(30), A2 => EN, ZN => n165);
   U64 : OAI21_X1 port map( B1 => n132, B2 => EN, A => n164, ZN => n100);
   U65 : NAND2_X1 port map( A1 => DIN(31), A2 => EN, ZN => n164);
   U66 : BUF_X1 port map( A => RST, Z => n97);
   U67 : BUF_X1 port map( A => RST, Z => n98);
   U68 : BUF_X1 port map( A => RST, Z => n99);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_6 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_6;

architecture SYN_bhv of mux21_NBIT32_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n15, ZN => n5);
   U2 : INV_X1 port map( A => n15, ZN => n4);
   U3 : BUF_X1 port map( A => n3, Z => n13);
   U4 : BUF_X1 port map( A => n2, Z => n12);
   U5 : BUF_X1 port map( A => n2, Z => n10);
   U6 : BUF_X1 port map( A => n1, Z => n9);
   U7 : BUF_X1 port map( A => n2, Z => n11);
   U8 : BUF_X1 port map( A => n3, Z => n15);
   U9 : BUF_X1 port map( A => n3, Z => n14);
   U10 : BUF_X1 port map( A => n1, Z => n8);
   U11 : BUF_X1 port map( A => n1, Z => n7);
   U12 : BUF_X1 port map( A => S, Z => n3);
   U13 : BUF_X1 port map( A => S, Z => n2);
   U14 : BUF_X1 port map( A => S, Z => n1);
   U15 : INV_X1 port map( A => n104, ZN => Z(31));
   U16 : INV_X1 port map( A => n105, ZN => Z(3));
   U17 : INV_X1 port map( A => n106, ZN => Z(4));
   U18 : INV_X1 port map( A => n107, ZN => Z(5));
   U19 : INV_X1 port map( A => n108, ZN => Z(6));
   U20 : INV_X1 port map( A => n110, ZN => Z(8));
   U21 : INV_X1 port map( A => n81, ZN => Z(10));
   U22 : INV_X1 port map( A => n109, ZN => Z(7));
   U23 : INV_X1 port map( A => n102, ZN => Z(2));
   U24 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => n8, ZN => 
                           n102);
   U25 : INV_X1 port map( A => n82, ZN => Z(11));
   U26 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => B(11), B2 => n14, ZN 
                           => n82);
   U27 : INV_X1 port map( A => n83, ZN => Z(12));
   U28 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => B(12), B2 => n13, ZN 
                           => n83);
   U29 : INV_X1 port map( A => n84, ZN => Z(13));
   U30 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n13, ZN 
                           => n84);
   U31 : INV_X1 port map( A => n85, ZN => Z(14));
   U32 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n13, ZN 
                           => n85);
   U33 : INV_X1 port map( A => n86, ZN => Z(15));
   U34 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n13, ZN 
                           => n86);
   U35 : INV_X1 port map( A => n87, ZN => Z(16));
   U36 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => B(16), B2 => n12, ZN 
                           => n87);
   U37 : INV_X1 port map( A => n88, ZN => Z(17));
   U38 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n12, ZN 
                           => n88);
   U39 : INV_X1 port map( A => n89, ZN => Z(18));
   U40 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => B(18), B2 => n12, ZN 
                           => n89);
   U41 : INV_X1 port map( A => n90, ZN => Z(19));
   U42 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => B(19), B2 => n12, ZN 
                           => n90);
   U43 : INV_X1 port map( A => n92, ZN => Z(20));
   U44 : AOI22_X1 port map( A1 => A(20), A2 => n5, B1 => B(20), B2 => n11, ZN 
                           => n92);
   U45 : INV_X1 port map( A => n93, ZN => Z(21));
   U46 : AOI22_X1 port map( A1 => A(21), A2 => n5, B1 => B(21), B2 => n11, ZN 
                           => n93);
   U47 : INV_X1 port map( A => n94, ZN => Z(22));
   U48 : AOI22_X1 port map( A1 => A(22), A2 => n5, B1 => B(22), B2 => n10, ZN 
                           => n94);
   U49 : INV_X1 port map( A => n95, ZN => Z(23));
   U50 : AOI22_X1 port map( A1 => A(23), A2 => n5, B1 => B(23), B2 => n10, ZN 
                           => n95);
   U51 : INV_X1 port map( A => n96, ZN => Z(24));
   U52 : AOI22_X1 port map( A1 => A(24), A2 => n5, B1 => B(24), B2 => n10, ZN 
                           => n96);
   U53 : INV_X1 port map( A => n97, ZN => Z(25));
   U54 : AOI22_X1 port map( A1 => A(25), A2 => n5, B1 => B(25), B2 => n10, ZN 
                           => n97);
   U55 : INV_X1 port map( A => n98, ZN => Z(26));
   U56 : AOI22_X1 port map( A1 => A(26), A2 => n5, B1 => B(26), B2 => n9, ZN =>
                           n98);
   U57 : INV_X1 port map( A => n99, ZN => Z(27));
   U58 : AOI22_X1 port map( A1 => A(27), A2 => n5, B1 => B(27), B2 => n9, ZN =>
                           n99);
   U59 : INV_X1 port map( A => n100, ZN => Z(28));
   U60 : AOI22_X1 port map( A1 => A(28), A2 => n5, B1 => B(28), B2 => n9, ZN =>
                           n100);
   U61 : INV_X1 port map( A => n101, ZN => Z(29));
   U62 : AOI22_X1 port map( A1 => A(29), A2 => n5, B1 => B(29), B2 => n9, ZN =>
                           n101);
   U63 : INV_X1 port map( A => n103, ZN => Z(30));
   U64 : AOI22_X1 port map( A1 => A(30), A2 => n5, B1 => B(30), B2 => n11, ZN 
                           => n103);
   U65 : INV_X1 port map( A => n91, ZN => Z(1));
   U66 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n11, ZN => 
                           n91);
   U67 : INV_X1 port map( A => n80, ZN => Z(0));
   U68 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => n14, ZN => 
                           n80);
   U69 : INV_X1 port map( A => n111, ZN => Z(9));
   U70 : AOI22_X1 port map( A1 => A(31), A2 => n6, B1 => B(31), B2 => n8, ZN =>
                           n104);
   U71 : AOI22_X1 port map( A1 => A(3), A2 => n6, B1 => B(3), B2 => n8, ZN => 
                           n105);
   U72 : AOI22_X1 port map( A1 => A(6), A2 => n6, B1 => B(6), B2 => n7, ZN => 
                           n108);
   U73 : AOI22_X1 port map( A1 => A(4), A2 => n6, B1 => B(4), B2 => n8, ZN => 
                           n106);
   U74 : AOI22_X1 port map( A1 => A(7), A2 => n6, B1 => B(7), B2 => n7, ZN => 
                           n109);
   U75 : AOI22_X1 port map( A1 => A(5), A2 => n6, B1 => B(5), B2 => n7, ZN => 
                           n107);
   U76 : AOI22_X1 port map( A1 => A(9), A2 => n6, B1 => n14, B2 => B(9), ZN => 
                           n111);
   U77 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => B(10), B2 => n14, ZN 
                           => n81);
   U78 : AOI22_X1 port map( A1 => A(8), A2 => n6, B1 => B(8), B2 => n7, ZN => 
                           n110);
   U79 : INV_X1 port map( A => n15, ZN => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_5;

architecture SYN_bhv of mux21_NBIT32_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => n4);
   U2 : INV_X1 port map( A => n14, ZN => n5);
   U3 : BUF_X1 port map( A => n1, Z => n6);
   U4 : BUF_X1 port map( A => n3, Z => n12);
   U5 : BUF_X1 port map( A => n2, Z => n11);
   U6 : BUF_X1 port map( A => n2, Z => n9);
   U7 : BUF_X1 port map( A => n3, Z => n14);
   U8 : BUF_X1 port map( A => n3, Z => n13);
   U9 : BUF_X1 port map( A => n1, Z => n7);
   U10 : BUF_X1 port map( A => n2, Z => n10);
   U11 : BUF_X1 port map( A => n1, Z => n8);
   U12 : BUF_X1 port map( A => S, Z => n3);
   U13 : BUF_X1 port map( A => S, Z => n1);
   U14 : BUF_X1 port map( A => S, Z => n2);
   U15 : INV_X1 port map( A => n98, ZN => Z(27));
   U16 : INV_X1 port map( A => n97, ZN => Z(26));
   U17 : INV_X1 port map( A => n100, ZN => Z(29));
   U18 : INV_X1 port map( A => n102, ZN => Z(30));
   U19 : INV_X1 port map( A => n103, ZN => Z(31));
   U20 : INV_X1 port map( A => n99, ZN => Z(28));
   U21 : INV_X1 port map( A => n90, ZN => Z(1));
   U22 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n10, ZN => 
                           n90);
   U23 : INV_X1 port map( A => n101, ZN => Z(2));
   U24 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           n101);
   U25 : INV_X1 port map( A => n104, ZN => Z(3));
   U26 : AOI22_X1 port map( A1 => A(3), A2 => n4, B1 => B(3), B2 => n7, ZN => 
                           n104);
   U27 : INV_X1 port map( A => n105, ZN => Z(4));
   U28 : AOI22_X1 port map( A1 => A(4), A2 => n5, B1 => B(4), B2 => n7, ZN => 
                           n105);
   U29 : INV_X1 port map( A => n106, ZN => Z(5));
   U30 : AOI22_X1 port map( A1 => A(5), A2 => n4, B1 => B(5), B2 => n6, ZN => 
                           n106);
   U31 : INV_X1 port map( A => n107, ZN => Z(6));
   U32 : AOI22_X1 port map( A1 => A(6), A2 => n5, B1 => B(6), B2 => n6, ZN => 
                           n107);
   U33 : INV_X1 port map( A => n108, ZN => Z(7));
   U34 : AOI22_X1 port map( A1 => A(7), A2 => n4, B1 => B(7), B2 => n6, ZN => 
                           n108);
   U35 : INV_X1 port map( A => n109, ZN => Z(8));
   U36 : AOI22_X1 port map( A1 => A(8), A2 => n5, B1 => B(8), B2 => n6, ZN => 
                           n109);
   U37 : INV_X1 port map( A => n80, ZN => Z(10));
   U38 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => B(10), B2 => n13, ZN 
                           => n80);
   U39 : INV_X1 port map( A => n81, ZN => Z(11));
   U40 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => B(11), B2 => n13, ZN 
                           => n81);
   U41 : INV_X1 port map( A => n82, ZN => Z(12));
   U42 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => B(12), B2 => n12, ZN 
                           => n82);
   U43 : INV_X1 port map( A => n83, ZN => Z(13));
   U44 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n12, ZN 
                           => n83);
   U45 : INV_X1 port map( A => n84, ZN => Z(14));
   U46 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n12, ZN 
                           => n84);
   U47 : INV_X1 port map( A => n85, ZN => Z(15));
   U48 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n12, ZN 
                           => n85);
   U49 : INV_X1 port map( A => n86, ZN => Z(16));
   U50 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => B(16), B2 => n11, ZN 
                           => n86);
   U51 : INV_X1 port map( A => n87, ZN => Z(17));
   U52 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n11, ZN 
                           => n87);
   U53 : INV_X1 port map( A => n88, ZN => Z(18));
   U54 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => B(18), B2 => n11, ZN 
                           => n88);
   U55 : INV_X1 port map( A => n89, ZN => Z(19));
   U56 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => B(19), B2 => n11, ZN 
                           => n89);
   U57 : INV_X1 port map( A => n91, ZN => Z(20));
   U58 : AOI22_X1 port map( A1 => A(20), A2 => n5, B1 => B(20), B2 => n10, ZN 
                           => n91);
   U59 : INV_X1 port map( A => n92, ZN => Z(21));
   U60 : AOI22_X1 port map( A1 => A(21), A2 => n5, B1 => B(21), B2 => n10, ZN 
                           => n92);
   U61 : INV_X1 port map( A => n93, ZN => Z(22));
   U62 : AOI22_X1 port map( A1 => A(22), A2 => n5, B1 => B(22), B2 => n9, ZN =>
                           n93);
   U63 : INV_X1 port map( A => n94, ZN => Z(23));
   U64 : AOI22_X1 port map( A1 => A(23), A2 => n5, B1 => B(23), B2 => n9, ZN =>
                           n94);
   U65 : INV_X1 port map( A => n95, ZN => Z(24));
   U66 : AOI22_X1 port map( A1 => A(24), A2 => n5, B1 => B(24), B2 => n9, ZN =>
                           n95);
   U67 : INV_X1 port map( A => n96, ZN => Z(25));
   U68 : AOI22_X1 port map( A1 => A(25), A2 => n5, B1 => B(25), B2 => n9, ZN =>
                           n96);
   U69 : INV_X1 port map( A => n110, ZN => Z(9));
   U70 : AOI22_X1 port map( A1 => A(9), A2 => n4, B1 => n13, B2 => B(9), ZN => 
                           n110);
   U71 : INV_X1 port map( A => n79, ZN => Z(0));
   U72 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => n13, ZN => 
                           n79);
   U73 : AOI22_X1 port map( A1 => A(29), A2 => n5, B1 => B(29), B2 => n8, ZN =>
                           n100);
   U74 : AOI22_X1 port map( A1 => A(26), A2 => n5, B1 => B(26), B2 => n8, ZN =>
                           n97);
   U75 : AOI22_X1 port map( A1 => A(30), A2 => n5, B1 => B(30), B2 => n10, ZN 
                           => n102);
   U76 : AOI22_X1 port map( A1 => A(27), A2 => n5, B1 => B(27), B2 => n8, ZN =>
                           n98);
   U77 : AOI22_X1 port map( A1 => A(28), A2 => n5, B1 => B(28), B2 => n8, ZN =>
                           n99);
   U78 : AOI22_X1 port map( A1 => A(31), A2 => n5, B1 => B(31), B2 => n7, ZN =>
                           n103);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_4;

architecture SYN_bhv of mux21_NBIT32_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n68, Z => n1);
   U2 : BUF_X1 port map( A => n68, Z => n2);
   U3 : BUF_X1 port map( A => n68, Z => n3);
   U4 : INV_X1 port map( A => n69, ZN => Z(0));
   U5 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => S, ZN => n69
                           );
   U6 : INV_X1 port map( A => n97, ZN => Z(6));
   U7 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => S, ZN => n97
                           );
   U8 : INV_X1 port map( A => n73, ZN => Z(13));
   U9 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => S, ZN => 
                           n73);
   U10 : INV_X1 port map( A => n77, ZN => Z(17));
   U11 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => S, ZN => 
                           n77);
   U12 : INV_X1 port map( A => n81, ZN => Z(20));
   U13 : AOI22_X1 port map( A1 => A(20), A2 => n2, B1 => B(20), B2 => S, ZN => 
                           n81);
   U14 : INV_X1 port map( A => n85, ZN => Z(24));
   U15 : AOI22_X1 port map( A1 => A(24), A2 => n2, B1 => B(24), B2 => S, ZN => 
                           n85);
   U16 : INV_X1 port map( A => n89, ZN => Z(28));
   U17 : AOI22_X1 port map( A1 => A(28), A2 => n2, B1 => B(28), B2 => S, ZN => 
                           n89);
   U18 : INV_X1 port map( A => n93, ZN => Z(31));
   U19 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => S, ZN => 
                           n93);
   U20 : INV_X1 port map( A => n94, ZN => Z(3));
   U21 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => S, ZN => 
                           n94);
   U22 : INV_X1 port map( A => n98, ZN => Z(7));
   U23 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => S, ZN => 
                           n98);
   U24 : INV_X1 port map( A => n70, ZN => Z(10));
   U25 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => S, ZN => 
                           n70);
   U26 : INV_X1 port map( A => n74, ZN => Z(14));
   U27 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => S, ZN => 
                           n74);
   U28 : INV_X1 port map( A => n78, ZN => Z(18));
   U29 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => S, ZN => 
                           n78);
   U30 : INV_X1 port map( A => n82, ZN => Z(21));
   U31 : AOI22_X1 port map( A1 => A(21), A2 => n2, B1 => B(21), B2 => S, ZN => 
                           n82);
   U32 : INV_X1 port map( A => n86, ZN => Z(25));
   U33 : AOI22_X1 port map( A1 => A(25), A2 => n2, B1 => B(25), B2 => S, ZN => 
                           n86);
   U34 : INV_X1 port map( A => n90, ZN => Z(29));
   U35 : AOI22_X1 port map( A1 => A(29), A2 => n2, B1 => B(29), B2 => S, ZN => 
                           n90);
   U36 : INV_X1 port map( A => n91, ZN => Z(2));
   U37 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => S, ZN => 
                           n91);
   U38 : INV_X1 port map( A => n95, ZN => Z(4));
   U39 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => S, ZN => 
                           n95);
   U40 : INV_X1 port map( A => n99, ZN => Z(8));
   U41 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => S, ZN => 
                           n99);
   U42 : INV_X1 port map( A => n71, ZN => Z(11));
   U43 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => S, ZN => 
                           n71);
   U44 : INV_X1 port map( A => n75, ZN => Z(15));
   U45 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => S, ZN => 
                           n75);
   U46 : INV_X1 port map( A => n79, ZN => Z(19));
   U47 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => S, ZN => 
                           n79);
   U48 : INV_X1 port map( A => n83, ZN => Z(22));
   U49 : AOI22_X1 port map( A1 => A(22), A2 => n2, B1 => B(22), B2 => S, ZN => 
                           n83);
   U50 : INV_X1 port map( A => n87, ZN => Z(26));
   U51 : AOI22_X1 port map( A1 => A(26), A2 => n2, B1 => B(26), B2 => S, ZN => 
                           n87);
   U52 : INV_X1 port map( A => n80, ZN => Z(1));
   U53 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => S, ZN => 
                           n80);
   U54 : INV_X1 port map( A => n96, ZN => Z(5));
   U55 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => S, ZN => 
                           n96);
   U56 : INV_X1 port map( A => n72, ZN => Z(12));
   U57 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => S, ZN => 
                           n72);
   U58 : INV_X1 port map( A => n76, ZN => Z(16));
   U59 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => S, ZN => 
                           n76);
   U60 : INV_X1 port map( A => n84, ZN => Z(23));
   U61 : AOI22_X1 port map( A1 => A(23), A2 => n2, B1 => B(23), B2 => S, ZN => 
                           n84);
   U62 : INV_X1 port map( A => n88, ZN => Z(27));
   U63 : AOI22_X1 port map( A1 => A(27), A2 => n2, B1 => B(27), B2 => S, ZN => 
                           n88);
   U64 : INV_X1 port map( A => n92, ZN => Z(30));
   U65 : AOI22_X1 port map( A1 => A(30), A2 => n2, B1 => B(30), B2 => S, ZN => 
                           n92);
   U66 : INV_X1 port map( A => n100, ZN => Z(9));
   U67 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => S, B2 => B(9), ZN => 
                           n100);
   U68 : INV_X1 port map( A => S, ZN => n68);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_3;

architecture SYN_bhv of mux21_NBIT32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n68, Z => n1);
   U2 : BUF_X1 port map( A => n68, Z => n2);
   U3 : BUF_X1 port map( A => n68, Z => n3);
   U4 : INV_X1 port map( A => n80, ZN => Z(1));
   U5 : AOI22_X1 port map( A1 => A(1), A2 => n1, B1 => B(1), B2 => S, ZN => n80
                           );
   U6 : INV_X1 port map( A => n69, ZN => Z(0));
   U7 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => S, ZN => n69
                           );
   U8 : INV_X1 port map( A => n94, ZN => Z(3));
   U9 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => S, ZN => n94
                           );
   U10 : INV_X1 port map( A => n81, ZN => Z(20));
   U11 : AOI22_X1 port map( A1 => A(20), A2 => n2, B1 => B(20), B2 => S, ZN => 
                           n81);
   U12 : INV_X1 port map( A => n82, ZN => Z(21));
   U13 : AOI22_X1 port map( A1 => A(21), A2 => n2, B1 => B(21), B2 => S, ZN => 
                           n82);
   U14 : INV_X1 port map( A => n83, ZN => Z(22));
   U15 : AOI22_X1 port map( A1 => A(22), A2 => n2, B1 => B(22), B2 => S, ZN => 
                           n83);
   U16 : INV_X1 port map( A => n84, ZN => Z(23));
   U17 : AOI22_X1 port map( A1 => A(23), A2 => n2, B1 => B(23), B2 => S, ZN => 
                           n84);
   U18 : INV_X1 port map( A => n77, ZN => Z(17));
   U19 : AOI22_X1 port map( A1 => A(17), A2 => n1, B1 => B(17), B2 => S, ZN => 
                           n77);
   U20 : INV_X1 port map( A => n78, ZN => Z(18));
   U21 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => S, ZN => 
                           n78);
   U22 : INV_X1 port map( A => n79, ZN => Z(19));
   U23 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => S, ZN => 
                           n79);
   U24 : INV_X1 port map( A => n73, ZN => Z(13));
   U25 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => S, ZN => 
                           n73);
   U26 : INV_X1 port map( A => n74, ZN => Z(14));
   U27 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => S, ZN => 
                           n74);
   U28 : INV_X1 port map( A => n75, ZN => Z(15));
   U29 : AOI22_X1 port map( A1 => A(15), A2 => n1, B1 => B(15), B2 => S, ZN => 
                           n75);
   U30 : INV_X1 port map( A => n76, ZN => Z(16));
   U31 : AOI22_X1 port map( A1 => A(16), A2 => n1, B1 => B(16), B2 => S, ZN => 
                           n76);
   U32 : INV_X1 port map( A => n70, ZN => Z(10));
   U33 : AOI22_X1 port map( A1 => A(10), A2 => n1, B1 => B(10), B2 => S, ZN => 
                           n70);
   U34 : INV_X1 port map( A => n71, ZN => Z(11));
   U35 : AOI22_X1 port map( A1 => A(11), A2 => n1, B1 => B(11), B2 => S, ZN => 
                           n71);
   U36 : INV_X1 port map( A => n72, ZN => Z(12));
   U37 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => S, ZN => 
                           n72);
   U38 : INV_X1 port map( A => n97, ZN => Z(6));
   U39 : AOI22_X1 port map( A1 => A(6), A2 => n3, B1 => B(6), B2 => S, ZN => 
                           n97);
   U40 : INV_X1 port map( A => n98, ZN => Z(7));
   U41 : AOI22_X1 port map( A1 => A(7), A2 => n3, B1 => B(7), B2 => S, ZN => 
                           n98);
   U42 : INV_X1 port map( A => n99, ZN => Z(8));
   U43 : AOI22_X1 port map( A1 => A(8), A2 => n3, B1 => B(8), B2 => S, ZN => 
                           n99);
   U44 : INV_X1 port map( A => n95, ZN => Z(4));
   U45 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => B(4), B2 => S, ZN => 
                           n95);
   U46 : INV_X1 port map( A => n96, ZN => Z(5));
   U47 : AOI22_X1 port map( A1 => A(5), A2 => n3, B1 => B(5), B2 => S, ZN => 
                           n96);
   U48 : INV_X1 port map( A => n89, ZN => Z(28));
   U49 : AOI22_X1 port map( A1 => A(28), A2 => n2, B1 => B(28), B2 => S, ZN => 
                           n89);
   U50 : INV_X1 port map( A => n90, ZN => Z(29));
   U51 : AOI22_X1 port map( A1 => A(29), A2 => n2, B1 => B(29), B2 => S, ZN => 
                           n90);
   U52 : INV_X1 port map( A => n91, ZN => Z(2));
   U53 : AOI22_X1 port map( A1 => A(2), A2 => n2, B1 => B(2), B2 => S, ZN => 
                           n91);
   U54 : INV_X1 port map( A => n92, ZN => Z(30));
   U55 : AOI22_X1 port map( A1 => A(30), A2 => n2, B1 => B(30), B2 => S, ZN => 
                           n92);
   U56 : INV_X1 port map( A => n85, ZN => Z(24));
   U57 : AOI22_X1 port map( A1 => A(24), A2 => n2, B1 => B(24), B2 => S, ZN => 
                           n85);
   U58 : INV_X1 port map( A => n86, ZN => Z(25));
   U59 : AOI22_X1 port map( A1 => A(25), A2 => n2, B1 => B(25), B2 => S, ZN => 
                           n86);
   U60 : INV_X1 port map( A => n87, ZN => Z(26));
   U61 : AOI22_X1 port map( A1 => A(26), A2 => n2, B1 => B(26), B2 => S, ZN => 
                           n87);
   U62 : INV_X1 port map( A => n88, ZN => Z(27));
   U63 : AOI22_X1 port map( A1 => A(27), A2 => n2, B1 => B(27), B2 => S, ZN => 
                           n88);
   U64 : INV_X1 port map( A => n93, ZN => Z(31));
   U65 : AOI22_X1 port map( A1 => A(31), A2 => n3, B1 => B(31), B2 => S, ZN => 
                           n93);
   U66 : INV_X1 port map( A => n100, ZN => Z(9));
   U67 : AOI22_X1 port map( A1 => A(9), A2 => n3, B1 => S, B2 => B(9), ZN => 
                           n100);
   U68 : INV_X1 port map( A => S, ZN => n68);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_2;

architecture SYN_bhv of mux21_NBIT32_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => n4);
   U2 : INV_X1 port map( A => n14, ZN => n5);
   U3 : BUF_X1 port map( A => n1, Z => n6);
   U4 : BUF_X1 port map( A => n3, Z => n12);
   U5 : BUF_X1 port map( A => n2, Z => n11);
   U6 : BUF_X1 port map( A => n2, Z => n9);
   U7 : BUF_X1 port map( A => n1, Z => n8);
   U8 : BUF_X1 port map( A => n2, Z => n10);
   U9 : BUF_X1 port map( A => n1, Z => n7);
   U10 : BUF_X1 port map( A => n3, Z => n14);
   U11 : BUF_X1 port map( A => n3, Z => n13);
   U12 : INV_X1 port map( A => n103, ZN => Z(31));
   U13 : AOI22_X1 port map( A1 => A(31), A2 => n4, B1 => B(31), B2 => n7, ZN =>
                           n103);
   U14 : BUF_X1 port map( A => S, Z => n3);
   U15 : BUF_X1 port map( A => S, Z => n2);
   U16 : BUF_X1 port map( A => S, Z => n1);
   U17 : INV_X1 port map( A => n79, ZN => Z(0));
   U18 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => n13, ZN => 
                           n79);
   U19 : INV_X1 port map( A => n104, ZN => Z(3));
   U20 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => B(3), B2 => n7, ZN => 
                           n104);
   U21 : INV_X1 port map( A => n105, ZN => Z(4));
   U22 : AOI22_X1 port map( A1 => A(4), A2 => n4, B1 => B(4), B2 => n7, ZN => 
                           n105);
   U23 : INV_X1 port map( A => n106, ZN => Z(5));
   U24 : AOI22_X1 port map( A1 => A(5), A2 => n5, B1 => B(5), B2 => n6, ZN => 
                           n106);
   U25 : INV_X1 port map( A => n107, ZN => Z(6));
   U26 : AOI22_X1 port map( A1 => A(6), A2 => n4, B1 => B(6), B2 => n6, ZN => 
                           n107);
   U27 : INV_X1 port map( A => n108, ZN => Z(7));
   U28 : AOI22_X1 port map( A1 => A(7), A2 => n5, B1 => B(7), B2 => n6, ZN => 
                           n108);
   U29 : INV_X1 port map( A => n109, ZN => Z(8));
   U30 : AOI22_X1 port map( A1 => A(8), A2 => n4, B1 => B(8), B2 => n6, ZN => 
                           n109);
   U31 : INV_X1 port map( A => n110, ZN => Z(9));
   U32 : AOI22_X1 port map( A1 => A(9), A2 => n5, B1 => n13, B2 => B(9), ZN => 
                           n110);
   U33 : INV_X1 port map( A => n85, ZN => Z(15));
   U34 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n12, ZN 
                           => n85);
   U35 : INV_X1 port map( A => n86, ZN => Z(16));
   U36 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => B(16), B2 => n11, ZN 
                           => n86);
   U37 : INV_X1 port map( A => n87, ZN => Z(17));
   U38 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n11, ZN 
                           => n87);
   U39 : INV_X1 port map( A => n88, ZN => Z(18));
   U40 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => B(18), B2 => n11, ZN 
                           => n88);
   U41 : INV_X1 port map( A => n89, ZN => Z(19));
   U42 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => B(19), B2 => n11, ZN 
                           => n89);
   U43 : INV_X1 port map( A => n91, ZN => Z(20));
   U44 : AOI22_X1 port map( A1 => A(20), A2 => n5, B1 => B(20), B2 => n10, ZN 
                           => n91);
   U45 : INV_X1 port map( A => n92, ZN => Z(21));
   U46 : AOI22_X1 port map( A1 => A(21), A2 => n5, B1 => B(21), B2 => n10, ZN 
                           => n92);
   U47 : INV_X1 port map( A => n93, ZN => Z(22));
   U48 : AOI22_X1 port map( A1 => A(22), A2 => n5, B1 => B(22), B2 => n9, ZN =>
                           n93);
   U49 : INV_X1 port map( A => n94, ZN => Z(23));
   U50 : AOI22_X1 port map( A1 => A(23), A2 => n5, B1 => B(23), B2 => n9, ZN =>
                           n94);
   U51 : INV_X1 port map( A => n95, ZN => Z(24));
   U52 : AOI22_X1 port map( A1 => A(24), A2 => n5, B1 => B(24), B2 => n9, ZN =>
                           n95);
   U53 : INV_X1 port map( A => n96, ZN => Z(25));
   U54 : AOI22_X1 port map( A1 => A(25), A2 => n5, B1 => B(25), B2 => n9, ZN =>
                           n96);
   U55 : INV_X1 port map( A => n97, ZN => Z(26));
   U56 : AOI22_X1 port map( A1 => A(26), A2 => n5, B1 => B(26), B2 => n8, ZN =>
                           n97);
   U57 : INV_X1 port map( A => n98, ZN => Z(27));
   U58 : AOI22_X1 port map( A1 => A(27), A2 => n5, B1 => B(27), B2 => n8, ZN =>
                           n98);
   U59 : INV_X1 port map( A => n99, ZN => Z(28));
   U60 : AOI22_X1 port map( A1 => A(28), A2 => n5, B1 => B(28), B2 => n8, ZN =>
                           n99);
   U61 : INV_X1 port map( A => n100, ZN => Z(29));
   U62 : AOI22_X1 port map( A1 => A(29), A2 => n5, B1 => B(29), B2 => n8, ZN =>
                           n100);
   U63 : INV_X1 port map( A => n102, ZN => Z(30));
   U64 : AOI22_X1 port map( A1 => A(30), A2 => n5, B1 => B(30), B2 => n10, ZN 
                           => n102);
   U65 : INV_X1 port map( A => n84, ZN => Z(14));
   U66 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n12, ZN 
                           => n84);
   U67 : INV_X1 port map( A => n90, ZN => Z(1));
   U68 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n10, ZN => 
                           n90);
   U69 : INV_X1 port map( A => n101, ZN => Z(2));
   U70 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           n101);
   U71 : INV_X1 port map( A => n80, ZN => Z(10));
   U72 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => B(10), B2 => n13, ZN 
                           => n80);
   U73 : INV_X1 port map( A => n81, ZN => Z(11));
   U74 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => B(11), B2 => n13, ZN 
                           => n81);
   U75 : INV_X1 port map( A => n82, ZN => Z(12));
   U76 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => B(12), B2 => n12, ZN 
                           => n82);
   U77 : INV_X1 port map( A => n83, ZN => Z(13));
   U78 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n12, ZN 
                           => n83);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_1;

architecture SYN_bhv of mux21_NBIT32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => n4);
   U2 : INV_X1 port map( A => n14, ZN => n5);
   U3 : BUF_X1 port map( A => n1, Z => n6);
   U4 : BUF_X1 port map( A => n3, Z => n12);
   U5 : BUF_X1 port map( A => n2, Z => n11);
   U6 : BUF_X1 port map( A => n2, Z => n9);
   U7 : BUF_X1 port map( A => n1, Z => n8);
   U8 : BUF_X1 port map( A => n2, Z => n10);
   U9 : BUF_X1 port map( A => n1, Z => n7);
   U10 : BUF_X1 port map( A => n3, Z => n14);
   U11 : BUF_X1 port map( A => n3, Z => n13);
   U12 : BUF_X1 port map( A => S, Z => n3);
   U13 : BUF_X1 port map( A => S, Z => n2);
   U14 : BUF_X1 port map( A => S, Z => n1);
   U15 : INV_X1 port map( A => n79, ZN => Z(0));
   U16 : AOI22_X1 port map( A1 => A(0), A2 => n4, B1 => B(0), B2 => n13, ZN => 
                           n79);
   U17 : INV_X1 port map( A => n90, ZN => Z(1));
   U18 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n10, ZN => 
                           n90);
   U19 : INV_X1 port map( A => n101, ZN => Z(2));
   U20 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => n7, ZN => 
                           n101);
   U21 : INV_X1 port map( A => n104, ZN => Z(3));
   U22 : AOI22_X1 port map( A1 => A(3), A2 => n4, B1 => B(3), B2 => n7, ZN => 
                           n104);
   U23 : INV_X1 port map( A => n105, ZN => Z(4));
   U24 : AOI22_X1 port map( A1 => A(4), A2 => n5, B1 => B(4), B2 => n7, ZN => 
                           n105);
   U25 : INV_X1 port map( A => n106, ZN => Z(5));
   U26 : AOI22_X1 port map( A1 => A(5), A2 => n4, B1 => B(5), B2 => n6, ZN => 
                           n106);
   U27 : INV_X1 port map( A => n107, ZN => Z(6));
   U28 : AOI22_X1 port map( A1 => A(6), A2 => n5, B1 => B(6), B2 => n6, ZN => 
                           n107);
   U29 : INV_X1 port map( A => n108, ZN => Z(7));
   U30 : AOI22_X1 port map( A1 => A(7), A2 => n4, B1 => B(7), B2 => n6, ZN => 
                           n108);
   U31 : INV_X1 port map( A => n109, ZN => Z(8));
   U32 : AOI22_X1 port map( A1 => A(8), A2 => n5, B1 => B(8), B2 => n6, ZN => 
                           n109);
   U33 : INV_X1 port map( A => n110, ZN => Z(9));
   U34 : AOI22_X1 port map( A1 => A(9), A2 => n4, B1 => n13, B2 => B(9), ZN => 
                           n110);
   U35 : INV_X1 port map( A => n80, ZN => Z(10));
   U36 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => B(10), B2 => n13, ZN 
                           => n80);
   U37 : INV_X1 port map( A => n81, ZN => Z(11));
   U38 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => B(11), B2 => n13, ZN 
                           => n81);
   U39 : INV_X1 port map( A => n82, ZN => Z(12));
   U40 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => B(12), B2 => n12, ZN 
                           => n82);
   U41 : INV_X1 port map( A => n83, ZN => Z(13));
   U42 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n12, ZN 
                           => n83);
   U43 : INV_X1 port map( A => n84, ZN => Z(14));
   U44 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n12, ZN 
                           => n84);
   U45 : INV_X1 port map( A => n85, ZN => Z(15));
   U46 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n12, ZN 
                           => n85);
   U47 : INV_X1 port map( A => n86, ZN => Z(16));
   U48 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => B(16), B2 => n11, ZN 
                           => n86);
   U49 : INV_X1 port map( A => n87, ZN => Z(17));
   U50 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => B(17), B2 => n11, ZN 
                           => n87);
   U51 : INV_X1 port map( A => n88, ZN => Z(18));
   U52 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => B(18), B2 => n11, ZN 
                           => n88);
   U53 : INV_X1 port map( A => n89, ZN => Z(19));
   U54 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => B(19), B2 => n11, ZN 
                           => n89);
   U55 : INV_X1 port map( A => n91, ZN => Z(20));
   U56 : AOI22_X1 port map( A1 => A(20), A2 => n5, B1 => B(20), B2 => n10, ZN 
                           => n91);
   U57 : INV_X1 port map( A => n92, ZN => Z(21));
   U58 : AOI22_X1 port map( A1 => A(21), A2 => n5, B1 => B(21), B2 => n10, ZN 
                           => n92);
   U59 : INV_X1 port map( A => n93, ZN => Z(22));
   U60 : AOI22_X1 port map( A1 => A(22), A2 => n5, B1 => B(22), B2 => n9, ZN =>
                           n93);
   U61 : INV_X1 port map( A => n94, ZN => Z(23));
   U62 : AOI22_X1 port map( A1 => A(23), A2 => n5, B1 => B(23), B2 => n9, ZN =>
                           n94);
   U63 : INV_X1 port map( A => n95, ZN => Z(24));
   U64 : AOI22_X1 port map( A1 => A(24), A2 => n5, B1 => B(24), B2 => n9, ZN =>
                           n95);
   U65 : INV_X1 port map( A => n96, ZN => Z(25));
   U66 : AOI22_X1 port map( A1 => A(25), A2 => n5, B1 => B(25), B2 => n9, ZN =>
                           n96);
   U67 : INV_X1 port map( A => n97, ZN => Z(26));
   U68 : AOI22_X1 port map( A1 => A(26), A2 => n5, B1 => B(26), B2 => n8, ZN =>
                           n97);
   U69 : INV_X1 port map( A => n98, ZN => Z(27));
   U70 : AOI22_X1 port map( A1 => A(27), A2 => n5, B1 => B(27), B2 => n8, ZN =>
                           n98);
   U71 : INV_X1 port map( A => n99, ZN => Z(28));
   U72 : AOI22_X1 port map( A1 => A(28), A2 => n5, B1 => B(28), B2 => n8, ZN =>
                           n99);
   U73 : INV_X1 port map( A => n100, ZN => Z(29));
   U74 : AOI22_X1 port map( A1 => A(29), A2 => n5, B1 => B(29), B2 => n8, ZN =>
                           n100);
   U75 : INV_X1 port map( A => n102, ZN => Z(30));
   U76 : AOI22_X1 port map( A1 => A(30), A2 => n5, B1 => B(30), B2 => n10, ZN 
                           => n102);
   U77 : INV_X1 port map( A => n103, ZN => Z(31));
   U78 : AOI22_X1 port map( A1 => A(31), A2 => n5, B1 => B(31), B2 => n7, ZN =>
                           n103);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ff_2 is

   port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);

end ff_2;

architecture SYN_bhv of ff_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CLK, RN => RST, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => EN, A => n6, ZN => n4);
   U3 : NAND2_X1 port map( A1 => EN, A2 => D, ZN => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ff_1 is

   port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);

end ff_1;

architecture SYN_bhv of ff_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CLK, RN => RST, Q => Q, QN => n5);
   U2 : OAI21_X1 port map( B1 => n5, B2 => EN, A => n6, ZN => n4);
   U3 : NAND2_X1 port map( A1 => EN, A2 => D, ZN => n6);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity RCA_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_0;

architecture SYN_STRUCTURAL of RCA_N4_0 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_select_basic_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_basic_N4_0;

architecture SYN_struct of carry_select_basic_N4_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, Y1_3_port, Y1_2_port, Y1_1_port, 
      Y1_0_port, Y2_3_port, Y2_2_port, Y2_1_port, Y2_0_port, n6, n7, n8, n9, n5
      , n_1155, n_1156 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => Y1_3_port, 
                           S(2) => Y1_2_port, S(1) => Y1_1_port, S(0) => 
                           Y1_0_port, Co => n_1155);
   RCA1 : RCA_N4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => Y2_3_port, 
                           S(2) => Y2_2_port, S(1) => Y2_1_port, S(0) => 
                           Y2_0_port, Co => n_1156);
   U3 : INV_X1 port map( A => C_i, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => S(3));
   U5 : AOI22_X1 port map( A1 => Y1_3_port, A2 => n5, B1 => Y2_3_port, B2 => 
                           C_i, ZN => n6);
   U6 : INV_X1 port map( A => n8, ZN => S(1));
   U7 : AOI22_X1 port map( A1 => Y1_1_port, A2 => n5, B1 => Y2_1_port, B2 => 
                           C_i, ZN => n8);
   U8 : INV_X1 port map( A => n7, ZN => S(2));
   U9 : AOI22_X1 port map( A1 => Y1_2_port, A2 => n5, B1 => Y2_2_port, B2 => 
                           C_i, ZN => n7);
   U10 : INV_X1 port map( A => n9, ZN => S(0));
   U11 : AOI22_X1 port map( A1 => Y1_0_port, A2 => n5, B1 => Y2_0_port, B2 => 
                           C_i, ZN => n9);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PGblock_0 is

   port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);

end PGblock_0;

architecture SYN_bhv of PGblock_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Gk_1j, B2 => Pik, A => Gik, ZN => n2);
   U3 : AND2_X1 port map( A1 => Pk_1j, A2 => Pik, ZN => Pij);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Gblock_0 is

   port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);

end Gblock_0;

architecture SYN_bhv of Gblock_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gk_1j, A => Gik, ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity PG_net_0 is

   port( a, b : in std_logic;  p, g : out std_logic);

end PG_net_0;

architecture SYN_bhv of PG_net_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity rca_bhv_numBit32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end rca_bhv_numBit32_0;

architecture SYN_BEHAVIORAL of rca_bhv_numBit32_0 is

   component rca_bhv_numBit32_0_DW01_add_0
      port( A, B : in std_logic_vector (32 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (32 downto 0);  CO : out std_logic);
   end component;
   
   signal n_1157 : std_logic;

begin
   
   add_1_root_add_35_2 : rca_bhv_numBit32_0_DW01_add_0 port map( A(32) => A(31)
                           , A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(32) => Co, SUM(31)
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1157);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux5to1_numBit32_0 is

   port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  SEL_in :
         in std_logic_vector (2 downto 0);  Z : out std_logic_vector (31 downto
         0));

end mux5to1_numBit32_0;

architecture SYN_bhv of mux5to1_numBit32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n1, n2
      , n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91 : std_logic;

begin
   
   U109 : OAI33_X1 port map( A1 => n91, A2 => SEL_in(2), A3 => SEL_in(1), B1 =>
                           n90, B2 => SEL_in(2), B3 => SEL_in(0), ZN => n8);
   U2 : BUF_X1 port map( A => n10, Z => n4);
   U3 : BUF_X1 port map( A => n10, Z => n77);
   U4 : BUF_X1 port map( A => n10, Z => n78);
   U5 : INV_X1 port map( A => SEL_in(1), ZN => n90);
   U6 : AOI222_X1 port map( A1 => IN4(2), A2 => n85, B1 => IN2(2), B2 => n82, 
                           C1 => IN5(2), C2 => n79, ZN => n68);
   U7 : AOI222_X1 port map( A1 => IN4(3), A2 => n85, B1 => IN2(3), B2 => n82, 
                           C1 => IN5(3), C2 => n79, ZN => n66);
   U8 : AOI222_X1 port map( A1 => IN4(4), A2 => n85, B1 => IN2(4), B2 => n82, 
                           C1 => IN5(4), C2 => n79, ZN => n64);
   U9 : AOI222_X1 port map( A1 => IN4(5), A2 => n85, B1 => IN2(5), B2 => n82, 
                           C1 => IN5(5), C2 => n79, ZN => n62);
   U10 : AOI222_X1 port map( A1 => IN4(6), A2 => n85, B1 => IN2(6), B2 => n82, 
                           C1 => IN5(6), C2 => n79, ZN => n60);
   U11 : AOI222_X1 port map( A1 => IN4(7), A2 => n85, B1 => IN2(7), B2 => n82, 
                           C1 => IN5(7), C2 => n79, ZN => n58);
   U12 : AOI222_X1 port map( A1 => IN4(8), A2 => n85, B1 => IN2(8), B2 => n82, 
                           C1 => IN5(8), C2 => n79, ZN => n56);
   U13 : AOI222_X1 port map( A1 => IN4(9), A2 => n85, B1 => IN2(9), B2 => n82, 
                           C1 => IN5(9), C2 => n79, ZN => n54);
   U14 : AOI222_X1 port map( A1 => IN4(10), A2 => n85, B1 => IN2(10), B2 => n82
                           , C1 => IN5(10), C2 => n79, ZN => n52);
   U15 : AOI222_X1 port map( A1 => IN4(11), A2 => n85, B1 => IN2(11), B2 => n82
                           , C1 => IN5(11), C2 => n79, ZN => n50);
   U16 : AOI222_X1 port map( A1 => IN4(12), A2 => n86, B1 => IN2(12), B2 => n83
                           , C1 => IN5(12), C2 => n80, ZN => n48);
   U17 : AOI222_X1 port map( A1 => IN4(13), A2 => n86, B1 => IN2(13), B2 => n83
                           , C1 => IN5(13), C2 => n80, ZN => n46);
   U18 : AOI222_X1 port map( A1 => IN4(14), A2 => n86, B1 => IN2(14), B2 => n83
                           , C1 => IN5(14), C2 => n80, ZN => n44);
   U19 : AOI222_X1 port map( A1 => IN4(15), A2 => n86, B1 => IN2(15), B2 => n83
                           , C1 => IN5(15), C2 => n80, ZN => n42);
   U20 : AOI222_X1 port map( A1 => IN4(25), A2 => n87, B1 => IN2(25), B2 => n84
                           , C1 => IN5(25), C2 => n81, ZN => n22);
   U21 : AOI222_X1 port map( A1 => IN4(26), A2 => n87, B1 => IN2(26), B2 => n84
                           , C1 => IN5(26), C2 => n81, ZN => n20);
   U22 : AOI222_X1 port map( A1 => IN4(27), A2 => n87, B1 => IN2(27), B2 => n84
                           , C1 => IN5(27), C2 => n81, ZN => n18);
   U23 : AOI222_X1 port map( A1 => IN4(28), A2 => n87, B1 => IN2(28), B2 => n84
                           , C1 => IN5(28), C2 => n81, ZN => n16);
   U24 : AOI222_X1 port map( A1 => IN4(29), A2 => n87, B1 => IN2(29), B2 => n84
                           , C1 => IN5(29), C2 => n81, ZN => n14);
   U25 : AOI222_X1 port map( A1 => IN4(30), A2 => n87, B1 => IN2(30), B2 => n84
                           , C1 => IN5(30), C2 => n81, ZN => n12);
   U26 : AOI222_X1 port map( A1 => IN4(1), A2 => n85, B1 => IN2(1), B2 => n82, 
                           C1 => IN5(1), C2 => n79, ZN => n70);
   U27 : AOI222_X1 port map( A1 => IN4(16), A2 => n86, B1 => IN2(16), B2 => n83
                           , C1 => IN5(16), C2 => n80, ZN => n40);
   U28 : AOI222_X1 port map( A1 => IN4(17), A2 => n86, B1 => IN2(17), B2 => n83
                           , C1 => IN5(17), C2 => n80, ZN => n38);
   U29 : AOI222_X1 port map( A1 => IN4(18), A2 => n86, B1 => IN2(18), B2 => n83
                           , C1 => IN5(18), C2 => n80, ZN => n36);
   U30 : AOI222_X1 port map( A1 => IN4(19), A2 => n86, B1 => IN2(19), B2 => n83
                           , C1 => IN5(19), C2 => n80, ZN => n34);
   U31 : AOI222_X1 port map( A1 => IN4(20), A2 => n86, B1 => IN2(20), B2 => n83
                           , C1 => IN5(20), C2 => n80, ZN => n32);
   U32 : AOI222_X1 port map( A1 => IN4(21), A2 => n86, B1 => IN2(21), B2 => n83
                           , C1 => IN5(21), C2 => n80, ZN => n30);
   U33 : AOI222_X1 port map( A1 => IN4(22), A2 => n86, B1 => IN2(22), B2 => n83
                           , C1 => IN5(22), C2 => n80, ZN => n28);
   U34 : AOI222_X1 port map( A1 => IN4(23), A2 => n86, B1 => IN2(23), B2 => n83
                           , C1 => IN5(23), C2 => n80, ZN => n26);
   U35 : AOI222_X1 port map( A1 => IN4(24), A2 => n86, B1 => IN2(24), B2 => n83
                           , C1 => IN5(24), C2 => n80, ZN => n24);
   U36 : BUF_X1 port map( A => n9, Z => n79);
   U37 : BUF_X1 port map( A => n9, Z => n80);
   U38 : BUF_X1 port map( A => n7, Z => n85);
   U39 : BUF_X1 port map( A => n7, Z => n86);
   U40 : BUF_X1 port map( A => n89, Z => n1);
   U41 : BUF_X1 port map( A => n89, Z => n2);
   U42 : NOR2_X1 port map( A1 => n88, A2 => n75, ZN => n10);
   U43 : INV_X1 port map( A => n74, ZN => n88);
   U44 : BUF_X1 port map( A => n89, Z => n3);
   U45 : BUF_X1 port map( A => n9, Z => n81);
   U46 : BUF_X1 port map( A => n7, Z => n87);
   U47 : NOR4_X1 port map( A1 => n76, A2 => n85, A3 => n79, A4 => n82, ZN => 
                           n74);
   U48 : NOR3_X1 port map( A1 => n90, A2 => SEL_in(2), A3 => n91, ZN => n7);
   U49 : BUF_X1 port map( A => n8, Z => n82);
   U50 : BUF_X1 port map( A => n8, Z => n83);
   U51 : BUF_X1 port map( A => n8, Z => n84);
   U52 : NOR2_X1 port map( A1 => n90, A2 => n91, ZN => n75);
   U53 : AND3_X1 port map( A1 => n91, A2 => n90, A3 => SEL_in(2), ZN => n9);
   U54 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => Z(3));
   U55 : INV_X1 port map( A => n73, ZN => n89);
   U56 : AOI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => n73);
   U57 : AOI22_X1 port map( A1 => IN3(1), A2 => n4, B1 => IN1(1), B2 => n1, ZN 
                           => n69);
   U58 : AOI22_X1 port map( A1 => IN3(2), A2 => n4, B1 => IN1(2), B2 => n1, ZN 
                           => n67);
   U59 : AOI22_X1 port map( A1 => IN3(3), A2 => n4, B1 => IN1(3), B2 => n1, ZN 
                           => n65);
   U60 : AOI22_X1 port map( A1 => IN3(4), A2 => n4, B1 => IN1(4), B2 => n1, ZN 
                           => n63);
   U61 : AOI22_X1 port map( A1 => IN3(5), A2 => n4, B1 => IN1(5), B2 => n1, ZN 
                           => n61);
   U62 : AOI22_X1 port map( A1 => IN3(6), A2 => n4, B1 => IN1(6), B2 => n1, ZN 
                           => n59);
   U63 : AOI22_X1 port map( A1 => IN3(7), A2 => n4, B1 => IN1(7), B2 => n1, ZN 
                           => n57);
   U64 : AOI22_X1 port map( A1 => IN3(8), A2 => n4, B1 => IN1(8), B2 => n1, ZN 
                           => n55);
   U65 : AOI22_X1 port map( A1 => IN3(9), A2 => n4, B1 => IN1(9), B2 => n1, ZN 
                           => n53);
   U66 : AOI22_X1 port map( A1 => IN3(10), A2 => n4, B1 => IN1(10), B2 => n1, 
                           ZN => n51);
   U67 : AOI22_X1 port map( A1 => IN3(11), A2 => n4, B1 => IN1(11), B2 => n1, 
                           ZN => n49);
   U68 : AOI22_X1 port map( A1 => IN3(12), A2 => n77, B1 => IN1(12), B2 => n2, 
                           ZN => n47);
   U69 : AOI22_X1 port map( A1 => IN3(13), A2 => n77, B1 => IN1(13), B2 => n2, 
                           ZN => n45);
   U70 : AOI22_X1 port map( A1 => IN3(14), A2 => n77, B1 => IN1(14), B2 => n2, 
                           ZN => n43);
   U71 : NOR3_X1 port map( A1 => SEL_in(1), A2 => SEL_in(2), A3 => SEL_in(0), 
                           ZN => n76);
   U72 : AOI222_X1 port map( A1 => IN4(0), A2 => n85, B1 => IN2(0), B2 => n82, 
                           C1 => IN5(0), C2 => n79, ZN => n72);
   U73 : AOI22_X1 port map( A1 => IN3(15), A2 => n77, B1 => IN1(15), B2 => n2, 
                           ZN => n41);
   U74 : AOI22_X1 port map( A1 => IN3(24), A2 => n78, B1 => IN1(24), B2 => n3, 
                           ZN => n23);
   U75 : AOI22_X1 port map( A1 => IN3(25), A2 => n78, B1 => IN1(25), B2 => n3, 
                           ZN => n21);
   U76 : AOI22_X1 port map( A1 => IN3(26), A2 => n78, B1 => IN1(26), B2 => n3, 
                           ZN => n19);
   U77 : AOI22_X1 port map( A1 => IN3(27), A2 => n78, B1 => IN1(27), B2 => n3, 
                           ZN => n17);
   U78 : AOI22_X1 port map( A1 => IN3(28), A2 => n78, B1 => IN1(28), B2 => n3, 
                           ZN => n15);
   U79 : AOI22_X1 port map( A1 => IN3(29), A2 => n78, B1 => IN1(29), B2 => n3, 
                           ZN => n13);
   U80 : AOI22_X1 port map( A1 => IN3(30), A2 => n78, B1 => IN1(30), B2 => n3, 
                           ZN => n11);
   U81 : AOI22_X1 port map( A1 => IN3(0), A2 => n4, B1 => IN1(0), B2 => n1, ZN 
                           => n71);
   U82 : AOI22_X1 port map( A1 => IN3(19), A2 => n77, B1 => IN1(19), B2 => n2, 
                           ZN => n33);
   U83 : AOI22_X1 port map( A1 => IN3(20), A2 => n77, B1 => IN1(20), B2 => n2, 
                           ZN => n31);
   U84 : AOI22_X1 port map( A1 => IN3(21), A2 => n77, B1 => IN1(21), B2 => n2, 
                           ZN => n29);
   U85 : AOI22_X1 port map( A1 => IN3(22), A2 => n77, B1 => IN1(22), B2 => n2, 
                           ZN => n27);
   U86 : AOI22_X1 port map( A1 => IN3(23), A2 => n77, B1 => IN1(23), B2 => n2, 
                           ZN => n25);
   U87 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => Z(4));
   U88 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => Z(5));
   U89 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => Z(6));
   U90 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => Z(7));
   U91 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => Z(8));
   U92 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => Z(9));
   U93 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => Z(10));
   U94 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => Z(11));
   U95 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => Z(12));
   U96 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => Z(13));
   U97 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => Z(14));
   U98 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => Z(15));
   U99 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => Z(16));
   U100 : AOI22_X1 port map( A1 => IN3(16), A2 => n77, B1 => IN1(16), B2 => n2,
                           ZN => n39);
   U101 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => Z(17));
   U102 : AOI22_X1 port map( A1 => IN3(17), A2 => n77, B1 => IN1(17), B2 => n2,
                           ZN => n37);
   U103 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => Z(18));
   U104 : AOI22_X1 port map( A1 => IN3(18), A2 => n77, B1 => IN1(18), B2 => n2,
                           ZN => n35);
   U105 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => Z(19));
   U106 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => Z(20));
   U107 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => Z(21));
   U108 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => Z(22));
   U110 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => Z(23));
   U111 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => Z(24));
   U112 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => Z(25));
   U113 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => Z(26));
   U114 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => Z(27));
   U115 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => Z(28));
   U116 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => Z(29));
   U117 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => Z(30));
   U118 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => Z(2));
   U119 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => Z(0));
   U120 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => Z(1));
   U121 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Z(31));
   U122 : AOI22_X1 port map( A1 => IN3(31), A2 => n78, B1 => IN1(31), B2 => n3,
                           ZN => n5);
   U123 : AOI222_X1 port map( A1 => IN4(31), A2 => n87, B1 => IN2(31), B2 => 
                           n84, C1 => IN5(31), C2 => n81, ZN => n6);
   U124 : INV_X1 port map( A => SEL_in(0), ZN => n91);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity booth_encoder_numBit16 is

   port( B : in std_logic_vector (15 downto 0);  SEL_out : out std_logic_vector
         (23 downto 0));

end booth_encoder_numBit16;

architecture SYN_structural of booth_encoder_numBit16 is

signal X_Logic0_port : std_logic;

begin
   SEL_out <= ( B(15), B(14), B(13), B(13), B(12), B(11), B(11), B(10), B(9), 
      B(9), B(8), B(7), B(7), B(6), B(5), B(5), B(4), B(3), B(3), B(2), B(1), 
      B(1), B(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8;

architecture SYN_structural of SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   component carry_select_basic_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_basic_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  C_i : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CSBI_1 : carry_select_basic_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) 
                           => A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), 
                           B(1) => B(1), B(0) => B(0), C_i => Ci(0), S(3) => 
                           S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CSBI_2 : carry_select_basic_N4_7 port map( A(3) => A(7), A(2) => A(6), A(1) 
                           => A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), 
                           B(1) => B(5), B(0) => B(4), C_i => Ci(1), S(3) => 
                           S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   CSBI_3 : carry_select_basic_N4_6 port map( A(3) => A(11), A(2) => A(10), 
                           A(1) => A(9), A(0) => A(8), B(3) => B(11), B(2) => 
                           B(10), B(1) => B(9), B(0) => B(8), C_i => Ci(2), 
                           S(3) => S(11), S(2) => S(10), S(1) => S(9), S(0) => 
                           S(8));
   CSBI_4 : carry_select_basic_N4_5 port map( A(3) => A(15), A(2) => A(14), 
                           A(1) => A(13), A(0) => A(12), B(3) => B(15), B(2) =>
                           B(14), B(1) => B(13), B(0) => B(12), C_i => Ci(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   CSBI_5 : carry_select_basic_N4_4 port map( A(3) => A(19), A(2) => A(18), 
                           A(1) => A(17), A(0) => A(16), B(3) => B(19), B(2) =>
                           B(18), B(1) => B(17), B(0) => B(16), C_i => Ci(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   CSBI_6 : carry_select_basic_N4_3 port map( A(3) => A(23), A(2) => A(22), 
                           A(1) => A(21), A(0) => A(20), B(3) => B(23), B(2) =>
                           B(22), B(1) => B(21), B(0) => B(20), C_i => Ci(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   CSBI_7 : carry_select_basic_N4_2 port map( A(3) => A(27), A(2) => A(26), 
                           A(1) => A(25), A(0) => A(24), B(3) => B(27), B(2) =>
                           B(26), B(1) => B(25), B(0) => B(24), C_i => Ci(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   CSBI_8 : carry_select_basic_N4_1 port map( A(3) => A(31), A(2) => A(30), 
                           A(1) => A(29), A(0) => A(28), B(3) => B(31), B(2) =>
                           B(30), B(1) => B(29), B(0) => B(28), C_i => Ci(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity carry_generator_NBIT32_NBIT_PER_BLOCK4 is

   port( A, B : in std_logic_vector (32 downto 1);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end carry_generator_NBIT32_NBIT_PER_BLOCK4;

architecture SYN_struct of carry_generator_NBIT32_NBIT_PER_BLOCK4 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component PGblock_1
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_2
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_3
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_4
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_5
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_6
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_7
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_8
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_9
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_10
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_11
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_12
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_13
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_14
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_15
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_16
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_17
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_18
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_19
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_20
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_21
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_22
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_23
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_24
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_25
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_26
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PGblock_0
      port( Pik, Gik, Pk_1j, Gk_1j : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component Gblock_1
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_2
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_3
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_4
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_5
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_6
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_7
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_8
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component Gblock_0
      port( Pik, Gik, Gk_1j : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_net_1
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_2
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_3
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_4
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_5
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_6
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_7
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_8
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_9
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_10
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_11
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_12
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_13
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_14
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_15
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_16
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_17
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_18
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_19
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_20
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_21
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_22
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_23
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_24
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_25
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_26
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_27
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_28
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_29
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_30
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component PG_net_0
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   signal Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port, G_16_16_port, G_16_15_port, G_16_13_port, 
      G_16_9_port, G_15_15_port, G_14_14_port, G_14_13_port, G_13_13_port, 
      G_12_12_port, G_12_11_port, G_12_9_port, G_11_11_port, G_10_10_port, 
      G_10_9_port, G_9_9_port, G_8_8_port, G_8_7_port, G_8_5_port, G_7_7_port, 
      G_6_6_port, G_6_5_port, G_5_5_port, G_4_4_port, G_4_3_port, G_3_3_port, 
      G_2_2_port, G_2_1_port, G_1_1_port, P_16_16_port, P_16_15_port, 
      P_16_13_port, P_16_9_port, P_15_15_port, P_14_14_port, P_14_13_port, 
      P_13_13_port, P_12_12_port, P_12_11_port, P_12_9_port, P_11_11_port, 
      P_10_10_port, P_10_9_port, P_9_9_port, P_8_8_port, P_8_7_port, P_8_5_port
      , P_7_7_port, P_6_6_port, P_6_5_port, P_5_5_port, P_4_4_port, P_4_3_port,
      P_3_3_port, P_2_2_port, G_32_32_port, G_32_31_port, G_32_29_port, 
      G_32_25_port, G_32_17_port, G_31_31_port, G_30_30_port, G_30_29_port, 
      G_29_29_port, G_28_28_port, G_28_27_port, G_28_25_port, G_28_17_port, 
      G_27_27_port, G_26_26_port, G_26_25_port, G_25_25_port, G_24_24_port, 
      G_24_23_port, G_24_21_port, G_24_17_port, G_23_23_port, G_22_22_port, 
      G_22_21_port, G_21_21_port, G_20_20_port, G_20_19_port, G_20_17_port, 
      G_19_19_port, G_18_18_port, G_18_17_port, G_17_17_port, P_32_32_port, 
      P_32_31_port, P_32_29_port, P_32_25_port, P_32_17_port, P_31_31_port, 
      P_30_30_port, P_30_29_port, P_29_29_port, P_28_28_port, P_28_27_port, 
      P_28_25_port, P_28_17_port, P_27_27_port, P_26_26_port, P_26_25_port, 
      P_25_25_port, P_24_24_port, P_24_23_port, P_24_21_port, P_24_17_port, 
      P_23_23_port, P_22_22_port, P_22_21_port, P_21_21_port, P_20_20_port, 
      P_20_19_port, P_20_17_port, P_19_19_port, P_18_18_port, P_18_17_port, 
      P_17_17_port, n3, n1, n2 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port );
   
   PGnetblock_2 : PG_net_0 port map( a => A(2), b => B(2), p => P_2_2_port, g 
                           => G_2_2_port);
   PGnetblock_3 : PG_net_30 port map( a => A(3), b => B(3), p => P_3_3_port, g 
                           => G_3_3_port);
   PGnetblock_4 : PG_net_29 port map( a => A(4), b => B(4), p => P_4_4_port, g 
                           => G_4_4_port);
   PGnetblock_5 : PG_net_28 port map( a => A(5), b => B(5), p => P_5_5_port, g 
                           => G_5_5_port);
   PGnetblock_6 : PG_net_27 port map( a => A(6), b => B(6), p => P_6_6_port, g 
                           => G_6_6_port);
   PGnetblock_7 : PG_net_26 port map( a => A(7), b => B(7), p => P_7_7_port, g 
                           => G_7_7_port);
   PGnetblock_8 : PG_net_25 port map( a => A(8), b => B(8), p => P_8_8_port, g 
                           => G_8_8_port);
   PGnetblock_9 : PG_net_24 port map( a => A(9), b => B(9), p => P_9_9_port, g 
                           => G_9_9_port);
   PGnetblock_10 : PG_net_23 port map( a => A(10), b => B(10), p => 
                           P_10_10_port, g => G_10_10_port);
   PGnetblock_11 : PG_net_22 port map( a => A(11), b => B(11), p => 
                           P_11_11_port, g => G_11_11_port);
   PGnetblock_12 : PG_net_21 port map( a => A(12), b => B(12), p => 
                           P_12_12_port, g => G_12_12_port);
   PGnetblock_13 : PG_net_20 port map( a => A(13), b => B(13), p => 
                           P_13_13_port, g => G_13_13_port);
   PGnetblock_14 : PG_net_19 port map( a => A(14), b => B(14), p => 
                           P_14_14_port, g => G_14_14_port);
   PGnetblock_15 : PG_net_18 port map( a => A(15), b => B(15), p => 
                           P_15_15_port, g => G_15_15_port);
   PGnetblock_16 : PG_net_17 port map( a => A(16), b => B(16), p => 
                           P_16_16_port, g => G_16_16_port);
   PGnetblock_17 : PG_net_16 port map( a => A(17), b => B(17), p => 
                           P_17_17_port, g => G_17_17_port);
   PGnetblock_18 : PG_net_15 port map( a => A(18), b => B(18), p => 
                           P_18_18_port, g => G_18_18_port);
   PGnetblock_19 : PG_net_14 port map( a => A(19), b => B(19), p => 
                           P_19_19_port, g => G_19_19_port);
   PGnetblock_20 : PG_net_13 port map( a => A(20), b => B(20), p => 
                           P_20_20_port, g => G_20_20_port);
   PGnetblock_21 : PG_net_12 port map( a => A(21), b => B(21), p => 
                           P_21_21_port, g => G_21_21_port);
   PGnetblock_22 : PG_net_11 port map( a => A(22), b => B(22), p => 
                           P_22_22_port, g => G_22_22_port);
   PGnetblock_23 : PG_net_10 port map( a => A(23), b => B(23), p => 
                           P_23_23_port, g => G_23_23_port);
   PGnetblock_24 : PG_net_9 port map( a => A(24), b => B(24), p => P_24_24_port
                           , g => G_24_24_port);
   PGnetblock_25 : PG_net_8 port map( a => A(25), b => B(25), p => P_25_25_port
                           , g => G_25_25_port);
   PGnetblock_26 : PG_net_7 port map( a => A(26), b => B(26), p => P_26_26_port
                           , g => G_26_26_port);
   PGnetblock_27 : PG_net_6 port map( a => A(27), b => B(27), p => P_27_27_port
                           , g => G_27_27_port);
   PGnetblock_28 : PG_net_5 port map( a => A(28), b => B(28), p => P_28_28_port
                           , g => G_28_28_port);
   PGnetblock_29 : PG_net_4 port map( a => A(29), b => B(29), p => P_29_29_port
                           , g => G_29_29_port);
   PGnetblock_30 : PG_net_3 port map( a => A(30), b => B(30), p => P_30_30_port
                           , g => G_30_30_port);
   PGnetblock_31 : PG_net_2 port map( a => A(31), b => B(31), p => P_31_31_port
                           , g => G_31_31_port);
   PGnetblock_32 : PG_net_1 port map( a => A(32), b => B(32), p => P_32_32_port
                           , g => G_32_32_port);
   GB_low_1_2 : Gblock_0 port map( Pik => P_2_2_port, Gik => G_2_2_port, Gk_1j 
                           => G_1_1_port, Gij => G_2_1_port);
   GB_low_2_4 : Gblock_8 port map( Pik => P_4_3_port, Gik => G_4_3_port, Gk_1j 
                           => G_2_1_port, Gij => Co_0_port);
   GB_low_3_8 : Gblock_7 port map( Pik => P_8_5_port, Gik => G_8_5_port, Gk_1j 
                           => Co_0_port, Gij => Co_1_port);
   GB_high_4_16_0 : Gblock_6 port map( Pik => P_16_9_port, Gik => G_16_9_port, 
                           Gk_1j => Co_1_port, Gij => Co_3_port);
   GB_high_4_16_1 : Gblock_5 port map( Pik => P_12_9_port, Gik => G_12_9_port, 
                           Gk_1j => Co_1_port, Gij => Co_2_port);
   GB_high_5_32_0 : Gblock_4 port map( Pik => P_32_17_port, Gik => G_32_17_port
                           , Gk_1j => Co_3_port, Gij => Co_7_port);
   GB_high_5_32_1 : Gblock_3 port map( Pik => P_28_17_port, Gik => G_28_17_port
                           , Gk_1j => Co_3_port, Gij => Co_6_port);
   GB_high_5_32_2 : Gblock_2 port map( Pik => P_24_17_port, Gik => G_24_17_port
                           , Gk_1j => Co_3_port, Gij => Co_5_port);
   GB_high_5_32_3 : Gblock_1 port map( Pik => P_20_17_port, Gik => G_20_17_port
                           , Gk_1j => Co_3_port, Gij => Co_4_port);
   PGB_low_1_4 : PGblock_0 port map( Pik => P_4_4_port, Gik => G_4_4_port, 
                           Pk_1j => P_3_3_port, Gk_1j => G_3_3_port, Pij => 
                           P_4_3_port, Gij => G_4_3_port);
   PGB_low_1_6 : PGblock_26 port map( Pik => P_6_6_port, Gik => G_6_6_port, 
                           Pk_1j => P_5_5_port, Gk_1j => G_5_5_port, Pij => 
                           P_6_5_port, Gij => G_6_5_port);
   PGB_low_1_8 : PGblock_25 port map( Pik => P_8_8_port, Gik => G_8_8_port, 
                           Pk_1j => P_7_7_port, Gk_1j => G_7_7_port, Pij => 
                           P_8_7_port, Gij => G_8_7_port);
   PGB_low_1_10 : PGblock_24 port map( Pik => P_10_10_port, Gik => G_10_10_port
                           , Pk_1j => P_9_9_port, Gk_1j => G_9_9_port, Pij => 
                           P_10_9_port, Gij => G_10_9_port);
   PGB_low_1_12 : PGblock_23 port map( Pik => P_12_12_port, Gik => G_12_12_port
                           , Pk_1j => P_11_11_port, Gk_1j => G_11_11_port, Pij 
                           => P_12_11_port, Gij => G_12_11_port);
   PGB_low_1_14 : PGblock_22 port map( Pik => P_14_14_port, Gik => G_14_14_port
                           , Pk_1j => P_13_13_port, Gk_1j => G_13_13_port, Pij 
                           => P_14_13_port, Gij => G_14_13_port);
   PGB_low_1_16 : PGblock_21 port map( Pik => P_16_16_port, Gik => G_16_16_port
                           , Pk_1j => P_15_15_port, Gk_1j => G_15_15_port, Pij 
                           => P_16_15_port, Gij => G_16_15_port);
   PGB_low_1_18 : PGblock_20 port map( Pik => P_18_18_port, Gik => G_18_18_port
                           , Pk_1j => P_17_17_port, Gk_1j => G_17_17_port, Pij 
                           => P_18_17_port, Gij => G_18_17_port);
   PGB_low_1_20 : PGblock_19 port map( Pik => P_20_20_port, Gik => G_20_20_port
                           , Pk_1j => P_19_19_port, Gk_1j => G_19_19_port, Pij 
                           => P_20_19_port, Gij => G_20_19_port);
   PGB_low_1_22 : PGblock_18 port map( Pik => P_22_22_port, Gik => G_22_22_port
                           , Pk_1j => P_21_21_port, Gk_1j => G_21_21_port, Pij 
                           => P_22_21_port, Gij => G_22_21_port);
   PGB_low_1_24 : PGblock_17 port map( Pik => P_24_24_port, Gik => G_24_24_port
                           , Pk_1j => P_23_23_port, Gk_1j => G_23_23_port, Pij 
                           => P_24_23_port, Gij => G_24_23_port);
   PGB_low_1_26 : PGblock_16 port map( Pik => P_26_26_port, Gik => G_26_26_port
                           , Pk_1j => P_25_25_port, Gk_1j => G_25_25_port, Pij 
                           => P_26_25_port, Gij => G_26_25_port);
   PGB_low_1_28 : PGblock_15 port map( Pik => P_28_28_port, Gik => G_28_28_port
                           , Pk_1j => P_27_27_port, Gk_1j => G_27_27_port, Pij 
                           => P_28_27_port, Gij => G_28_27_port);
   PGB_low_1_30 : PGblock_14 port map( Pik => P_30_30_port, Gik => G_30_30_port
                           , Pk_1j => P_29_29_port, Gk_1j => G_29_29_port, Pij 
                           => P_30_29_port, Gij => G_30_29_port);
   PGB_low_1_32 : PGblock_13 port map( Pik => P_32_32_port, Gik => G_32_32_port
                           , Pk_1j => P_31_31_port, Gk_1j => G_31_31_port, Pij 
                           => P_32_31_port, Gij => G_32_31_port);
   PGB_low_2_8 : PGblock_12 port map( Pik => P_8_7_port, Gik => G_8_7_port, 
                           Pk_1j => P_6_5_port, Gk_1j => G_6_5_port, Pij => 
                           P_8_5_port, Gij => G_8_5_port);
   PGB_low_2_12 : PGblock_11 port map( Pik => P_12_11_port, Gik => G_12_11_port
                           , Pk_1j => P_10_9_port, Gk_1j => G_10_9_port, Pij =>
                           P_12_9_port, Gij => G_12_9_port);
   PGB_low_2_16 : PGblock_10 port map( Pik => P_16_15_port, Gik => G_16_15_port
                           , Pk_1j => P_14_13_port, Gk_1j => G_14_13_port, Pij 
                           => P_16_13_port, Gij => G_16_13_port);
   PGB_low_2_20 : PGblock_9 port map( Pik => P_20_19_port, Gik => G_20_19_port,
                           Pk_1j => P_18_17_port, Gk_1j => G_18_17_port, Pij =>
                           P_20_17_port, Gij => G_20_17_port);
   PGB_low_2_24 : PGblock_8 port map( Pik => P_24_23_port, Gik => G_24_23_port,
                           Pk_1j => P_22_21_port, Gk_1j => G_22_21_port, Pij =>
                           P_24_21_port, Gij => G_24_21_port);
   PGB_low_2_28 : PGblock_7 port map( Pik => P_28_27_port, Gik => G_28_27_port,
                           Pk_1j => P_26_25_port, Gk_1j => G_26_25_port, Pij =>
                           P_28_25_port, Gij => G_28_25_port);
   PGB_low_2_32 : PGblock_6 port map( Pik => P_32_31_port, Gik => G_32_31_port,
                           Pk_1j => P_30_29_port, Gk_1j => G_30_29_port, Pij =>
                           P_32_29_port, Gij => G_32_29_port);
   PGB_low_3_16 : PGblock_5 port map( Pik => P_16_13_port, Gik => G_16_13_port,
                           Pk_1j => P_12_9_port, Gk_1j => G_12_9_port, Pij => 
                           P_16_9_port, Gij => G_16_9_port);
   PGB_low_3_24 : PGblock_4 port map( Pik => P_24_21_port, Gik => G_24_21_port,
                           Pk_1j => P_20_17_port, Gk_1j => G_20_17_port, Pij =>
                           P_24_17_port, Gij => G_24_17_port);
   PGB_low_3_32 : PGblock_3 port map( Pik => P_32_29_port, Gik => G_32_29_port,
                           Pk_1j => P_28_25_port, Gk_1j => G_28_25_port, Pij =>
                           P_32_25_port, Gij => G_32_25_port);
   PGB_high_4_32_0 : PGblock_2 port map( Pik => P_32_25_port, Gik => 
                           G_32_25_port, Pk_1j => P_24_17_port, Gk_1j => 
                           G_24_17_port, Pij => P_32_17_port, Gij => 
                           G_32_17_port);
   PGB_high_4_32_1 : PGblock_1 port map( Pik => P_28_25_port, Gik => 
                           G_28_25_port, Pk_1j => P_24_17_port, Gk_1j => 
                           G_24_17_port, Pij => P_28_17_port, Gij => 
                           G_28_17_port);
   U1 : INV_X1 port map( A => A(1), ZN => n1);
   U2 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => G_1_1_port);
   U3 : INV_X1 port map( A => B(1), ZN => n2);
   U4 : OAI21_X1 port map( B1 => A(1), B2 => B(1), A => Cin, ZN => n3);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity BOOTHMUL_numBit16 is

   port( A, B : in std_logic_vector (15 downto 0);  P : out std_logic_vector 
         (31 downto 0));

end BOOTHMUL_numBit16;

architecture SYN_mixed of BOOTHMUL_numBit16 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component rca_bhv_numBit32_1
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component rca_bhv_numBit32_2
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component rca_bhv_numBit32_3
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component rca_bhv_numBit32_4
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component rca_bhv_numBit32_5
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component rca_bhv_numBit32_6
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component rca_bhv_numBit32_0
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   component mux5to1_numBit32_1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux5to1_numBit32_2
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux5to1_numBit32_3
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux5to1_numBit32_4
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux5to1_numBit32_5
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux5to1_numBit32_6
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux5to1_numBit32_7
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux5to1_numBit32_0
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic_vector (31 downto 0);  
            SEL_in : in std_logic_vector (2 downto 0);  Z : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component booth_encoder_numBit16
      port( B : in std_logic_vector (15 downto 0);  SEL_out : out 
            std_logic_vector (23 downto 0));
   end component;
   
   signal X_Logic0_port, encoder_out_23_port, encoder_out_22_port, 
      encoder_out_21_port, encoder_out_20_port, encoder_out_19_port, 
      encoder_out_18_port, encoder_out_17_port, encoder_out_16_port, 
      encoder_out_15_port, encoder_out_14_port, encoder_out_13_port, 
      encoder_out_12_port, encoder_out_11_port, encoder_out_10_port, 
      encoder_out_9_port, encoder_out_8_port, encoder_out_7_port, 
      encoder_out_6_port, encoder_out_5_port, encoder_out_4_port, 
      encoder_out_3_port, encoder_out_2_port, encoder_out_1_port, 
      encoder_out_0_port, A_minus_31_port, A_minus_15_port, A_minus_14_port, 
      A_minus_13_port, A_minus_12_port, A_minus_11_port, A_minus_10_port, 
      A_minus_9_port, A_minus_8_port, A_minus_7_port, A_minus_6_port, 
      A_minus_5_port, A_minus_4_port, A_minus_3_port, A_minus_2_port, 
      A_minus_1_port, A_minus_0_port, sum_op_7_31_port, sum_op_7_30_port, 
      sum_op_7_29_port, sum_op_7_28_port, sum_op_7_27_port, sum_op_7_26_port, 
      sum_op_7_25_port, sum_op_7_24_port, sum_op_7_23_port, sum_op_7_22_port, 
      sum_op_7_21_port, sum_op_7_20_port, sum_op_7_19_port, sum_op_7_18_port, 
      sum_op_7_17_port, sum_op_7_16_port, sum_op_7_15_port, sum_op_7_14_port, 
      sum_op_7_13_port, sum_op_7_12_port, sum_op_7_11_port, sum_op_7_10_port, 
      sum_op_7_9_port, sum_op_7_8_port, sum_op_7_7_port, sum_op_7_6_port, 
      sum_op_7_5_port, sum_op_7_4_port, sum_op_7_3_port, sum_op_7_2_port, 
      sum_op_7_1_port, sum_op_7_0_port, sum_op_6_31_port, sum_op_6_30_port, 
      sum_op_6_29_port, sum_op_6_28_port, sum_op_6_27_port, sum_op_6_26_port, 
      sum_op_6_25_port, sum_op_6_24_port, sum_op_6_23_port, sum_op_6_22_port, 
      sum_op_6_21_port, sum_op_6_20_port, sum_op_6_19_port, sum_op_6_18_port, 
      sum_op_6_17_port, sum_op_6_16_port, sum_op_6_15_port, sum_op_6_14_port, 
      sum_op_6_13_port, sum_op_6_12_port, sum_op_6_11_port, sum_op_6_10_port, 
      sum_op_6_9_port, sum_op_6_8_port, sum_op_6_7_port, sum_op_6_6_port, 
      sum_op_6_5_port, sum_op_6_4_port, sum_op_6_3_port, sum_op_6_2_port, 
      sum_op_6_1_port, sum_op_6_0_port, sum_op_5_31_port, sum_op_5_30_port, 
      sum_op_5_29_port, sum_op_5_28_port, sum_op_5_27_port, sum_op_5_26_port, 
      sum_op_5_25_port, sum_op_5_24_port, sum_op_5_23_port, sum_op_5_22_port, 
      sum_op_5_21_port, sum_op_5_20_port, sum_op_5_19_port, sum_op_5_18_port, 
      sum_op_5_17_port, sum_op_5_16_port, sum_op_5_15_port, sum_op_5_14_port, 
      sum_op_5_13_port, sum_op_5_12_port, sum_op_5_11_port, sum_op_5_10_port, 
      sum_op_5_9_port, sum_op_5_8_port, sum_op_5_7_port, sum_op_5_6_port, 
      sum_op_5_5_port, sum_op_5_4_port, sum_op_5_3_port, sum_op_5_2_port, 
      sum_op_5_1_port, sum_op_5_0_port, sum_op_4_31_port, sum_op_4_30_port, 
      sum_op_4_29_port, sum_op_4_28_port, sum_op_4_27_port, sum_op_4_26_port, 
      sum_op_4_25_port, sum_op_4_24_port, sum_op_4_23_port, sum_op_4_22_port, 
      sum_op_4_21_port, sum_op_4_20_port, sum_op_4_19_port, sum_op_4_18_port, 
      sum_op_4_17_port, sum_op_4_16_port, sum_op_4_15_port, sum_op_4_14_port, 
      sum_op_4_13_port, sum_op_4_12_port, sum_op_4_11_port, sum_op_4_10_port, 
      sum_op_4_9_port, sum_op_4_8_port, sum_op_4_7_port, sum_op_4_6_port, 
      sum_op_4_5_port, sum_op_4_4_port, sum_op_4_3_port, sum_op_4_2_port, 
      sum_op_4_1_port, sum_op_4_0_port, sum_op_3_31_port, sum_op_3_30_port, 
      sum_op_3_29_port, sum_op_3_28_port, sum_op_3_27_port, sum_op_3_26_port, 
      sum_op_3_25_port, sum_op_3_24_port, sum_op_3_23_port, sum_op_3_22_port, 
      sum_op_3_21_port, sum_op_3_20_port, sum_op_3_19_port, sum_op_3_18_port, 
      sum_op_3_17_port, sum_op_3_16_port, sum_op_3_15_port, sum_op_3_14_port, 
      sum_op_3_13_port, sum_op_3_12_port, sum_op_3_11_port, sum_op_3_10_port, 
      sum_op_3_9_port, sum_op_3_8_port, sum_op_3_7_port, sum_op_3_6_port, 
      sum_op_3_5_port, sum_op_3_4_port, sum_op_3_3_port, sum_op_3_2_port, 
      sum_op_3_1_port, sum_op_3_0_port, sum_op_2_31_port, sum_op_2_30_port, 
      sum_op_2_29_port, sum_op_2_28_port, sum_op_2_27_port, sum_op_2_26_port, 
      sum_op_2_25_port, sum_op_2_24_port, sum_op_2_23_port, sum_op_2_22_port, 
      sum_op_2_21_port, sum_op_2_20_port, sum_op_2_19_port, sum_op_2_18_port, 
      sum_op_2_17_port, sum_op_2_16_port, sum_op_2_15_port, sum_op_2_14_port, 
      sum_op_2_13_port, sum_op_2_12_port, sum_op_2_11_port, sum_op_2_10_port, 
      sum_op_2_9_port, sum_op_2_8_port, sum_op_2_7_port, sum_op_2_6_port, 
      sum_op_2_5_port, sum_op_2_4_port, sum_op_2_3_port, sum_op_2_2_port, 
      sum_op_2_1_port, sum_op_2_0_port, sum_op_1_31_port, sum_op_1_30_port, 
      sum_op_1_29_port, sum_op_1_28_port, sum_op_1_27_port, sum_op_1_26_port, 
      sum_op_1_25_port, sum_op_1_24_port, sum_op_1_23_port, sum_op_1_22_port, 
      sum_op_1_21_port, sum_op_1_20_port, sum_op_1_19_port, sum_op_1_18_port, 
      sum_op_1_17_port, sum_op_1_16_port, sum_op_1_15_port, sum_op_1_14_port, 
      sum_op_1_13_port, sum_op_1_12_port, sum_op_1_11_port, sum_op_1_10_port, 
      sum_op_1_9_port, sum_op_1_8_port, sum_op_1_7_port, sum_op_1_6_port, 
      sum_op_1_5_port, sum_op_1_4_port, sum_op_1_3_port, sum_op_1_2_port, 
      sum_op_1_1_port, sum_op_1_0_port, sum_op_0_31_port, sum_op_0_30_port, 
      sum_op_0_29_port, sum_op_0_28_port, sum_op_0_27_port, sum_op_0_26_port, 
      sum_op_0_25_port, sum_op_0_24_port, sum_op_0_23_port, sum_op_0_22_port, 
      sum_op_0_21_port, sum_op_0_20_port, sum_op_0_19_port, sum_op_0_18_port, 
      sum_op_0_17_port, sum_op_0_16_port, sum_op_0_15_port, sum_op_0_14_port, 
      sum_op_0_13_port, sum_op_0_12_port, sum_op_0_11_port, sum_op_0_10_port, 
      sum_op_0_9_port, sum_op_0_8_port, sum_op_0_7_port, sum_op_0_6_port, 
      sum_op_0_5_port, sum_op_0_4_port, sum_op_0_3_port, sum_op_0_2_port, 
      sum_op_0_1_port, sum_op_0_0_port, rca_out_5_31_port, rca_out_5_30_port, 
      rca_out_5_29_port, rca_out_5_28_port, rca_out_5_27_port, 
      rca_out_5_26_port, rca_out_5_25_port, rca_out_5_24_port, 
      rca_out_5_23_port, rca_out_5_22_port, rca_out_5_21_port, 
      rca_out_5_20_port, rca_out_5_19_port, rca_out_5_18_port, 
      rca_out_5_17_port, rca_out_5_16_port, rca_out_5_15_port, 
      rca_out_5_14_port, rca_out_5_13_port, rca_out_5_12_port, 
      rca_out_5_11_port, rca_out_5_10_port, rca_out_5_9_port, rca_out_5_8_port,
      rca_out_5_7_port, rca_out_5_6_port, rca_out_5_5_port, rca_out_5_4_port, 
      rca_out_5_3_port, rca_out_5_2_port, rca_out_5_1_port, rca_out_5_0_port, 
      rca_out_4_31_port, rca_out_4_30_port, rca_out_4_29_port, 
      rca_out_4_28_port, rca_out_4_27_port, rca_out_4_26_port, 
      rca_out_4_25_port, rca_out_4_24_port, rca_out_4_23_port, 
      rca_out_4_22_port, rca_out_4_21_port, rca_out_4_20_port, 
      rca_out_4_19_port, rca_out_4_18_port, rca_out_4_17_port, 
      rca_out_4_16_port, rca_out_4_15_port, rca_out_4_14_port, 
      rca_out_4_13_port, rca_out_4_12_port, rca_out_4_11_port, 
      rca_out_4_10_port, rca_out_4_9_port, rca_out_4_8_port, rca_out_4_7_port, 
      rca_out_4_6_port, rca_out_4_5_port, rca_out_4_4_port, rca_out_4_3_port, 
      rca_out_4_2_port, rca_out_4_1_port, rca_out_4_0_port, rca_out_3_31_port, 
      rca_out_3_30_port, rca_out_3_29_port, rca_out_3_28_port, 
      rca_out_3_27_port, rca_out_3_26_port, rca_out_3_25_port, 
      rca_out_3_24_port, rca_out_3_23_port, rca_out_3_22_port, 
      rca_out_3_21_port, rca_out_3_20_port, rca_out_3_19_port, 
      rca_out_3_18_port, rca_out_3_17_port, rca_out_3_16_port, 
      rca_out_3_15_port, rca_out_3_14_port, rca_out_3_13_port, 
      rca_out_3_12_port, rca_out_3_11_port, rca_out_3_10_port, rca_out_3_9_port
      , rca_out_3_8_port, rca_out_3_7_port, rca_out_3_6_port, rca_out_3_5_port,
      rca_out_3_4_port, rca_out_3_3_port, rca_out_3_2_port, rca_out_3_1_port, 
      rca_out_3_0_port, rca_out_2_31_port, rca_out_2_30_port, rca_out_2_29_port
      , rca_out_2_28_port, rca_out_2_27_port, rca_out_2_26_port, 
      rca_out_2_25_port, rca_out_2_24_port, rca_out_2_23_port, 
      rca_out_2_22_port, rca_out_2_21_port, rca_out_2_20_port, 
      rca_out_2_19_port, rca_out_2_18_port, rca_out_2_17_port, 
      rca_out_2_16_port, rca_out_2_15_port, rca_out_2_14_port, 
      rca_out_2_13_port, rca_out_2_12_port, rca_out_2_11_port, 
      rca_out_2_10_port, rca_out_2_9_port, rca_out_2_8_port, rca_out_2_7_port, 
      rca_out_2_6_port, rca_out_2_5_port, rca_out_2_4_port, rca_out_2_3_port, 
      rca_out_2_2_port, rca_out_2_1_port, rca_out_2_0_port, rca_out_1_31_port, 
      rca_out_1_30_port, rca_out_1_29_port, rca_out_1_28_port, 
      rca_out_1_27_port, rca_out_1_26_port, rca_out_1_25_port, 
      rca_out_1_24_port, rca_out_1_23_port, rca_out_1_22_port, 
      rca_out_1_21_port, rca_out_1_20_port, rca_out_1_19_port, 
      rca_out_1_18_port, rca_out_1_17_port, rca_out_1_16_port, 
      rca_out_1_15_port, rca_out_1_14_port, rca_out_1_13_port, 
      rca_out_1_12_port, rca_out_1_11_port, rca_out_1_10_port, rca_out_1_9_port
      , rca_out_1_8_port, rca_out_1_7_port, rca_out_1_6_port, rca_out_1_5_port,
      rca_out_1_4_port, rca_out_1_3_port, rca_out_1_2_port, rca_out_1_1_port, 
      rca_out_1_0_port, rca_out_0_31_port, rca_out_0_30_port, rca_out_0_29_port
      , rca_out_0_28_port, rca_out_0_27_port, rca_out_0_26_port, 
      rca_out_0_25_port, rca_out_0_24_port, rca_out_0_23_port, 
      rca_out_0_22_port, rca_out_0_21_port, rca_out_0_20_port, 
      rca_out_0_19_port, rca_out_0_18_port, rca_out_0_17_port, 
      rca_out_0_16_port, rca_out_0_15_port, rca_out_0_14_port, 
      rca_out_0_13_port, rca_out_0_12_port, rca_out_0_11_port, 
      rca_out_0_10_port, rca_out_0_9_port, rca_out_0_8_port, rca_out_0_7_port, 
      rca_out_0_6_port, rca_out_0_5_port, rca_out_0_4_port, rca_out_0_3_port, 
      rca_out_0_2_port, rca_out_0_1_port, rca_out_0_0_port, add_65_carry_2_port
      , add_65_carry_3_port, add_65_carry_4_port, add_65_carry_5_port, 
      add_65_carry_6_port, add_65_carry_7_port, add_65_carry_8_port, 
      add_65_carry_9_port, add_65_carry_10_port, add_65_carry_11_port, 
      add_65_carry_12_port, add_65_carry_13_port, add_65_carry_14_port, 
      add_65_carry_15_port, add_65_A_0_port, add_65_A_1_port, add_65_A_2_port, 
      add_65_A_3_port, add_65_A_4_port, add_65_A_5_port, add_65_A_6_port, 
      add_65_A_7_port, add_65_A_8_port, add_65_A_9_port, add_65_A_10_port, 
      add_65_A_11_port, add_65_A_12_port, add_65_A_13_port, add_65_A_14_port, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n_1158, n_1159, n_1160, 
      n_1161, n_1162, n_1163, n_1164, n_1165 : std_logic;

begin
   
   X_Logic0_port <= '0';
   encode : booth_encoder_numBit16 port map( B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           SEL_out(23) => encoder_out_23_port, SEL_out(22) => 
                           encoder_out_22_port, SEL_out(21) => 
                           encoder_out_21_port, SEL_out(20) => 
                           encoder_out_20_port, SEL_out(19) => 
                           encoder_out_19_port, SEL_out(18) => 
                           encoder_out_18_port, SEL_out(17) => 
                           encoder_out_17_port, SEL_out(16) => 
                           encoder_out_16_port, SEL_out(15) => 
                           encoder_out_15_port, SEL_out(14) => 
                           encoder_out_14_port, SEL_out(13) => 
                           encoder_out_13_port, SEL_out(12) => 
                           encoder_out_12_port, SEL_out(11) => 
                           encoder_out_11_port, SEL_out(10) => 
                           encoder_out_10_port, SEL_out(9) => 
                           encoder_out_9_port, SEL_out(8) => encoder_out_8_port
                           , SEL_out(7) => encoder_out_7_port, SEL_out(6) => 
                           encoder_out_6_port, SEL_out(5) => encoder_out_5_port
                           , SEL_out(4) => encoder_out_4_port, SEL_out(3) => 
                           encoder_out_3_port, SEL_out(2) => encoder_out_2_port
                           , SEL_out(1) => encoder_out_1_port, SEL_out(0) => 
                           n_1158);
   mux0_0 : mux5to1_numBit32_0 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => n48, IN2(30) => n48, 
                           IN2(29) => n49, IN2(28) => n48, IN2(27) => n48, 
                           IN2(26) => n49, IN2(25) => n48, IN2(24) => n49, 
                           IN2(23) => n48, IN2(22) => n48, IN2(21) => n48, 
                           IN2(20) => n49, IN2(19) => n48, IN2(18) => n49, 
                           IN2(17) => n48, IN2(16) => n49, IN2(15) => n48, 
                           IN2(14) => A(14), IN2(13) => A(13), IN2(12) => A(12)
                           , IN2(11) => A(11), IN2(10) => A(10), IN2(9) => A(9)
                           , IN2(8) => A(8), IN2(7) => A(7), IN2(6) => A(6), 
                           IN2(5) => A(5), IN2(4) => A(4), IN2(3) => A(3), 
                           IN2(2) => A(2), IN2(1) => A(1), IN2(0) => A(0), 
                           IN3(31) => n35, IN3(30) => n31, IN3(29) => n31, 
                           IN3(28) => n36, IN3(27) => n31, IN3(26) => n35, 
                           IN3(25) => n31, IN3(24) => n36, IN3(23) => n31, 
                           IN3(22) => n36, IN3(21) => n32, IN3(20) => n35, 
                           IN3(19) => n32, IN3(18) => n35, IN3(17) => n33, 
                           IN3(16) => n34, IN3(15) => A_minus_15_port, IN3(14) 
                           => n2, IN3(13) => n4, IN3(12) => n6, IN3(11) => n8, 
                           IN3(10) => n10, IN3(9) => n12, IN3(8) => n14, IN3(7)
                           => n16, IN3(6) => n18, IN3(5) => n20, IN3(4) => n22,
                           IN3(3) => n24, IN3(2) => n26, IN3(1) => n28, IN3(0) 
                           => A_minus_0_port, IN4(31) => n42, IN4(30) => n42, 
                           IN4(29) => n42, IN4(28) => n42, IN4(27) => n42, 
                           IN4(26) => n42, IN4(25) => n42, IN4(24) => n42, 
                           IN4(23) => n42, IN4(22) => n42, IN4(21) => n42, 
                           IN4(20) => n43, IN4(19) => n43, IN4(18) => n43, 
                           IN4(17) => n43, IN4(16) => n43, IN4(15) => A(14), 
                           IN4(14) => A(13), IN4(13) => A(12), IN4(12) => A(11)
                           , IN4(11) => A(10), IN4(10) => A(9), IN4(9) => A(8),
                           IN4(8) => A(7), IN4(7) => A(6), IN4(6) => A(5), 
                           IN4(5) => A(4), IN4(4) => A(3), IN4(3) => A(2), 
                           IN4(2) => A(1), IN4(1) => A(0), IN4(0) => 
                           X_Logic0_port, IN5(31) => n41, IN5(30) => n41, 
                           IN5(29) => n41, IN5(28) => n41, IN5(27) => n41, 
                           IN5(26) => n41, IN5(25) => n40, IN5(24) => n40, 
                           IN5(23) => n39, IN5(22) => n40, IN5(21) => n38, 
                           IN5(20) => n39, IN5(19) => n38, IN5(18) => n38, 
                           IN5(17) => n39, IN5(16) => A_minus_15_port, IN5(15) 
                           => n2, IN5(14) => n4, IN5(13) => n6, IN5(12) => n8, 
                           IN5(11) => n10, IN5(10) => n12, IN5(9) => n14, 
                           IN5(8) => n16, IN5(7) => n18, IN5(6) => n20, IN5(5) 
                           => n22, IN5(4) => n24, IN5(3) => n26, IN5(2) => n28,
                           IN5(1) => A_minus_0_port, IN5(0) => X_Logic0_port, 
                           SEL_in(2) => encoder_out_2_port, SEL_in(1) => 
                           encoder_out_1_port, SEL_in(0) => encoder_out_0_port,
                           Z(31) => sum_op_0_31_port, Z(30) => sum_op_0_30_port
                           , Z(29) => sum_op_0_29_port, Z(28) => 
                           sum_op_0_28_port, Z(27) => sum_op_0_27_port, Z(26) 
                           => sum_op_0_26_port, Z(25) => sum_op_0_25_port, 
                           Z(24) => sum_op_0_24_port, Z(23) => sum_op_0_23_port
                           , Z(22) => sum_op_0_22_port, Z(21) => 
                           sum_op_0_21_port, Z(20) => sum_op_0_20_port, Z(19) 
                           => sum_op_0_19_port, Z(18) => sum_op_0_18_port, 
                           Z(17) => sum_op_0_17_port, Z(16) => sum_op_0_16_port
                           , Z(15) => sum_op_0_15_port, Z(14) => 
                           sum_op_0_14_port, Z(13) => sum_op_0_13_port, Z(12) 
                           => sum_op_0_12_port, Z(11) => sum_op_0_11_port, 
                           Z(10) => sum_op_0_10_port, Z(9) => sum_op_0_9_port, 
                           Z(8) => sum_op_0_8_port, Z(7) => sum_op_0_7_port, 
                           Z(6) => sum_op_0_6_port, Z(5) => sum_op_0_5_port, 
                           Z(4) => sum_op_0_4_port, Z(3) => sum_op_0_3_port, 
                           Z(2) => sum_op_0_2_port, Z(1) => sum_op_0_1_port, 
                           Z(0) => sum_op_0_0_port);
   mux_i_1 : mux5to1_numBit32_7 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => n52, IN2(30) => n51, 
                           IN2(29) => n51, IN2(28) => n51, IN2(27) => n51, 
                           IN2(26) => n51, IN2(25) => n50, IN2(24) => n50, 
                           IN2(23) => n50, IN2(22) => n50, IN2(21) => n50, 
                           IN2(20) => n49, IN2(19) => n49, IN2(18) => n49, 
                           IN2(17) => n49, IN2(16) => A(14), IN2(15) => A(13), 
                           IN2(14) => A(12), IN2(13) => A(11), IN2(12) => A(10)
                           , IN2(11) => A(9), IN2(10) => A(8), IN2(9) => A(7), 
                           IN2(8) => A(6), IN2(7) => A(5), IN2(6) => A(4), 
                           IN2(5) => A(3), IN2(4) => A(2), IN2(3) => A(1), 
                           IN2(2) => A(0), IN2(1) => X_Logic0_port, IN2(0) => 
                           X_Logic0_port, IN3(31) => n31, IN3(30) => n36, 
                           IN3(29) => n31, IN3(28) => n35, IN3(27) => n31, 
                           IN3(26) => n35, IN3(25) => n32, IN3(24) => n36, 
                           IN3(23) => n32, IN3(22) => n35, IN3(21) => n33, 
                           IN3(20) => n34, IN3(19) => n33, IN3(18) => n34, 
                           IN3(17) => A_minus_15_port, IN3(16) => n2, IN3(15) 
                           => n4, IN3(14) => n6, IN3(13) => n8, IN3(12) => n10,
                           IN3(11) => n12, IN3(10) => n14, IN3(9) => n16, 
                           IN3(8) => n18, IN3(7) => n20, IN3(6) => n22, IN3(5) 
                           => n24, IN3(4) => n26, IN3(3) => n28, IN3(2) => 
                           A_minus_0_port, IN3(1) => X_Logic0_port, IN3(0) => 
                           X_Logic0_port, IN4(31) => n47, IN4(30) => n47, 
                           IN4(29) => n47, IN4(28) => n47, IN4(27) => n46, 
                           IN4(26) => n47, IN4(25) => n47, IN4(24) => n47, 
                           IN4(23) => n46, IN4(22) => n46, IN4(21) => n46, 
                           IN4(20) => n46, IN4(19) => n46, IN4(18) => n42, 
                           IN4(17) => A(14), IN4(16) => A(13), IN4(15) => A(12)
                           , IN4(14) => A(11), IN4(13) => A(10), IN4(12) => 
                           A(9), IN4(11) => A(8), IN4(10) => A(7), IN4(9) => 
                           A(6), IN4(8) => A(5), IN4(7) => A(4), IN4(6) => A(3)
                           , IN4(5) => A(2), IN4(4) => A(1), IN4(3) => A(0), 
                           IN4(2) => X_Logic0_port, IN4(1) => X_Logic0_port, 
                           IN4(0) => X_Logic0_port, IN5(31) => n41, IN5(30) => 
                           n41, IN5(29) => n40, IN5(28) => n40, IN5(27) => n40,
                           IN5(26) => n40, IN5(25) => n40, IN5(24) => n41, 
                           IN5(23) => n37, IN5(22) => n39, IN5(21) => n37, 
                           IN5(20) => n39, IN5(19) => n37, IN5(18) => 
                           A_minus_15_port, IN5(17) => n2, IN5(16) => n4, 
                           IN5(15) => n6, IN5(14) => n8, IN5(13) => n10, 
                           IN5(12) => n12, IN5(11) => n14, IN5(10) => n16, 
                           IN5(9) => n18, IN5(8) => n20, IN5(7) => n22, IN5(6) 
                           => n24, IN5(5) => n26, IN5(4) => n28, IN5(3) => 
                           A_minus_0_port, IN5(2) => X_Logic0_port, IN5(1) => 
                           X_Logic0_port, IN5(0) => X_Logic0_port, SEL_in(2) =>
                           encoder_out_5_port, SEL_in(1) => encoder_out_4_port,
                           SEL_in(0) => encoder_out_3_port, Z(31) => 
                           sum_op_1_31_port, Z(30) => sum_op_1_30_port, Z(29) 
                           => sum_op_1_29_port, Z(28) => sum_op_1_28_port, 
                           Z(27) => sum_op_1_27_port, Z(26) => sum_op_1_26_port
                           , Z(25) => sum_op_1_25_port, Z(24) => 
                           sum_op_1_24_port, Z(23) => sum_op_1_23_port, Z(22) 
                           => sum_op_1_22_port, Z(21) => sum_op_1_21_port, 
                           Z(20) => sum_op_1_20_port, Z(19) => sum_op_1_19_port
                           , Z(18) => sum_op_1_18_port, Z(17) => 
                           sum_op_1_17_port, Z(16) => sum_op_1_16_port, Z(15) 
                           => sum_op_1_15_port, Z(14) => sum_op_1_14_port, 
                           Z(13) => sum_op_1_13_port, Z(12) => sum_op_1_12_port
                           , Z(11) => sum_op_1_11_port, Z(10) => 
                           sum_op_1_10_port, Z(9) => sum_op_1_9_port, Z(8) => 
                           sum_op_1_8_port, Z(7) => sum_op_1_7_port, Z(6) => 
                           sum_op_1_6_port, Z(5) => sum_op_1_5_port, Z(4) => 
                           sum_op_1_4_port, Z(3) => sum_op_1_3_port, Z(2) => 
                           sum_op_1_2_port, Z(1) => sum_op_1_1_port, Z(0) => 
                           sum_op_1_0_port);
   mux_i_2 : mux5to1_numBit32_6 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => A(15), IN2(30) => A(15), 
                           IN2(29) => A(15), IN2(28) => A(15), IN2(27) => A(15)
                           , IN2(26) => A(15), IN2(25) => n48, IN2(24) => A(15)
                           , IN2(23) => A(15), IN2(22) => n53, IN2(21) => n53, 
                           IN2(20) => n53, IN2(19) => n53, IN2(18) => A(14), 
                           IN2(17) => A(13), IN2(16) => A(12), IN2(15) => A(11)
                           , IN2(14) => A(10), IN2(13) => A(9), IN2(12) => A(8)
                           , IN2(11) => A(7), IN2(10) => A(6), IN2(9) => A(5), 
                           IN2(8) => A(4), IN2(7) => A(3), IN2(6) => A(2), 
                           IN2(5) => A(1), IN2(4) => A(0), IN2(3) => 
                           X_Logic0_port, IN2(2) => X_Logic0_port, IN2(1) => 
                           X_Logic0_port, IN2(0) => X_Logic0_port, IN3(31) => 
                           n31, IN3(30) => n36, IN3(29) => n31, IN3(28) => n36,
                           IN3(27) => n32, IN3(26) => n36, IN3(25) => n32, 
                           IN3(24) => n36, IN3(23) => n33, IN3(22) => n34, 
                           IN3(21) => n33, IN3(20) => n34, IN3(19) => 
                           A_minus_15_port, IN3(18) => n2, IN3(17) => n4, 
                           IN3(16) => n6, IN3(15) => n8, IN3(14) => n10, 
                           IN3(13) => n12, IN3(12) => n14, IN3(11) => n16, 
                           IN3(10) => n18, IN3(9) => n20, IN3(8) => n22, IN3(7)
                           => n24, IN3(6) => n26, IN3(5) => n28, IN3(4) => 
                           A_minus_0_port, IN3(3) => X_Logic0_port, IN3(2) => 
                           X_Logic0_port, IN3(1) => X_Logic0_port, IN3(0) => 
                           X_Logic0_port, IN4(31) => n46, IN4(30) => n46, 
                           IN4(29) => n46, IN4(28) => n46, IN4(27) => n46, 
                           IN4(26) => n47, IN4(25) => n46, IN4(24) => n47, 
                           IN4(23) => n45, IN4(22) => n47, IN4(21) => n47, 
                           IN4(20) => n47, IN4(19) => A(14), IN4(18) => A(13), 
                           IN4(17) => A(12), IN4(16) => A(11), IN4(15) => A(10)
                           , IN4(14) => A(9), IN4(13) => A(8), IN4(12) => A(7),
                           IN4(11) => A(6), IN4(10) => A(5), IN4(9) => A(4), 
                           IN4(8) => A(3), IN4(7) => A(2), IN4(6) => A(1), 
                           IN4(5) => A(0), IN4(4) => X_Logic0_port, IN4(3) => 
                           X_Logic0_port, IN4(2) => X_Logic0_port, IN4(1) => 
                           X_Logic0_port, IN4(0) => X_Logic0_port, IN5(31) => 
                           n41, IN5(30) => n41, IN5(29) => n40, IN5(28) => n40,
                           IN5(27) => n39, IN5(26) => n39, IN5(25) => n38, 
                           IN5(24) => n38, IN5(23) => n37, IN5(22) => n37, 
                           IN5(21) => n38, IN5(20) => A_minus_15_port, IN5(19) 
                           => n2, IN5(18) => n4, IN5(17) => n6, IN5(16) => n8, 
                           IN5(15) => n10, IN5(14) => n12, IN5(13) => n14, 
                           IN5(12) => n16, IN5(11) => n18, IN5(10) => n20, 
                           IN5(9) => n22, IN5(8) => n24, IN5(7) => n26, IN5(6) 
                           => n28, IN5(5) => A_minus_0_port, IN5(4) => 
                           X_Logic0_port, IN5(3) => X_Logic0_port, IN5(2) => 
                           X_Logic0_port, IN5(1) => X_Logic0_port, IN5(0) => 
                           X_Logic0_port, SEL_in(2) => encoder_out_8_port, 
                           SEL_in(1) => encoder_out_7_port, SEL_in(0) => 
                           encoder_out_6_port, Z(31) => sum_op_2_31_port, Z(30)
                           => sum_op_2_30_port, Z(29) => sum_op_2_29_port, 
                           Z(28) => sum_op_2_28_port, Z(27) => sum_op_2_27_port
                           , Z(26) => sum_op_2_26_port, Z(25) => 
                           sum_op_2_25_port, Z(24) => sum_op_2_24_port, Z(23) 
                           => sum_op_2_23_port, Z(22) => sum_op_2_22_port, 
                           Z(21) => sum_op_2_21_port, Z(20) => sum_op_2_20_port
                           , Z(19) => sum_op_2_19_port, Z(18) => 
                           sum_op_2_18_port, Z(17) => sum_op_2_17_port, Z(16) 
                           => sum_op_2_16_port, Z(15) => sum_op_2_15_port, 
                           Z(14) => sum_op_2_14_port, Z(13) => sum_op_2_13_port
                           , Z(12) => sum_op_2_12_port, Z(11) => 
                           sum_op_2_11_port, Z(10) => sum_op_2_10_port, Z(9) =>
                           sum_op_2_9_port, Z(8) => sum_op_2_8_port, Z(7) => 
                           sum_op_2_7_port, Z(6) => sum_op_2_6_port, Z(5) => 
                           sum_op_2_5_port, Z(4) => sum_op_2_4_port, Z(3) => 
                           sum_op_2_3_port, Z(2) => sum_op_2_2_port, Z(1) => 
                           sum_op_2_1_port, Z(0) => sum_op_2_0_port);
   mux_i_3 : mux5to1_numBit32_5 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => n52, IN2(30) => n52, 
                           IN2(29) => n50, IN2(28) => n53, IN2(27) => n53, 
                           IN2(26) => n53, IN2(25) => n53, IN2(24) => n53, 
                           IN2(23) => n53, IN2(22) => n53, IN2(21) => n53, 
                           IN2(20) => A(14), IN2(19) => A(13), IN2(18) => A(12)
                           , IN2(17) => A(11), IN2(16) => A(10), IN2(15) => 
                           A(9), IN2(14) => A(8), IN2(13) => A(7), IN2(12) => 
                           A(6), IN2(11) => A(5), IN2(10) => A(4), IN2(9) => 
                           A(3), IN2(8) => A(2), IN2(7) => A(1), IN2(6) => A(0)
                           , IN2(5) => X_Logic0_port, IN2(4) => X_Logic0_port, 
                           IN2(3) => X_Logic0_port, IN2(2) => X_Logic0_port, 
                           IN2(1) => X_Logic0_port, IN2(0) => X_Logic0_port, 
                           IN3(31) => n31, IN3(30) => n35, IN3(29) => n32, 
                           IN3(28) => n35, IN3(27) => n32, IN3(26) => n36, 
                           IN3(25) => n33, IN3(24) => n34, IN3(23) => n33, 
                           IN3(22) => n34, IN3(21) => A_minus_15_port, IN3(20) 
                           => n2, IN3(19) => n4, IN3(18) => n6, IN3(17) => n8, 
                           IN3(16) => n10, IN3(15) => n12, IN3(14) => n14, 
                           IN3(13) => n16, IN3(12) => n18, IN3(11) => n20, 
                           IN3(10) => n22, IN3(9) => n24, IN3(8) => n26, IN3(7)
                           => n28, IN3(6) => A_minus_0_port, IN3(5) => 
                           X_Logic0_port, IN3(4) => X_Logic0_port, IN3(3) => 
                           X_Logic0_port, IN3(2) => X_Logic0_port, IN3(1) => 
                           X_Logic0_port, IN3(0) => X_Logic0_port, IN4(31) => 
                           n45, IN4(30) => n45, IN4(29) => n45, IN4(28) => n45,
                           IN4(27) => n45, IN4(26) => n45, IN4(25) => n45, 
                           IN4(24) => n45, IN4(23) => n45, IN4(22) => n45, 
                           IN4(21) => A(14), IN4(20) => A(13), IN4(19) => A(12)
                           , IN4(18) => A(11), IN4(17) => A(10), IN4(16) => 
                           A(9), IN4(15) => A(8), IN4(14) => A(7), IN4(13) => 
                           A(6), IN4(12) => A(5), IN4(11) => A(4), IN4(10) => 
                           A(3), IN4(9) => A(2), IN4(8) => A(1), IN4(7) => A(0)
                           , IN4(6) => X_Logic0_port, IN4(5) => X_Logic0_port, 
                           IN4(4) => X_Logic0_port, IN4(3) => X_Logic0_port, 
                           IN4(2) => X_Logic0_port, IN4(1) => X_Logic0_port, 
                           IN4(0) => X_Logic0_port, IN5(31) => n40, IN5(30) => 
                           n40, IN5(29) => n39, IN5(28) => n39, IN5(27) => n37,
                           IN5(26) => n38, IN5(25) => n38, IN5(24) => n37, 
                           IN5(23) => n38, IN5(22) => A_minus_15_port, IN5(21) 
                           => n2, IN5(20) => n4, IN5(19) => n6, IN5(18) => n8, 
                           IN5(17) => n10, IN5(16) => n12, IN5(15) => n14, 
                           IN5(14) => n16, IN5(13) => n18, IN5(12) => n20, 
                           IN5(11) => n22, IN5(10) => n24, IN5(9) => n26, 
                           IN5(8) => n28, IN5(7) => A_minus_0_port, IN5(6) => 
                           X_Logic0_port, IN5(5) => X_Logic0_port, IN5(4) => 
                           X_Logic0_port, IN5(3) => X_Logic0_port, IN5(2) => 
                           X_Logic0_port, IN5(1) => X_Logic0_port, IN5(0) => 
                           X_Logic0_port, SEL_in(2) => encoder_out_11_port, 
                           SEL_in(1) => encoder_out_10_port, SEL_in(0) => 
                           encoder_out_9_port, Z(31) => sum_op_3_31_port, Z(30)
                           => sum_op_3_30_port, Z(29) => sum_op_3_29_port, 
                           Z(28) => sum_op_3_28_port, Z(27) => sum_op_3_27_port
                           , Z(26) => sum_op_3_26_port, Z(25) => 
                           sum_op_3_25_port, Z(24) => sum_op_3_24_port, Z(23) 
                           => sum_op_3_23_port, Z(22) => sum_op_3_22_port, 
                           Z(21) => sum_op_3_21_port, Z(20) => sum_op_3_20_port
                           , Z(19) => sum_op_3_19_port, Z(18) => 
                           sum_op_3_18_port, Z(17) => sum_op_3_17_port, Z(16) 
                           => sum_op_3_16_port, Z(15) => sum_op_3_15_port, 
                           Z(14) => sum_op_3_14_port, Z(13) => sum_op_3_13_port
                           , Z(12) => sum_op_3_12_port, Z(11) => 
                           sum_op_3_11_port, Z(10) => sum_op_3_10_port, Z(9) =>
                           sum_op_3_9_port, Z(8) => sum_op_3_8_port, Z(7) => 
                           sum_op_3_7_port, Z(6) => sum_op_3_6_port, Z(5) => 
                           sum_op_3_5_port, Z(4) => sum_op_3_4_port, Z(3) => 
                           sum_op_3_3_port, Z(2) => sum_op_3_2_port, Z(1) => 
                           sum_op_3_1_port, Z(0) => sum_op_3_0_port);
   mux_i_4 : mux5to1_numBit32_4 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => n52, IN2(30) => n52, 
                           IN2(29) => n52, IN2(28) => n52, IN2(27) => n52, 
                           IN2(26) => n52, IN2(25) => n52, IN2(24) => n52, 
                           IN2(23) => n52, IN2(22) => A(14), IN2(21) => A(13), 
                           IN2(20) => A(12), IN2(19) => A(11), IN2(18) => A(10)
                           , IN2(17) => A(9), IN2(16) => A(8), IN2(15) => A(7),
                           IN2(14) => A(6), IN2(13) => A(5), IN2(12) => A(4), 
                           IN2(11) => A(3), IN2(10) => A(2), IN2(9) => A(1), 
                           IN2(8) => A(0), IN2(7) => X_Logic0_port, IN2(6) => 
                           X_Logic0_port, IN2(5) => X_Logic0_port, IN2(4) => 
                           X_Logic0_port, IN2(3) => X_Logic0_port, IN2(2) => 
                           X_Logic0_port, IN2(1) => X_Logic0_port, IN2(0) => 
                           X_Logic0_port, IN3(31) => n31, IN3(30) => n36, 
                           IN3(29) => n32, IN3(28) => n36, IN3(27) => n33, 
                           IN3(26) => n34, IN3(25) => n33, IN3(24) => n34, 
                           IN3(23) => A_minus_15_port, IN3(22) => n2, IN3(21) 
                           => n4, IN3(20) => n6, IN3(19) => n8, IN3(18) => n10,
                           IN3(17) => n12, IN3(16) => n14, IN3(15) => n16, 
                           IN3(14) => n18, IN3(13) => n20, IN3(12) => n22, 
                           IN3(11) => n24, IN3(10) => n26, IN3(9) => n28, 
                           IN3(8) => A_minus_0_port, IN3(7) => X_Logic0_port, 
                           IN3(6) => X_Logic0_port, IN3(5) => X_Logic0_port, 
                           IN3(4) => X_Logic0_port, IN3(3) => X_Logic0_port, 
                           IN3(2) => X_Logic0_port, IN3(1) => X_Logic0_port, 
                           IN3(0) => X_Logic0_port, IN4(31) => n44, IN4(30) => 
                           n44, IN4(29) => n44, IN4(28) => n44, IN4(27) => n44,
                           IN4(26) => n44, IN4(25) => n44, IN4(24) => n44, 
                           IN4(23) => A(14), IN4(22) => A(13), IN4(21) => A(12)
                           , IN4(20) => A(11), IN4(19) => A(10), IN4(18) => 
                           A(9), IN4(17) => A(8), IN4(16) => A(7), IN4(15) => 
                           A(6), IN4(14) => A(5), IN4(13) => A(4), IN4(12) => 
                           A(3), IN4(11) => A(2), IN4(10) => A(1), IN4(9) => 
                           A(0), IN4(8) => X_Logic0_port, IN4(7) => 
                           X_Logic0_port, IN4(6) => X_Logic0_port, IN4(5) => 
                           X_Logic0_port, IN4(4) => X_Logic0_port, IN4(3) => 
                           X_Logic0_port, IN4(2) => X_Logic0_port, IN4(1) => 
                           X_Logic0_port, IN4(0) => X_Logic0_port, IN5(31) => 
                           n39, IN5(30) => n39, IN5(29) => n38, IN5(28) => n41,
                           IN5(27) => n37, IN5(26) => n38, IN5(25) => n39, 
                           IN5(24) => A_minus_15_port, IN5(23) => n2, IN5(22) 
                           => n4, IN5(21) => n6, IN5(20) => n8, IN5(19) => n10,
                           IN5(18) => n12, IN5(17) => n14, IN5(16) => n16, 
                           IN5(15) => n18, IN5(14) => n20, IN5(13) => n22, 
                           IN5(12) => n24, IN5(11) => n26, IN5(10) => n28, 
                           IN5(9) => A_minus_0_port, IN5(8) => X_Logic0_port, 
                           IN5(7) => X_Logic0_port, IN5(6) => X_Logic0_port, 
                           IN5(5) => X_Logic0_port, IN5(4) => X_Logic0_port, 
                           IN5(3) => X_Logic0_port, IN5(2) => X_Logic0_port, 
                           IN5(1) => X_Logic0_port, IN5(0) => X_Logic0_port, 
                           SEL_in(2) => encoder_out_14_port, SEL_in(1) => 
                           encoder_out_13_port, SEL_in(0) => 
                           encoder_out_12_port, Z(31) => sum_op_4_31_port, 
                           Z(30) => sum_op_4_30_port, Z(29) => sum_op_4_29_port
                           , Z(28) => sum_op_4_28_port, Z(27) => 
                           sum_op_4_27_port, Z(26) => sum_op_4_26_port, Z(25) 
                           => sum_op_4_25_port, Z(24) => sum_op_4_24_port, 
                           Z(23) => sum_op_4_23_port, Z(22) => sum_op_4_22_port
                           , Z(21) => sum_op_4_21_port, Z(20) => 
                           sum_op_4_20_port, Z(19) => sum_op_4_19_port, Z(18) 
                           => sum_op_4_18_port, Z(17) => sum_op_4_17_port, 
                           Z(16) => sum_op_4_16_port, Z(15) => sum_op_4_15_port
                           , Z(14) => sum_op_4_14_port, Z(13) => 
                           sum_op_4_13_port, Z(12) => sum_op_4_12_port, Z(11) 
                           => sum_op_4_11_port, Z(10) => sum_op_4_10_port, Z(9)
                           => sum_op_4_9_port, Z(8) => sum_op_4_8_port, Z(7) =>
                           sum_op_4_7_port, Z(6) => sum_op_4_6_port, Z(5) => 
                           sum_op_4_5_port, Z(4) => sum_op_4_4_port, Z(3) => 
                           sum_op_4_3_port, Z(2) => sum_op_4_2_port, Z(1) => 
                           sum_op_4_1_port, Z(0) => sum_op_4_0_port);
   mux_i_5 : mux5to1_numBit32_3 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => n51, IN2(30) => n51, 
                           IN2(29) => n51, IN2(28) => n51, IN2(27) => n51, 
                           IN2(26) => n51, IN2(25) => n51, IN2(24) => A(14), 
                           IN2(23) => A(13), IN2(22) => A(12), IN2(21) => A(11)
                           , IN2(20) => A(10), IN2(19) => A(9), IN2(18) => A(8)
                           , IN2(17) => A(7), IN2(16) => A(6), IN2(15) => A(5),
                           IN2(14) => A(4), IN2(13) => A(3), IN2(12) => A(2), 
                           IN2(11) => A(1), IN2(10) => A(0), IN2(9) => 
                           X_Logic0_port, IN2(8) => X_Logic0_port, IN2(7) => 
                           X_Logic0_port, IN2(6) => X_Logic0_port, IN2(5) => 
                           X_Logic0_port, IN2(4) => X_Logic0_port, IN2(3) => 
                           X_Logic0_port, IN2(2) => X_Logic0_port, IN2(1) => 
                           X_Logic0_port, IN2(0) => X_Logic0_port, IN3(31) => 
                           n32, IN3(30) => n35, IN3(29) => n32, IN3(28) => n35,
                           IN3(27) => n33, IN3(26) => n34, IN3(25) => 
                           A_minus_15_port, IN3(24) => n2, IN3(23) => n4, 
                           IN3(22) => n6, IN3(21) => n8, IN3(20) => n10, 
                           IN3(19) => n12, IN3(18) => n14, IN3(17) => n16, 
                           IN3(16) => n18, IN3(15) => n20, IN3(14) => n22, 
                           IN3(13) => n24, IN3(12) => n26, IN3(11) => n28, 
                           IN3(10) => A_minus_0_port, IN3(9) => X_Logic0_port, 
                           IN3(8) => X_Logic0_port, IN3(7) => X_Logic0_port, 
                           IN3(6) => X_Logic0_port, IN3(5) => X_Logic0_port, 
                           IN3(4) => X_Logic0_port, IN3(3) => X_Logic0_port, 
                           IN3(2) => X_Logic0_port, IN3(1) => X_Logic0_port, 
                           IN3(0) => X_Logic0_port, IN4(31) => n43, IN4(30) => 
                           n43, IN4(29) => n44, IN4(28) => n44, IN4(27) => n44,
                           IN4(26) => n44, IN4(25) => A(14), IN4(24) => A(13), 
                           IN4(23) => A(12), IN4(22) => A(11), IN4(21) => A(10)
                           , IN4(20) => A(9), IN4(19) => A(8), IN4(18) => A(7),
                           IN4(17) => A(6), IN4(16) => A(5), IN4(15) => A(4), 
                           IN4(14) => A(3), IN4(13) => A(2), IN4(12) => A(1), 
                           IN4(11) => A(0), IN4(10) => X_Logic0_port, IN4(9) =>
                           X_Logic0_port, IN4(8) => X_Logic0_port, IN4(7) => 
                           X_Logic0_port, IN4(6) => X_Logic0_port, IN4(5) => 
                           X_Logic0_port, IN4(4) => X_Logic0_port, IN4(3) => 
                           X_Logic0_port, IN4(2) => X_Logic0_port, IN4(1) => 
                           X_Logic0_port, IN4(0) => X_Logic0_port, IN5(31) => 
                           n40, IN5(30) => n39, IN5(29) => n37, IN5(28) => n38,
                           IN5(27) => n37, IN5(26) => A_minus_15_port, IN5(25) 
                           => n2, IN5(24) => n4, IN5(23) => n6, IN5(22) => n8, 
                           IN5(21) => n10, IN5(20) => n12, IN5(19) => n14, 
                           IN5(18) => n16, IN5(17) => n18, IN5(16) => n20, 
                           IN5(15) => n22, IN5(14) => n24, IN5(13) => n26, 
                           IN5(12) => n28, IN5(11) => A_minus_0_port, IN5(10) 
                           => X_Logic0_port, IN5(9) => X_Logic0_port, IN5(8) =>
                           X_Logic0_port, IN5(7) => X_Logic0_port, IN5(6) => 
                           X_Logic0_port, IN5(5) => X_Logic0_port, IN5(4) => 
                           X_Logic0_port, IN5(3) => X_Logic0_port, IN5(2) => 
                           X_Logic0_port, IN5(1) => X_Logic0_port, IN5(0) => 
                           X_Logic0_port, SEL_in(2) => encoder_out_17_port, 
                           SEL_in(1) => encoder_out_16_port, SEL_in(0) => 
                           encoder_out_15_port, Z(31) => sum_op_5_31_port, 
                           Z(30) => sum_op_5_30_port, Z(29) => sum_op_5_29_port
                           , Z(28) => sum_op_5_28_port, Z(27) => 
                           sum_op_5_27_port, Z(26) => sum_op_5_26_port, Z(25) 
                           => sum_op_5_25_port, Z(24) => sum_op_5_24_port, 
                           Z(23) => sum_op_5_23_port, Z(22) => sum_op_5_22_port
                           , Z(21) => sum_op_5_21_port, Z(20) => 
                           sum_op_5_20_port, Z(19) => sum_op_5_19_port, Z(18) 
                           => sum_op_5_18_port, Z(17) => sum_op_5_17_port, 
                           Z(16) => sum_op_5_16_port, Z(15) => sum_op_5_15_port
                           , Z(14) => sum_op_5_14_port, Z(13) => 
                           sum_op_5_13_port, Z(12) => sum_op_5_12_port, Z(11) 
                           => sum_op_5_11_port, Z(10) => sum_op_5_10_port, Z(9)
                           => sum_op_5_9_port, Z(8) => sum_op_5_8_port, Z(7) =>
                           sum_op_5_7_port, Z(6) => sum_op_5_6_port, Z(5) => 
                           sum_op_5_5_port, Z(4) => sum_op_5_4_port, Z(3) => 
                           sum_op_5_3_port, Z(2) => sum_op_5_2_port, Z(1) => 
                           sum_op_5_1_port, Z(0) => sum_op_5_0_port);
   mux_i_6 : mux5to1_numBit32_2 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => n50, IN2(30) => n50, 
                           IN2(29) => n50, IN2(28) => n50, IN2(27) => n50, 
                           IN2(26) => A(14), IN2(25) => A(13), IN2(24) => A(12)
                           , IN2(23) => A(11), IN2(22) => A(10), IN2(21) => 
                           A(9), IN2(20) => A(8), IN2(19) => A(7), IN2(18) => 
                           A(6), IN2(17) => A(5), IN2(16) => A(4), IN2(15) => 
                           A(3), IN2(14) => A(2), IN2(13) => A(1), IN2(12) => 
                           A(0), IN2(11) => X_Logic0_port, IN2(10) => 
                           X_Logic0_port, IN2(9) => X_Logic0_port, IN2(8) => 
                           X_Logic0_port, IN2(7) => X_Logic0_port, IN2(6) => 
                           X_Logic0_port, IN2(5) => X_Logic0_port, IN2(4) => 
                           X_Logic0_port, IN2(3) => X_Logic0_port, IN2(2) => 
                           X_Logic0_port, IN2(1) => X_Logic0_port, IN2(0) => 
                           X_Logic0_port, IN3(31) => n32, IN3(30) => n35, 
                           IN3(29) => n33, IN3(28) => n34, IN3(27) => 
                           A_minus_15_port, IN3(26) => n2, IN3(25) => n4, 
                           IN3(24) => n6, IN3(23) => n8, IN3(22) => n10, 
                           IN3(21) => n12, IN3(20) => n14, IN3(19) => n16, 
                           IN3(18) => n18, IN3(17) => n20, IN3(16) => n22, 
                           IN3(15) => n24, IN3(14) => n26, IN3(13) => n28, 
                           IN3(12) => A_minus_0_port, IN3(11) => X_Logic0_port,
                           IN3(10) => X_Logic0_port, IN3(9) => X_Logic0_port, 
                           IN3(8) => X_Logic0_port, IN3(7) => X_Logic0_port, 
                           IN3(6) => X_Logic0_port, IN3(5) => X_Logic0_port, 
                           IN3(4) => X_Logic0_port, IN3(3) => X_Logic0_port, 
                           IN3(2) => X_Logic0_port, IN3(1) => X_Logic0_port, 
                           IN3(0) => X_Logic0_port, IN4(31) => n43, IN4(30) => 
                           n43, IN4(29) => n43, IN4(28) => n43, IN4(27) => 
                           A(14), IN4(26) => A(13), IN4(25) => A(12), IN4(24) 
                           => A(11), IN4(23) => A(10), IN4(22) => A(9), IN4(21)
                           => A(8), IN4(20) => A(7), IN4(19) => A(6), IN4(18) 
                           => A(5), IN4(17) => A(4), IN4(16) => A(3), IN4(15) 
                           => A(2), IN4(14) => A(1), IN4(13) => A(0), IN4(12) 
                           => X_Logic0_port, IN4(11) => X_Logic0_port, IN4(10) 
                           => X_Logic0_port, IN4(9) => X_Logic0_port, IN4(8) =>
                           X_Logic0_port, IN4(7) => X_Logic0_port, IN4(6) => 
                           X_Logic0_port, IN4(5) => X_Logic0_port, IN4(4) => 
                           X_Logic0_port, IN4(3) => X_Logic0_port, IN4(2) => 
                           X_Logic0_port, IN4(1) => X_Logic0_port, IN4(0) => 
                           X_Logic0_port, IN5(31) => n37, IN5(30) => n38, 
                           IN5(29) => n37, IN5(28) => A_minus_15_port, IN5(27) 
                           => n2, IN5(26) => n4, IN5(25) => n6, IN5(24) => n8, 
                           IN5(23) => n10, IN5(22) => n12, IN5(21) => n14, 
                           IN5(20) => n16, IN5(19) => n18, IN5(18) => n20, 
                           IN5(17) => n22, IN5(16) => n24, IN5(15) => n26, 
                           IN5(14) => n28, IN5(13) => A_minus_0_port, IN5(12) 
                           => X_Logic0_port, IN5(11) => X_Logic0_port, IN5(10) 
                           => X_Logic0_port, IN5(9) => X_Logic0_port, IN5(8) =>
                           X_Logic0_port, IN5(7) => X_Logic0_port, IN5(6) => 
                           X_Logic0_port, IN5(5) => X_Logic0_port, IN5(4) => 
                           X_Logic0_port, IN5(3) => X_Logic0_port, IN5(2) => 
                           X_Logic0_port, IN5(1) => X_Logic0_port, IN5(0) => 
                           X_Logic0_port, SEL_in(2) => encoder_out_20_port, 
                           SEL_in(1) => encoder_out_19_port, SEL_in(0) => 
                           encoder_out_18_port, Z(31) => sum_op_6_31_port, 
                           Z(30) => sum_op_6_30_port, Z(29) => sum_op_6_29_port
                           , Z(28) => sum_op_6_28_port, Z(27) => 
                           sum_op_6_27_port, Z(26) => sum_op_6_26_port, Z(25) 
                           => sum_op_6_25_port, Z(24) => sum_op_6_24_port, 
                           Z(23) => sum_op_6_23_port, Z(22) => sum_op_6_22_port
                           , Z(21) => sum_op_6_21_port, Z(20) => 
                           sum_op_6_20_port, Z(19) => sum_op_6_19_port, Z(18) 
                           => sum_op_6_18_port, Z(17) => sum_op_6_17_port, 
                           Z(16) => sum_op_6_16_port, Z(15) => sum_op_6_15_port
                           , Z(14) => sum_op_6_14_port, Z(13) => 
                           sum_op_6_13_port, Z(12) => sum_op_6_12_port, Z(11) 
                           => sum_op_6_11_port, Z(10) => sum_op_6_10_port, Z(9)
                           => sum_op_6_9_port, Z(8) => sum_op_6_8_port, Z(7) =>
                           sum_op_6_7_port, Z(6) => sum_op_6_6_port, Z(5) => 
                           sum_op_6_5_port, Z(4) => sum_op_6_4_port, Z(3) => 
                           sum_op_6_3_port, Z(2) => sum_op_6_2_port, Z(1) => 
                           sum_op_6_1_port, Z(0) => sum_op_6_0_port);
   mux_i_7 : mux5to1_numBit32_1 port map( IN1(31) => X_Logic0_port, IN1(30) => 
                           X_Logic0_port, IN1(29) => X_Logic0_port, IN1(28) => 
                           X_Logic0_port, IN1(27) => X_Logic0_port, IN1(26) => 
                           X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) => 
                           X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) => 
                           X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) => 
                           X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(31) => n49, IN2(30) => n49, 
                           IN2(29) => n50, IN2(28) => A(14), IN2(27) => A(13), 
                           IN2(26) => A(12), IN2(25) => A(11), IN2(24) => A(10)
                           , IN2(23) => A(9), IN2(22) => A(8), IN2(21) => A(7),
                           IN2(20) => A(6), IN2(19) => A(5), IN2(18) => A(4), 
                           IN2(17) => A(3), IN2(16) => A(2), IN2(15) => A(1), 
                           IN2(14) => A(0), IN2(13) => X_Logic0_port, IN2(12) 
                           => X_Logic0_port, IN2(11) => X_Logic0_port, IN2(10) 
                           => X_Logic0_port, IN2(9) => X_Logic0_port, IN2(8) =>
                           X_Logic0_port, IN2(7) => X_Logic0_port, IN2(6) => 
                           X_Logic0_port, IN2(5) => X_Logic0_port, IN2(4) => 
                           X_Logic0_port, IN2(3) => X_Logic0_port, IN2(2) => 
                           X_Logic0_port, IN2(1) => X_Logic0_port, IN2(0) => 
                           X_Logic0_port, IN3(31) => n33, IN3(30) => n34, 
                           IN3(29) => A_minus_15_port, IN3(28) => n2, IN3(27) 
                           => n4, IN3(26) => n6, IN3(25) => n8, IN3(24) => n10,
                           IN3(23) => n12, IN3(22) => n14, IN3(21) => n16, 
                           IN3(20) => n18, IN3(19) => n20, IN3(18) => n22, 
                           IN3(17) => n24, IN3(16) => n26, IN3(15) => n28, 
                           IN3(14) => A_minus_0_port, IN3(13) => X_Logic0_port,
                           IN3(12) => X_Logic0_port, IN3(11) => X_Logic0_port, 
                           IN3(10) => X_Logic0_port, IN3(9) => X_Logic0_port, 
                           IN3(8) => X_Logic0_port, IN3(7) => X_Logic0_port, 
                           IN3(6) => X_Logic0_port, IN3(5) => X_Logic0_port, 
                           IN3(4) => X_Logic0_port, IN3(3) => X_Logic0_port, 
                           IN3(2) => X_Logic0_port, IN3(1) => X_Logic0_port, 
                           IN3(0) => X_Logic0_port, IN4(31) => n43, IN4(30) => 
                           n45, IN4(29) => A(14), IN4(28) => A(13), IN4(27) => 
                           A(12), IN4(26) => A(11), IN4(25) => A(10), IN4(24) 
                           => A(9), IN4(23) => A(8), IN4(22) => A(7), IN4(21) 
                           => A(6), IN4(20) => A(5), IN4(19) => A(4), IN4(18) 
                           => A(3), IN4(17) => A(2), IN4(16) => A(1), IN4(15) 
                           => A(0), IN4(14) => X_Logic0_port, IN4(13) => 
                           X_Logic0_port, IN4(12) => X_Logic0_port, IN4(11) => 
                           X_Logic0_port, IN4(10) => X_Logic0_port, IN4(9) => 
                           X_Logic0_port, IN4(8) => X_Logic0_port, IN4(7) => 
                           X_Logic0_port, IN4(6) => X_Logic0_port, IN4(5) => 
                           X_Logic0_port, IN4(4) => X_Logic0_port, IN4(3) => 
                           X_Logic0_port, IN4(2) => X_Logic0_port, IN4(1) => 
                           X_Logic0_port, IN4(0) => X_Logic0_port, IN5(31) => 
                           n37, IN5(30) => A_minus_15_port, IN5(29) => n2, 
                           IN5(28) => n4, IN5(27) => n6, IN5(26) => n8, IN5(25)
                           => n10, IN5(24) => n12, IN5(23) => n14, IN5(22) => 
                           n16, IN5(21) => n18, IN5(20) => n20, IN5(19) => n22,
                           IN5(18) => n24, IN5(17) => n26, IN5(16) => n28, 
                           IN5(15) => A_minus_0_port, IN5(14) => X_Logic0_port,
                           IN5(13) => X_Logic0_port, IN5(12) => X_Logic0_port, 
                           IN5(11) => X_Logic0_port, IN5(10) => X_Logic0_port, 
                           IN5(9) => X_Logic0_port, IN5(8) => X_Logic0_port, 
                           IN5(7) => X_Logic0_port, IN5(6) => X_Logic0_port, 
                           IN5(5) => X_Logic0_port, IN5(4) => X_Logic0_port, 
                           IN5(3) => X_Logic0_port, IN5(2) => X_Logic0_port, 
                           IN5(1) => X_Logic0_port, IN5(0) => X_Logic0_port, 
                           SEL_in(2) => encoder_out_23_port, SEL_in(1) => 
                           encoder_out_22_port, SEL_in(0) => 
                           encoder_out_21_port, Z(31) => sum_op_7_31_port, 
                           Z(30) => sum_op_7_30_port, Z(29) => sum_op_7_29_port
                           , Z(28) => sum_op_7_28_port, Z(27) => 
                           sum_op_7_27_port, Z(26) => sum_op_7_26_port, Z(25) 
                           => sum_op_7_25_port, Z(24) => sum_op_7_24_port, 
                           Z(23) => sum_op_7_23_port, Z(22) => sum_op_7_22_port
                           , Z(21) => sum_op_7_21_port, Z(20) => 
                           sum_op_7_20_port, Z(19) => sum_op_7_19_port, Z(18) 
                           => sum_op_7_18_port, Z(17) => sum_op_7_17_port, 
                           Z(16) => sum_op_7_16_port, Z(15) => sum_op_7_15_port
                           , Z(14) => sum_op_7_14_port, Z(13) => 
                           sum_op_7_13_port, Z(12) => sum_op_7_12_port, Z(11) 
                           => sum_op_7_11_port, Z(10) => sum_op_7_10_port, Z(9)
                           => sum_op_7_9_port, Z(8) => sum_op_7_8_port, Z(7) =>
                           sum_op_7_7_port, Z(6) => sum_op_7_6_port, Z(5) => 
                           sum_op_7_5_port, Z(4) => sum_op_7_4_port, Z(3) => 
                           sum_op_7_3_port, Z(2) => sum_op_7_2_port, Z(1) => 
                           sum_op_7_1_port, Z(0) => sum_op_7_0_port);
   rca0_0 : rca_bhv_numBit32_0 port map( A(31) => sum_op_0_31_port, A(30) => 
                           sum_op_0_30_port, A(29) => sum_op_0_29_port, A(28) 
                           => sum_op_0_28_port, A(27) => sum_op_0_27_port, 
                           A(26) => sum_op_0_26_port, A(25) => sum_op_0_25_port
                           , A(24) => sum_op_0_24_port, A(23) => 
                           sum_op_0_23_port, A(22) => sum_op_0_22_port, A(21) 
                           => sum_op_0_21_port, A(20) => sum_op_0_20_port, 
                           A(19) => sum_op_0_19_port, A(18) => sum_op_0_18_port
                           , A(17) => sum_op_0_17_port, A(16) => 
                           sum_op_0_16_port, A(15) => sum_op_0_15_port, A(14) 
                           => sum_op_0_14_port, A(13) => sum_op_0_13_port, 
                           A(12) => sum_op_0_12_port, A(11) => sum_op_0_11_port
                           , A(10) => sum_op_0_10_port, A(9) => sum_op_0_9_port
                           , A(8) => sum_op_0_8_port, A(7) => sum_op_0_7_port, 
                           A(6) => sum_op_0_6_port, A(5) => sum_op_0_5_port, 
                           A(4) => sum_op_0_4_port, A(3) => sum_op_0_3_port, 
                           A(2) => sum_op_0_2_port, A(1) => sum_op_0_1_port, 
                           A(0) => sum_op_0_0_port, B(31) => sum_op_1_31_port, 
                           B(30) => sum_op_1_30_port, B(29) => sum_op_1_29_port
                           , B(28) => sum_op_1_28_port, B(27) => 
                           sum_op_1_27_port, B(26) => sum_op_1_26_port, B(25) 
                           => sum_op_1_25_port, B(24) => sum_op_1_24_port, 
                           B(23) => sum_op_1_23_port, B(22) => sum_op_1_22_port
                           , B(21) => sum_op_1_21_port, B(20) => 
                           sum_op_1_20_port, B(19) => sum_op_1_19_port, B(18) 
                           => sum_op_1_18_port, B(17) => sum_op_1_17_port, 
                           B(16) => sum_op_1_16_port, B(15) => sum_op_1_15_port
                           , B(14) => sum_op_1_14_port, B(13) => 
                           sum_op_1_13_port, B(12) => sum_op_1_12_port, B(11) 
                           => sum_op_1_11_port, B(10) => sum_op_1_10_port, B(9)
                           => sum_op_1_9_port, B(8) => sum_op_1_8_port, B(7) =>
                           sum_op_1_7_port, B(6) => sum_op_1_6_port, B(5) => 
                           sum_op_1_5_port, B(4) => sum_op_1_4_port, B(3) => 
                           sum_op_1_3_port, B(2) => sum_op_1_2_port, B(1) => 
                           sum_op_1_1_port, B(0) => sum_op_1_0_port, Ci => 
                           X_Logic0_port, S(31) => rca_out_0_31_port, S(30) => 
                           rca_out_0_30_port, S(29) => rca_out_0_29_port, S(28)
                           => rca_out_0_28_port, S(27) => rca_out_0_27_port, 
                           S(26) => rca_out_0_26_port, S(25) => 
                           rca_out_0_25_port, S(24) => rca_out_0_24_port, S(23)
                           => rca_out_0_23_port, S(22) => rca_out_0_22_port, 
                           S(21) => rca_out_0_21_port, S(20) => 
                           rca_out_0_20_port, S(19) => rca_out_0_19_port, S(18)
                           => rca_out_0_18_port, S(17) => rca_out_0_17_port, 
                           S(16) => rca_out_0_16_port, S(15) => 
                           rca_out_0_15_port, S(14) => rca_out_0_14_port, S(13)
                           => rca_out_0_13_port, S(12) => rca_out_0_12_port, 
                           S(11) => rca_out_0_11_port, S(10) => 
                           rca_out_0_10_port, S(9) => rca_out_0_9_port, S(8) =>
                           rca_out_0_8_port, S(7) => rca_out_0_7_port, S(6) => 
                           rca_out_0_6_port, S(5) => rca_out_0_5_port, S(4) => 
                           rca_out_0_4_port, S(3) => rca_out_0_3_port, S(2) => 
                           rca_out_0_2_port, S(1) => rca_out_0_1_port, S(0) => 
                           rca_out_0_0_port, Co => n_1159);
   rca_i_1 : rca_bhv_numBit32_6 port map( A(31) => rca_out_0_31_port, A(30) => 
                           rca_out_0_30_port, A(29) => rca_out_0_29_port, A(28)
                           => rca_out_0_28_port, A(27) => rca_out_0_27_port, 
                           A(26) => rca_out_0_26_port, A(25) => 
                           rca_out_0_25_port, A(24) => rca_out_0_24_port, A(23)
                           => rca_out_0_23_port, A(22) => rca_out_0_22_port, 
                           A(21) => rca_out_0_21_port, A(20) => 
                           rca_out_0_20_port, A(19) => rca_out_0_19_port, A(18)
                           => rca_out_0_18_port, A(17) => rca_out_0_17_port, 
                           A(16) => rca_out_0_16_port, A(15) => 
                           rca_out_0_15_port, A(14) => rca_out_0_14_port, A(13)
                           => rca_out_0_13_port, A(12) => rca_out_0_12_port, 
                           A(11) => rca_out_0_11_port, A(10) => 
                           rca_out_0_10_port, A(9) => rca_out_0_9_port, A(8) =>
                           rca_out_0_8_port, A(7) => rca_out_0_7_port, A(6) => 
                           rca_out_0_6_port, A(5) => rca_out_0_5_port, A(4) => 
                           rca_out_0_4_port, A(3) => rca_out_0_3_port, A(2) => 
                           rca_out_0_2_port, A(1) => rca_out_0_1_port, A(0) => 
                           rca_out_0_0_port, B(31) => sum_op_2_31_port, B(30) 
                           => sum_op_2_30_port, B(29) => sum_op_2_29_port, 
                           B(28) => sum_op_2_28_port, B(27) => sum_op_2_27_port
                           , B(26) => sum_op_2_26_port, B(25) => 
                           sum_op_2_25_port, B(24) => sum_op_2_24_port, B(23) 
                           => sum_op_2_23_port, B(22) => sum_op_2_22_port, 
                           B(21) => sum_op_2_21_port, B(20) => sum_op_2_20_port
                           , B(19) => sum_op_2_19_port, B(18) => 
                           sum_op_2_18_port, B(17) => sum_op_2_17_port, B(16) 
                           => sum_op_2_16_port, B(15) => sum_op_2_15_port, 
                           B(14) => sum_op_2_14_port, B(13) => sum_op_2_13_port
                           , B(12) => sum_op_2_12_port, B(11) => 
                           sum_op_2_11_port, B(10) => sum_op_2_10_port, B(9) =>
                           sum_op_2_9_port, B(8) => sum_op_2_8_port, B(7) => 
                           sum_op_2_7_port, B(6) => sum_op_2_6_port, B(5) => 
                           sum_op_2_5_port, B(4) => sum_op_2_4_port, B(3) => 
                           sum_op_2_3_port, B(2) => sum_op_2_2_port, B(1) => 
                           sum_op_2_1_port, B(0) => sum_op_2_0_port, Ci => 
                           X_Logic0_port, S(31) => rca_out_1_31_port, S(30) => 
                           rca_out_1_30_port, S(29) => rca_out_1_29_port, S(28)
                           => rca_out_1_28_port, S(27) => rca_out_1_27_port, 
                           S(26) => rca_out_1_26_port, S(25) => 
                           rca_out_1_25_port, S(24) => rca_out_1_24_port, S(23)
                           => rca_out_1_23_port, S(22) => rca_out_1_22_port, 
                           S(21) => rca_out_1_21_port, S(20) => 
                           rca_out_1_20_port, S(19) => rca_out_1_19_port, S(18)
                           => rca_out_1_18_port, S(17) => rca_out_1_17_port, 
                           S(16) => rca_out_1_16_port, S(15) => 
                           rca_out_1_15_port, S(14) => rca_out_1_14_port, S(13)
                           => rca_out_1_13_port, S(12) => rca_out_1_12_port, 
                           S(11) => rca_out_1_11_port, S(10) => 
                           rca_out_1_10_port, S(9) => rca_out_1_9_port, S(8) =>
                           rca_out_1_8_port, S(7) => rca_out_1_7_port, S(6) => 
                           rca_out_1_6_port, S(5) => rca_out_1_5_port, S(4) => 
                           rca_out_1_4_port, S(3) => rca_out_1_3_port, S(2) => 
                           rca_out_1_2_port, S(1) => rca_out_1_1_port, S(0) => 
                           rca_out_1_0_port, Co => n_1160);
   rca_i_2 : rca_bhv_numBit32_5 port map( A(31) => rca_out_1_31_port, A(30) => 
                           rca_out_1_30_port, A(29) => rca_out_1_29_port, A(28)
                           => rca_out_1_28_port, A(27) => rca_out_1_27_port, 
                           A(26) => rca_out_1_26_port, A(25) => 
                           rca_out_1_25_port, A(24) => rca_out_1_24_port, A(23)
                           => rca_out_1_23_port, A(22) => rca_out_1_22_port, 
                           A(21) => rca_out_1_21_port, A(20) => 
                           rca_out_1_20_port, A(19) => rca_out_1_19_port, A(18)
                           => rca_out_1_18_port, A(17) => rca_out_1_17_port, 
                           A(16) => rca_out_1_16_port, A(15) => 
                           rca_out_1_15_port, A(14) => rca_out_1_14_port, A(13)
                           => rca_out_1_13_port, A(12) => rca_out_1_12_port, 
                           A(11) => rca_out_1_11_port, A(10) => 
                           rca_out_1_10_port, A(9) => rca_out_1_9_port, A(8) =>
                           rca_out_1_8_port, A(7) => rca_out_1_7_port, A(6) => 
                           rca_out_1_6_port, A(5) => rca_out_1_5_port, A(4) => 
                           rca_out_1_4_port, A(3) => rca_out_1_3_port, A(2) => 
                           rca_out_1_2_port, A(1) => rca_out_1_1_port, A(0) => 
                           rca_out_1_0_port, B(31) => sum_op_3_31_port, B(30) 
                           => sum_op_3_30_port, B(29) => sum_op_3_29_port, 
                           B(28) => sum_op_3_28_port, B(27) => sum_op_3_27_port
                           , B(26) => sum_op_3_26_port, B(25) => 
                           sum_op_3_25_port, B(24) => sum_op_3_24_port, B(23) 
                           => sum_op_3_23_port, B(22) => sum_op_3_22_port, 
                           B(21) => sum_op_3_21_port, B(20) => sum_op_3_20_port
                           , B(19) => sum_op_3_19_port, B(18) => 
                           sum_op_3_18_port, B(17) => sum_op_3_17_port, B(16) 
                           => sum_op_3_16_port, B(15) => sum_op_3_15_port, 
                           B(14) => sum_op_3_14_port, B(13) => sum_op_3_13_port
                           , B(12) => sum_op_3_12_port, B(11) => 
                           sum_op_3_11_port, B(10) => sum_op_3_10_port, B(9) =>
                           sum_op_3_9_port, B(8) => sum_op_3_8_port, B(7) => 
                           sum_op_3_7_port, B(6) => sum_op_3_6_port, B(5) => 
                           sum_op_3_5_port, B(4) => sum_op_3_4_port, B(3) => 
                           sum_op_3_3_port, B(2) => sum_op_3_2_port, B(1) => 
                           sum_op_3_1_port, B(0) => sum_op_3_0_port, Ci => 
                           X_Logic0_port, S(31) => rca_out_2_31_port, S(30) => 
                           rca_out_2_30_port, S(29) => rca_out_2_29_port, S(28)
                           => rca_out_2_28_port, S(27) => rca_out_2_27_port, 
                           S(26) => rca_out_2_26_port, S(25) => 
                           rca_out_2_25_port, S(24) => rca_out_2_24_port, S(23)
                           => rca_out_2_23_port, S(22) => rca_out_2_22_port, 
                           S(21) => rca_out_2_21_port, S(20) => 
                           rca_out_2_20_port, S(19) => rca_out_2_19_port, S(18)
                           => rca_out_2_18_port, S(17) => rca_out_2_17_port, 
                           S(16) => rca_out_2_16_port, S(15) => 
                           rca_out_2_15_port, S(14) => rca_out_2_14_port, S(13)
                           => rca_out_2_13_port, S(12) => rca_out_2_12_port, 
                           S(11) => rca_out_2_11_port, S(10) => 
                           rca_out_2_10_port, S(9) => rca_out_2_9_port, S(8) =>
                           rca_out_2_8_port, S(7) => rca_out_2_7_port, S(6) => 
                           rca_out_2_6_port, S(5) => rca_out_2_5_port, S(4) => 
                           rca_out_2_4_port, S(3) => rca_out_2_3_port, S(2) => 
                           rca_out_2_2_port, S(1) => rca_out_2_1_port, S(0) => 
                           rca_out_2_0_port, Co => n_1161);
   rca_i_3 : rca_bhv_numBit32_4 port map( A(31) => rca_out_2_31_port, A(30) => 
                           rca_out_2_30_port, A(29) => rca_out_2_29_port, A(28)
                           => rca_out_2_28_port, A(27) => rca_out_2_27_port, 
                           A(26) => rca_out_2_26_port, A(25) => 
                           rca_out_2_25_port, A(24) => rca_out_2_24_port, A(23)
                           => rca_out_2_23_port, A(22) => rca_out_2_22_port, 
                           A(21) => rca_out_2_21_port, A(20) => 
                           rca_out_2_20_port, A(19) => rca_out_2_19_port, A(18)
                           => rca_out_2_18_port, A(17) => rca_out_2_17_port, 
                           A(16) => rca_out_2_16_port, A(15) => 
                           rca_out_2_15_port, A(14) => rca_out_2_14_port, A(13)
                           => rca_out_2_13_port, A(12) => rca_out_2_12_port, 
                           A(11) => rca_out_2_11_port, A(10) => 
                           rca_out_2_10_port, A(9) => rca_out_2_9_port, A(8) =>
                           rca_out_2_8_port, A(7) => rca_out_2_7_port, A(6) => 
                           rca_out_2_6_port, A(5) => rca_out_2_5_port, A(4) => 
                           rca_out_2_4_port, A(3) => rca_out_2_3_port, A(2) => 
                           rca_out_2_2_port, A(1) => rca_out_2_1_port, A(0) => 
                           rca_out_2_0_port, B(31) => sum_op_4_31_port, B(30) 
                           => sum_op_4_30_port, B(29) => sum_op_4_29_port, 
                           B(28) => sum_op_4_28_port, B(27) => sum_op_4_27_port
                           , B(26) => sum_op_4_26_port, B(25) => 
                           sum_op_4_25_port, B(24) => sum_op_4_24_port, B(23) 
                           => sum_op_4_23_port, B(22) => sum_op_4_22_port, 
                           B(21) => sum_op_4_21_port, B(20) => sum_op_4_20_port
                           , B(19) => sum_op_4_19_port, B(18) => 
                           sum_op_4_18_port, B(17) => sum_op_4_17_port, B(16) 
                           => sum_op_4_16_port, B(15) => sum_op_4_15_port, 
                           B(14) => sum_op_4_14_port, B(13) => sum_op_4_13_port
                           , B(12) => sum_op_4_12_port, B(11) => 
                           sum_op_4_11_port, B(10) => sum_op_4_10_port, B(9) =>
                           sum_op_4_9_port, B(8) => sum_op_4_8_port, B(7) => 
                           sum_op_4_7_port, B(6) => sum_op_4_6_port, B(5) => 
                           sum_op_4_5_port, B(4) => sum_op_4_4_port, B(3) => 
                           sum_op_4_3_port, B(2) => sum_op_4_2_port, B(1) => 
                           sum_op_4_1_port, B(0) => sum_op_4_0_port, Ci => 
                           X_Logic0_port, S(31) => rca_out_3_31_port, S(30) => 
                           rca_out_3_30_port, S(29) => rca_out_3_29_port, S(28)
                           => rca_out_3_28_port, S(27) => rca_out_3_27_port, 
                           S(26) => rca_out_3_26_port, S(25) => 
                           rca_out_3_25_port, S(24) => rca_out_3_24_port, S(23)
                           => rca_out_3_23_port, S(22) => rca_out_3_22_port, 
                           S(21) => rca_out_3_21_port, S(20) => 
                           rca_out_3_20_port, S(19) => rca_out_3_19_port, S(18)
                           => rca_out_3_18_port, S(17) => rca_out_3_17_port, 
                           S(16) => rca_out_3_16_port, S(15) => 
                           rca_out_3_15_port, S(14) => rca_out_3_14_port, S(13)
                           => rca_out_3_13_port, S(12) => rca_out_3_12_port, 
                           S(11) => rca_out_3_11_port, S(10) => 
                           rca_out_3_10_port, S(9) => rca_out_3_9_port, S(8) =>
                           rca_out_3_8_port, S(7) => rca_out_3_7_port, S(6) => 
                           rca_out_3_6_port, S(5) => rca_out_3_5_port, S(4) => 
                           rca_out_3_4_port, S(3) => rca_out_3_3_port, S(2) => 
                           rca_out_3_2_port, S(1) => rca_out_3_1_port, S(0) => 
                           rca_out_3_0_port, Co => n_1162);
   rca_i_4 : rca_bhv_numBit32_3 port map( A(31) => rca_out_3_31_port, A(30) => 
                           rca_out_3_30_port, A(29) => rca_out_3_29_port, A(28)
                           => rca_out_3_28_port, A(27) => rca_out_3_27_port, 
                           A(26) => rca_out_3_26_port, A(25) => 
                           rca_out_3_25_port, A(24) => rca_out_3_24_port, A(23)
                           => rca_out_3_23_port, A(22) => rca_out_3_22_port, 
                           A(21) => rca_out_3_21_port, A(20) => 
                           rca_out_3_20_port, A(19) => rca_out_3_19_port, A(18)
                           => rca_out_3_18_port, A(17) => rca_out_3_17_port, 
                           A(16) => rca_out_3_16_port, A(15) => 
                           rca_out_3_15_port, A(14) => rca_out_3_14_port, A(13)
                           => rca_out_3_13_port, A(12) => rca_out_3_12_port, 
                           A(11) => rca_out_3_11_port, A(10) => 
                           rca_out_3_10_port, A(9) => rca_out_3_9_port, A(8) =>
                           rca_out_3_8_port, A(7) => rca_out_3_7_port, A(6) => 
                           rca_out_3_6_port, A(5) => rca_out_3_5_port, A(4) => 
                           rca_out_3_4_port, A(3) => rca_out_3_3_port, A(2) => 
                           rca_out_3_2_port, A(1) => rca_out_3_1_port, A(0) => 
                           rca_out_3_0_port, B(31) => sum_op_5_31_port, B(30) 
                           => sum_op_5_30_port, B(29) => sum_op_5_29_port, 
                           B(28) => sum_op_5_28_port, B(27) => sum_op_5_27_port
                           , B(26) => sum_op_5_26_port, B(25) => 
                           sum_op_5_25_port, B(24) => sum_op_5_24_port, B(23) 
                           => sum_op_5_23_port, B(22) => sum_op_5_22_port, 
                           B(21) => sum_op_5_21_port, B(20) => sum_op_5_20_port
                           , B(19) => sum_op_5_19_port, B(18) => 
                           sum_op_5_18_port, B(17) => sum_op_5_17_port, B(16) 
                           => sum_op_5_16_port, B(15) => sum_op_5_15_port, 
                           B(14) => sum_op_5_14_port, B(13) => sum_op_5_13_port
                           , B(12) => sum_op_5_12_port, B(11) => 
                           sum_op_5_11_port, B(10) => sum_op_5_10_port, B(9) =>
                           sum_op_5_9_port, B(8) => sum_op_5_8_port, B(7) => 
                           sum_op_5_7_port, B(6) => sum_op_5_6_port, B(5) => 
                           sum_op_5_5_port, B(4) => sum_op_5_4_port, B(3) => 
                           sum_op_5_3_port, B(2) => sum_op_5_2_port, B(1) => 
                           sum_op_5_1_port, B(0) => sum_op_5_0_port, Ci => 
                           X_Logic0_port, S(31) => rca_out_4_31_port, S(30) => 
                           rca_out_4_30_port, S(29) => rca_out_4_29_port, S(28)
                           => rca_out_4_28_port, S(27) => rca_out_4_27_port, 
                           S(26) => rca_out_4_26_port, S(25) => 
                           rca_out_4_25_port, S(24) => rca_out_4_24_port, S(23)
                           => rca_out_4_23_port, S(22) => rca_out_4_22_port, 
                           S(21) => rca_out_4_21_port, S(20) => 
                           rca_out_4_20_port, S(19) => rca_out_4_19_port, S(18)
                           => rca_out_4_18_port, S(17) => rca_out_4_17_port, 
                           S(16) => rca_out_4_16_port, S(15) => 
                           rca_out_4_15_port, S(14) => rca_out_4_14_port, S(13)
                           => rca_out_4_13_port, S(12) => rca_out_4_12_port, 
                           S(11) => rca_out_4_11_port, S(10) => 
                           rca_out_4_10_port, S(9) => rca_out_4_9_port, S(8) =>
                           rca_out_4_8_port, S(7) => rca_out_4_7_port, S(6) => 
                           rca_out_4_6_port, S(5) => rca_out_4_5_port, S(4) => 
                           rca_out_4_4_port, S(3) => rca_out_4_3_port, S(2) => 
                           rca_out_4_2_port, S(1) => rca_out_4_1_port, S(0) => 
                           rca_out_4_0_port, Co => n_1163);
   rca_i_5 : rca_bhv_numBit32_2 port map( A(31) => rca_out_4_31_port, A(30) => 
                           rca_out_4_30_port, A(29) => rca_out_4_29_port, A(28)
                           => rca_out_4_28_port, A(27) => rca_out_4_27_port, 
                           A(26) => rca_out_4_26_port, A(25) => 
                           rca_out_4_25_port, A(24) => rca_out_4_24_port, A(23)
                           => rca_out_4_23_port, A(22) => rca_out_4_22_port, 
                           A(21) => rca_out_4_21_port, A(20) => 
                           rca_out_4_20_port, A(19) => rca_out_4_19_port, A(18)
                           => rca_out_4_18_port, A(17) => rca_out_4_17_port, 
                           A(16) => rca_out_4_16_port, A(15) => 
                           rca_out_4_15_port, A(14) => rca_out_4_14_port, A(13)
                           => rca_out_4_13_port, A(12) => rca_out_4_12_port, 
                           A(11) => rca_out_4_11_port, A(10) => 
                           rca_out_4_10_port, A(9) => rca_out_4_9_port, A(8) =>
                           rca_out_4_8_port, A(7) => rca_out_4_7_port, A(6) => 
                           rca_out_4_6_port, A(5) => rca_out_4_5_port, A(4) => 
                           rca_out_4_4_port, A(3) => rca_out_4_3_port, A(2) => 
                           rca_out_4_2_port, A(1) => rca_out_4_1_port, A(0) => 
                           rca_out_4_0_port, B(31) => sum_op_6_31_port, B(30) 
                           => sum_op_6_30_port, B(29) => sum_op_6_29_port, 
                           B(28) => sum_op_6_28_port, B(27) => sum_op_6_27_port
                           , B(26) => sum_op_6_26_port, B(25) => 
                           sum_op_6_25_port, B(24) => sum_op_6_24_port, B(23) 
                           => sum_op_6_23_port, B(22) => sum_op_6_22_port, 
                           B(21) => sum_op_6_21_port, B(20) => sum_op_6_20_port
                           , B(19) => sum_op_6_19_port, B(18) => 
                           sum_op_6_18_port, B(17) => sum_op_6_17_port, B(16) 
                           => sum_op_6_16_port, B(15) => sum_op_6_15_port, 
                           B(14) => sum_op_6_14_port, B(13) => sum_op_6_13_port
                           , B(12) => sum_op_6_12_port, B(11) => 
                           sum_op_6_11_port, B(10) => sum_op_6_10_port, B(9) =>
                           sum_op_6_9_port, B(8) => sum_op_6_8_port, B(7) => 
                           sum_op_6_7_port, B(6) => sum_op_6_6_port, B(5) => 
                           sum_op_6_5_port, B(4) => sum_op_6_4_port, B(3) => 
                           sum_op_6_3_port, B(2) => sum_op_6_2_port, B(1) => 
                           sum_op_6_1_port, B(0) => sum_op_6_0_port, Ci => 
                           X_Logic0_port, S(31) => rca_out_5_31_port, S(30) => 
                           rca_out_5_30_port, S(29) => rca_out_5_29_port, S(28)
                           => rca_out_5_28_port, S(27) => rca_out_5_27_port, 
                           S(26) => rca_out_5_26_port, S(25) => 
                           rca_out_5_25_port, S(24) => rca_out_5_24_port, S(23)
                           => rca_out_5_23_port, S(22) => rca_out_5_22_port, 
                           S(21) => rca_out_5_21_port, S(20) => 
                           rca_out_5_20_port, S(19) => rca_out_5_19_port, S(18)
                           => rca_out_5_18_port, S(17) => rca_out_5_17_port, 
                           S(16) => rca_out_5_16_port, S(15) => 
                           rca_out_5_15_port, S(14) => rca_out_5_14_port, S(13)
                           => rca_out_5_13_port, S(12) => rca_out_5_12_port, 
                           S(11) => rca_out_5_11_port, S(10) => 
                           rca_out_5_10_port, S(9) => rca_out_5_9_port, S(8) =>
                           rca_out_5_8_port, S(7) => rca_out_5_7_port, S(6) => 
                           rca_out_5_6_port, S(5) => rca_out_5_5_port, S(4) => 
                           rca_out_5_4_port, S(3) => rca_out_5_3_port, S(2) => 
                           rca_out_5_2_port, S(1) => rca_out_5_1_port, S(0) => 
                           rca_out_5_0_port, Co => n_1164);
   rca_i_6 : rca_bhv_numBit32_1 port map( A(31) => rca_out_5_31_port, A(30) => 
                           rca_out_5_30_port, A(29) => rca_out_5_29_port, A(28)
                           => rca_out_5_28_port, A(27) => rca_out_5_27_port, 
                           A(26) => rca_out_5_26_port, A(25) => 
                           rca_out_5_25_port, A(24) => rca_out_5_24_port, A(23)
                           => rca_out_5_23_port, A(22) => rca_out_5_22_port, 
                           A(21) => rca_out_5_21_port, A(20) => 
                           rca_out_5_20_port, A(19) => rca_out_5_19_port, A(18)
                           => rca_out_5_18_port, A(17) => rca_out_5_17_port, 
                           A(16) => rca_out_5_16_port, A(15) => 
                           rca_out_5_15_port, A(14) => rca_out_5_14_port, A(13)
                           => rca_out_5_13_port, A(12) => rca_out_5_12_port, 
                           A(11) => rca_out_5_11_port, A(10) => 
                           rca_out_5_10_port, A(9) => rca_out_5_9_port, A(8) =>
                           rca_out_5_8_port, A(7) => rca_out_5_7_port, A(6) => 
                           rca_out_5_6_port, A(5) => rca_out_5_5_port, A(4) => 
                           rca_out_5_4_port, A(3) => rca_out_5_3_port, A(2) => 
                           rca_out_5_2_port, A(1) => rca_out_5_1_port, A(0) => 
                           rca_out_5_0_port, B(31) => sum_op_7_31_port, B(30) 
                           => sum_op_7_30_port, B(29) => sum_op_7_29_port, 
                           B(28) => sum_op_7_28_port, B(27) => sum_op_7_27_port
                           , B(26) => sum_op_7_26_port, B(25) => 
                           sum_op_7_25_port, B(24) => sum_op_7_24_port, B(23) 
                           => sum_op_7_23_port, B(22) => sum_op_7_22_port, 
                           B(21) => sum_op_7_21_port, B(20) => sum_op_7_20_port
                           , B(19) => sum_op_7_19_port, B(18) => 
                           sum_op_7_18_port, B(17) => sum_op_7_17_port, B(16) 
                           => sum_op_7_16_port, B(15) => sum_op_7_15_port, 
                           B(14) => sum_op_7_14_port, B(13) => sum_op_7_13_port
                           , B(12) => sum_op_7_12_port, B(11) => 
                           sum_op_7_11_port, B(10) => sum_op_7_10_port, B(9) =>
                           sum_op_7_9_port, B(8) => sum_op_7_8_port, B(7) => 
                           sum_op_7_7_port, B(6) => sum_op_7_6_port, B(5) => 
                           sum_op_7_5_port, B(4) => sum_op_7_4_port, B(3) => 
                           sum_op_7_3_port, B(2) => sum_op_7_2_port, B(1) => 
                           sum_op_7_1_port, B(0) => sum_op_7_0_port, Ci => 
                           X_Logic0_port, S(31) => P(31), S(30) => P(30), S(29)
                           => P(29), S(28) => P(28), S(27) => P(27), S(26) => 
                           P(26), S(25) => P(25), S(24) => P(24), S(23) => 
                           P(23), S(22) => P(22), S(21) => P(21), S(20) => 
                           P(20), S(19) => P(19), S(18) => P(18), S(17) => 
                           P(17), S(16) => P(16), S(15) => P(15), S(14) => 
                           P(14), S(13) => P(13), S(12) => P(12), S(11) => 
                           P(11), S(10) => P(10), S(9) => P(9), S(8) => P(8), 
                           S(7) => P(7), S(6) => P(6), S(5) => P(5), S(4) => 
                           P(4), S(3) => P(3), S(2) => P(2), S(1) => P(1), S(0)
                           => P(0), Co => n_1165);
   add_65_U1_1_1 : HA_X1 port map( A => add_65_A_1_port, B => add_65_A_0_port, 
                           CO => add_65_carry_2_port, S => A_minus_1_port);
   add_65_U1_1_2 : HA_X1 port map( A => add_65_A_2_port, B => 
                           add_65_carry_2_port, CO => add_65_carry_3_port, S =>
                           A_minus_2_port);
   add_65_U1_1_3 : HA_X1 port map( A => add_65_A_3_port, B => 
                           add_65_carry_3_port, CO => add_65_carry_4_port, S =>
                           A_minus_3_port);
   add_65_U1_1_4 : HA_X1 port map( A => add_65_A_4_port, B => 
                           add_65_carry_4_port, CO => add_65_carry_5_port, S =>
                           A_minus_4_port);
   add_65_U1_1_5 : HA_X1 port map( A => add_65_A_5_port, B => 
                           add_65_carry_5_port, CO => add_65_carry_6_port, S =>
                           A_minus_5_port);
   add_65_U1_1_6 : HA_X1 port map( A => add_65_A_6_port, B => 
                           add_65_carry_6_port, CO => add_65_carry_7_port, S =>
                           A_minus_6_port);
   add_65_U1_1_7 : HA_X1 port map( A => add_65_A_7_port, B => 
                           add_65_carry_7_port, CO => add_65_carry_8_port, S =>
                           A_minus_7_port);
   add_65_U1_1_8 : HA_X1 port map( A => add_65_A_8_port, B => 
                           add_65_carry_8_port, CO => add_65_carry_9_port, S =>
                           A_minus_8_port);
   add_65_U1_1_9 : HA_X1 port map( A => add_65_A_9_port, B => 
                           add_65_carry_9_port, CO => add_65_carry_10_port, S 
                           => A_minus_9_port);
   add_65_U1_1_10 : HA_X1 port map( A => add_65_A_10_port, B => 
                           add_65_carry_10_port, CO => add_65_carry_11_port, S 
                           => A_minus_10_port);
   add_65_U1_1_11 : HA_X1 port map( A => add_65_A_11_port, B => 
                           add_65_carry_11_port, CO => add_65_carry_12_port, S 
                           => A_minus_11_port);
   add_65_U1_1_12 : HA_X1 port map( A => add_65_A_12_port, B => 
                           add_65_carry_12_port, CO => add_65_carry_13_port, S 
                           => A_minus_12_port);
   add_65_U1_1_13 : HA_X1 port map( A => add_65_A_13_port, B => 
                           add_65_carry_13_port, CO => add_65_carry_14_port, S 
                           => A_minus_13_port);
   add_65_U1_1_14 : HA_X1 port map( A => add_65_A_14_port, B => 
                           add_65_carry_14_port, CO => add_65_carry_15_port, S 
                           => A_minus_14_port);
   U3 : INV_X1 port map( A => A_minus_14_port, ZN => n1);
   U4 : INV_X1 port map( A => n1, ZN => n2);
   U5 : INV_X1 port map( A => A_minus_13_port, ZN => n3);
   U6 : INV_X1 port map( A => n3, ZN => n4);
   U7 : INV_X1 port map( A => A_minus_12_port, ZN => n5);
   U8 : INV_X1 port map( A => n5, ZN => n6);
   U9 : INV_X1 port map( A => A_minus_11_port, ZN => n7);
   U10 : INV_X1 port map( A => n7, ZN => n8);
   U11 : INV_X1 port map( A => A_minus_10_port, ZN => n9);
   U12 : INV_X1 port map( A => n9, ZN => n10);
   U13 : INV_X1 port map( A => A_minus_9_port, ZN => n11);
   U14 : INV_X1 port map( A => n11, ZN => n12);
   U15 : INV_X1 port map( A => A_minus_8_port, ZN => n13);
   U16 : INV_X1 port map( A => n13, ZN => n14);
   U17 : INV_X1 port map( A => A_minus_7_port, ZN => n15);
   U18 : INV_X1 port map( A => n15, ZN => n16);
   U19 : INV_X1 port map( A => A_minus_6_port, ZN => n17);
   U20 : INV_X1 port map( A => n17, ZN => n18);
   U21 : INV_X1 port map( A => A_minus_5_port, ZN => n19);
   U22 : INV_X1 port map( A => n19, ZN => n20);
   U23 : INV_X1 port map( A => A_minus_4_port, ZN => n21);
   U24 : INV_X1 port map( A => n21, ZN => n22);
   U25 : INV_X1 port map( A => A_minus_3_port, ZN => n23);
   U26 : INV_X1 port map( A => n23, ZN => n24);
   U27 : INV_X1 port map( A => A_minus_2_port, ZN => n25);
   U28 : INV_X1 port map( A => n25, ZN => n26);
   U29 : INV_X1 port map( A => A_minus_1_port, ZN => n27);
   U30 : INV_X1 port map( A => n27, ZN => n28);
   U31 : BUF_X1 port map( A => n30, Z => n40);
   U32 : BUF_X1 port map( A => n30, Z => n39);
   U33 : BUF_X1 port map( A => n30, Z => n37);
   U34 : BUF_X1 port map( A => n30, Z => n38);
   U35 : BUF_X1 port map( A => n29, Z => n36);
   U36 : BUF_X1 port map( A => n29, Z => n31);
   U37 : BUF_X1 port map( A => n29, Z => n33);
   U38 : BUF_X1 port map( A => n29, Z => n35);
   U39 : BUF_X1 port map( A => n29, Z => n32);
   U40 : BUF_X1 port map( A => n29, Z => n34);
   U41 : BUF_X1 port map( A => n30, Z => n41);
   U42 : BUF_X1 port map( A => A_minus_31_port, Z => n29);
   U43 : BUF_X1 port map( A => A_minus_31_port, Z => n30);
   U44 : INV_X1 port map( A => n54, ZN => n42);
   U45 : INV_X1 port map( A => n54, ZN => n43);
   U46 : INV_X1 port map( A => n54, ZN => n47);
   U47 : INV_X1 port map( A => n54, ZN => n46);
   U48 : INV_X1 port map( A => n54, ZN => n44);
   U49 : INV_X1 port map( A => n54, ZN => n45);
   U50 : INV_X1 port map( A => n54, ZN => n48);
   U51 : INV_X1 port map( A => n54, ZN => n53);
   U52 : INV_X1 port map( A => n54, ZN => n52);
   U53 : INV_X1 port map( A => n54, ZN => n51);
   U54 : INV_X1 port map( A => n54, ZN => n50);
   U55 : INV_X1 port map( A => n54, ZN => n49);
   U56 : INV_X1 port map( A => add_65_A_0_port, ZN => A_minus_0_port);
   U57 : INV_X1 port map( A => A(0), ZN => add_65_A_0_port);
   U58 : INV_X1 port map( A => A(14), ZN => add_65_A_14_port);
   U59 : INV_X1 port map( A => A(1), ZN => add_65_A_1_port);
   U60 : INV_X1 port map( A => A(2), ZN => add_65_A_2_port);
   U61 : INV_X1 port map( A => A(3), ZN => add_65_A_3_port);
   U62 : INV_X1 port map( A => A(4), ZN => add_65_A_4_port);
   U63 : INV_X1 port map( A => A(5), ZN => add_65_A_5_port);
   U64 : INV_X1 port map( A => A(6), ZN => add_65_A_6_port);
   U65 : INV_X1 port map( A => A(7), ZN => add_65_A_7_port);
   U66 : INV_X1 port map( A => A(8), ZN => add_65_A_8_port);
   U67 : INV_X1 port map( A => A(9), ZN => add_65_A_9_port);
   U68 : INV_X1 port map( A => A(10), ZN => add_65_A_10_port);
   U69 : INV_X1 port map( A => A(11), ZN => add_65_A_11_port);
   U70 : INV_X1 port map( A => A(12), ZN => add_65_A_12_port);
   U71 : INV_X1 port map( A => A(13), ZN => add_65_A_13_port);
   U72 : XOR2_X2 port map( A => add_65_carry_15_port, B => n54, Z => 
                           A_minus_15_port);
   U73 : INV_X1 port map( A => A(15), ZN => n54);
   U74 : NOR2_X1 port map( A1 => add_65_carry_15_port, A2 => A(15), ZN => 
                           A_minus_31_port);
   encoder_out_0_port <= '0';

end SYN_mixed;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity P4Adder_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (31 downto 0);  Cout : out std_logic);

end P4Adder_NBIT32;

architecture SYN_struct of P4Adder_NBIT32 is

   component SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component carry_generator_NBIT32_NBIT_PER_BLOCK4
      port( A, B : in std_logic_vector (32 downto 1);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal Csum_7_port, Csum_6_port, Csum_5_port, Csum_4_port, Csum_3_port, 
      Csum_2_port, Csum_1_port : std_logic;

begin
   
   Carrygen0 : carry_generator_NBIT32_NBIT_PER_BLOCK4 port map( A(32) => A(31),
                           A(31) => A(30), A(30) => A(29), A(29) => A(28), 
                           A(28) => A(27), A(27) => A(26), A(26) => A(25), 
                           A(25) => A(24), A(24) => A(23), A(23) => A(22), 
                           A(22) => A(21), A(21) => A(20), A(20) => A(19), 
                           A(19) => A(18), A(18) => A(17), A(17) => A(16), 
                           A(16) => A(15), A(15) => A(14), A(14) => A(13), 
                           A(13) => A(12), A(12) => A(11), A(11) => A(10), 
                           A(10) => A(9), A(9) => A(8), A(8) => A(7), A(7) => 
                           A(6), A(6) => A(5), A(5) => A(4), A(4) => A(3), A(3)
                           => A(2), A(2) => A(1), A(1) => A(0), B(32) => B(31),
                           B(31) => B(30), B(30) => B(29), B(29) => B(28), 
                           B(28) => B(27), B(27) => B(26), B(26) => B(25), 
                           B(25) => B(24), B(24) => B(23), B(23) => B(22), 
                           B(22) => B(21), B(21) => B(20), B(20) => B(19), 
                           B(19) => B(18), B(18) => B(17), B(17) => B(16), 
                           B(16) => B(15), B(15) => B(14), B(14) => B(13), 
                           B(13) => B(12), B(12) => B(11), B(11) => B(10), 
                           B(10) => B(9), B(9) => B(8), B(8) => B(7), B(7) => 
                           B(6), B(6) => B(5), B(5) => B(4), B(4) => B(3), B(3)
                           => B(2), B(2) => B(1), B(1) => B(0), Cin => Cin, 
                           Co(7) => Cout, Co(6) => Csum_7_port, Co(5) => 
                           Csum_6_port, Co(4) => Csum_5_port, Co(3) => 
                           Csum_4_port, Co(2) => Csum_3_port, Co(1) => 
                           Csum_2_port, Co(0) => Csum_1_port);
   Sumgen0 : SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), Ci(7) => 
                           Csum_7_port, Ci(6) => Csum_6_port, Ci(5) => 
                           Csum_5_port, Ci(4) => Csum_4_port, Ci(3) => 
                           Csum_3_port, Ci(2) => Csum_2_port, Ci(1) => 
                           Csum_1_port, Ci(0) => Cin, S(31) => S(31), S(30) => 
                           S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           S(21), S(20) => S(20), S(19) => S(19), S(18) => 
                           S(18), S(17) => S(17), S(16) => S(16), S(15) => 
                           S(15), S(14) => S(14), S(13) => S(13), S(12) => 
                           S(12), S(11) => S(11), S(10) => S(10), S(9) => S(9),
                           S(8) => S(8), S(7) => S(7), S(6) => S(6), S(5) => 
                           S(5), S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1)
                           => S(1), S(0) => S(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity shifter_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  LOGIC_ARITH, LEFT_RIGHT : 
         in std_logic;  RES : out std_logic_vector (31 downto 0));

end shifter_NBIT32;

architecture SYN_bhv of shifter_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X4
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X2
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, 
      n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
      n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, 
      n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, 
      n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n1, n2, n3, n4, n5, n6, 
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n266, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649 : std_logic;

begin
   
   U264 : AOI21_X2 port map( B1 => A(31), B2 => B(18), A => n483, ZN => n282);
   U267 : OAI21_X2 port map( B1 => n613, B2 => n629, A => n486, ZN => n285);
   U269 : AOI21_X2 port map( B1 => A(31), B2 => n39, A => n487, ZN => n288);
   U388 : AOI221_X2 port map( B1 => n31, B2 => A(18), C1 => n21, C2 => A(17), A
                           => n568, ZN => n196);
   U428 : NOR2_X2 port map( A1 => n639, A2 => n39, ZN => n165);
   U461 : NOR2_X2 port map( A1 => n643, A2 => n39, ZN => n199);
   U637 : NAND3_X1 port map( A1 => n227, A2 => n647, A3 => n228, ZN => n226);
   U638 : NAND3_X1 port map( A1 => n227, A2 => n647, A3 => B(4), ZN => n428);
   U639 : NAND3_X1 port map( A1 => n445, A2 => n199, A3 => LEFT_RIGHT, ZN => 
                           n240);
   U641 : NAND3_X1 port map( A1 => n489, A2 => n629, A3 => n579, ZN => n255);
   U642 : NAND3_X1 port map( A1 => n267, A2 => n199, A3 => n445, ZN => n138);
   U2 : NOR4_X1 port map( A1 => B(20), A2 => B(21), A3 => B(19), A4 => n594, ZN
                           => n484);
   U3 : NOR2_X2 port map( A1 => n640, A2 => B(3), ZN => n262);
   U4 : NOR2_X2 port map( A1 => n490, A2 => B(11), ZN => n283);
   U5 : NAND3_X1 port map( A1 => n445, A2 => n35, A3 => LEFT_RIGHT, ZN => n269)
                           ;
   U6 : INV_X1 port map( A => n167, ZN => n636);
   U7 : NOR2_X1 port map( A1 => n637, A2 => B(4), ZN => n167);
   U8 : INV_X1 port map( A => n169, ZN => n645);
   U9 : INV_X1 port map( A => n165, ZN => n638);
   U10 : INV_X1 port map( A => n199, ZN => n642);
   U11 : INV_X1 port map( A => n32, ZN => n28);
   U12 : INV_X1 port map( A => n32, ZN => n26);
   U13 : INV_X1 port map( A => n32, ZN => n27);
   U14 : INV_X1 port map( A => n22, ZN => n14);
   U15 : INV_X1 port map( A => n22, ZN => n15);
   U16 : INV_X1 port map( A => n21, ZN => n16);
   U17 : INV_X1 port map( A => n505, ZN => n644);
   U18 : INV_X1 port map( A => n31, ZN => n29);
   U19 : INV_X1 port map( A => n493, ZN => n641);
   U20 : NOR2_X1 port map( A1 => n646, A2 => n39, ZN => n169);
   U21 : NAND2_X1 port map( A1 => n488, A2 => n454, ZN => n161);
   U22 : INV_X1 port map( A => n42, ZN => n39);
   U23 : OAI222_X1 port map( A1 => n79, A2 => n645, B1 => n63, B2 => n636, C1 
                           => n91, C2 => n638, ZN => n371);
   U24 : OAI222_X1 port map( A1 => n82, A2 => n645, B1 => n62, B2 => n636, C1 
                           => n95, C2 => n638, ZN => n360);
   U25 : OAI222_X1 port map( A1 => n85, A2 => n645, B1 => n73, B2 => n636, C1 
                           => n99, C2 => n638, ZN => n349);
   U26 : OAI222_X1 port map( A1 => n87, A2 => n645, B1 => n76, B2 => n636, C1 
                           => n104, C2 => n638, ZN => n338);
   U27 : NOR2_X1 port map( A1 => n41, A2 => n643, ZN => n493);
   U28 : OAI22_X1 port map( A1 => n116, A2 => n643, B1 => n127, B2 => n639, ZN 
                           => n383);
   U29 : INV_X1 port map( A => n454, ZN => n637);
   U30 : AOI21_X1 port map( B1 => n135, B2 => n2, A => n519, ZN => n286);
   U31 : AOI21_X1 port map( B1 => n130, B2 => n3, A => n519, ZN => n312);
   U32 : BUF_X1 port map( A => n138, Z => n34);
   U33 : BUF_X1 port map( A => n138, Z => n33);
   U34 : NOR2_X1 port map( A1 => n383, A2 => n359, ZN => n197);
   U35 : NOR2_X1 port map( A1 => n119, A2 => n359, ZN => n181);
   U36 : BUF_X1 port map( A => n138, Z => n35);
   U37 : NAND2_X1 port map( A1 => n488, A2 => n5, ZN => n505);
   U38 : INV_X1 port map( A => n182, ZN => n119);
   U39 : INV_X1 port map( A => n238, ZN => n107);
   U40 : INV_X1 port map( A => n214, ZN => n56);
   U41 : INV_X1 port map( A => n202, ZN => n50);
   U42 : INV_X1 port map( A => n188, ZN => n48);
   U43 : NOR2_X1 port map( A1 => n613, A2 => n148, ZN => n150);
   U44 : OAI21_X2 port map( B1 => n612, B2 => n633, A => n481, ZN => n279);
   U45 : NOR2_X1 port map( A1 => n640, A2 => n647, ZN => n454);
   U46 : NAND2_X1 port map( A1 => n484, A2 => n631, ZN => n281);
   U47 : AOI222_X1 port map( A1 => n370, A2 => n262, B1 => n320, B2 => n260, C1
                           => n185, C2 => n3, ZN => n238);
   U48 : INV_X1 port map( A => n356, ZN => n643);
   U49 : AOI222_X1 port map( A1 => n168, A2 => n262, B1 => n355, B2 => n260, C1
                           => n170, C2 => n3, ZN => n471);
   U50 : AOI222_X1 port map( A1 => n402, A2 => n262, B1 => n403, B2 => n260, C1
                           => n464, C2 => n2, ZN => n461);
   U51 : NAND2_X1 port map( A1 => n488, A2 => n262, ZN => n157);
   U52 : NAND2_X1 port map( A1 => n488, A2 => n260, ZN => n158);
   U53 : OAI222_X1 port map( A1 => n374, A2 => n639, B1 => n646, B2 => n375, C1
                           => n376, C2 => n643, ZN => n172);
   U54 : OAI222_X1 port map( A1 => n132, A2 => n639, B1 => n362, B2 => n646, C1
                           => n363, C2 => n643, ZN => n139);
   U55 : OAI222_X1 port map( A1 => n614, A2 => n639, B1 => n293, B2 => n646, C1
                           => n405, C2 => n643, ZN => n348);
   U56 : OAI222_X1 port map( A1 => n616, A2 => n639, B1 => n46, B2 => n646, C1 
                           => n387, C2 => n643, ZN => n337);
   U57 : AOI221_X1 port map( B1 => n130, B2 => n262, C1 => n355, C2 => n2, A =>
                           n359, ZN => n159);
   U58 : AOI221_X1 port map( B1 => n135, B2 => n262, C1 => n403, C2 => n3, A =>
                           n359, ZN => n347);
   U59 : OAI221_X1 port map( B1 => n106, B2 => n639, C1 => n90, C2 => n643, A 
                           => n607, ZN => n480);
   U60 : AOI22_X1 port map( A1 => n454, A2 => n320, B1 => n260, B2 => n370, ZN 
                           => n607);
   U61 : AOI222_X1 port map( A1 => n169, A2 => n185, B1 => n493, B2 => n320, C1
                           => n167, C2 => n370, ZN => n550);
   U62 : OAI222_X1 port map( A1 => n62, A2 => n645, B1 => n363, B2 => n636, C1 
                           => n82, C2 => n638, ZN => n418);
   U63 : OAI222_X1 port map( A1 => n73, A2 => n645, B1 => n405, B2 => n636, C1 
                           => n85, C2 => n638, ZN => n404);
   U64 : OAI222_X1 port map( A1 => n76, A2 => n645, B1 => n387, B2 => n636, C1 
                           => n87, C2 => n638, ZN => n386);
   U65 : INV_X1 port map( A => n260, ZN => n646);
   U66 : NOR2_X1 port map( A1 => n648, A2 => B(4), ZN => n488);
   U67 : INV_X1 port map( A => n262, ZN => n639);
   U68 : INV_X1 port map( A => n332, ZN => n628);
   U69 : OAI222_X1 port map( A1 => n133, A2 => n14, B1 => n29, B2 => n615, C1 
                           => n1, C2 => n103, ZN => n602);
   U70 : OAI221_X1 port map( B1 => n363, B2 => n639, C1 => n62, C2 => n643, A 
                           => n522, ZN => n314);
   U71 : AOI22_X1 port map( A1 => n454, A2 => n58, B1 => n260, B2 => n420, ZN 
                           => n522);
   U72 : OAI221_X1 port map( B1 => n405, B2 => n639, C1 => n73, C2 => n643, A 
                           => n509, ZN => n290);
   U73 : AOI22_X1 port map( A1 => n454, A2 => n52, B1 => n260, B2 => n407, ZN 
                           => n509);
   U74 : OAI221_X1 port map( B1 => n387, B2 => n639, C1 => n76, C2 => n643, A 
                           => n496, ZN => n271);
   U75 : AOI22_X1 port map( A1 => n454, A2 => n390, B1 => n260, B2 => n389, ZN 
                           => n496);
   U76 : OAI21_X1 port map( B1 => n613, B2 => n631, A => n486, ZN => n253);
   U77 : NOR2_X1 port map( A1 => n613, A2 => n647, ZN => n359);
   U78 : NOR2_X1 port map( A1 => n613, A2 => n2, ZN => n519);
   U79 : AOI221_X1 port map( B1 => n219, B2 => n199, C1 => n223, C2 => n39, A 
                           => n224, ZN => n222);
   U80 : OAI222_X1 port map( A1 => n638, A2 => n71, B1 => n636, B2 => n93, C1 
                           => n645, C2 => n81, ZN => n224);
   U81 : AOI221_X1 port map( B1 => n207, B2 => n199, C1 => n211, C2 => n39, A 
                           => n212, ZN => n210);
   U82 : OAI222_X1 port map( A1 => n638, A2 => n68, B1 => n636, B2 => n97, C1 
                           => n645, C2 => n84, ZN => n212);
   U83 : AOI221_X1 port map( B1 => n193, B2 => n199, C1 => n115, C2 => n39, A 
                           => n200, ZN => n198);
   U84 : OAI222_X1 port map( A1 => n638, A2 => n75, B1 => n636, B2 => n101, C1 
                           => n645, C2 => n196, ZN => n200);
   U85 : OAI22_X1 port map( A1 => n8, A2 => n131, B1 => n1, B2 => n266, ZN => 
                           n533);
   U86 : OAI221_X1 port map( B1 => n618, B2 => n642, C1 => n238, C2 => n41, A 
                           => n239, ZN => n229);
   U87 : AOI222_X1 port map( A1 => n165, A2 => n178, B1 => n167, B2 => n186, C1
                           => n169, C2 => n184, ZN => n239);
   U88 : OAI221_X1 port map( B1 => n65, B2 => n642, C1 => n182, C2 => n41, A =>
                           n183, ZN => n173);
   U89 : AOI222_X1 port map( A1 => n165, A2 => n184, B1 => n167, B2 => n185, C1
                           => n169, C2 => n186, ZN => n183);
   U90 : OAI221_X1 port map( B1 => n71, B2 => n642, C1 => n163, C2 => n42, A =>
                           n164, ZN => n141);
   U91 : AOI222_X1 port map( A1 => n165, A2 => n166, B1 => n167, B2 => n168, C1
                           => n169, C2 => n170, ZN => n164);
   U92 : OAI221_X1 port map( B1 => n68, B2 => n642, C1 => n344, C2 => n42, A =>
                           n581, ZN => n572);
   U93 : AOI222_X1 port map( A1 => n165, A2 => n516, B1 => n167, B2 => n402, C1
                           => n169, C2 => n464, ZN => n581);
   U94 : OAI221_X1 port map( B1 => n93, B2 => n638, C1 => n81, C2 => n642, A =>
                           n534, ZN => n526);
   U95 : AOI222_X1 port map( A1 => n169, A2 => n168, B1 => n493, B2 => n129, C1
                           => n167, C2 => n355, ZN => n534);
   U96 : OAI221_X1 port map( B1 => n97, B2 => n638, C1 => n84, C2 => n642, A =>
                           n520, ZN => n511);
   U97 : AOI222_X1 port map( A1 => n169, A2 => n402, B1 => n493, B2 => n134, C1
                           => n167, C2 => n403, ZN => n520);
   U98 : OAI221_X1 port map( B1 => n101, B2 => n638, C1 => n196, C2 => n642, A 
                           => n507, ZN => n498);
   U99 : AOI222_X1 port map( A1 => n169, A2 => n453, B1 => n493, B2 => n382, C1
                           => n167, C2 => n506, ZN => n507);
   U100 : NOR2_X1 port map( A1 => n613, A2 => n8, ZN => n382);
   U101 : OAI221_X1 port map( B1 => n127, B2 => n161, C1 => n116, C2 => n158, A
                           => n162, ZN => n503);
   U102 : OAI221_X1 port map( B1 => n237, B2 => n160, C1 => n90, C2 => n161, A 
                           => n162, ZN => n235);
   U103 : OAI221_X1 port map( B1 => n110, B2 => n160, C1 => n93, C2 => n161, A 
                           => n162, ZN => n220);
   U104 : OAI221_X1 port map( B1 => n113, B2 => n160, C1 => n97, C2 => n161, A 
                           => n162, ZN => n208);
   U105 : OAI221_X1 port map( B1 => n197, B2 => n160, C1 => n101, C2 => n161, A
                           => n162, ZN => n194);
   U106 : OAI221_X1 port map( B1 => n181, B2 => n160, C1 => n106, C2 => n161, A
                           => n162, ZN => n179);
   U107 : OAI221_X1 port map( B1 => n159, B2 => n160, C1 => n109, C2 => n161, A
                           => n162, ZN => n155);
   U108 : OAI221_X1 port map( B1 => n347, B2 => n160, C1 => n112, C2 => n161, A
                           => n162, ZN => n577);
   U109 : OAI221_X1 port map( B1 => n336, B2 => n160, C1 => n116, C2 => n161, A
                           => n162, ZN => n560);
   U110 : OAI221_X1 port map( B1 => n323, B2 => n160, C1 => n118, C2 => n161, A
                           => n162, ZN => n548);
   U111 : INV_X1 port map( A => n370, ZN => n118);
   U112 : OAI221_X1 port map( B1 => n312, B2 => n160, C1 => n121, C2 => n161, A
                           => n162, ZN => n531);
   U113 : INV_X1 port map( A => n355, ZN => n121);
   U114 : OAI221_X1 port map( B1 => n286, B2 => n160, C1 => n124, C2 => n161, A
                           => n162, ZN => n517);
   U115 : INV_X1 port map( A => n403, ZN => n124);
   U116 : AND2_X1 port map( A1 => n491, A2 => n633, ZN => n276);
   U117 : AOI22_X1 port map( A1 => n480, A2 => n39, B1 => n43, B2 => n64, ZN =>
                           n587);
   U118 : INV_X1 port map( A => n601, ZN => n64);
   U119 : AOI221_X1 port map( B1 => n4, B2 => n602, C1 => n454, C2 => n184, A 
                           => n603, ZN => n601);
   U120 : OAI22_X1 port map( A1 => n618, A2 => n639, B1 => n65, B2 => n646, ZN 
                           => n603);
   U121 : AOI22_X1 port map( A1 => n420, A2 => n2, B1 => n58, B2 => n262, ZN =>
                           n214);
   U122 : AOI22_X1 port map( A1 => n407, A2 => n5, B1 => n52, B2 => n262, ZN =>
                           n202);
   U123 : AOI22_X1 port map( A1 => n389, A2 => n3, B1 => n390, B2 => n262, ZN 
                           => n188);
   U124 : AOI22_X1 port map( A1 => n168, A2 => n3, B1 => n355, B2 => n262, ZN 
                           => n413);
   U125 : AOI22_X1 port map( A1 => n402, A2 => n5, B1 => n403, B2 => n262, ZN 
                           => n396);
   U126 : AOI22_X1 port map( A1 => n452, A2 => n4, B1 => n453, B2 => n262, ZN 
                           => n449);
   U127 : AOI22_X1 port map( A1 => n370, A2 => n4, B1 => n320, B2 => n262, ZN 
                           => n182);
   U128 : AOI22_X1 port map( A1 => n355, A2 => n2, B1 => n129, B2 => n262, ZN 
                           => n163);
   U129 : AOI22_X1 port map( A1 => n403, A2 => n4, B1 => n134, B2 => n262, ZN 
                           => n344);
   U130 : AOI21_X1 port map( B1 => n148, B2 => n232, A => n150, ZN => n231);
   U131 : OAI21_X1 port map( B1 => n233, B2 => n152, A => n153, ZN => n232);
   U132 : AOI211_X1 port map( C1 => n644, C2 => n234, A => n235, B => n236, ZN 
                           => n233);
   U133 : OAI22_X1 port map( A1 => n65, A2 => n157, B1 => n78, B2 => n158, ZN 
                           => n236);
   U134 : AOI21_X1 port map( B1 => n148, B2 => n217, A => n150, ZN => n216);
   U135 : OAI21_X1 port map( B1 => n218, B2 => n152, A => n153, ZN => n217);
   U136 : AOI211_X1 port map( C1 => n644, C2 => n219, A => n220, B => n221, ZN 
                           => n218);
   U137 : OAI22_X1 port map( A1 => n71, A2 => n157, B1 => n81, B2 => n158, ZN 
                           => n221);
   U138 : AOI21_X1 port map( B1 => n148, B2 => n205, A => n150, ZN => n204);
   U139 : OAI21_X1 port map( B1 => n206, B2 => n152, A => n153, ZN => n205);
   U140 : AOI211_X1 port map( C1 => n644, C2 => n207, A => n208, B => n209, ZN 
                           => n206);
   U141 : OAI22_X1 port map( A1 => n68, A2 => n157, B1 => n84, B2 => n158, ZN 
                           => n209);
   U142 : AOI21_X1 port map( B1 => n148, B2 => n191, A => n150, ZN => n190);
   U143 : OAI21_X1 port map( B1 => n192, B2 => n152, A => n153, ZN => n191);
   U144 : AOI211_X1 port map( C1 => n644, C2 => n193, A => n194, B => n195, ZN 
                           => n192);
   U145 : OAI22_X1 port map( A1 => n75, A2 => n157, B1 => n196, B2 => n158, ZN 
                           => n195);
   U146 : AOI21_X1 port map( B1 => n148, B2 => n176, A => n150, ZN => n175);
   U147 : OAI21_X1 port map( B1 => n177, B2 => n152, A => n153, ZN => n176);
   U148 : AOI211_X1 port map( C1 => n644, C2 => n178, A => n179, B => n180, ZN 
                           => n177);
   U149 : OAI22_X1 port map( A1 => n78, A2 => n157, B1 => n90, B2 => n158, ZN 
                           => n180);
   U150 : AOI21_X1 port map( B1 => n148, B2 => n149, A => n150, ZN => n145);
   U151 : OAI21_X1 port map( B1 => n151, B2 => n152, A => n153, ZN => n149);
   U152 : AOI211_X1 port map( C1 => n644, C2 => n154, A => n155, B => n156, ZN 
                           => n151);
   U153 : OAI22_X1 port map( A1 => n81, A2 => n157, B1 => n93, B2 => n158, ZN 
                           => n156);
   U154 : AOI21_X1 port map( B1 => n148, B2 => n575, A => n150, ZN => n574);
   U155 : OAI21_X1 port map( B1 => n576, B2 => n152, A => n153, ZN => n575);
   U156 : AOI211_X1 port map( C1 => n644, C2 => n305, A => n577, B => n578, ZN 
                           => n576);
   U157 : OAI22_X1 port map( A1 => n84, A2 => n157, B1 => n97, B2 => n158, ZN 
                           => n578);
   U158 : AOI21_X1 port map( B1 => n148, B2 => n558, A => n150, ZN => n557);
   U159 : OAI21_X1 port map( B1 => n559, B2 => n152, A => n153, ZN => n558);
   U160 : AOI211_X1 port map( C1 => n644, C2 => n261, A => n560, B => n561, ZN 
                           => n559);
   U161 : OAI22_X1 port map( A1 => n196, A2 => n157, B1 => n101, B2 => n158, ZN
                           => n561);
   U162 : AOI21_X1 port map( B1 => n148, B2 => n546, A => n150, ZN => n545);
   U163 : OAI21_X1 port map( B1 => n547, B2 => n152, A => n153, ZN => n546);
   U164 : AOI211_X1 port map( C1 => n644, C2 => n184, A => n548, B => n549, ZN 
                           => n547);
   U165 : OAI22_X1 port map( A1 => n90, A2 => n157, B1 => n106, B2 => n158, ZN 
                           => n549);
   U166 : AOI21_X1 port map( B1 => n148, B2 => n529, A => n150, ZN => n528);
   U167 : OAI21_X1 port map( B1 => n530, B2 => n152, A => n153, ZN => n529);
   U168 : AOI211_X1 port map( C1 => n644, C2 => n166, A => n531, B => n532, ZN 
                           => n530);
   U169 : OAI22_X1 port map( A1 => n93, A2 => n157, B1 => n109, B2 => n158, ZN 
                           => n532);
   U170 : AOI21_X1 port map( B1 => n148, B2 => n514, A => n150, ZN => n513);
   U171 : OAI21_X1 port map( B1 => n515, B2 => n152, A => n153, ZN => n514);
   U172 : AOI211_X1 port map( C1 => n644, C2 => n516, A => n517, B => n518, ZN 
                           => n515);
   U173 : OAI22_X1 port map( A1 => n97, A2 => n157, B1 => n112, B2 => n158, ZN 
                           => n518);
   U174 : AOI21_X1 port map( B1 => n283, B2 => n415, A => n285, ZN => n414);
   U175 : OAI21_X1 port map( B1 => n110, B2 => n287, A => n288, ZN => n415);
   U176 : AOI21_X1 port map( B1 => n283, B2 => n398, A => n285, ZN => n397);
   U177 : OAI21_X1 port map( B1 => n113, B2 => n287, A => n288, ZN => n398);
   U178 : AOI21_X1 port map( B1 => n283, B2 => n385, A => n285, ZN => n384);
   U179 : OAI21_X1 port map( B1 => n197, B2 => n287, A => n288, ZN => n385);
   U180 : AOI21_X1 port map( B1 => n283, B2 => n369, A => n285, ZN => n368);
   U181 : OAI21_X1 port map( B1 => n181, B2 => n287, A => n288, ZN => n369);
   U182 : AOI21_X1 port map( B1 => n283, B2 => n335, A => n285, ZN => n334);
   U183 : OAI21_X1 port map( B1 => n336, B2 => n287, A => n288, ZN => n335);
   U184 : OAI211_X1 port map( C1 => n127, C2 => n646, A => n401, B => n449, ZN 
                           => n257);
   U185 : AOI21_X1 port map( B1 => n320, B2 => n4, A => n519, ZN => n323);
   U186 : AOI21_X1 port map( B1 => n506, B2 => n5, A => n519, ZN => n336);
   U187 : NAND2_X1 port map( A1 => n484, A2 => n633, ZN => n249);
   U188 : OAI21_X1 port map( B1 => n417, B2 => n637, A => n471, ZN => n440);
   U189 : OAI21_X1 port map( B1 => n400, B2 => n637, A => n461, ZN => n302);
   U190 : NOR2_X1 port map( A1 => n613, A2 => n484, ZN => n483);
   U191 : OAI21_X1 port map( B1 => n412, B2 => n637, A => n471, ZN => n434);
   U192 : OAI21_X1 port map( B1 => n395, B2 => n637, A => n461, ZN => n297);
   U193 : OAI21_X1 port map( B1 => n412, B2 => n646, A => n413, ZN => n223);
   U194 : OAI21_X1 port map( B1 => n395, B2 => n646, A => n396, ZN => n211);
   U195 : OAI21_X1 port map( B1 => n333, B2 => n647, A => n449, ZN => n246);
   U196 : OAI21_X1 port map( B1 => n482, B2 => n281, A => n282, ZN => n479);
   U197 : AOI21_X1 port map( B1 => n283, B2 => n485, A => n285, ZN => n482);
   U198 : OAI21_X1 port map( B1 => n89, B2 => n287, A => n288, ZN => n485);
   U199 : INV_X1 port map( A => n480, ZN => n89);
   U200 : OAI21_X1 port map( B1 => n472, B2 => n281, A => n282, ZN => n470);
   U201 : AOI21_X1 port map( B1 => n283, B2 => n473, A => n285, ZN => n472);
   U202 : OAI21_X1 port map( B1 => n94, B2 => n287, A => n288, ZN => n473);
   U203 : INV_X1 port map( A => n440, ZN => n94);
   U204 : OAI21_X1 port map( B1 => n462, B2 => n281, A => n282, ZN => n460);
   U205 : AOI21_X1 port map( B1 => n283, B2 => n463, A => n285, ZN => n462);
   U206 : OAI21_X1 port map( B1 => n98, B2 => n287, A => n288, ZN => n463);
   U207 : INV_X1 port map( A => n302, ZN => n98);
   U208 : OAI21_X1 port map( B1 => n450, B2 => n281, A => n282, ZN => n448);
   U209 : AOI21_X1 port map( B1 => n283, B2 => n451, A => n285, ZN => n450);
   U210 : OAI21_X1 port map( B1 => n102, B2 => n287, A => n288, ZN => n451);
   U211 : INV_X1 port map( A => n257, ZN => n102);
   U212 : OAI21_X1 port map( B1 => n425, B2 => n281, A => n282, ZN => n424);
   U213 : AOI21_X1 port map( B1 => n283, B2 => n426, A => n285, ZN => n425);
   U214 : OAI21_X1 port map( B1 => n237, B2 => n287, A => n288, ZN => n426);
   U215 : OAI21_X1 port map( B1 => n357, B2 => n281, A => n282, ZN => n354);
   U216 : AOI21_X1 port map( B1 => n283, B2 => n358, A => n285, ZN => n357);
   U217 : OAI21_X1 port map( B1 => n159, B2 => n287, A => n288, ZN => n358);
   U218 : OAI21_X1 port map( B1 => n345, B2 => n281, A => n282, ZN => n343);
   U219 : AOI21_X1 port map( B1 => n283, B2 => n346, A => n285, ZN => n345);
   U220 : OAI21_X1 port map( B1 => n347, B2 => n287, A => n288, ZN => n346);
   U221 : OAI21_X1 port map( B1 => n321, B2 => n281, A => n282, ZN => n319);
   U222 : AOI21_X1 port map( B1 => n283, B2 => n322, A => n285, ZN => n321);
   U223 : OAI21_X1 port map( B1 => n323, B2 => n287, A => n288, ZN => n322);
   U224 : OAI21_X1 port map( B1 => n310, B2 => n281, A => n282, ZN => n309);
   U225 : AOI21_X1 port map( B1 => n283, B2 => n311, A => n285, ZN => n310);
   U226 : OAI21_X1 port map( B1 => n312, B2 => n287, A => n288, ZN => n311);
   U227 : OAI21_X1 port map( B1 => n280, B2 => n281, A => n282, ZN => n277);
   U228 : AOI21_X1 port map( B1 => n283, B2 => n284, A => n285, ZN => n280);
   U229 : OAI21_X1 port map( B1 => n286, B2 => n287, A => n288, ZN => n284);
   U230 : AOI22_X1 port map( A1 => n246, A2 => n39, B1 => n43, B2 => n247, ZN 
                           => n245);
   U231 : AOI22_X1 port map( A1 => n434, A2 => n39, B1 => n42, B2 => n435, ZN 
                           => n433);
   U232 : AOI22_X1 port map( A1 => n297, A2 => n39, B1 => n42, B2 => n298, ZN 
                           => n296);
   U233 : INV_X1 port map( A => n452, ZN => n101);
   U234 : INV_X1 port map( A => n464, ZN => n97);
   U235 : INV_X1 port map( A => n170, ZN => n93);
   U236 : INV_X1 port map( A => n186, ZN => n90);
   U237 : INV_X1 port map( A => n516, ZN => n84);
   U238 : INV_X1 port map( A => n166, ZN => n81);
   U239 : NOR2_X1 port map( A1 => n266, A2 => n8, ZN => n580);
   U240 : AOI21_X1 port map( B1 => n251, B2 => n438, A => n253, ZN => n437);
   U241 : OAI21_X1 port map( B1 => n439, B2 => n255, A => n256, ZN => n438);
   U242 : AOI22_X1 port map( A1 => n435, A2 => n40, B1 => B(4), B2 => n440, ZN 
                           => n439);
   U243 : AOI21_X1 port map( B1 => n251, B2 => n300, A => n253, ZN => n299);
   U244 : OAI21_X1 port map( B1 => n301, B2 => n255, A => n256, ZN => n300);
   U245 : AOI22_X1 port map( A1 => n298, A2 => n40, B1 => B(4), B2 => n302, ZN 
                           => n301);
   U246 : AOI21_X1 port map( B1 => n251, B2 => n252, A => n253, ZN => n248);
   U247 : OAI21_X1 port map( B1 => n254, B2 => n255, A => n256, ZN => n252);
   U248 : AOI22_X1 port map( A1 => n247, A2 => n40, B1 => B(4), B2 => n257, ZN 
                           => n254);
   U249 : BUF_X1 port map( A => n356, Z => n2);
   U250 : BUF_X1 port map( A => n356, Z => n3);
   U251 : INV_X1 port map( A => n293, ZN => n52);
   U252 : INV_X1 port map( A => n184, ZN => n78);
   U253 : INV_X1 port map( A => n506, ZN => n127);
   U254 : INV_X1 port map( A => n185, ZN => n106);
   U255 : INV_X1 port map( A => n412, ZN => n129);
   U256 : INV_X1 port map( A => n395, ZN => n134);
   U257 : INV_X1 port map( A => n390, ZN => n46);
   U258 : BUF_X1 port map( A => n356, Z => n4);
   U259 : BUF_X1 port map( A => n356, Z => n5);
   U260 : INV_X1 port map( A => n453, ZN => n116);
   U261 : INV_X1 port map( A => n154, ZN => n71);
   U262 : INV_X1 port map( A => n305, ZN => n68);
   U263 : INV_X1 port map( A => n178, ZN => n65);
   U265 : INV_X1 port map( A => n168, ZN => n109);
   U266 : INV_X1 port map( A => n402, ZN => n112);
   U268 : INV_X1 port map( A => n261, ZN => n75);
   U270 : INV_X1 port map( A => n419, ZN => n82);
   U271 : INV_X1 port map( A => n406, ZN => n85);
   U272 : INV_X1 port map( A => n388, ZN => n87);
   U273 : BUF_X1 port map( A => n44, Z => n42);
   U274 : INV_X1 port map( A => n362, ZN => n58);
   U275 : INV_X1 port map( A => n474, ZN => n62);
   U276 : INV_X1 port map( A => n465, ZN => n73);
   U277 : INV_X1 port map( A => n455, ZN => n76);
   U278 : INV_X1 port map( A => n267, ZN => n8);
   U279 : BUF_X1 port map( A => n44, Z => n43);
   U280 : BUF_X1 port map( A => n44, Z => n40);
   U281 : INV_X1 port map( A => n417, ZN => n130);
   U282 : INV_X1 port map( A => n400, ZN => n135);
   U283 : BUF_X1 port map( A => n44, Z => n41);
   U284 : INV_X1 port map( A => n373, ZN => n79);
   U285 : INV_X1 port map( A => n420, ZN => n132);
   U286 : INV_X1 port map( A => n407, ZN => n614);
   U287 : INV_X1 port map( A => n389, ZN => n616);
   U288 : INV_X1 port map( A => n429, ZN => n63);
   U289 : INV_X1 port map( A => n372, ZN => n91);
   U290 : INV_X1 port map( A => n361, ZN => n95);
   U291 : INV_X1 port map( A => n350, ZN => n99);
   U292 : INV_X1 port map( A => n339, ZN => n104);
   U293 : AND2_X1 port map( A1 => n238, A2 => n401, ZN => n237);
   U294 : INV_X1 port map( A => n234, ZN => n618);
   U295 : INV_X1 port map( A => n416, ZN => n110);
   U296 : OAI211_X1 port map( C1 => n417, C2 => n646, A => n401, B => n413, ZN 
                           => n416);
   U297 : INV_X1 port map( A => n399, ZN => n113);
   U298 : OAI211_X1 port map( C1 => n400, C2 => n646, A => n401, B => n396, ZN 
                           => n399);
   U299 : INV_X1 port map( A => n381, ZN => n115);
   U300 : AOI21_X1 port map( B1 => n260, B2 => n382, A => n383, ZN => n381);
   U301 : OR4_X1 port map( A1 => B(21), A2 => B(20), A3 => B(19), A4 => B(18), 
                           ZN => n598);
   U302 : OAI22_X1 port map( A1 => n88, A2 => n1, B1 => n86, B2 => n8, ZN => 
                           n568);
   U303 : AOI222_X1 port map( A1 => n11, A2 => A(1), B1 => A(0), B2 => n18, C1 
                           => n7, C2 => A(2), ZN => n293);
   U304 : AOI221_X1 port map( B1 => n31, B2 => A(6), C1 => n20, C2 => A(7), A 
                           => n525, ZN => n363);
   U305 : OAI22_X1 port map( A1 => n623, A2 => n1, B1 => n624, B2 => n8, ZN => 
                           n525);
   U306 : AOI221_X1 port map( B1 => n30, B2 => A(7), C1 => n20, C2 => A(8), A 
                           => n570, ZN => n405);
   U307 : OAI22_X1 port map( A1 => n624, A2 => n1, B1 => n66, B2 => n8, ZN => 
                           n570);
   U308 : AOI221_X1 port map( B1 => n31, B2 => A(8), C1 => n21, C2 => A(9), A 
                           => n552, ZN => n387);
   U309 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n74, B2 => n8, ZN => 
                           n552);
   U310 : AOI221_X1 port map( B1 => n30, B2 => A(5), C1 => n20, C2 => A(6), A 
                           => n541, ZN => n376);
   U311 : OAI22_X1 port map( A1 => n622, A2 => n1, B1 => n623, B2 => n8, ZN => 
                           n541);
   U312 : OAI221_X1 port map( B1 => n29, B2 => n613, C1 => n17, C2 => n266, A 
                           => n609, ZN => n320);
   U313 : AOI22_X1 port map( A1 => A(29), A2 => n10, B1 => A(28), B2 => n267, 
                           ZN => n609);
   U314 : OAI221_X1 port map( B1 => n27, B2 => n128, C1 => n15, C2 => n126, A 
                           => n535, ZN => n355);
   U315 : AOI22_X1 port map( A1 => A(26), A2 => n11, B1 => A(25), B2 => n6, ZN 
                           => n535);
   U316 : OAI221_X1 port map( B1 => n28, B2 => n131, C1 => n16, C2 => n128, A 
                           => n585, ZN => n403);
   U317 : AOI22_X1 port map( A1 => A(27), A2 => n9, B1 => A(26), B2 => n267, ZN
                           => n585);
   U318 : OR3_X1 port map( A1 => B(22), A2 => B(24), A3 => B(23), ZN => n594);
   U319 : NAND3_X1 port map( A1 => n489, A2 => n629, A3 => n600, ZN => n152);
   U320 : NOR3_X1 port map( A1 => B(12), A2 => B(14), A3 => B(13), ZN => n600);
   U321 : NAND3_X1 port map( A1 => n592, A2 => n632, A3 => n599, ZN => n146);
   U322 : INV_X1 port map( A => B(22), ZN => n632);
   U323 : NOR3_X1 port map( A1 => B(23), A2 => B(25), A3 => B(24), ZN => n599);
   U324 : NAND2_X1 port map( A1 => A(31), A2 => n648, ZN => n162);
   U325 : OAI221_X1 port map( B1 => n29, B2 => n86, C1 => n17, C2 => n83, A => 
                           n606, ZN => n184);
   U326 : AOI22_X1 port map( A1 => A(13), A2 => n10, B1 => A(12), B2 => n267, 
                           ZN => n606);
   U327 : OAI221_X1 port map( B1 => n29, B2 => n126, C1 => n17, C2 => n123, A 
                           => n608, ZN => n370);
   U328 : AOI22_X1 port map( A1 => A(25), A2 => n10, B1 => A(24), B2 => n267, 
                           ZN => n608);
   U329 : NAND2_X1 port map( A1 => n488, A2 => n489, ZN => n287);
   U330 : OAI221_X1 port map( B1 => n27, B2 => n117, C1 => n15, C2 => n114, A 
                           => n536, ZN => n168);
   U331 : AOI22_X1 port map( A1 => A(22), A2 => n9, B1 => A(21), B2 => n7, ZN 
                           => n536);
   U332 : OAI221_X1 port map( B1 => n28, B2 => n120, C1 => n16, C2 => n117, A 
                           => n583, ZN => n402);
   U333 : AOI22_X1 port map( A1 => A(23), A2 => n9, B1 => A(22), B2 => n267, ZN
                           => n583);
   U334 : AOI221_X1 port map( B1 => A(1), B2 => n32, C1 => A(2), C2 => n18, A 
                           => n540, ZN => n374);
   U335 : OAI22_X1 port map( A1 => n615, A2 => n1, B1 => n617, B2 => n8, ZN => 
                           n540);
   U336 : NAND2_X1 port map( A1 => A(31), A2 => n152, ZN => n153);
   U337 : NAND2_X1 port map( A1 => A(31), A2 => n146, ZN => n147);
   U338 : NOR2_X2 port map( A1 => n612, A2 => n591, ZN => n144);
   U339 : OAI221_X1 port map( B1 => n28, B2 => n266, C1 => n16, C2 => n131, A 
                           => n564, ZN => n506);
   U340 : AOI22_X1 port map( A1 => A(28), A2 => n9, B1 => A(27), B2 => n7, ZN 
                           => n564);
   U341 : OAI221_X1 port map( B1 => n28, B2 => n123, C1 => n16, C2 => n120, A 
                           => n565, ZN => n453);
   U342 : AOI22_X1 port map( A1 => A(24), A2 => n9, B1 => A(23), B2 => n7, ZN 
                           => n565);
   U343 : NOR2_X2 port map( A1 => n647, A2 => B(2), ZN => n260);
   U344 : OAI221_X1 port map( B1 => n26, B2 => n114, C1 => n14, C2 => n111, A 
                           => n611, ZN => n185);
   U345 : AOI22_X1 port map( A1 => A(21), A2 => n11, B1 => A(20), B2 => n6, ZN 
                           => n611);
   U346 : AOI222_X1 port map( A1 => n429, A2 => n5, B1 => n620, B2 => n262, C1 
                           => n227, C2 => B(3), ZN => n327);
   U347 : INV_X1 port map( A => n376, ZN => n620);
   U348 : OAI221_X1 port map( B1 => n26, B2 => n77, C1 => n15, C2 => n74, A => 
                           n444, ZN => n154);
   U349 : AOI22_X1 port map( A1 => A(10), A2 => n11, B1 => A(9), B2 => n6, ZN 
                           => n444);
   U350 : OAI221_X1 port map( B1 => n29, B2 => n80, C1 => n16, C2 => n77, A => 
                           n586, ZN => n305);
   U351 : AOI22_X1 port map( A1 => A(11), A2 => n10, B1 => A(10), B2 => n267, 
                           ZN => n586);
   U352 : OAI221_X1 port map( B1 => n28, B2 => n83, C1 => n16, C2 => n80, A => 
                           n567, ZN => n261);
   U353 : AOI22_X1 port map( A1 => A(12), A2 => n9, B1 => A(11), B2 => n7, ZN 
                           => n567);
   U354 : OAI221_X1 port map( B1 => n26, B2 => n623, C1 => n14, C2 => n622, A 
                           => n443, ZN => n219);
   U355 : AOI22_X1 port map( A1 => A(6), A2 => n11, B1 => A(5), B2 => n7, ZN =>
                           n443);
   U356 : OAI221_X1 port map( B1 => n26, B2 => n624, C1 => n14, C2 => n623, A 
                           => n306, ZN => n207);
   U357 : AOI22_X1 port map( A1 => A(7), A2 => n11, B1 => A(6), B2 => n6, ZN =>
                           n306);
   U358 : OAI221_X1 port map( B1 => n27, B2 => n66, C1 => n15, C2 => n624, A =>
                           n265, ZN => n193);
   U359 : AOI22_X1 port map( A1 => A(8), A2 => n10, B1 => A(7), B2 => n6, ZN =>
                           n265);
   U360 : OAI221_X1 port map( B1 => n29, B2 => n100, C1 => n17, C2 => n96, A =>
                           n610, ZN => n186);
   U361 : AOI22_X1 port map( A1 => A(17), A2 => n10, B1 => A(16), B2 => n267, 
                           ZN => n610);
   U362 : OAI221_X1 port map( B1 => n29, B2 => n74, C1 => n17, C2 => n66, A => 
                           n604, ZN => n178);
   U363 : AOI22_X1 port map( A1 => A(9), A2 => n10, B1 => A(8), B2 => n267, ZN 
                           => n604);
   U364 : OAI221_X1 port map( B1 => n27, B2 => n88, C1 => n15, C2 => n86, A => 
                           n537, ZN => n166);
   U365 : AOI22_X1 port map( A1 => A(14), A2 => n11, B1 => A(13), B2 => n7, ZN 
                           => n537);
   U366 : OAI221_X1 port map( B1 => n28, B2 => n92, C1 => n16, C2 => n88, A => 
                           n584, ZN => n516);
   U367 : AOI22_X1 port map( A1 => A(15), A2 => n9, B1 => A(14), B2 => n7, ZN 
                           => n584);
   U368 : OAI221_X1 port map( B1 => n27, B2 => n80, C1 => n15, C2 => n83, A => 
                           n494, ZN => n373);
   U369 : AOI22_X1 port map( A1 => A(15), A2 => n9, B1 => A(16), B2 => n6, ZN 
                           => n494);
   U370 : OAI221_X1 port map( B1 => n27, B2 => n133, C1 => n15, C2 => n615, A 
                           => n523, ZN => n420);
   U371 : AOI22_X1 port map( A1 => A(4), A2 => n10, B1 => A(5), B2 => n7, ZN =>
                           n523);
   U372 : OAI221_X1 port map( B1 => n28, B2 => n615, C1 => n16, C2 => n617, A 
                           => n571, ZN => n407);
   U373 : AOI22_X1 port map( A1 => A(5), A2 => n9, B1 => A(6), B2 => n7, ZN => 
                           n571);
   U374 : OAI221_X1 port map( B1 => n28, B2 => n617, C1 => n16, C2 => n619, A 
                           => n554, ZN => n389);
   U375 : AOI22_X1 port map( A1 => A(6), A2 => n9, B1 => A(7), B2 => n7, ZN => 
                           n554);
   U376 : OAI221_X1 port map( B1 => n49, B2 => n29, C1 => n103, C2 => n14, A =>
                           n553, ZN => n390);
   U377 : AOI22_X1 port map( A1 => A(2), A2 => n9, B1 => A(3), B2 => n7, ZN => 
                           n553);
   U378 : OAI221_X1 port map( B1 => n28, B2 => n624, C1 => n16, C2 => n66, A =>
                           n542, ZN => n429);
   U379 : AOI22_X1 port map( A1 => A(11), A2 => n9, B1 => A(12), B2 => n7, ZN 
                           => n542);
   U380 : OAI221_X1 port map( B1 => n28, B2 => n111, C1 => n16, C2 => n108, A 
                           => n566, ZN => n452);
   U381 : AOI22_X1 port map( A1 => A(20), A2 => n9, B1 => A(19), B2 => n7, ZN 
                           => n566);
   U382 : OAI221_X1 port map( B1 => n28, B2 => n105, C1 => n16, C2 => n100, A 
                           => n538, ZN => n170);
   U383 : AOI22_X1 port map( A1 => A(18), A2 => n9, B1 => A(17), B2 => n7, ZN 
                           => n538);
   U384 : OAI221_X1 port map( B1 => n28, B2 => n108, C1 => n16, C2 => n105, A 
                           => n582, ZN => n464);
   U385 : AOI22_X1 port map( A1 => A(19), A2 => n10, B1 => A(18), B2 => n7, ZN 
                           => n582);
   U386 : INV_X1 port map( A => A(31), ZN => n613);
   U387 : AOI22_X1 port map( A1 => n267, A2 => A(1), B1 => n11, B2 => A(0), ZN 
                           => n362);
   U389 : NAND2_X1 port map( A1 => B(4), A2 => n579, ZN => n160);
   U390 : OAI222_X1 port map( A1 => n79, A2 => n636, B1 => n326, B2 => n642, C1
                           => n91, C2 => n645, ZN => n325);
   U391 : AOI222_X1 port map( A1 => A(27), A2 => n10, B1 => A(25), B2 => n30, 
                           C1 => A(26), C2 => n18, ZN => n326);
   U392 : AOI222_X1 port map( A1 => A(28), A2 => n10, B1 => A(26), B2 => n30, 
                           C1 => A(27), C2 => n19, ZN => n316);
   U393 : AOI222_X1 port map( A1 => A(29), A2 => n11, B1 => A(27), B2 => n32, 
                           C1 => A(28), C2 => n18, ZN => n292);
   U394 : AOI222_X1 port map( A1 => A(30), A2 => n11, B1 => A(28), B2 => n30, 
                           C1 => A(29), C2 => n22, ZN => n273);
   U395 : AOI21_X1 port map( B1 => A(31), B2 => B(11), A => n487, ZN => n256);
   U396 : AOI21_X1 port map( B1 => A(31), B2 => B(25), A => n483, ZN => n250);
   U397 : OAI222_X1 port map( A1 => n171, A2 => n36, B1 => n55, B2 => n626, C1 
                           => n623, C2 => n33, ZN => RES(8));
   U398 : INV_X1 port map( A => n172, ZN => n55);
   U399 : AOI221_X1 port map( B1 => n140, B2 => n173, C1 => n142, C2 => n174, A
                           => n144, ZN => n171);
   U400 : OAI21_X1 port map( B1 => n175, B2 => n146, A => n147, ZN => n174);
   U401 : OAI222_X1 port map( A1 => n187, A2 => n36, B1 => n188, B2 => n626, C1
                           => n622, C2 => n33, ZN => RES(7));
   U402 : AOI221_X1 port map( B1 => n140, B2 => n61, C1 => n142, C2 => n189, A 
                           => n144, ZN => n187);
   U403 : INV_X1 port map( A => n198, ZN => n61);
   U404 : OAI21_X1 port map( B1 => n190, B2 => n146, A => n147, ZN => n189);
   U405 : OAI222_X1 port map( A1 => n136, A2 => n36, B1 => n59, B2 => n626, C1 
                           => n624, C2 => n33, ZN => RES(9));
   U406 : INV_X1 port map( A => n139, ZN => n59);
   U407 : AOI221_X1 port map( B1 => n140, B2 => n141, C1 => n142, C2 => n143, A
                           => n144, ZN => n136);
   U408 : OAI21_X1 port map( B1 => n145, B2 => n146, A => n147, ZN => n143);
   U409 : OAI222_X1 port map( A1 => n539, A2 => n36, B1 => n327, B2 => n626, C1
                           => n77, C2 => n35, ZN => RES(12));
   U410 : AOI221_X1 port map( B1 => n140, B2 => n543, C1 => n142, C2 => n544, A
                           => n144, ZN => n539);
   U411 : OAI21_X1 port map( B1 => n545, B2 => n146, A => n147, ZN => n544);
   U412 : OAI221_X1 port map( B1 => n90, B2 => n638, C1 => n78, C2 => n642, A 
                           => n550, ZN => n543);
   U413 : OAI222_X1 port map( A1 => n521, A2 => n36, B1 => n57, B2 => n626, C1 
                           => n80, C2 => n35, ZN => RES(13));
   U414 : INV_X1 port map( A => n314, ZN => n57);
   U415 : AOI221_X1 port map( B1 => n140, B2 => n526, C1 => n142, C2 => n527, A
                           => n144, ZN => n521);
   U416 : OAI21_X1 port map( B1 => n528, B2 => n146, A => n147, ZN => n527);
   U417 : OAI222_X1 port map( A1 => n508, A2 => n36, B1 => n51, B2 => n626, C1 
                           => n83, C2 => n35, ZN => RES(14));
   U418 : INV_X1 port map( A => n290, ZN => n51);
   U419 : AOI221_X1 port map( B1 => n140, B2 => n511, C1 => n142, C2 => n512, A
                           => n144, ZN => n508);
   U420 : OAI21_X1 port map( B1 => n513, B2 => n146, A => n147, ZN => n512);
   U421 : OAI222_X1 port map( A1 => n551, A2 => n36, B1 => n45, B2 => n626, C1 
                           => n74, C2 => n35, ZN => RES(11));
   U422 : INV_X1 port map( A => n337, ZN => n45);
   U423 : AOI221_X1 port map( B1 => n140, B2 => n555, C1 => n142, C2 => n556, A
                           => n144, ZN => n551);
   U424 : OAI21_X1 port map( B1 => n557, B2 => n146, A => n147, ZN => n556);
   U425 : OAI222_X1 port map( A1 => n495, A2 => n36, B1 => n47, B2 => n626, C1 
                           => n86, C2 => n35, ZN => RES(15));
   U426 : INV_X1 port map( A => n271, ZN => n47);
   U427 : AOI221_X1 port map( B1 => n140, B2 => n498, C1 => n142, C2 => n499, A
                           => n144, ZN => n495);
   U429 : OAI21_X1 port map( B1 => n500, B2 => n146, A => n147, ZN => n499);
   U430 : OAI222_X1 port map( A1 => n569, A2 => n36, B1 => n53, B2 => n626, C1 
                           => n66, C2 => n35, ZN => RES(10));
   U431 : INV_X1 port map( A => n348, ZN => n53);
   U432 : AOI221_X1 port map( B1 => n140, B2 => n572, C1 => n142, C2 => n573, A
                           => n144, ZN => n569);
   U433 : OAI21_X1 port map( B1 => n574, B2 => n146, A => n147, ZN => n573);
   U434 : OAI222_X1 port map( A1 => n201, A2 => n36, B1 => n202, B2 => n626, C1
                           => n621, C2 => n33, ZN => RES(6));
   U435 : AOI221_X1 port map( B1 => n140, B2 => n67, C1 => n142, C2 => n203, A 
                           => n144, ZN => n201);
   U436 : INV_X1 port map( A => n210, ZN => n67);
   U437 : OAI21_X1 port map( B1 => n204, B2 => n146, A => n147, ZN => n203);
   U438 : OAI222_X1 port map( A1 => n213, A2 => n36, B1 => n214, B2 => n626, C1
                           => n619, C2 => n33, ZN => RES(5));
   U439 : AOI221_X1 port map( B1 => n140, B2 => n70, C1 => n142, C2 => n215, A 
                           => n144, ZN => n213);
   U440 : INV_X1 port map( A => n222, ZN => n70);
   U441 : OAI21_X1 port map( B1 => n216, B2 => n146, A => n147, ZN => n215);
   U442 : OAI221_X1 port map( B1 => n27, B2 => n83, C1 => n15, C2 => n86, A => 
                           n476, ZN => n419);
   U443 : AOI22_X1 port map( A1 => A(16), A2 => n11, B1 => A(17), B2 => n6, ZN 
                           => n476);
   U444 : OAI221_X1 port map( B1 => n27, B2 => n86, C1 => n15, C2 => n88, A => 
                           n467, ZN => n406);
   U445 : AOI22_X1 port map( A1 => A(17), A2 => n9, B1 => A(18), B2 => n7, ZN 
                           => n467);
   U446 : OAI221_X1 port map( B1 => n27, B2 => n88, C1 => n15, C2 => n92, A => 
                           n457, ZN => n388);
   U447 : AOI22_X1 port map( A1 => A(18), A2 => n10, B1 => A(19), B2 => n6, ZN 
                           => n457);
   U448 : OAI221_X1 port map( B1 => n26, B2 => n92, C1 => n14, C2 => n96, A => 
                           n430, ZN => n372);
   U449 : AOI22_X1 port map( A1 => A(19), A2 => n11, B1 => A(20), B2 => n6, ZN 
                           => n430);
   U450 : OAI221_X1 port map( B1 => n29, B2 => n622, C1 => n17, C2 => n621, A 
                           => n605, ZN => n234);
   U451 : AOI22_X1 port map( A1 => A(5), A2 => n10, B1 => A(4), B2 => n267, ZN 
                           => n605);
   U452 : OAI221_X1 port map( B1 => n258, B2 => n643, C1 => n196, C2 => n637, A
                           => n259, ZN => n247);
   U453 : AOI22_X1 port map( A1 => n260, A2 => n261, B1 => n262, B2 => n193, ZN
                           => n259);
   U454 : AOI222_X1 port map( A1 => A(4), A2 => n11, B1 => A(6), B2 => n31, C1 
                           => A(5), C2 => n19, ZN => n258);
   U455 : OAI221_X1 port map( B1 => n303, B2 => n643, C1 => n84, C2 => n637, A 
                           => n304, ZN => n298);
   U456 : AOI22_X1 port map( A1 => n260, A2 => n305, B1 => n262, B2 => n207, ZN
                           => n304);
   U457 : AOI222_X1 port map( A1 => A(3), A2 => n10, B1 => A(5), B2 => n32, C1 
                           => A(4), C2 => n19, ZN => n303);
   U458 : OAI221_X1 port map( B1 => n441, B2 => n643, C1 => n81, C2 => n637, A 
                           => n442, ZN => n435);
   U459 : AOI22_X1 port map( A1 => n260, A2 => n154, B1 => n262, B2 => n219, ZN
                           => n442);
   U460 : AOI222_X1 port map( A1 => A(2), A2 => n10, B1 => A(4), B2 => n30, C1 
                           => A(3), C2 => n20, ZN => n441);
   U462 : INV_X1 port map( A => n228, ZN => n626);
   U463 : OAI221_X1 port map( B1 => n27, B2 => n66, C1 => n15, C2 => n74, A => 
                           n524, ZN => n474);
   U464 : AOI22_X1 port map( A1 => A(12), A2 => n11, B1 => A(13), B2 => n7, ZN 
                           => n524);
   U465 : OAI221_X1 port map( B1 => n27, B2 => n74, C1 => n15, C2 => n77, A => 
                           n510, ZN => n465);
   U466 : AOI22_X1 port map( A1 => A(13), A2 => n9, B1 => A(14), B2 => n6, ZN 
                           => n510);
   U467 : OAI221_X1 port map( B1 => n27, B2 => n77, C1 => n15, C2 => n80, A => 
                           n497, ZN => n455);
   U468 : AOI22_X1 port map( A1 => A(14), A2 => n10, B1 => A(15), B2 => n7, ZN 
                           => n497);
   U469 : OAI221_X1 port map( B1 => n26, B2 => n96, C1 => n14, C2 => n100, A =>
                           n421, ZN => n361);
   U470 : AOI22_X1 port map( A1 => A(20), A2 => n11, B1 => A(21), B2 => n6, ZN 
                           => n421);
   U471 : OAI221_X1 port map( B1 => n26, B2 => n100, C1 => n14, C2 => n105, A 
                           => n408, ZN => n350);
   U472 : AOI22_X1 port map( A1 => A(21), A2 => n11, B1 => A(22), B2 => n6, ZN 
                           => n408);
   U473 : OAI221_X1 port map( B1 => n26, B2 => n105, C1 => n14, C2 => n108, A 
                           => n391, ZN => n339);
   U474 : AOI22_X1 port map( A1 => A(22), A2 => n9, B1 => A(23), B2 => n6, ZN 
                           => n391);
   U475 : OAI221_X1 port map( B1 => n26, B2 => n108, C1 => n14, C2 => n111, A 
                           => n377, ZN => n324);
   U476 : AOI22_X1 port map( A1 => A(23), A2 => n9, B1 => A(24), B2 => n6, ZN 
                           => n377);
   U477 : OAI221_X1 port map( B1 => n26, B2 => n111, C1 => n14, C2 => n114, A 
                           => n364, ZN => n313);
   U478 : AOI22_X1 port map( A1 => A(24), A2 => n10, B1 => A(25), B2 => n6, ZN 
                           => n364);
   U479 : OAI221_X1 port map( B1 => n26, B2 => n114, C1 => n14, C2 => n117, A 
                           => n351, ZN => n289);
   U480 : AOI22_X1 port map( A1 => A(25), A2 => n11, B1 => A(26), B2 => n6, ZN 
                           => n351);
   U481 : OAI221_X1 port map( B1 => n26, B2 => n117, C1 => n14, C2 => n120, A 
                           => n340, ZN => n270);
   U482 : AOI22_X1 port map( A1 => A(26), A2 => n10, B1 => A(27), B2 => n6, ZN 
                           => n340);
   U483 : AOI22_X1 port map( A1 => n640, A2 => n506, B1 => B(2), B2 => n382, ZN
                           => n333);
   U484 : AOI21_X1 port map( B1 => n22, B2 => A(31), A => n533, ZN => n412);
   U485 : AOI21_X1 port map( B1 => n11, B2 => A(31), A => n580, ZN => n395);
   U486 : AOI21_X1 port map( B1 => B(1), B2 => A(31), A => n533, ZN => n417);
   U487 : AOI21_X1 port map( B1 => n8, B2 => A(31), A => n580, ZN => n400);
   U488 : NOR2_X1 port map( A1 => n490, A2 => B(18), ZN => n251);
   U489 : OAI22_X1 port map( A1 => B(2), A2 => n374, B1 => n640, B2 => n375, ZN
                           => n227);
   U490 : OAI221_X1 port map( B1 => n196, B2 => n638, C1 => n75, C2 => n642, A 
                           => n562, ZN => n555);
   U491 : AOI221_X1 port map( B1 => n169, B2 => n452, C1 => n167, C2 => n453, A
                           => n563, ZN => n562);
   U492 : NOR3_X1 port map( A1 => n41, A2 => B(3), A3 => n333, ZN => n563);
   U493 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n267);
   U494 : AOI21_X1 port map( B1 => n634, B2 => n590, A => n144, ZN => n481);
   U495 : INV_X1 port map( A => n592, ZN => n634);
   U496 : NAND2_X1 port map( A1 => A(31), A2 => n490, ZN => n486);
   U497 : OAI221_X1 port map( B1 => n225, B2 => n36, C1 => n617, C2 => n33, A 
                           => n226, ZN => RES(4));
   U498 : AOI221_X1 port map( B1 => n140, B2 => n229, C1 => n142, C2 => n230, A
                           => n144, ZN => n225);
   U499 : OAI21_X1 port map( B1 => n231, B2 => n146, A => n147, ZN => n230);
   U500 : NAND2_X1 port map( A1 => n454, A2 => A(31), ZN => n401);
   U501 : NOR2_X1 port map( A1 => B(2), A2 => B(3), ZN => n356);
   U502 : AOI21_X1 port map( B1 => n148, B2 => n501, A => n150, ZN => n500);
   U503 : OAI21_X1 port map( B1 => n502, B2 => n152, A => n153, ZN => n501);
   U504 : AOI211_X1 port map( C1 => B(4), C2 => A(31), A => n503, B => n504, ZN
                           => n502);
   U505 : OAI22_X1 port map( A1 => n196, A2 => n505, B1 => n101, B2 => n157, ZN
                           => n504);
   U506 : INV_X1 port map( A => A(10), ZN => n66);
   U507 : OAI21_X1 port map( B1 => n489, B2 => n613, A => n162, ZN => n487);
   U508 : NOR3_X1 port map( A1 => n332, A2 => B(3), A3 => n333, ZN => n331);
   U509 : INV_X1 port map( A => B(3), ZN => n647);
   U510 : INV_X1 port map( A => A(11), ZN => n74);
   U511 : INV_X1 port map( A => A(15), ZN => n86);
   U512 : INV_X1 port map( A => A(9), ZN => n624);
   U513 : INV_X1 port map( A => A(16), ZN => n88);
   U514 : BUF_X1 port map( A => n137, Z => n36);
   U515 : BUF_X1 port map( A => n137, Z => n37);
   U516 : NAND2_X1 port map( A1 => A(0), A2 => n6, ZN => n375);
   U517 : INV_X1 port map( A => A(23), ZN => n114);
   U518 : INV_X1 port map( A => A(19), ZN => n100);
   U519 : INV_X1 port map( A => A(24), ZN => n117);
   U520 : INV_X1 port map( A => A(20), ZN => n105);
   U521 : INV_X1 port map( A => A(21), ZN => n108);
   U522 : INV_X1 port map( A => A(22), ZN => n111);
   U523 : INV_X1 port map( A => A(8), ZN => n623);
   U524 : INV_X1 port map( A => A(12), ZN => n77);
   U525 : INV_X1 port map( A => A(13), ZN => n80);
   U526 : INV_X1 port map( A => A(14), ZN => n83);
   U527 : INV_X1 port map( A => A(30), ZN => n266);
   U528 : INV_X1 port map( A => A(3), ZN => n615);
   U529 : OR4_X1 port map( A1 => B(13), A2 => B(14), A3 => B(12), A4 => n596, 
                           ZN => n490);
   U530 : OR3_X1 port map( A1 => B(15), A2 => B(17), A3 => B(16), ZN => n596);
   U531 : INV_X1 port map( A => B(2), ZN => n640);
   U532 : INV_X1 port map( A => A(17), ZN => n92);
   U533 : INV_X1 port map( A => A(7), ZN => n622);
   U534 : INV_X1 port map( A => A(18), ZN => n96);
   U535 : INV_X1 port map( A => A(25), ZN => n120);
   U536 : AND3_X1 port map( A1 => n579, A2 => n591, A3 => n597, ZN => n445);
   U537 : NOR3_X1 port map( A1 => n152, A2 => n146, A3 => n630, ZN => n597);
   U538 : INV_X1 port map( A => n148, ZN => n630);
   U539 : INV_X1 port map( A => A(4), ZN => n617);
   U540 : INV_X1 port map( A => n590, ZN => n612);
   U541 : INV_X1 port map( A => A(27), ZN => n126);
   U542 : INV_X1 port map( A => A(26), ZN => n123);
   U543 : INV_X1 port map( A => A(6), ZN => n621);
   U544 : INV_X1 port map( A => A(5), ZN => n619);
   U545 : INV_X1 port map( A => A(28), ZN => n128);
   U546 : INV_X1 port map( A => A(29), ZN => n131);
   U547 : INV_X1 port map( A => B(25), ZN => n633);
   U548 : INV_X1 port map( A => A(2), ZN => n133);
   U549 : AND2_X1 port map( A1 => n140, A2 => n199, ZN => n278);
   U550 : INV_X1 port map( A => A(1), ZN => n103);
   U551 : INV_X1 port map( A => n579, ZN => n648);
   U552 : INV_X1 port map( A => A(0), ZN => n49);
   U553 : OR2_X1 port map( A1 => n625, A2 => B(1), ZN => n1);
   U554 : NAND2_X1 port map( A1 => n140, A2 => n40, ZN => n332);
   U555 : INV_X1 port map( A => n436, ZN => n627);
   U556 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n263);
   U557 : NAND2_X1 port map( A1 => B(1), A2 => n625, ZN => n264);
   U558 : INV_X1 port map( A => B(11), ZN => n629);
   U559 : INV_X1 port map( A => B(18), ZN => n631);
   U560 : AND2_X1 port map( A1 => n142, A2 => n592, ZN => n491);
   U561 : BUF_X1 port map( A => n137, Z => n38);
   U562 : INV_X1 port map( A => B(0), ZN => n625);
   U563 : INV_X1 port map( A => B(4), ZN => n44);
   U564 : NOR2_X2 port map( A1 => n635, A2 => LOGIC_ARITH, ZN => n142);
   U565 : INV_X1 port map( A => n591, ZN => n635);
   U566 : NOR3_X1 port map( A1 => B(9), A2 => B(8), A3 => B(10), ZN => n489);
   U567 : NOR3_X1 port map( A1 => B(7), A2 => B(6), A3 => B(5), ZN => n579);
   U568 : NOR3_X1 port map( A1 => B(28), A2 => B(27), A3 => B(26), ZN => n592);
   U569 : OAI222_X1 port map( A1 => n468, A2 => n269, B1 => n469, B2 => n37, C1
                           => n92, C2 => n34, ZN => RES(17));
   U570 : AOI221_X1 port map( B1 => n165, B2 => n474, C1 => n199, C2 => n419, A
                           => n475, ZN => n468);
   U571 : AOI221_X1 port map( B1 => n276, B2 => n470, C1 => n628, C2 => n434, A
                           => n279, ZN => n469);
   U572 : OAI222_X1 port map( A1 => n132, A2 => n636, B1 => n362, B2 => n641, 
                           C1 => n363, C2 => n645, ZN => n475);
   U573 : OAI222_X1 port map( A1 => n458, A2 => n269, B1 => n459, B2 => n38, C1
                           => n96, C2 => n34, ZN => RES(18));
   U574 : AOI221_X1 port map( B1 => n165, B2 => n465, C1 => n199, C2 => n406, A
                           => n466, ZN => n458);
   U575 : AOI221_X1 port map( B1 => n276, B2 => n460, C1 => n628, C2 => n297, A
                           => n279, ZN => n459);
   U576 : OAI222_X1 port map( A1 => n614, A2 => n636, B1 => n293, B2 => n641, 
                           C1 => n405, C2 => n645, ZN => n466);
   U577 : OAI222_X1 port map( A1 => n446, A2 => n269, B1 => n447, B2 => n37, C1
                           => n100, C2 => n34, ZN => RES(19));
   U578 : AOI221_X1 port map( B1 => n165, B2 => n455, C1 => n199, C2 => n388, A
                           => n456, ZN => n446);
   U579 : AOI221_X1 port map( B1 => n276, B2 => n448, C1 => n628, C2 => n246, A
                           => n279, ZN => n447);
   U580 : OAI222_X1 port map( A1 => n616, A2 => n636, B1 => n46, B2 => n641, C1
                           => n387, C2 => n645, ZN => n456);
   U581 : OAI222_X1 port map( A1 => n422, A2 => n269, B1 => n423, B2 => n37, C1
                           => n105, C2 => n34, ZN => RES(20));
   U582 : AOI221_X1 port map( B1 => n165, B2 => n373, C1 => n199, C2 => n372, A
                           => n427, ZN => n422);
   U583 : AOI221_X1 port map( B1 => n276, B2 => n424, C1 => n628, C2 => n107, A
                           => n279, ZN => n423);
   U584 : OAI221_X1 port map( B1 => n376, B2 => n636, C1 => n63, C2 => n645, A 
                           => n428, ZN => n427);
   U585 : OAI222_X1 port map( A1 => n409, A2 => n269, B1 => n410, B2 => n37, C1
                           => n108, C2 => n34, ZN => RES(21));
   U586 : AOI221_X1 port map( B1 => n276, B2 => n411, C1 => n628, C2 => n223, A
                           => n279, ZN => n410);
   U587 : AOI221_X1 port map( B1 => n199, B2 => n361, C1 => B(4), C2 => n56, A 
                           => n418, ZN => n409);
   U588 : OAI21_X1 port map( B1 => n414, B2 => n281, A => n282, ZN => n411);
   U589 : OAI222_X1 port map( A1 => n392, A2 => n269, B1 => n393, B2 => n37, C1
                           => n111, C2 => n34, ZN => RES(22));
   U590 : AOI221_X1 port map( B1 => n276, B2 => n394, C1 => n628, C2 => n211, A
                           => n279, ZN => n393);
   U591 : AOI221_X1 port map( B1 => n199, B2 => n350, C1 => B(4), C2 => n50, A 
                           => n404, ZN => n392);
   U592 : OAI21_X1 port map( B1 => n397, B2 => n281, A => n282, ZN => n394);
   U593 : OAI222_X1 port map( A1 => n378, A2 => n269, B1 => n379, B2 => n37, C1
                           => n114, C2 => n34, ZN => RES(23));
   U594 : AOI221_X1 port map( B1 => n276, B2 => n380, C1 => n628, C2 => n115, A
                           => n279, ZN => n379);
   U595 : AOI221_X1 port map( B1 => n199, B2 => n339, C1 => B(4), C2 => n48, A 
                           => n386, ZN => n378);
   U596 : OAI21_X1 port map( B1 => n384, B2 => n281, A => n282, ZN => n380);
   U597 : OAI222_X1 port map( A1 => n365, A2 => n269, B1 => n366, B2 => n37, C1
                           => n117, C2 => n34, ZN => RES(24));
   U598 : AOI221_X1 port map( B1 => n276, B2 => n367, C1 => n628, C2 => n119, A
                           => n279, ZN => n366);
   U599 : AOI221_X1 port map( B1 => n199, B2 => n324, C1 => n39, C2 => n172, A 
                           => n371, ZN => n365);
   U600 : OAI21_X1 port map( B1 => n368, B2 => n281, A => n282, ZN => n367);
   U601 : OAI222_X1 port map( A1 => n352, A2 => n269, B1 => n353, B2 => n37, C1
                           => n120, C2 => n34, ZN => RES(25));
   U602 : AOI221_X1 port map( B1 => n276, B2 => n354, C1 => n628, C2 => n122, A
                           => n279, ZN => n353);
   U603 : AOI221_X1 port map( B1 => n199, B2 => n313, C1 => n39, C2 => n139, A 
                           => n360, ZN => n352);
   U604 : INV_X1 port map( A => n163, ZN => n122);
   U605 : OAI222_X1 port map( A1 => n477, A2 => n269, B1 => n478, B2 => n38, C1
                           => n88, C2 => n35, ZN => RES(16));
   U606 : AOI221_X1 port map( B1 => n165, B2 => n429, C1 => n199, C2 => n373, A
                           => n492, ZN => n477);
   U607 : AOI221_X1 port map( B1 => n276, B2 => n479, C1 => n628, C2 => n480, A
                           => n279, ZN => n478);
   U608 : OAI222_X1 port map( A1 => n374, A2 => n636, B1 => n375, B2 => n641, 
                           C1 => n376, C2 => n645, ZN => n492);
   U609 : OAI222_X1 port map( A1 => n341, A2 => n269, B1 => n342, B2 => n37, C1
                           => n123, C2 => n34, ZN => RES(26));
   U610 : AOI221_X1 port map( B1 => n276, B2 => n343, C1 => n628, C2 => n125, A
                           => n279, ZN => n342);
   U611 : AOI221_X1 port map( B1 => n199, B2 => n289, C1 => n39, C2 => n348, A 
                           => n349, ZN => n341);
   U612 : INV_X1 port map( A => n344, ZN => n125);
   U613 : OAI222_X1 port map( A1 => n328, A2 => n269, B1 => n329, B2 => n37, C1
                           => n126, C2 => n34, ZN => RES(27));
   U614 : AOI211_X1 port map( C1 => n276, C2 => n330, A => n279, B => n331, ZN 
                           => n329);
   U615 : AOI221_X1 port map( B1 => n199, B2 => n270, C1 => n39, C2 => n337, A 
                           => n338, ZN => n328);
   U616 : OAI21_X1 port map( B1 => n334, B2 => n281, A => n282, ZN => n330);
   U617 : OAI222_X1 port map( A1 => n317, A2 => n269, B1 => n318, B2 => n37, C1
                           => n128, C2 => n34, ZN => RES(28));
   U618 : AOI221_X1 port map( B1 => n165, B2 => n324, C1 => n39, C2 => n54, A 
                           => n325, ZN => n317);
   U619 : AOI221_X1 port map( B1 => n276, B2 => n319, C1 => n278, C2 => n320, A
                           => n279, ZN => n318);
   U620 : INV_X1 port map( A => n327, ZN => n54);
   U621 : OAI222_X1 port map( A1 => n307, A2 => n269, B1 => n308, B2 => n37, C1
                           => n131, C2 => n33, ZN => RES(29));
   U622 : AOI221_X1 port map( B1 => n165, B2 => n313, C1 => n39, C2 => n314, A 
                           => n315, ZN => n307);
   U623 : AOI221_X1 port map( B1 => n276, B2 => n309, C1 => n278, C2 => n129, A
                           => n279, ZN => n308);
   U624 : OAI222_X1 port map( A1 => n82, A2 => n636, B1 => n316, B2 => n642, C1
                           => n95, C2 => n645, ZN => n315);
   U625 : OAI222_X1 port map( A1 => n274, A2 => n269, B1 => n275, B2 => n38, C1
                           => n266, C2 => n33, ZN => RES(30));
   U626 : AOI221_X1 port map( B1 => n165, B2 => n289, C1 => n39, C2 => n290, A 
                           => n291, ZN => n274);
   U627 : AOI221_X1 port map( B1 => n276, B2 => n277, C1 => n278, C2 => n134, A
                           => n279, ZN => n275);
   U628 : OAI222_X1 port map( A1 => n85, A2 => n636, B1 => n292, B2 => n642, C1
                           => n99, C2 => n645, ZN => n291);
   U629 : OAI221_X1 port map( B1 => n293, B2 => n240, C1 => n133, C2 => n33, A 
                           => n294, ZN => RES(2));
   U630 : AOI221_X1 port map( B1 => n242, B2 => n295, C1 => n627, C2 => n69, A 
                           => n244, ZN => n294);
   U631 : INV_X1 port map( A => n296, ZN => n69);
   U632 : OAI21_X1 port map( B1 => n299, B2 => n249, A => n250, ZN => n295);
   U633 : OAI221_X1 port map( B1 => n362, B2 => n240, C1 => n103, C2 => n33, A 
                           => n431, ZN => RES(1));
   U634 : AOI221_X1 port map( B1 => n242, B2 => n432, C1 => n627, C2 => n72, A 
                           => n244, ZN => n431);
   U635 : INV_X1 port map( A => n433, ZN => n72);
   U636 : OAI21_X1 port map( B1 => n437, B2 => n249, A => n250, ZN => n432);
   U640 : OAI221_X1 port map( B1 => n46, B2 => n240, C1 => n615, C2 => n33, A 
                           => n241, ZN => RES(3));
   U643 : AOI221_X1 port map( B1 => n242, B2 => n243, C1 => n627, C2 => n60, A 
                           => n244, ZN => n241);
   U644 : INV_X1 port map( A => n245, ZN => n60);
   U645 : OAI21_X1 port map( B1 => n248, B2 => n249, A => n250, ZN => n243);
   U646 : NOR2_X1 port map( A1 => B(29), A2 => B(30), ZN => n591);
   U647 : AND2_X1 port map( A1 => LOGIC_ARITH, A2 => n445, ZN => n140);
   U648 : NOR2_X1 port map( A1 => n613, A2 => LOGIC_ARITH, ZN => n590);
   U649 : OAI221_X1 port map( B1 => n587, B2 => n436, C1 => n49, C2 => n33, A 
                           => n588, ZN => RES(0));
   U650 : NOR2_X1 port map( A1 => n269, A2 => n39, ZN => n228);
   U651 : AOI21_X1 port map( B1 => n242, B2 => n589, A => n244, ZN => n588);
   U652 : OAI21_X1 port map( B1 => n593, B2 => n249, A => n250, ZN => n589);
   U653 : AOI21_X1 port map( B1 => n251, B2 => n595, A => n253, ZN => n593);
   U654 : OAI21_X1 port map( B1 => n587, B2 => n255, A => n256, ZN => n595);
   U655 : AND2_X1 port map( A1 => n491, A2 => n649, ZN => n242);
   U656 : NAND2_X1 port map( A1 => n35, A2 => n649, ZN => n137);
   U657 : NAND2_X1 port map( A1 => n140, A2 => n649, ZN => n436);
   U658 : NOR2_X1 port map( A1 => n481, A2 => LEFT_RIGHT, ZN => n244);
   U659 : INV_X1 port map( A => LEFT_RIGHT, ZN => n649);
   U660 : OAI222_X1 port map( A1 => n268, A2 => n269, B1 => LEFT_RIGHT, B2 => 
                           n612, C1 => n613, C2 => n34, ZN => RES(31));
   U661 : AOI221_X1 port map( B1 => n165, B2 => n270, C1 => n39, C2 => n271, A 
                           => n272, ZN => n268);
   U662 : OAI222_X1 port map( A1 => n87, A2 => n636, B1 => n273, B2 => n642, C1
                           => n104, C2 => n645, ZN => n272);
   U663 : NOR4_X4 port map( A1 => B(16), A2 => B(17), A3 => B(15), A4 => n598, 
                           ZN => n148);
   U664 : INV_X1 port map( A => n8, ZN => n6);
   U665 : INV_X1 port map( A => n8, ZN => n7);
   U666 : INV_X1 port map( A => n1, ZN => n9);
   U667 : INV_X1 port map( A => n1, ZN => n10);
   U668 : INV_X1 port map( A => n1, ZN => n11);
   U669 : CLKBUF_X1 port map( A => n264, Z => n12);
   U670 : CLKBUF_X1 port map( A => n264, Z => n13);
   U671 : INV_X1 port map( A => n19, ZN => n17);
   U672 : INV_X1 port map( A => n12, ZN => n18);
   U673 : INV_X1 port map( A => n12, ZN => n19);
   U674 : INV_X1 port map( A => n264, ZN => n20);
   U675 : INV_X1 port map( A => n13, ZN => n21);
   U676 : INV_X1 port map( A => n13, ZN => n22);
   U677 : CLKBUF_X1 port map( A => n263, Z => n23);
   U678 : CLKBUF_X1 port map( A => n263, Z => n24);
   U679 : CLKBUF_X1 port map( A => n263, Z => n25);
   U680 : INV_X1 port map( A => n23, ZN => n30);
   U681 : INV_X1 port map( A => n24, ZN => n31);
   U682 : INV_X1 port map( A => n25, ZN => n32);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity comparator_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  OPSel : in std_logic_vector
         (0 to 2);  RES : out std_logic_vector (31 downto 0));

end comparator_NBIT32;

architecture SYN_bhv of comparator_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component comparator_NBIT32_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   signal X_Logic0_port, N26, N27, N28, N29, N30, N31, n10, n15, n16, n17, n18,
      n19, n20, RES_0_port, n2, n3, n4 : std_logic;

begin
   RES <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, RES_0_port 
      );
   
   X_Logic0_port <= '0';
   n10 <= '0';
   r57 : comparator_NBIT32_DW01_cmp6_0 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), TC => n10, LT => N30, GT => N28,
                           EQ => N26, LE => N31, GE => N29, NE => N27);
   U3 : INV_X1 port map( A => n15, ZN => RES_0_port);
   U4 : AOI21_X1 port map( B1 => n16, B2 => n4, A => n17, ZN => n15);
   U5 : INV_X1 port map( A => OPSel(2), ZN => n3);
   U6 : OAI22_X1 port map( A1 => n19, A2 => n2, B1 => OPSel(1), B2 => n20, ZN 
                           => n16);
   U7 : INV_X1 port map( A => OPSel(1), ZN => n2);
   U8 : AOI22_X1 port map( A1 => N28, A2 => n3, B1 => N29, B2 => OPSel(2), ZN 
                           => n19);
   U9 : AOI22_X1 port map( A1 => N26, A2 => n3, B1 => N27, B2 => OPSel(2), ZN 
                           => n20);
   U10 : NOR3_X1 port map( A1 => n4, A2 => OPSel(1), A3 => n18, ZN => n17);
   U11 : AOI22_X1 port map( A1 => N30, A2 => n3, B1 => OPSel(2), B2 => N31, ZN 
                           => n18);
   U12 : INV_X1 port map( A => OPSel(0), ZN => n4);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ALU_NBIT32 is

   port( OP1, OP2 : in std_logic_vector (31 downto 0);  ALU_OPC : in 
         std_logic_vector (0 to 4);  ALU_RES : out std_logic_vector (31 downto 
         0));

end ALU_NBIT32;

architecture SYN_struct of ALU_NBIT32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux21_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux41_NBIT32_1
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component BOOTHMUL_numBit16
      port( A, B : in std_logic_vector (15 downto 0);  P : out std_logic_vector
            (31 downto 0));
   end component;
   
   component P4Adder_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component shifter_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  LOGIC_ARITH, LEFT_RIGHT 
            : in std_logic;  RES : out std_logic_vector (31 downto 0));
   end component;
   
   component comparator_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  OPSel : in 
            std_logic_vector (0 to 2);  RES : out std_logic_vector (31 downto 
            0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, select_type_sig_1_port, select_type_sig_0_port, 
      select_zero_sig, A_CMP_31_port, A_CMP_30_port, A_CMP_29_port, 
      A_CMP_28_port, A_CMP_27_port, A_CMP_26_port, A_CMP_25_port, A_CMP_24_port
      , A_CMP_23_port, A_CMP_22_port, A_CMP_21_port, A_CMP_20_port, 
      A_CMP_19_port, A_CMP_18_port, A_CMP_17_port, A_CMP_16_port, A_CMP_15_port
      , A_CMP_14_port, A_CMP_13_port, A_CMP_12_port, A_CMP_11_port, 
      A_CMP_10_port, A_CMP_9_port, A_CMP_8_port, A_CMP_7_port, A_CMP_6_port, 
      A_CMP_5_port, A_CMP_4_port, A_CMP_3_port, A_CMP_2_port, A_CMP_1_port, 
      A_CMP_0_port, B_CMP_31_port, B_CMP_30_port, B_CMP_29_port, B_CMP_28_port,
      B_CMP_27_port, B_CMP_26_port, B_CMP_25_port, B_CMP_24_port, B_CMP_23_port
      , B_CMP_22_port, B_CMP_21_port, B_CMP_20_port, B_CMP_19_port, 
      B_CMP_18_port, B_CMP_17_port, B_CMP_16_port, B_CMP_15_port, B_CMP_14_port
      , B_CMP_13_port, B_CMP_12_port, B_CMP_11_port, B_CMP_10_port, 
      B_CMP_9_port, B_CMP_8_port, B_CMP_7_port, B_CMP_6_port, B_CMP_5_port, 
      B_CMP_4_port, B_CMP_3_port, B_CMP_2_port, B_CMP_1_port, B_CMP_0_port, 
      A_SHF_31_port, A_SHF_30_port, A_SHF_29_port, A_SHF_28_port, A_SHF_27_port
      , A_SHF_26_port, A_SHF_25_port, A_SHF_24_port, A_SHF_23_port, 
      A_SHF_22_port, A_SHF_21_port, A_SHF_20_port, A_SHF_19_port, A_SHF_18_port
      , A_SHF_17_port, A_SHF_16_port, A_SHF_15_port, A_SHF_14_port, 
      A_SHF_13_port, A_SHF_12_port, A_SHF_11_port, A_SHF_10_port, A_SHF_9_port,
      A_SHF_8_port, A_SHF_7_port, A_SHF_6_port, A_SHF_5_port, A_SHF_4_port, 
      A_SHF_3_port, A_SHF_2_port, A_SHF_1_port, A_SHF_0_port, B_SHF_31_port, 
      B_SHF_30_port, B_SHF_29_port, B_SHF_28_port, B_SHF_27_port, B_SHF_26_port
      , B_SHF_25_port, B_SHF_24_port, B_SHF_23_port, B_SHF_22_port, 
      B_SHF_21_port, B_SHF_20_port, B_SHF_19_port, B_SHF_18_port, B_SHF_17_port
      , B_SHF_16_port, B_SHF_15_port, B_SHF_14_port, B_SHF_13_port, 
      B_SHF_12_port, B_SHF_11_port, B_SHF_10_port, B_SHF_9_port, B_SHF_8_port, 
      B_SHF_7_port, B_SHF_6_port, B_SHF_5_port, B_SHF_4_port, B_SHF_3_port, 
      B_SHF_2_port, B_SHF_1_port, B_SHF_0_port, A_ADD_31_port, A_ADD_30_port, 
      A_ADD_29_port, A_ADD_28_port, A_ADD_27_port, A_ADD_26_port, A_ADD_25_port
      , A_ADD_24_port, A_ADD_23_port, A_ADD_22_port, A_ADD_21_port, 
      A_ADD_20_port, A_ADD_19_port, A_ADD_18_port, A_ADD_17_port, A_ADD_16_port
      , A_ADD_15_port, A_ADD_14_port, A_ADD_13_port, A_ADD_12_port, 
      A_ADD_11_port, A_ADD_10_port, A_ADD_9_port, A_ADD_8_port, A_ADD_7_port, 
      A_ADD_6_port, A_ADD_5_port, A_ADD_4_port, A_ADD_3_port, A_ADD_2_port, 
      A_ADD_1_port, A_ADD_0_port, B_ADD_31_port, B_ADD_30_port, B_ADD_29_port, 
      B_ADD_28_port, B_ADD_27_port, B_ADD_26_port, B_ADD_25_port, B_ADD_24_port
      , B_ADD_23_port, B_ADD_22_port, B_ADD_21_port, B_ADD_20_port, 
      B_ADD_19_port, B_ADD_18_port, B_ADD_17_port, B_ADD_16_port, B_ADD_15_port
      , B_ADD_14_port, B_ADD_13_port, B_ADD_12_port, B_ADD_11_port, 
      B_ADD_10_port, B_ADD_9_port, B_ADD_8_port, B_ADD_7_port, B_ADD_6_port, 
      B_ADD_5_port, B_ADD_4_port, B_ADD_3_port, B_ADD_2_port, B_ADD_1_port, 
      B_ADD_0_port, A_MUL_15_port, A_MUL_14_port, A_MUL_13_port, A_MUL_12_port,
      A_MUL_11_port, A_MUL_10_port, A_MUL_9_port, A_MUL_8_port, A_MUL_7_port, 
      A_MUL_6_port, A_MUL_5_port, A_MUL_4_port, A_MUL_3_port, A_MUL_2_port, 
      A_MUL_1_port, A_MUL_0_port, B_MUL_15_port, B_MUL_14_port, B_MUL_13_port, 
      B_MUL_12_port, B_MUL_11_port, B_MUL_10_port, B_MUL_9_port, B_MUL_8_port, 
      B_MUL_7_port, B_MUL_6_port, B_MUL_5_port, B_MUL_4_port, B_MUL_3_port, 
      B_MUL_2_port, B_MUL_1_port, B_MUL_0_port, LOGIC_ARITH, LEFT_RIGHT, 
      OPSel_1_port, OPSel_0_port, ADD_SUB, LOGIC_RES_31_port, LOGIC_RES_30_port
      , LOGIC_RES_29_port, LOGIC_RES_28_port, LOGIC_RES_27_port, 
      LOGIC_RES_26_port, LOGIC_RES_25_port, LOGIC_RES_24_port, 
      LOGIC_RES_23_port, LOGIC_RES_22_port, LOGIC_RES_21_port, 
      LOGIC_RES_20_port, LOGIC_RES_19_port, LOGIC_RES_18_port, 
      LOGIC_RES_17_port, LOGIC_RES_16_port, LOGIC_RES_15_port, 
      LOGIC_RES_14_port, LOGIC_RES_13_port, LOGIC_RES_12_port, 
      LOGIC_RES_11_port, LOGIC_RES_10_port, LOGIC_RES_9_port, LOGIC_RES_8_port,
      LOGIC_RES_7_port, LOGIC_RES_6_port, LOGIC_RES_5_port, LOGIC_RES_4_port, 
      LOGIC_RES_3_port, LOGIC_RES_2_port, LOGIC_RES_1_port, LOGIC_RES_0_port, 
      COMP_RES_31_port, COMP_RES_30_port, COMP_RES_29_port, COMP_RES_28_port, 
      COMP_RES_27_port, COMP_RES_26_port, COMP_RES_25_port, COMP_RES_24_port, 
      COMP_RES_23_port, COMP_RES_22_port, COMP_RES_21_port, COMP_RES_20_port, 
      COMP_RES_19_port, COMP_RES_18_port, COMP_RES_17_port, COMP_RES_16_port, 
      COMP_RES_15_port, COMP_RES_14_port, COMP_RES_13_port, COMP_RES_12_port, 
      COMP_RES_11_port, COMP_RES_10_port, COMP_RES_9_port, COMP_RES_8_port, 
      COMP_RES_7_port, COMP_RES_6_port, COMP_RES_5_port, COMP_RES_4_port, 
      COMP_RES_3_port, COMP_RES_2_port, COMP_RES_1_port, COMP_RES_0_port, 
      SHIFT_RES_31_port, SHIFT_RES_30_port, SHIFT_RES_29_port, 
      SHIFT_RES_28_port, SHIFT_RES_27_port, SHIFT_RES_26_port, 
      SHIFT_RES_25_port, SHIFT_RES_24_port, SHIFT_RES_23_port, 
      SHIFT_RES_22_port, SHIFT_RES_21_port, SHIFT_RES_20_port, 
      SHIFT_RES_19_port, SHIFT_RES_18_port, SHIFT_RES_17_port, 
      SHIFT_RES_16_port, SHIFT_RES_15_port, SHIFT_RES_14_port, 
      SHIFT_RES_13_port, SHIFT_RES_12_port, SHIFT_RES_11_port, 
      SHIFT_RES_10_port, SHIFT_RES_9_port, SHIFT_RES_8_port, SHIFT_RES_7_port, 
      SHIFT_RES_6_port, SHIFT_RES_5_port, SHIFT_RES_4_port, SHIFT_RES_3_port, 
      SHIFT_RES_2_port, SHIFT_RES_1_port, SHIFT_RES_0_port, ADD_SUB_RES_31_port
      , ADD_SUB_RES_30_port, ADD_SUB_RES_29_port, ADD_SUB_RES_28_port, 
      ADD_SUB_RES_27_port, ADD_SUB_RES_26_port, ADD_SUB_RES_25_port, 
      ADD_SUB_RES_24_port, ADD_SUB_RES_23_port, ADD_SUB_RES_22_port, 
      ADD_SUB_RES_21_port, ADD_SUB_RES_20_port, ADD_SUB_RES_19_port, 
      ADD_SUB_RES_18_port, ADD_SUB_RES_17_port, ADD_SUB_RES_16_port, 
      ADD_SUB_RES_15_port, ADD_SUB_RES_14_port, ADD_SUB_RES_13_port, 
      ADD_SUB_RES_12_port, ADD_SUB_RES_11_port, ADD_SUB_RES_10_port, 
      ADD_SUB_RES_9_port, ADD_SUB_RES_8_port, ADD_SUB_RES_7_port, 
      ADD_SUB_RES_6_port, ADD_SUB_RES_5_port, ADD_SUB_RES_4_port, 
      ADD_SUB_RES_3_port, ADD_SUB_RES_2_port, ADD_SUB_RES_1_port, 
      ADD_SUB_RES_0_port, MUL_RES_31_port, MUL_RES_30_port, MUL_RES_29_port, 
      MUL_RES_28_port, MUL_RES_27_port, MUL_RES_26_port, MUL_RES_25_port, 
      MUL_RES_24_port, MUL_RES_23_port, MUL_RES_22_port, MUL_RES_21_port, 
      MUL_RES_20_port, MUL_RES_19_port, MUL_RES_18_port, MUL_RES_17_port, 
      MUL_RES_16_port, MUL_RES_15_port, MUL_RES_14_port, MUL_RES_13_port, 
      MUL_RES_12_port, MUL_RES_11_port, MUL_RES_10_port, MUL_RES_9_port, 
      MUL_RES_8_port, MUL_RES_7_port, MUL_RES_6_port, MUL_RES_5_port, 
      MUL_RES_4_port, MUL_RES_3_port, MUL_RES_2_port, MUL_RES_1_port, 
      MUL_RES_0_port, sig_intraMux_31_port, sig_intraMux_30_port, 
      sig_intraMux_29_port, sig_intraMux_28_port, sig_intraMux_27_port, 
      sig_intraMux_26_port, sig_intraMux_25_port, sig_intraMux_24_port, 
      sig_intraMux_23_port, sig_intraMux_22_port, sig_intraMux_21_port, 
      sig_intraMux_20_port, sig_intraMux_19_port, sig_intraMux_18_port, 
      sig_intraMux_17_port, sig_intraMux_16_port, sig_intraMux_15_port, 
      sig_intraMux_14_port, sig_intraMux_13_port, sig_intraMux_12_port, 
      sig_intraMux_11_port, sig_intraMux_10_port, sig_intraMux_9_port, 
      sig_intraMux_8_port, sig_intraMux_7_port, sig_intraMux_6_port, 
      sig_intraMux_5_port, sig_intraMux_4_port, sig_intraMux_3_port, 
      sig_intraMux_2_port, sig_intraMux_1_port, sig_intraMux_0_port, 
      sig_ALU_RES_31_port, sig_ALU_RES_30_port, sig_ALU_RES_29_port, 
      sig_ALU_RES_28_port, sig_ALU_RES_27_port, sig_ALU_RES_26_port, 
      sig_ALU_RES_25_port, sig_ALU_RES_24_port, sig_ALU_RES_23_port, 
      sig_ALU_RES_22_port, sig_ALU_RES_21_port, sig_ALU_RES_20_port, 
      sig_ALU_RES_19_port, sig_ALU_RES_18_port, sig_ALU_RES_17_port, 
      sig_ALU_RES_16_port, sig_ALU_RES_15_port, sig_ALU_RES_14_port, 
      sig_ALU_RES_13_port, sig_ALU_RES_12_port, sig_ALU_RES_11_port, 
      sig_ALU_RES_10_port, sig_ALU_RES_9_port, sig_ALU_RES_8_port, 
      sig_ALU_RES_7_port, sig_ALU_RES_6_port, sig_ALU_RES_5_port, 
      sig_ALU_RES_4_port, sig_ALU_RES_3_port, sig_ALU_RES_2_port, 
      sig_ALU_RES_1_port, sig_ALU_RES_0_port, n78, n79, n80, n81, n82, n83, n84
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n85, n86, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n_1166, n_1167, n_1168, n_1169, n_1170, 
      n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, 
      n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, 
      n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   U227 : OAI22_X2 port map( A1 => n191, A2 => n35, B1 => n41, B2 => n68, ZN =>
                           A_SHF_31_port);
   U257 : NOR2_X2 port map( A1 => n75, A2 => n26, ZN => A_MUL_9_port);
   U258 : NOR2_X2 port map( A1 => n74, A2 => n26, ZN => A_MUL_8_port);
   U259 : NOR2_X2 port map( A1 => n73, A2 => n26, ZN => A_MUL_7_port);
   U260 : NOR2_X2 port map( A1 => n72, A2 => n26, ZN => A_MUL_6_port);
   U261 : NOR2_X2 port map( A1 => n71, A2 => n25, ZN => A_MUL_5_port);
   U262 : NOR2_X2 port map( A1 => n70, A2 => n25, ZN => A_MUL_4_port);
   U263 : NOR2_X2 port map( A1 => n69, A2 => n25, ZN => A_MUL_3_port);
   U264 : NOR2_X2 port map( A1 => n66, A2 => n25, ZN => A_MUL_2_port);
   U265 : NOR2_X2 port map( A1 => n55, A2 => n25, ZN => A_MUL_1_port);
   U267 : NOR2_X2 port map( A1 => n49, A2 => n25, ZN => A_MUL_14_port);
   U268 : NOR2_X2 port map( A1 => n48, A2 => n25, ZN => A_MUL_13_port);
   U269 : NOR2_X2 port map( A1 => n47, A2 => n25, ZN => A_MUL_12_port);
   U270 : NOR2_X2 port map( A1 => n46, A2 => n25, ZN => A_MUL_11_port);
   U271 : NOR2_X2 port map( A1 => n45, A2 => n25, ZN => A_MUL_10_port);
   U272 : NOR2_X2 port map( A1 => n44, A2 => n25, ZN => A_MUL_0_port);
   U427 : NAND3_X1 port map( A1 => n209, A2 => n208, A3 => n80, ZN => n79);
   U428 : NAND3_X1 port map( A1 => n43, A2 => n37, A3 => n34, ZN => 
                           select_type_sig_1_port);
   U429 : NAND3_X1 port map( A1 => n84, A2 => n3, A3 => n34, ZN => 
                           select_type_sig_0_port);
   U430 : NAND3_X1 port map( A1 => ALU_OPC(1), A2 => n209, A3 => n156, ZN => 
                           n84);
   U431 : NAND3_X1 port map( A1 => ALU_OPC(4), A2 => ALU_OPC(1), A3 => n156, ZN
                           => n158);
   U432 : NAND3_X1 port map( A1 => ALU_OPC(0), A2 => ALU_OPC(3), A3 => n162, ZN
                           => n82);
   U434 : NAND3_X1 port map( A1 => n208, A2 => n206, A3 => ALU_OPC(0), ZN => 
                           n164);
   U435 : OAI33_X1 port map( A1 => n208, A2 => n202, A3 => n209, B1 => n170, B2
                           => ALU_OPC(4), B3 => n207, ZN => ADD_SUB);
   U436 : NAND3_X1 port map( A1 => n206, A2 => n201, A3 => n208, ZN => n170);
   Comp : comparator_NBIT32 port map( A(31) => A_CMP_31_port, A(30) => 
                           A_CMP_30_port, A(29) => A_CMP_29_port, A(28) => 
                           A_CMP_28_port, A(27) => A_CMP_27_port, A(26) => 
                           A_CMP_26_port, A(25) => A_CMP_25_port, A(24) => 
                           A_CMP_24_port, A(23) => A_CMP_23_port, A(22) => 
                           A_CMP_22_port, A(21) => A_CMP_21_port, A(20) => 
                           A_CMP_20_port, A(19) => A_CMP_19_port, A(18) => 
                           A_CMP_18_port, A(17) => A_CMP_17_port, A(16) => 
                           A_CMP_16_port, A(15) => A_CMP_15_port, A(14) => 
                           A_CMP_14_port, A(13) => A_CMP_13_port, A(12) => 
                           A_CMP_12_port, A(11) => A_CMP_11_port, A(10) => 
                           A_CMP_10_port, A(9) => A_CMP_9_port, A(8) => 
                           A_CMP_8_port, A(7) => A_CMP_7_port, A(6) => 
                           A_CMP_6_port, A(5) => A_CMP_5_port, A(4) => 
                           A_CMP_4_port, A(3) => A_CMP_3_port, A(2) => 
                           A_CMP_2_port, A(1) => A_CMP_1_port, A(0) => 
                           A_CMP_0_port, B(31) => B_CMP_31_port, B(30) => 
                           B_CMP_30_port, B(29) => B_CMP_29_port, B(28) => 
                           B_CMP_28_port, B(27) => B_CMP_27_port, B(26) => 
                           B_CMP_26_port, B(25) => B_CMP_25_port, B(24) => 
                           B_CMP_24_port, B(23) => B_CMP_23_port, B(22) => 
                           B_CMP_22_port, B(21) => B_CMP_21_port, B(20) => 
                           B_CMP_20_port, B(19) => B_CMP_19_port, B(18) => 
                           B_CMP_18_port, B(17) => B_CMP_17_port, B(16) => 
                           B_CMP_16_port, B(15) => B_CMP_15_port, B(14) => 
                           B_CMP_14_port, B(13) => B_CMP_13_port, B(12) => 
                           B_CMP_12_port, B(11) => B_CMP_11_port, B(10) => 
                           B_CMP_10_port, B(9) => B_CMP_9_port, B(8) => 
                           B_CMP_8_port, B(7) => B_CMP_7_port, B(6) => 
                           B_CMP_6_port, B(5) => B_CMP_5_port, B(4) => 
                           B_CMP_4_port, B(3) => B_CMP_3_port, B(2) => 
                           B_CMP_2_port, B(1) => B_CMP_1_port, B(0) => 
                           B_CMP_0_port, OPSel(0) => n203, OPSel(1) => 
                           OPSel_1_port, OPSel(2) => OPSel_0_port, RES(31) => 
                           n_1166, RES(30) => n_1167, RES(29) => n_1168, 
                           RES(28) => n_1169, RES(27) => n_1170, RES(26) => 
                           n_1171, RES(25) => n_1172, RES(24) => n_1173, 
                           RES(23) => n_1174, RES(22) => n_1175, RES(21) => 
                           n_1176, RES(20) => n_1177, RES(19) => n_1178, 
                           RES(18) => n_1179, RES(17) => n_1180, RES(16) => 
                           n_1181, RES(15) => n_1182, RES(14) => n_1183, 
                           RES(13) => n_1184, RES(12) => n_1185, RES(11) => 
                           n_1186, RES(10) => n_1187, RES(9) => n_1188, RES(8) 
                           => n_1189, RES(7) => n_1190, RES(6) => n_1191, 
                           RES(5) => n_1192, RES(4) => n_1193, RES(3) => n_1194
                           , RES(2) => n_1195, RES(1) => n_1196, RES(0) => 
                           COMP_RES_0_port);
   Shift : shifter_NBIT32 port map( A(31) => A_SHF_31_port, A(30) => 
                           A_SHF_30_port, A(29) => A_SHF_29_port, A(28) => 
                           A_SHF_28_port, A(27) => A_SHF_27_port, A(26) => 
                           A_SHF_26_port, A(25) => A_SHF_25_port, A(24) => 
                           A_SHF_24_port, A(23) => A_SHF_23_port, A(22) => 
                           A_SHF_22_port, A(21) => A_SHF_21_port, A(20) => 
                           A_SHF_20_port, A(19) => A_SHF_19_port, A(18) => 
                           A_SHF_18_port, A(17) => A_SHF_17_port, A(16) => 
                           A_SHF_16_port, A(15) => A_SHF_15_port, A(14) => 
                           A_SHF_14_port, A(13) => A_SHF_13_port, A(12) => 
                           A_SHF_12_port, A(11) => A_SHF_11_port, A(10) => 
                           A_SHF_10_port, A(9) => A_SHF_9_port, A(8) => 
                           A_SHF_8_port, A(7) => A_SHF_7_port, A(6) => 
                           A_SHF_6_port, A(5) => A_SHF_5_port, A(4) => 
                           A_SHF_4_port, A(3) => A_SHF_3_port, A(2) => 
                           A_SHF_2_port, A(1) => A_SHF_1_port, A(0) => 
                           A_SHF_0_port, B(31) => B_SHF_31_port, B(30) => 
                           B_SHF_30_port, B(29) => B_SHF_29_port, B(28) => 
                           B_SHF_28_port, B(27) => B_SHF_27_port, B(26) => 
                           B_SHF_26_port, B(25) => B_SHF_25_port, B(24) => 
                           B_SHF_24_port, B(23) => B_SHF_23_port, B(22) => 
                           B_SHF_22_port, B(21) => B_SHF_21_port, B(20) => 
                           B_SHF_20_port, B(19) => B_SHF_19_port, B(18) => 
                           B_SHF_18_port, B(17) => B_SHF_17_port, B(16) => 
                           B_SHF_16_port, B(15) => B_SHF_15_port, B(14) => 
                           B_SHF_14_port, B(13) => B_SHF_13_port, B(12) => 
                           B_SHF_12_port, B(11) => B_SHF_11_port, B(10) => 
                           B_SHF_10_port, B(9) => B_SHF_9_port, B(8) => 
                           B_SHF_8_port, B(7) => B_SHF_7_port, B(6) => 
                           B_SHF_6_port, B(5) => B_SHF_5_port, B(4) => 
                           B_SHF_4_port, B(3) => B_SHF_3_port, B(2) => 
                           B_SHF_2_port, B(1) => B_SHF_1_port, B(0) => 
                           B_SHF_0_port, LOGIC_ARITH => LOGIC_ARITH, LEFT_RIGHT
                           => LEFT_RIGHT, RES(31) => SHIFT_RES_31_port, RES(30)
                           => SHIFT_RES_30_port, RES(29) => SHIFT_RES_29_port, 
                           RES(28) => SHIFT_RES_28_port, RES(27) => 
                           SHIFT_RES_27_port, RES(26) => SHIFT_RES_26_port, 
                           RES(25) => SHIFT_RES_25_port, RES(24) => 
                           SHIFT_RES_24_port, RES(23) => SHIFT_RES_23_port, 
                           RES(22) => SHIFT_RES_22_port, RES(21) => 
                           SHIFT_RES_21_port, RES(20) => SHIFT_RES_20_port, 
                           RES(19) => SHIFT_RES_19_port, RES(18) => 
                           SHIFT_RES_18_port, RES(17) => SHIFT_RES_17_port, 
                           RES(16) => SHIFT_RES_16_port, RES(15) => 
                           SHIFT_RES_15_port, RES(14) => SHIFT_RES_14_port, 
                           RES(13) => SHIFT_RES_13_port, RES(12) => 
                           SHIFT_RES_12_port, RES(11) => SHIFT_RES_11_port, 
                           RES(10) => SHIFT_RES_10_port, RES(9) => 
                           SHIFT_RES_9_port, RES(8) => SHIFT_RES_8_port, RES(7)
                           => SHIFT_RES_7_port, RES(6) => SHIFT_RES_6_port, 
                           RES(5) => SHIFT_RES_5_port, RES(4) => 
                           SHIFT_RES_4_port, RES(3) => SHIFT_RES_3_port, RES(2)
                           => SHIFT_RES_2_port, RES(1) => SHIFT_RES_1_port, 
                           RES(0) => SHIFT_RES_0_port);
   Add_Sub_unit : P4Adder_NBIT32 port map( A(31) => A_ADD_31_port, A(30) => 
                           A_ADD_30_port, A(29) => A_ADD_29_port, A(28) => 
                           A_ADD_28_port, A(27) => A_ADD_27_port, A(26) => 
                           A_ADD_26_port, A(25) => A_ADD_25_port, A(24) => 
                           A_ADD_24_port, A(23) => A_ADD_23_port, A(22) => 
                           A_ADD_22_port, A(21) => A_ADD_21_port, A(20) => 
                           A_ADD_20_port, A(19) => A_ADD_19_port, A(18) => 
                           A_ADD_18_port, A(17) => A_ADD_17_port, A(16) => 
                           A_ADD_16_port, A(15) => A_ADD_15_port, A(14) => 
                           A_ADD_14_port, A(13) => A_ADD_13_port, A(12) => 
                           A_ADD_12_port, A(11) => A_ADD_11_port, A(10) => 
                           A_ADD_10_port, A(9) => A_ADD_9_port, A(8) => 
                           A_ADD_8_port, A(7) => A_ADD_7_port, A(6) => 
                           A_ADD_6_port, A(5) => A_ADD_5_port, A(4) => 
                           A_ADD_4_port, A(3) => A_ADD_3_port, A(2) => 
                           A_ADD_2_port, A(1) => A_ADD_1_port, A(0) => 
                           A_ADD_0_port, B(31) => B_ADD_31_port, B(30) => 
                           B_ADD_30_port, B(29) => B_ADD_29_port, B(28) => 
                           B_ADD_28_port, B(27) => B_ADD_27_port, B(26) => 
                           B_ADD_26_port, B(25) => B_ADD_25_port, B(24) => 
                           B_ADD_24_port, B(23) => B_ADD_23_port, B(22) => 
                           B_ADD_22_port, B(21) => B_ADD_21_port, B(20) => 
                           B_ADD_20_port, B(19) => B_ADD_19_port, B(18) => 
                           B_ADD_18_port, B(17) => B_ADD_17_port, B(16) => 
                           B_ADD_16_port, B(15) => B_ADD_15_port, B(14) => 
                           B_ADD_14_port, B(13) => B_ADD_13_port, B(12) => 
                           B_ADD_12_port, B(11) => B_ADD_11_port, B(10) => 
                           B_ADD_10_port, B(9) => B_ADD_9_port, B(8) => 
                           B_ADD_8_port, B(7) => B_ADD_7_port, B(6) => 
                           B_ADD_6_port, B(5) => B_ADD_5_port, B(4) => 
                           B_ADD_4_port, B(3) => B_ADD_3_port, B(2) => 
                           B_ADD_2_port, B(1) => B_ADD_1_port, B(0) => 
                           B_ADD_0_port, Cin => n2, S(31) => 
                           ADD_SUB_RES_31_port, S(30) => ADD_SUB_RES_30_port, 
                           S(29) => ADD_SUB_RES_29_port, S(28) => 
                           ADD_SUB_RES_28_port, S(27) => ADD_SUB_RES_27_port, 
                           S(26) => ADD_SUB_RES_26_port, S(25) => 
                           ADD_SUB_RES_25_port, S(24) => ADD_SUB_RES_24_port, 
                           S(23) => ADD_SUB_RES_23_port, S(22) => 
                           ADD_SUB_RES_22_port, S(21) => ADD_SUB_RES_21_port, 
                           S(20) => ADD_SUB_RES_20_port, S(19) => 
                           ADD_SUB_RES_19_port, S(18) => ADD_SUB_RES_18_port, 
                           S(17) => ADD_SUB_RES_17_port, S(16) => 
                           ADD_SUB_RES_16_port, S(15) => ADD_SUB_RES_15_port, 
                           S(14) => ADD_SUB_RES_14_port, S(13) => 
                           ADD_SUB_RES_13_port, S(12) => ADD_SUB_RES_12_port, 
                           S(11) => ADD_SUB_RES_11_port, S(10) => 
                           ADD_SUB_RES_10_port, S(9) => ADD_SUB_RES_9_port, 
                           S(8) => ADD_SUB_RES_8_port, S(7) => 
                           ADD_SUB_RES_7_port, S(6) => ADD_SUB_RES_6_port, S(5)
                           => ADD_SUB_RES_5_port, S(4) => ADD_SUB_RES_4_port, 
                           S(3) => ADD_SUB_RES_3_port, S(2) => 
                           ADD_SUB_RES_2_port, S(1) => ADD_SUB_RES_1_port, S(0)
                           => ADD_SUB_RES_0_port, Cout => n_1197);
   Booth_mul : BOOTHMUL_numBit16 port map( A(15) => A_MUL_15_port, A(14) => 
                           A_MUL_14_port, A(13) => A_MUL_13_port, A(12) => 
                           A_MUL_12_port, A(11) => A_MUL_11_port, A(10) => 
                           A_MUL_10_port, A(9) => A_MUL_9_port, A(8) => 
                           A_MUL_8_port, A(7) => A_MUL_7_port, A(6) => 
                           A_MUL_6_port, A(5) => A_MUL_5_port, A(4) => 
                           A_MUL_4_port, A(3) => A_MUL_3_port, A(2) => 
                           A_MUL_2_port, A(1) => A_MUL_1_port, A(0) => 
                           A_MUL_0_port, B(15) => B_MUL_15_port, B(14) => 
                           B_MUL_14_port, B(13) => B_MUL_13_port, B(12) => 
                           B_MUL_12_port, B(11) => B_MUL_11_port, B(10) => 
                           B_MUL_10_port, B(9) => B_MUL_9_port, B(8) => 
                           B_MUL_8_port, B(7) => B_MUL_7_port, B(6) => 
                           B_MUL_6_port, B(5) => B_MUL_5_port, B(4) => 
                           B_MUL_4_port, B(3) => B_MUL_3_port, B(2) => 
                           B_MUL_2_port, B(1) => B_MUL_1_port, B(0) => 
                           B_MUL_0_port, P(31) => MUL_RES_31_port, P(30) => 
                           MUL_RES_30_port, P(29) => MUL_RES_29_port, P(28) => 
                           MUL_RES_28_port, P(27) => MUL_RES_27_port, P(26) => 
                           MUL_RES_26_port, P(25) => MUL_RES_25_port, P(24) => 
                           MUL_RES_24_port, P(23) => MUL_RES_23_port, P(22) => 
                           MUL_RES_22_port, P(21) => MUL_RES_21_port, P(20) => 
                           MUL_RES_20_port, P(19) => MUL_RES_19_port, P(18) => 
                           MUL_RES_18_port, P(17) => MUL_RES_17_port, P(16) => 
                           MUL_RES_16_port, P(15) => MUL_RES_15_port, P(14) => 
                           MUL_RES_14_port, P(13) => MUL_RES_13_port, P(12) => 
                           MUL_RES_12_port, P(11) => MUL_RES_11_port, P(10) => 
                           MUL_RES_10_port, P(9) => MUL_RES_9_port, P(8) => 
                           MUL_RES_8_port, P(7) => MUL_RES_7_port, P(6) => 
                           MUL_RES_6_port, P(5) => MUL_RES_5_port, P(4) => 
                           MUL_RES_4_port, P(3) => MUL_RES_3_port, P(2) => 
                           MUL_RES_2_port, P(1) => MUL_RES_1_port, P(0) => 
                           MUL_RES_0_port);
   Res_mux : mux41_NBIT32_1 port map( A(31) => ADD_SUB_RES_31_port, A(30) => 
                           ADD_SUB_RES_30_port, A(29) => ADD_SUB_RES_29_port, 
                           A(28) => ADD_SUB_RES_28_port, A(27) => 
                           ADD_SUB_RES_27_port, A(26) => ADD_SUB_RES_26_port, 
                           A(25) => ADD_SUB_RES_25_port, A(24) => 
                           ADD_SUB_RES_24_port, A(23) => ADD_SUB_RES_23_port, 
                           A(22) => ADD_SUB_RES_22_port, A(21) => 
                           ADD_SUB_RES_21_port, A(20) => ADD_SUB_RES_20_port, 
                           A(19) => ADD_SUB_RES_19_port, A(18) => 
                           ADD_SUB_RES_18_port, A(17) => ADD_SUB_RES_17_port, 
                           A(16) => ADD_SUB_RES_16_port, A(15) => 
                           ADD_SUB_RES_15_port, A(14) => ADD_SUB_RES_14_port, 
                           A(13) => ADD_SUB_RES_13_port, A(12) => 
                           ADD_SUB_RES_12_port, A(11) => ADD_SUB_RES_11_port, 
                           A(10) => ADD_SUB_RES_10_port, A(9) => 
                           ADD_SUB_RES_9_port, A(8) => ADD_SUB_RES_8_port, A(7)
                           => ADD_SUB_RES_7_port, A(6) => ADD_SUB_RES_6_port, 
                           A(5) => ADD_SUB_RES_5_port, A(4) => 
                           ADD_SUB_RES_4_port, A(3) => ADD_SUB_RES_3_port, A(2)
                           => ADD_SUB_RES_2_port, A(1) => ADD_SUB_RES_1_port, 
                           A(0) => ADD_SUB_RES_0_port, B(31) => 
                           LOGIC_RES_31_port, B(30) => LOGIC_RES_30_port, B(29)
                           => LOGIC_RES_29_port, B(28) => LOGIC_RES_28_port, 
                           B(27) => LOGIC_RES_27_port, B(26) => 
                           LOGIC_RES_26_port, B(25) => LOGIC_RES_25_port, B(24)
                           => LOGIC_RES_24_port, B(23) => LOGIC_RES_23_port, 
                           B(22) => LOGIC_RES_22_port, B(21) => 
                           LOGIC_RES_21_port, B(20) => LOGIC_RES_20_port, B(19)
                           => LOGIC_RES_19_port, B(18) => LOGIC_RES_18_port, 
                           B(17) => LOGIC_RES_17_port, B(16) => 
                           LOGIC_RES_16_port, B(15) => LOGIC_RES_15_port, B(14)
                           => LOGIC_RES_14_port, B(13) => LOGIC_RES_13_port, 
                           B(12) => LOGIC_RES_12_port, B(11) => 
                           LOGIC_RES_11_port, B(10) => LOGIC_RES_10_port, B(9) 
                           => LOGIC_RES_9_port, B(8) => LOGIC_RES_8_port, B(7) 
                           => LOGIC_RES_7_port, B(6) => LOGIC_RES_6_port, B(5) 
                           => LOGIC_RES_5_port, B(4) => LOGIC_RES_4_port, B(3) 
                           => LOGIC_RES_3_port, B(2) => LOGIC_RES_2_port, B(1) 
                           => LOGIC_RES_1_port, B(0) => LOGIC_RES_0_port, C(31)
                           => SHIFT_RES_31_port, C(30) => SHIFT_RES_30_port, 
                           C(29) => SHIFT_RES_29_port, C(28) => 
                           SHIFT_RES_28_port, C(27) => SHIFT_RES_27_port, C(26)
                           => SHIFT_RES_26_port, C(25) => SHIFT_RES_25_port, 
                           C(24) => SHIFT_RES_24_port, C(23) => 
                           SHIFT_RES_23_port, C(22) => SHIFT_RES_22_port, C(21)
                           => SHIFT_RES_21_port, C(20) => SHIFT_RES_20_port, 
                           C(19) => SHIFT_RES_19_port, C(18) => 
                           SHIFT_RES_18_port, C(17) => SHIFT_RES_17_port, C(16)
                           => SHIFT_RES_16_port, C(15) => SHIFT_RES_15_port, 
                           C(14) => SHIFT_RES_14_port, C(13) => 
                           SHIFT_RES_13_port, C(12) => SHIFT_RES_12_port, C(11)
                           => SHIFT_RES_11_port, C(10) => SHIFT_RES_10_port, 
                           C(9) => SHIFT_RES_9_port, C(8) => SHIFT_RES_8_port, 
                           C(7) => SHIFT_RES_7_port, C(6) => SHIFT_RES_6_port, 
                           C(5) => SHIFT_RES_5_port, C(4) => SHIFT_RES_4_port, 
                           C(3) => SHIFT_RES_3_port, C(2) => SHIFT_RES_2_port, 
                           C(1) => SHIFT_RES_1_port, C(0) => SHIFT_RES_0_port, 
                           D(31) => COMP_RES_31_port, D(30) => COMP_RES_30_port
                           , D(29) => COMP_RES_29_port, D(28) => 
                           COMP_RES_28_port, D(27) => COMP_RES_27_port, D(26) 
                           => COMP_RES_26_port, D(25) => COMP_RES_25_port, 
                           D(24) => COMP_RES_24_port, D(23) => COMP_RES_23_port
                           , D(22) => COMP_RES_22_port, D(21) => 
                           COMP_RES_21_port, D(20) => COMP_RES_20_port, D(19) 
                           => COMP_RES_19_port, D(18) => COMP_RES_18_port, 
                           D(17) => COMP_RES_17_port, D(16) => COMP_RES_16_port
                           , D(15) => COMP_RES_15_port, D(14) => 
                           COMP_RES_14_port, D(13) => COMP_RES_13_port, D(12) 
                           => COMP_RES_12_port, D(11) => COMP_RES_11_port, 
                           D(10) => COMP_RES_10_port, D(9) => COMP_RES_9_port, 
                           D(8) => COMP_RES_8_port, D(7) => COMP_RES_7_port, 
                           D(6) => COMP_RES_6_port, D(5) => COMP_RES_5_port, 
                           D(4) => COMP_RES_4_port, D(3) => COMP_RES_3_port, 
                           D(2) => COMP_RES_2_port, D(1) => COMP_RES_1_port, 
                           D(0) => COMP_RES_0_port, S(1) => 
                           select_type_sig_1_port, S(0) => 
                           select_type_sig_0_port, Z(31) => 
                           sig_intraMux_31_port, Z(30) => sig_intraMux_30_port,
                           Z(29) => sig_intraMux_29_port, Z(28) => 
                           sig_intraMux_28_port, Z(27) => sig_intraMux_27_port,
                           Z(26) => sig_intraMux_26_port, Z(25) => 
                           sig_intraMux_25_port, Z(24) => sig_intraMux_24_port,
                           Z(23) => sig_intraMux_23_port, Z(22) => 
                           sig_intraMux_22_port, Z(21) => sig_intraMux_21_port,
                           Z(20) => sig_intraMux_20_port, Z(19) => 
                           sig_intraMux_19_port, Z(18) => sig_intraMux_18_port,
                           Z(17) => sig_intraMux_17_port, Z(16) => 
                           sig_intraMux_16_port, Z(15) => sig_intraMux_15_port,
                           Z(14) => sig_intraMux_14_port, Z(13) => 
                           sig_intraMux_13_port, Z(12) => sig_intraMux_12_port,
                           Z(11) => sig_intraMux_11_port, Z(10) => 
                           sig_intraMux_10_port, Z(9) => sig_intraMux_9_port, 
                           Z(8) => sig_intraMux_8_port, Z(7) => 
                           sig_intraMux_7_port, Z(6) => sig_intraMux_6_port, 
                           Z(5) => sig_intraMux_5_port, Z(4) => 
                           sig_intraMux_4_port, Z(3) => sig_intraMux_3_port, 
                           Z(2) => sig_intraMux_2_port, Z(1) => 
                           sig_intraMux_1_port, Z(0) => sig_intraMux_0_port);
   Mul_mux : mux21_NBIT32_2 port map( A(31) => sig_intraMux_31_port, A(30) => 
                           sig_intraMux_30_port, A(29) => sig_intraMux_29_port,
                           A(28) => sig_intraMux_28_port, A(27) => 
                           sig_intraMux_27_port, A(26) => sig_intraMux_26_port,
                           A(25) => sig_intraMux_25_port, A(24) => 
                           sig_intraMux_24_port, A(23) => sig_intraMux_23_port,
                           A(22) => sig_intraMux_22_port, A(21) => 
                           sig_intraMux_21_port, A(20) => sig_intraMux_20_port,
                           A(19) => sig_intraMux_19_port, A(18) => 
                           sig_intraMux_18_port, A(17) => sig_intraMux_17_port,
                           A(16) => sig_intraMux_16_port, A(15) => 
                           sig_intraMux_15_port, A(14) => sig_intraMux_14_port,
                           A(13) => sig_intraMux_13_port, A(12) => 
                           sig_intraMux_12_port, A(11) => sig_intraMux_11_port,
                           A(10) => sig_intraMux_10_port, A(9) => 
                           sig_intraMux_9_port, A(8) => sig_intraMux_8_port, 
                           A(7) => sig_intraMux_7_port, A(6) => 
                           sig_intraMux_6_port, A(5) => sig_intraMux_5_port, 
                           A(4) => sig_intraMux_4_port, A(3) => 
                           sig_intraMux_3_port, A(2) => sig_intraMux_2_port, 
                           A(1) => sig_intraMux_1_port, A(0) => 
                           sig_intraMux_0_port, B(31) => MUL_RES_31_port, B(30)
                           => MUL_RES_30_port, B(29) => MUL_RES_29_port, B(28) 
                           => MUL_RES_28_port, B(27) => MUL_RES_27_port, B(26) 
                           => MUL_RES_26_port, B(25) => MUL_RES_25_port, B(24) 
                           => MUL_RES_24_port, B(23) => MUL_RES_23_port, B(22) 
                           => MUL_RES_22_port, B(21) => MUL_RES_21_port, B(20) 
                           => MUL_RES_20_port, B(19) => MUL_RES_19_port, B(18) 
                           => MUL_RES_18_port, B(17) => MUL_RES_17_port, B(16) 
                           => MUL_RES_16_port, B(15) => MUL_RES_15_port, B(14) 
                           => MUL_RES_14_port, B(13) => MUL_RES_13_port, B(12) 
                           => MUL_RES_12_port, B(11) => MUL_RES_11_port, B(10) 
                           => MUL_RES_10_port, B(9) => MUL_RES_9_port, B(8) => 
                           MUL_RES_8_port, B(7) => MUL_RES_7_port, B(6) => 
                           MUL_RES_6_port, B(5) => MUL_RES_5_port, B(4) => 
                           MUL_RES_4_port, B(3) => MUL_RES_3_port, B(2) => 
                           MUL_RES_2_port, B(1) => MUL_RES_1_port, B(0) => 
                           MUL_RES_0_port, S => n1, Z(31) => 
                           sig_ALU_RES_31_port, Z(30) => sig_ALU_RES_30_port, 
                           Z(29) => sig_ALU_RES_29_port, Z(28) => 
                           sig_ALU_RES_28_port, Z(27) => sig_ALU_RES_27_port, 
                           Z(26) => sig_ALU_RES_26_port, Z(25) => 
                           sig_ALU_RES_25_port, Z(24) => sig_ALU_RES_24_port, 
                           Z(23) => sig_ALU_RES_23_port, Z(22) => 
                           sig_ALU_RES_22_port, Z(21) => sig_ALU_RES_21_port, 
                           Z(20) => sig_ALU_RES_20_port, Z(19) => 
                           sig_ALU_RES_19_port, Z(18) => sig_ALU_RES_18_port, 
                           Z(17) => sig_ALU_RES_17_port, Z(16) => 
                           sig_ALU_RES_16_port, Z(15) => sig_ALU_RES_15_port, 
                           Z(14) => sig_ALU_RES_14_port, Z(13) => 
                           sig_ALU_RES_13_port, Z(12) => sig_ALU_RES_12_port, 
                           Z(11) => sig_ALU_RES_11_port, Z(10) => 
                           sig_ALU_RES_10_port, Z(9) => sig_ALU_RES_9_port, 
                           Z(8) => sig_ALU_RES_8_port, Z(7) => 
                           sig_ALU_RES_7_port, Z(6) => sig_ALU_RES_6_port, Z(5)
                           => sig_ALU_RES_5_port, Z(4) => sig_ALU_RES_4_port, 
                           Z(3) => sig_ALU_RES_3_port, Z(2) => 
                           sig_ALU_RES_2_port, Z(1) => sig_ALU_RES_1_port, Z(0)
                           => sig_ALU_RES_0_port);
   Zeros_mux : mux21_NBIT32_1 port map( A(31) => sig_ALU_RES_31_port, A(30) => 
                           sig_ALU_RES_30_port, A(29) => sig_ALU_RES_29_port, 
                           A(28) => sig_ALU_RES_28_port, A(27) => 
                           sig_ALU_RES_27_port, A(26) => sig_ALU_RES_26_port, 
                           A(25) => sig_ALU_RES_25_port, A(24) => 
                           sig_ALU_RES_24_port, A(23) => sig_ALU_RES_23_port, 
                           A(22) => sig_ALU_RES_22_port, A(21) => 
                           sig_ALU_RES_21_port, A(20) => sig_ALU_RES_20_port, 
                           A(19) => sig_ALU_RES_19_port, A(18) => 
                           sig_ALU_RES_18_port, A(17) => sig_ALU_RES_17_port, 
                           A(16) => sig_ALU_RES_16_port, A(15) => 
                           sig_ALU_RES_15_port, A(14) => sig_ALU_RES_14_port, 
                           A(13) => sig_ALU_RES_13_port, A(12) => 
                           sig_ALU_RES_12_port, A(11) => sig_ALU_RES_11_port, 
                           A(10) => sig_ALU_RES_10_port, A(9) => 
                           sig_ALU_RES_9_port, A(8) => sig_ALU_RES_8_port, A(7)
                           => sig_ALU_RES_7_port, A(6) => sig_ALU_RES_6_port, 
                           A(5) => sig_ALU_RES_5_port, A(4) => 
                           sig_ALU_RES_4_port, A(3) => sig_ALU_RES_3_port, A(2)
                           => sig_ALU_RES_2_port, A(1) => sig_ALU_RES_1_port, 
                           A(0) => sig_ALU_RES_0_port, B(31) => X_Logic0_port, 
                           B(30) => X_Logic0_port, B(29) => X_Logic0_port, 
                           B(28) => X_Logic0_port, B(27) => X_Logic0_port, 
                           B(26) => X_Logic0_port, B(25) => X_Logic0_port, 
                           B(24) => X_Logic0_port, B(23) => X_Logic0_port, 
                           B(22) => X_Logic0_port, B(21) => X_Logic0_port, 
                           B(20) => X_Logic0_port, B(19) => X_Logic0_port, 
                           B(18) => X_Logic0_port, B(17) => X_Logic0_port, 
                           B(16) => X_Logic0_port, B(15) => X_Logic0_port, 
                           B(14) => X_Logic0_port, B(13) => X_Logic0_port, 
                           B(12) => X_Logic0_port, B(11) => X_Logic0_port, 
                           B(10) => X_Logic0_port, B(9) => X_Logic0_port, B(8) 
                           => X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, S => select_zero_sig, Z(31) => 
                           ALU_RES(31), Z(30) => ALU_RES(30), Z(29) => 
                           ALU_RES(29), Z(28) => ALU_RES(28), Z(27) => 
                           ALU_RES(27), Z(26) => ALU_RES(26), Z(25) => 
                           ALU_RES(25), Z(24) => ALU_RES(24), Z(23) => 
                           ALU_RES(23), Z(22) => ALU_RES(22), Z(21) => 
                           ALU_RES(21), Z(20) => ALU_RES(20), Z(19) => 
                           ALU_RES(19), Z(18) => ALU_RES(18), Z(17) => 
                           ALU_RES(17), Z(16) => ALU_RES(16), Z(15) => 
                           ALU_RES(15), Z(14) => ALU_RES(14), Z(13) => 
                           ALU_RES(13), Z(12) => ALU_RES(12), Z(11) => 
                           ALU_RES(11), Z(10) => ALU_RES(10), Z(9) => 
                           ALU_RES(9), Z(8) => ALU_RES(8), Z(7) => ALU_RES(7), 
                           Z(6) => ALU_RES(6), Z(5) => ALU_RES(5), Z(4) => 
                           ALU_RES(4), Z(3) => ALU_RES(3), Z(2) => ALU_RES(2), 
                           Z(1) => ALU_RES(1), Z(0) => ALU_RES(0));
   U3 : OAI22_X1 port map( A1 => n194, A2 => n35, B1 => n40, B2 => n71, ZN => 
                           A_SHF_5_port);
   U4 : OAI22_X1 port map( A1 => n195, A2 => n35, B1 => n40, B2 => n72, ZN => 
                           A_SHF_6_port);
   U5 : OAI22_X1 port map( A1 => n185, A2 => n36, B1 => n41, B2 => n62, ZN => 
                           A_SHF_26_port);
   U6 : OAI22_X1 port map( A1 => n186, A2 => n36, B1 => n41, B2 => n63, ZN => 
                           A_SHF_27_port);
   U7 : AND3_X1 port map( A1 => ALU_OPC(4), A2 => ALU_OPC(2), A3 => n163, ZN =>
                           n1);
   U8 : INV_X1 port map( A => n199, ZN => n2);
   U9 : BUF_X1 port map( A => n168, Z => n13);
   U10 : BUF_X1 port map( A => n168, Z => n14);
   U11 : BUF_X1 port map( A => n168, Z => n15);
   U12 : OAI22_X1 port map( A1 => n175, A2 => n37, B1 => n42, B2 => n52, ZN => 
                           A_SHF_17_port);
   U13 : OAI22_X1 port map( A1 => n196, A2 => n35, B1 => n40, B2 => n73, ZN => 
                           A_SHF_7_port);
   U14 : OAI22_X1 port map( A1 => n176, A2 => n37, B1 => n42, B2 => n53, ZN => 
                           A_SHF_18_port);
   U15 : OAI22_X1 port map( A1 => n184, A2 => n36, B1 => n41, B2 => n61, ZN => 
                           A_SHF_25_port);
   U16 : OAI22_X1 port map( A1 => n187, A2 => n36, B1 => n41, B2 => n64, ZN => 
                           A_SHF_28_port);
   U17 : OAI22_X1 port map( A1 => n193, A2 => n36, B1 => n41, B2 => n70, ZN => 
                           A_SHF_4_port);
   U18 : NOR2_X1 port map( A1 => n38, A2 => n192, ZN => B_SHF_3_port);
   U19 : OAI22_X1 port map( A1 => n197, A2 => n35, B1 => n40, B2 => n74, ZN => 
                           A_SHF_8_port);
   U20 : OAI22_X1 port map( A1 => n189, A2 => n35, B1 => n41, B2 => n66, ZN => 
                           A_SHF_2_port);
   U21 : OAI22_X1 port map( A1 => n182, A2 => n36, B1 => n41, B2 => n59, ZN => 
                           A_SHF_23_port);
   U22 : OAI22_X1 port map( A1 => n183, A2 => n36, B1 => n41, B2 => n60, ZN => 
                           A_SHF_24_port);
   U23 : OAI22_X1 port map( A1 => n177, A2 => n36, B1 => n42, B2 => n54, ZN => 
                           A_SHF_19_port);
   U24 : OAI22_X1 port map( A1 => n179, A2 => n36, B1 => n42, B2 => n56, ZN => 
                           A_SHF_20_port);
   U25 : OAI22_X1 port map( A1 => n180, A2 => n36, B1 => n42, B2 => n57, ZN => 
                           A_SHF_21_port);
   U26 : OAI22_X1 port map( A1 => n181, A2 => n36, B1 => n42, B2 => n58, ZN => 
                           A_SHF_22_port);
   U27 : OAI22_X1 port map( A1 => n86, A2 => n37, B1 => n43, B2 => n47, ZN => 
                           A_SHF_12_port);
   U28 : OAI22_X1 port map( A1 => n171, A2 => n37, B1 => n42, B2 => n48, ZN => 
                           A_SHF_13_port);
   U29 : OAI22_X1 port map( A1 => n172, A2 => n37, B1 => n42, B2 => n49, ZN => 
                           A_SHF_14_port);
   U30 : NOR2_X1 port map( A1 => n192, A2 => n26, ZN => B_MUL_3_port);
   U31 : NOR2_X1 port map( A1 => n194, A2 => n26, ZN => B_MUL_5_port);
   U32 : NOR2_X1 port map( A1 => n196, A2 => n26, ZN => B_MUL_7_port);
   U33 : NOR2_X1 port map( A1 => n198, A2 => n26, ZN => B_MUL_9_port);
   U34 : NOR2_X1 port map( A1 => n178, A2 => n26, ZN => B_MUL_1_port);
   U35 : NOR2_X1 port map( A1 => n85, A2 => n26, ZN => B_MUL_11_port);
   U36 : NOR2_X1 port map( A1 => n171, A2 => n26, ZN => B_MUL_13_port);
   U37 : NOR2_X1 port map( A1 => n38, A2 => n198, ZN => B_SHF_9_port);
   U38 : NOR2_X1 port map( A1 => n38, A2 => n197, ZN => B_SHF_8_port);
   U39 : NOR2_X1 port map( A1 => n40, A2 => n77, ZN => B_SHF_10_port);
   U40 : OAI22_X1 port map( A1 => n178, A2 => n36, B1 => n42, B2 => n55, ZN => 
                           A_SHF_1_port);
   U41 : NOR2_X1 port map( A1 => n38, A2 => n189, ZN => B_SHF_2_port);
   U42 : OAI22_X1 port map( A1 => n198, A2 => n35, B1 => n40, B2 => n75, ZN => 
                           A_SHF_9_port);
   U43 : OAI22_X1 port map( A1 => n76, A2 => n35, B1 => n42, B2 => n44, ZN => 
                           A_SHF_0_port);
   U44 : NOR2_X1 port map( A1 => n38, A2 => n196, ZN => B_SHF_7_port);
   U45 : NOR2_X1 port map( A1 => n38, A2 => n195, ZN => B_SHF_6_port);
   U46 : NOR2_X1 port map( A1 => n38, A2 => n194, ZN => B_SHF_5_port);
   U47 : OAI22_X1 port map( A1 => n85, A2 => n37, B1 => n43, B2 => n46, ZN => 
                           A_SHF_11_port);
   U48 : OAI22_X1 port map( A1 => n173, A2 => n37, B1 => n42, B2 => n50, ZN => 
                           A_SHF_15_port);
   U49 : OAI22_X1 port map( A1 => n188, A2 => n35, B1 => n41, B2 => n65, ZN => 
                           A_SHF_29_port);
   U50 : OAI22_X1 port map( A1 => n174, A2 => n37, B1 => n42, B2 => n51, ZN => 
                           A_SHF_16_port);
   U51 : OAI22_X1 port map( A1 => n192, A2 => n35, B1 => n41, B2 => n69, ZN => 
                           A_SHF_3_port);
   U52 : NOR2_X1 port map( A1 => n13, A2 => n44, ZN => A_ADD_0_port);
   U53 : NOR2_X1 port map( A1 => n15, A2 => n70, ZN => A_ADD_4_port);
   U54 : NOR2_X1 port map( A1 => n15, A2 => n74, ZN => A_ADD_8_port);
   U55 : NOR2_X1 port map( A1 => n15, A2 => n71, ZN => A_ADD_5_port);
   U56 : NOR2_X1 port map( A1 => n15, A2 => n75, ZN => A_ADD_9_port);
   U57 : NOR2_X1 port map( A1 => n15, A2 => n72, ZN => A_ADD_6_port);
   U58 : NOR2_X1 port map( A1 => n15, A2 => n69, ZN => A_ADD_3_port);
   U59 : NOR2_X1 port map( A1 => n15, A2 => n73, ZN => A_ADD_7_port);
   U60 : NOR2_X1 port map( A1 => n15, A2 => n68, ZN => A_ADD_31_port);
   U61 : NOR2_X1 port map( A1 => n13, A2 => n47, ZN => A_ADD_12_port);
   U62 : NOR2_X1 port map( A1 => n13, A2 => n51, ZN => A_ADD_16_port);
   U63 : NOR2_X1 port map( A1 => n14, A2 => n60, ZN => A_ADD_24_port);
   U64 : NOR2_X1 port map( A1 => n13, A2 => n55, ZN => A_ADD_1_port);
   U65 : NOR2_X1 port map( A1 => n13, A2 => n48, ZN => A_ADD_13_port);
   U66 : NOR2_X1 port map( A1 => n13, A2 => n52, ZN => A_ADD_17_port);
   U67 : NOR2_X1 port map( A1 => n14, A2 => n61, ZN => A_ADD_25_port);
   U68 : NOR2_X1 port map( A1 => n14, A2 => n66, ZN => A_ADD_2_port);
   U69 : NOR2_X1 port map( A1 => n13, A2 => n45, ZN => A_ADD_10_port);
   U70 : NOR2_X1 port map( A1 => n13, A2 => n49, ZN => A_ADD_14_port);
   U71 : NOR2_X1 port map( A1 => n13, A2 => n53, ZN => A_ADD_18_port);
   U72 : NOR2_X1 port map( A1 => n14, A2 => n62, ZN => A_ADD_26_port);
   U73 : NOR2_X1 port map( A1 => n14, A2 => n58, ZN => A_ADD_22_port);
   U74 : NOR2_X1 port map( A1 => n14, A2 => n57, ZN => A_ADD_21_port);
   U75 : NOR2_X1 port map( A1 => n14, A2 => n56, ZN => A_ADD_20_port);
   U76 : NOR2_X1 port map( A1 => n14, A2 => n67, ZN => A_ADD_30_port);
   U77 : NOR2_X1 port map( A1 => n14, A2 => n65, ZN => A_ADD_29_port);
   U78 : NOR2_X1 port map( A1 => n14, A2 => n64, ZN => A_ADD_28_port);
   U79 : NOR2_X1 port map( A1 => n13, A2 => n46, ZN => A_ADD_11_port);
   U80 : NOR2_X1 port map( A1 => n13, A2 => n50, ZN => A_ADD_15_port);
   U81 : NOR2_X1 port map( A1 => n13, A2 => n54, ZN => A_ADD_19_port);
   U82 : NOR2_X1 port map( A1 => n14, A2 => n59, ZN => A_ADD_23_port);
   U83 : NOR2_X1 port map( A1 => n14, A2 => n63, ZN => A_ADD_27_port);
   U84 : NOR2_X1 port map( A1 => n39, A2 => n178, ZN => B_SHF_1_port);
   U85 : NOR2_X1 port map( A1 => n38, A2 => n187, ZN => B_SHF_28_port);
   U86 : NOR2_X1 port map( A1 => n38, A2 => n186, ZN => B_SHF_27_port);
   U87 : NOR2_X1 port map( A1 => n39, A2 => n185, ZN => B_SHF_26_port);
   U88 : OAI22_X1 port map( A1 => n77, A2 => n37, B1 => n43, B2 => n45, ZN => 
                           A_SHF_10_port);
   U89 : NOR2_X1 port map( A1 => n40, A2 => n85, ZN => B_SHF_11_port);
   U90 : NOR2_X1 port map( A1 => n173, A2 => n26, ZN => B_MUL_15_port);
   U91 : OAI22_X1 port map( A1 => n190, A2 => n35, B1 => n41, B2 => n67, ZN => 
                           A_SHF_30_port);
   U92 : NOR2_X1 port map( A1 => n39, A2 => n176, ZN => B_SHF_18_port);
   U93 : NOR2_X1 port map( A1 => n38, A2 => n188, ZN => B_SHF_29_port);
   U94 : NOR2_X1 port map( A1 => n38, A2 => n190, ZN => B_SHF_30_port);
   U95 : BUF_X1 port map( A => n205, Z => n7);
   U96 : BUF_X1 port map( A => n205, Z => n8);
   U97 : BUF_X1 port map( A => n205, Z => n9);
   U98 : BUF_X1 port map( A => n205, Z => n11);
   U99 : BUF_X1 port map( A => n205, Z => n10);
   U100 : NOR2_X1 port map( A1 => n39, A2 => n184, ZN => B_SHF_25_port);
   U101 : NOR2_X1 port map( A1 => n40, A2 => n76, ZN => B_SHF_0_port);
   U102 : NOR2_X1 port map( A1 => n39, A2 => n174, ZN => B_SHF_16_port);
   U103 : NOR2_X1 port map( A1 => n39, A2 => n175, ZN => B_SHF_17_port);
   U104 : NOR2_X1 port map( A1 => n40, A2 => n173, ZN => B_SHF_15_port);
   U105 : NOR2_X1 port map( A1 => n50, A2 => n25, ZN => A_MUL_15_port);
   U106 : NOR2_X1 port map( A1 => n189, A2 => n26, ZN => B_MUL_2_port);
   U107 : NOR2_X1 port map( A1 => n193, A2 => n25, ZN => B_MUL_4_port);
   U108 : NOR2_X1 port map( A1 => n195, A2 => n26, ZN => B_MUL_6_port);
   U109 : NOR2_X1 port map( A1 => n197, A2 => n25, ZN => B_MUL_8_port);
   U110 : NOR2_X1 port map( A1 => n76, A2 => n26, ZN => B_MUL_0_port);
   U111 : NOR2_X1 port map( A1 => n77, A2 => n26, ZN => B_MUL_10_port);
   U112 : NOR2_X1 port map( A1 => n86, A2 => n26, ZN => B_MUL_12_port);
   U113 : NOR2_X1 port map( A1 => n172, A2 => n26, ZN => B_MUL_14_port);
   U114 : BUF_X1 port map( A => n199, Z => n5);
   U115 : BUF_X1 port map( A => n199, Z => n4);
   U116 : OAI21_X1 port map( B1 => n43, B2 => n193, A => n37, ZN => 
                           B_SHF_4_port);
   U117 : BUF_X1 port map( A => n199, Z => n6);
   U118 : NOR2_X1 port map( A1 => n39, A2 => n183, ZN => B_SHF_24_port);
   U119 : NOR2_X1 port map( A1 => n39, A2 => n182, ZN => B_SHF_23_port);
   U120 : NOR2_X1 port map( A1 => n39, A2 => n181, ZN => B_SHF_22_port);
   U121 : NOR2_X1 port map( A1 => n30, A2 => n67, ZN => A_CMP_30_port);
   U122 : OAI22_X1 port map( A1 => n99, A2 => n194, B1 => n100, B2 => n71, ZN 
                           => LOGIC_RES_5_port);
   U123 : OAI22_X1 port map( A1 => n97, A2 => n195, B1 => n98, B2 => n72, ZN =>
                           LOGIC_RES_6_port);
   U124 : OAI22_X1 port map( A1 => n95, A2 => n196, B1 => n96, B2 => n73, ZN =>
                           LOGIC_RES_7_port);
   U125 : OAI22_X1 port map( A1 => n90, A2 => n198, B1 => n91, B2 => n75, ZN =>
                           LOGIC_RES_9_port);
   U126 : OAI22_X1 port map( A1 => n105, A2 => n191, B1 => n106, B2 => n68, ZN 
                           => LOGIC_RES_31_port);
   U127 : NOR2_X1 port map( A1 => n29, A2 => n55, ZN => A_CMP_1_port);
   U128 : OAI22_X1 port map( A1 => n151, A2 => n77, B1 => n152, B2 => n45, ZN 
                           => LOGIC_RES_10_port);
   U129 : OAI22_X1 port map( A1 => n149, A2 => n85, B1 => n150, B2 => n46, ZN 
                           => LOGIC_RES_11_port);
   U130 : OAI22_X1 port map( A1 => n145, A2 => n171, B1 => n146, B2 => n48, ZN 
                           => LOGIC_RES_13_port);
   U131 : OAI22_X1 port map( A1 => n143, A2 => n172, B1 => n144, B2 => n49, ZN 
                           => LOGIC_RES_14_port);
   U132 : OAI22_X1 port map( A1 => n141, A2 => n173, B1 => n142, B2 => n50, ZN 
                           => LOGIC_RES_15_port);
   U133 : OAI22_X1 port map( A1 => n137, A2 => n175, B1 => n138, B2 => n52, ZN 
                           => LOGIC_RES_17_port);
   U134 : OAI22_X1 port map( A1 => n135, A2 => n176, B1 => n136, B2 => n53, ZN 
                           => LOGIC_RES_18_port);
   U135 : OAI22_X1 port map( A1 => n133, A2 => n177, B1 => n134, B2 => n54, ZN 
                           => LOGIC_RES_19_port);
   U136 : OAI22_X1 port map( A1 => n127, A2 => n180, B1 => n128, B2 => n57, ZN 
                           => LOGIC_RES_21_port);
   U137 : OAI22_X1 port map( A1 => n125, A2 => n181, B1 => n126, B2 => n58, ZN 
                           => LOGIC_RES_22_port);
   U138 : OAI22_X1 port map( A1 => n123, A2 => n182, B1 => n124, B2 => n59, ZN 
                           => LOGIC_RES_23_port);
   U139 : OAI22_X1 port map( A1 => n119, A2 => n184, B1 => n120, B2 => n61, ZN 
                           => LOGIC_RES_25_port);
   U140 : OAI22_X1 port map( A1 => n117, A2 => n185, B1 => n118, B2 => n62, ZN 
                           => LOGIC_RES_26_port);
   U141 : OAI22_X1 port map( A1 => n115, A2 => n186, B1 => n116, B2 => n63, ZN 
                           => LOGIC_RES_27_port);
   U142 : OAI22_X1 port map( A1 => n111, A2 => n188, B1 => n112, B2 => n65, ZN 
                           => LOGIC_RES_29_port);
   U143 : OAI22_X1 port map( A1 => n107, A2 => n190, B1 => n108, B2 => n67, ZN 
                           => LOGIC_RES_30_port);
   U144 : NOR2_X1 port map( A1 => n39, A2 => n177, ZN => B_SHF_19_port);
   U145 : NOR2_X1 port map( A1 => n39, A2 => n180, ZN => B_SHF_21_port);
   U146 : NOR2_X1 port map( A1 => n40, A2 => n171, ZN => B_SHF_13_port);
   U147 : NOR2_X1 port map( A1 => n39, A2 => n179, ZN => B_SHF_20_port);
   U148 : NOR2_X1 port map( A1 => n40, A2 => n172, ZN => B_SHF_14_port);
   U149 : NOR2_X1 port map( A1 => n40, A2 => n86, ZN => B_SHF_12_port);
   U150 : NOR2_X1 port map( A1 => n34, A2 => n196, ZN => B_CMP_7_port);
   U151 : NOR2_X1 port map( A1 => n34, A2 => n198, ZN => B_CMP_9_port);
   U152 : AOI21_X1 port map( B1 => n9, B2 => n194, A => n21, ZN => n100);
   U153 : AOI21_X1 port map( B1 => n9, B2 => n195, A => n21, ZN => n98);
   U154 : AOI21_X1 port map( B1 => n9, B2 => n197, A => n21, ZN => n94);
   U155 : AOI21_X1 port map( B1 => n11, B2 => n178, A => n23, ZN => n132);
   U156 : AOI21_X1 port map( B1 => n10, B2 => n189, A => n22, ZN => n110);
   U157 : AOI21_X1 port map( B1 => n10, B2 => n192, A => n22, ZN => n104);
   U158 : AOI21_X1 port map( B1 => n10, B2 => n193, A => n22, ZN => n102);
   U159 : AOI21_X1 port map( B1 => n10, B2 => n196, A => n22, ZN => n96);
   U160 : AOI21_X1 port map( B1 => n10, B2 => n198, A => n22, ZN => n91);
   U161 : AOI21_X1 port map( B1 => n11, B2 => n172, A => n23, ZN => n144);
   U162 : AOI21_X1 port map( B1 => n11, B2 => n173, A => n23, ZN => n142);
   U163 : AOI21_X1 port map( B1 => n11, B2 => n174, A => n23, ZN => n140);
   U164 : AOI21_X1 port map( B1 => n11, B2 => n175, A => n23, ZN => n138);
   U165 : AOI21_X1 port map( B1 => n11, B2 => n176, A => n23, ZN => n136);
   U166 : AOI21_X1 port map( B1 => n11, B2 => n177, A => n23, ZN => n134);
   U167 : AOI21_X1 port map( B1 => n11, B2 => n179, A => n23, ZN => n130);
   U168 : AOI21_X1 port map( B1 => n11, B2 => n180, A => n23, ZN => n128);
   U169 : AOI21_X1 port map( B1 => n11, B2 => n181, A => n23, ZN => n126);
   U170 : AOI21_X1 port map( B1 => n11, B2 => n182, A => n23, ZN => n124);
   U171 : AOI21_X1 port map( B1 => n11, B2 => n183, A => n22, ZN => n122);
   U172 : AOI21_X1 port map( B1 => n10, B2 => n184, A => n22, ZN => n120);
   U173 : AOI21_X1 port map( B1 => n10, B2 => n185, A => n22, ZN => n118);
   U174 : AOI21_X1 port map( B1 => n10, B2 => n186, A => n22, ZN => n116);
   U175 : AOI21_X1 port map( B1 => n10, B2 => n187, A => n22, ZN => n114);
   U176 : AOI21_X1 port map( B1 => n10, B2 => n188, A => n22, ZN => n112);
   U177 : AOI21_X1 port map( B1 => n10, B2 => n190, A => n22, ZN => n108);
   U178 : AOI21_X1 port map( B1 => n10, B2 => n191, A => n22, ZN => n106);
   U179 : AOI21_X1 port map( B1 => n12, B2 => n77, A => n24, ZN => n152);
   U180 : AOI21_X1 port map( B1 => n12, B2 => n85, A => n24, ZN => n150);
   U181 : AOI21_X1 port map( B1 => n12, B2 => n86, A => n23, ZN => n148);
   U182 : AOI21_X1 port map( B1 => n12, B2 => n171, A => n23, ZN => n146);
   U183 : NOR2_X1 port map( A1 => n34, A2 => n197, ZN => B_CMP_8_port);
   U184 : NOR2_X1 port map( A1 => n34, A2 => n195, ZN => B_CMP_6_port);
   U185 : NOR2_X1 port map( A1 => n33, A2 => n190, ZN => B_CMP_30_port);
   U186 : NOR2_X1 port map( A1 => n31, A2 => n76, ZN => B_CMP_0_port);
   U187 : NOR2_X1 port map( A1 => n33, A2 => n192, ZN => B_CMP_3_port);
   U188 : NOR2_X1 port map( A1 => n33, A2 => n194, ZN => B_CMP_5_port);
   U189 : NOR2_X1 port map( A1 => n31, A2 => n85, ZN => B_CMP_11_port);
   U190 : NOR2_X1 port map( A1 => n32, A2 => n171, ZN => B_CMP_13_port);
   U191 : NOR2_X1 port map( A1 => n32, A2 => n173, ZN => B_CMP_15_port);
   U192 : NOR2_X1 port map( A1 => n32, A2 => n175, ZN => B_CMP_17_port);
   U193 : NOR2_X1 port map( A1 => n32, A2 => n177, ZN => B_CMP_19_port);
   U194 : NOR2_X1 port map( A1 => n32, A2 => n180, ZN => B_CMP_21_port);
   U195 : NOR2_X1 port map( A1 => n32, A2 => n182, ZN => B_CMP_23_port);
   U196 : NOR2_X1 port map( A1 => n33, A2 => n184, ZN => B_CMP_25_port);
   U197 : NOR2_X1 port map( A1 => n33, A2 => n186, ZN => B_CMP_27_port);
   U198 : NOR2_X1 port map( A1 => n33, A2 => n188, ZN => B_CMP_29_port);
   U199 : NOR2_X1 port map( A1 => n31, A2 => n68, ZN => A_CMP_31_port);
   U200 : NOR2_X1 port map( A1 => n33, A2 => n193, ZN => B_CMP_4_port);
   U201 : NOR2_X1 port map( A1 => n31, A2 => n86, ZN => B_CMP_12_port);
   U202 : NOR2_X1 port map( A1 => n32, A2 => n174, ZN => B_CMP_16_port);
   U203 : NOR2_X1 port map( A1 => n32, A2 => n179, ZN => B_CMP_20_port);
   U204 : NOR2_X1 port map( A1 => n33, A2 => n183, ZN => B_CMP_24_port);
   U205 : NOR2_X1 port map( A1 => n33, A2 => n187, ZN => B_CMP_28_port);
   U206 : NOR2_X1 port map( A1 => n33, A2 => n189, ZN => B_CMP_2_port);
   U207 : NOR2_X1 port map( A1 => n31, A2 => n77, ZN => B_CMP_10_port);
   U208 : NOR2_X1 port map( A1 => n32, A2 => n172, ZN => B_CMP_14_port);
   U209 : NOR2_X1 port map( A1 => n32, A2 => n176, ZN => B_CMP_18_port);
   U210 : NOR2_X1 port map( A1 => n32, A2 => n181, ZN => B_CMP_22_port);
   U211 : NOR2_X1 port map( A1 => n33, A2 => n185, ZN => B_CMP_26_port);
   U212 : AND2_X1 port map( A1 => n18, A2 => n6, ZN => n168);
   U213 : NOR2_X1 port map( A1 => n38, A2 => n191, ZN => B_SHF_31_port);
   U214 : NOR2_X1 port map( A1 => n32, A2 => n178, ZN => B_CMP_1_port);
   U215 : NOR2_X1 port map( A1 => n29, A2 => n44, ZN => A_CMP_0_port);
   U216 : NOR2_X1 port map( A1 => n31, A2 => n69, ZN => A_CMP_3_port);
   U217 : NOR2_X1 port map( A1 => n31, A2 => n71, ZN => A_CMP_5_port);
   U218 : NOR2_X1 port map( A1 => n31, A2 => n73, ZN => A_CMP_7_port);
   U219 : NOR2_X1 port map( A1 => n31, A2 => n75, ZN => A_CMP_9_port);
   U220 : NOR2_X1 port map( A1 => n29, A2 => n46, ZN => A_CMP_11_port);
   U221 : NOR2_X1 port map( A1 => n29, A2 => n48, ZN => A_CMP_13_port);
   U222 : NOR2_X1 port map( A1 => n29, A2 => n50, ZN => A_CMP_15_port);
   U223 : NOR2_X1 port map( A1 => n33, A2 => n191, ZN => B_CMP_31_port);
   U224 : NOR2_X1 port map( A1 => n29, A2 => n52, ZN => A_CMP_17_port);
   U225 : NOR2_X1 port map( A1 => n29, A2 => n54, ZN => A_CMP_19_port);
   U226 : NOR2_X1 port map( A1 => n30, A2 => n57, ZN => A_CMP_21_port);
   U228 : NOR2_X1 port map( A1 => n30, A2 => n59, ZN => A_CMP_23_port);
   U229 : NOR2_X1 port map( A1 => n30, A2 => n61, ZN => A_CMP_25_port);
   U230 : NOR2_X1 port map( A1 => n30, A2 => n63, ZN => A_CMP_27_port);
   U231 : NOR2_X1 port map( A1 => n30, A2 => n65, ZN => A_CMP_29_port);
   U232 : NOR2_X1 port map( A1 => n31, A2 => n70, ZN => A_CMP_4_port);
   U233 : NOR2_X1 port map( A1 => n31, A2 => n74, ZN => A_CMP_8_port);
   U234 : NOR2_X1 port map( A1 => n29, A2 => n47, ZN => A_CMP_12_port);
   U235 : NOR2_X1 port map( A1 => n30, A2 => n66, ZN => A_CMP_2_port);
   U236 : NOR2_X1 port map( A1 => n31, A2 => n72, ZN => A_CMP_6_port);
   U237 : NOR2_X1 port map( A1 => n29, A2 => n45, ZN => A_CMP_10_port);
   U238 : NOR2_X1 port map( A1 => n29, A2 => n49, ZN => A_CMP_14_port);
   U239 : NOR2_X1 port map( A1 => n29, A2 => n51, ZN => A_CMP_16_port);
   U240 : NOR2_X1 port map( A1 => n30, A2 => n56, ZN => A_CMP_20_port);
   U241 : NOR2_X1 port map( A1 => n30, A2 => n60, ZN => A_CMP_24_port);
   U242 : NOR2_X1 port map( A1 => n30, A2 => n64, ZN => A_CMP_28_port);
   U243 : NOR2_X1 port map( A1 => n29, A2 => n53, ZN => A_CMP_18_port);
   U244 : NOR2_X1 port map( A1 => n30, A2 => n58, ZN => A_CMP_22_port);
   U245 : NOR2_X1 port map( A1 => n30, A2 => n62, ZN => A_CMP_26_port);
   U246 : OAI22_X1 port map( A1 => OP2(0), A2 => n6, B1 => n76, B2 => n18, ZN 
                           => B_ADD_0_port);
   U247 : OAI22_X1 port map( A1 => OP2(4), A2 => n4, B1 => n193, B2 => n16, ZN 
                           => B_ADD_4_port);
   U248 : OAI22_X1 port map( A1 => OP2(8), A2 => n4, B1 => n197, B2 => n16, ZN 
                           => B_ADD_8_port);
   U249 : OAI22_X1 port map( A1 => OP2(12), A2 => n6, B1 => n86, B2 => n18, ZN 
                           => B_ADD_12_port);
   U250 : OAI22_X1 port map( A1 => OP2(16), A2 => n6, B1 => n174, B2 => n18, ZN
                           => B_ADD_16_port);
   U251 : OAI22_X1 port map( A1 => OP2(24), A2 => n5, B1 => n183, B2 => n17, ZN
                           => B_ADD_24_port);
   U252 : OAI22_X1 port map( A1 => OP2(5), A2 => n4, B1 => n194, B2 => n16, ZN 
                           => B_ADD_5_port);
   U253 : OAI22_X1 port map( A1 => OP2(1), A2 => n5, B1 => n178, B2 => n17, ZN 
                           => B_ADD_1_port);
   U254 : OAI22_X1 port map( A1 => OP2(9), A2 => n4, B1 => n198, B2 => n16, ZN 
                           => B_ADD_9_port);
   U255 : OAI22_X1 port map( A1 => OP2(13), A2 => n6, B1 => n171, B2 => n18, ZN
                           => B_ADD_13_port);
   U256 : OAI22_X1 port map( A1 => OP2(17), A2 => n5, B1 => n175, B2 => n17, ZN
                           => B_ADD_17_port);
   U266 : OAI22_X1 port map( A1 => OP2(25), A2 => n5, B1 => n184, B2 => n17, ZN
                           => B_ADD_25_port);
   U273 : OAI22_X1 port map( A1 => OP2(2), A2 => n4, B1 => n189, B2 => n16, ZN 
                           => B_ADD_2_port);
   U274 : OAI22_X1 port map( A1 => OP2(6), A2 => n4, B1 => n195, B2 => n16, ZN 
                           => B_ADD_6_port);
   U275 : OAI22_X1 port map( A1 => OP2(10), A2 => n6, B1 => n77, B2 => n18, ZN 
                           => B_ADD_10_port);
   U276 : OAI22_X1 port map( A1 => OP2(14), A2 => n6, B1 => n172, B2 => n18, ZN
                           => B_ADD_14_port);
   U277 : OAI22_X1 port map( A1 => OP2(18), A2 => n5, B1 => n176, B2 => n17, ZN
                           => B_ADD_18_port);
   U278 : OAI22_X1 port map( A1 => OP2(26), A2 => n5, B1 => n185, B2 => n17, ZN
                           => B_ADD_26_port);
   U279 : OAI22_X1 port map( A1 => OP2(22), A2 => n5, B1 => n181, B2 => n17, ZN
                           => B_ADD_22_port);
   U280 : OAI22_X1 port map( A1 => OP2(21), A2 => n5, B1 => n180, B2 => n17, ZN
                           => B_ADD_21_port);
   U281 : OAI22_X1 port map( A1 => OP2(20), A2 => n5, B1 => n179, B2 => n17, ZN
                           => B_ADD_20_port);
   U282 : OAI22_X1 port map( A1 => OP2(30), A2 => n4, B1 => n190, B2 => n16, ZN
                           => B_ADD_30_port);
   U283 : OAI22_X1 port map( A1 => OP2(29), A2 => n4, B1 => n188, B2 => n16, ZN
                           => B_ADD_29_port);
   U284 : OAI22_X1 port map( A1 => OP2(28), A2 => n4, B1 => n187, B2 => n16, ZN
                           => B_ADD_28_port);
   U285 : OAI22_X1 port map( A1 => OP2(3), A2 => n4, B1 => n192, B2 => n16, ZN 
                           => B_ADD_3_port);
   U286 : OAI22_X1 port map( A1 => OP2(7), A2 => n4, B1 => n196, B2 => n16, ZN 
                           => B_ADD_7_port);
   U287 : OAI22_X1 port map( A1 => OP2(11), A2 => n6, B1 => n85, B2 => n18, ZN 
                           => B_ADD_11_port);
   U288 : OAI22_X1 port map( A1 => OP2(15), A2 => n6, B1 => n173, B2 => n18, ZN
                           => B_ADD_15_port);
   U289 : OAI22_X1 port map( A1 => OP2(19), A2 => n5, B1 => n177, B2 => n17, ZN
                           => B_ADD_19_port);
   U290 : OAI22_X1 port map( A1 => OP2(23), A2 => n5, B1 => n182, B2 => n17, ZN
                           => B_ADD_23_port);
   U291 : OAI22_X1 port map( A1 => OP2(27), A2 => n5, B1 => n186, B2 => n17, ZN
                           => B_ADD_27_port);
   U292 : OAI22_X1 port map( A1 => OP2(31), A2 => n4, B1 => n191, B2 => n16, ZN
                           => B_ADD_31_port);
   U293 : INV_X1 port map( A => n1, ZN => n26);
   U294 : INV_X1 port map( A => n1, ZN => n25);
   U295 : INV_X1 port map( A => n3, ZN => n27);
   U296 : INV_X1 port map( A => n3, ZN => n28);
   U297 : INV_X1 port map( A => ADD_SUB, ZN => n199);
   U298 : AOI221_X1 port map( B1 => OP1(10), B2 => n27, C1 => n7, C2 => n45, A 
                           => n19, ZN => n151);
   U299 : AOI221_X1 port map( B1 => OP1(11), B2 => n28, C1 => n7, C2 => n46, A 
                           => n19, ZN => n149);
   U300 : AOI221_X1 port map( B1 => OP1(12), B2 => n27, C1 => n7, C2 => n47, A 
                           => n19, ZN => n147);
   U301 : AOI221_X1 port map( B1 => OP1(13), B2 => n28, C1 => n7, C2 => n48, A 
                           => n19, ZN => n145);
   U302 : AOI221_X1 port map( B1 => OP1(14), B2 => n27, C1 => n7, C2 => n49, A 
                           => n19, ZN => n143);
   U303 : AOI221_X1 port map( B1 => OP1(15), B2 => n28, C1 => n7, C2 => n50, A 
                           => n19, ZN => n141);
   U304 : AOI221_X1 port map( B1 => OP1(16), B2 => n27, C1 => n7, C2 => n51, A 
                           => n19, ZN => n139);
   U305 : AOI221_X1 port map( B1 => OP1(1), B2 => n28, C1 => n8, C2 => n55, A 
                           => n20, ZN => n131);
   U306 : AOI221_X1 port map( B1 => OP1(2), B2 => n27, C1 => n9, C2 => n66, A 
                           => n21, ZN => n109);
   U307 : AOI221_X1 port map( B1 => OP1(3), B2 => n27, C1 => n8, C2 => n69, A 
                           => n20, ZN => n103);
   U308 : AOI221_X1 port map( B1 => OP1(4), B2 => n27, C1 => n8, C2 => n70, A 
                           => n20, ZN => n101);
   U309 : AOI221_X1 port map( B1 => OP1(5), B2 => n27, C1 => n8, C2 => n71, A 
                           => n20, ZN => n99);
   U310 : AOI221_X1 port map( B1 => OP1(6), B2 => n27, C1 => n7, C2 => n72, A 
                           => n19, ZN => n97);
   U311 : AOI221_X1 port map( B1 => OP1(7), B2 => n27, C1 => n7, C2 => n73, A 
                           => n19, ZN => n95);
   U312 : AOI221_X1 port map( B1 => OP1(8), B2 => n27, C1 => n7, C2 => n74, A 
                           => n19, ZN => n93);
   U313 : AOI221_X1 port map( B1 => OP1(17), B2 => n28, C1 => n8, C2 => n52, A 
                           => n20, ZN => n137);
   U314 : AOI221_X1 port map( B1 => OP1(18), B2 => n28, C1 => n8, C2 => n53, A 
                           => n20, ZN => n135);
   U315 : AOI221_X1 port map( B1 => OP1(19), B2 => n28, C1 => n8, C2 => n54, A 
                           => n20, ZN => n133);
   U316 : AOI221_X1 port map( B1 => OP1(20), B2 => n28, C1 => n8, C2 => n56, A 
                           => n20, ZN => n129);
   U317 : AOI221_X1 port map( B1 => OP1(21), B2 => n28, C1 => n8, C2 => n57, A 
                           => n20, ZN => n127);
   U318 : AOI221_X1 port map( B1 => OP1(22), B2 => n28, C1 => n8, C2 => n58, A 
                           => n20, ZN => n125);
   U319 : AOI221_X1 port map( B1 => OP1(23), B2 => n28, C1 => n8, C2 => n59, A 
                           => n20, ZN => n123);
   U320 : AOI221_X1 port map( B1 => OP1(24), B2 => n28, C1 => n9, C2 => n60, A 
                           => n21, ZN => n121);
   U321 : AOI221_X1 port map( B1 => OP1(25), B2 => n28, C1 => n9, C2 => n61, A 
                           => n21, ZN => n119);
   U322 : AOI221_X1 port map( B1 => OP1(26), B2 => n28, C1 => n8, C2 => n62, A 
                           => n20, ZN => n117);
   U323 : AOI221_X1 port map( B1 => OP1(27), B2 => n28, C1 => n9, C2 => n63, A 
                           => n21, ZN => n115);
   U324 : AOI221_X1 port map( B1 => OP1(28), B2 => n27, C1 => n9, C2 => n64, A 
                           => n21, ZN => n113);
   U325 : AOI221_X1 port map( B1 => OP1(29), B2 => n27, C1 => n9, C2 => n65, A 
                           => n21, ZN => n111);
   U326 : AOI221_X1 port map( B1 => OP1(30), B2 => n27, C1 => n9, C2 => n67, A 
                           => n21, ZN => n107);
   U327 : AOI221_X1 port map( B1 => OP1(31), B2 => n27, C1 => n9, C2 => n68, A 
                           => n21, ZN => n105);
   U328 : AOI221_X1 port map( B1 => n27, B2 => OP1(9), C1 => n7, C2 => n75, A 
                           => n19, ZN => n90);
   U329 : BUF_X1 port map( A => n81, Z => n39);
   U330 : BUF_X1 port map( A => n81, Z => n40);
   U331 : BUF_X1 port map( A => n81, Z => n41);
   U332 : BUF_X1 port map( A => n81, Z => n42);
   U333 : INV_X1 port map( A => OP2(0), ZN => n76);
   U334 : INV_X1 port map( A => OP2(1), ZN => n178);
   U335 : INV_X1 port map( A => OP2(2), ZN => n189);
   U336 : INV_X1 port map( A => OP2(3), ZN => n192);
   U337 : INV_X1 port map( A => OP2(5), ZN => n194);
   U338 : INV_X1 port map( A => OP2(6), ZN => n195);
   U339 : INV_X1 port map( A => OP2(7), ZN => n196);
   U340 : INV_X1 port map( A => OP2(8), ZN => n197);
   U341 : INV_X1 port map( A => OP2(9), ZN => n198);
   U342 : INV_X1 port map( A => OP2(10), ZN => n77);
   U343 : INV_X1 port map( A => OP2(11), ZN => n85);
   U344 : INV_X1 port map( A => OP2(12), ZN => n86);
   U345 : INV_X1 port map( A => OP2(13), ZN => n171);
   U346 : INV_X1 port map( A => OP2(14), ZN => n172);
   U347 : INV_X1 port map( A => OP2(15), ZN => n173);
   U348 : INV_X1 port map( A => OP2(4), ZN => n193);
   U349 : BUF_X1 port map( A => n92, Z => n19);
   U350 : BUF_X1 port map( A => n92, Z => n20);
   U351 : OAI22_X1 port map( A1 => n153, A2 => n76, B1 => n154, B2 => n44, ZN 
                           => LOGIC_RES_0_port);
   U352 : AOI21_X1 port map( B1 => n9, B2 => n76, A => n21, ZN => n154);
   U353 : AOI221_X1 port map( B1 => OP1(0), B2 => n28, C1 => n7, C2 => n44, A 
                           => n19, ZN => n153);
   U354 : BUF_X1 port map( A => n92, Z => n23);
   U355 : BUF_X1 port map( A => n92, Z => n22);
   U356 : BUF_X1 port map( A => n82, Z => n35);
   U357 : BUF_X1 port map( A => n82, Z => n36);
   U358 : BUF_X1 port map( A => n92, Z => n21);
   U359 : BUF_X1 port map( A => n159, Z => n17);
   U360 : BUF_X1 port map( A => n159, Z => n16);
   U361 : BUF_X1 port map( A => n83, Z => n33);
   U362 : BUF_X1 port map( A => n83, Z => n31);
   U363 : BUF_X1 port map( A => n83, Z => n29);
   U364 : BUF_X1 port map( A => n83, Z => n32);
   U365 : BUF_X1 port map( A => n83, Z => n30);
   U366 : BUF_X1 port map( A => n81, Z => n38);
   U367 : INV_X1 port map( A => OP1(0), ZN => n44);
   U368 : INV_X1 port map( A => OP1(1), ZN => n55);
   U369 : INV_X1 port map( A => OP1(2), ZN => n66);
   U370 : INV_X1 port map( A => OP1(3), ZN => n69);
   U371 : INV_X1 port map( A => OP1(4), ZN => n70);
   U372 : INV_X1 port map( A => OP1(5), ZN => n71);
   U373 : INV_X1 port map( A => OP1(6), ZN => n72);
   U374 : INV_X1 port map( A => OP1(7), ZN => n73);
   U375 : INV_X1 port map( A => OP1(8), ZN => n74);
   U376 : INV_X1 port map( A => OP1(9), ZN => n75);
   U377 : INV_X1 port map( A => OP1(10), ZN => n45);
   U378 : INV_X1 port map( A => OP1(11), ZN => n46);
   U379 : INV_X1 port map( A => OP1(12), ZN => n47);
   U380 : INV_X1 port map( A => OP1(13), ZN => n48);
   U381 : INV_X1 port map( A => OP1(14), ZN => n49);
   U382 : INV_X1 port map( A => OP1(15), ZN => n50);
   U383 : BUF_X1 port map( A => n159, Z => n18);
   U384 : INV_X1 port map( A => OP2(16), ZN => n174);
   U385 : INV_X1 port map( A => OP2(17), ZN => n175);
   U386 : INV_X1 port map( A => OP2(18), ZN => n176);
   U387 : INV_X1 port map( A => OP2(19), ZN => n177);
   U388 : INV_X1 port map( A => OP2(20), ZN => n179);
   U389 : INV_X1 port map( A => OP2(21), ZN => n180);
   U390 : INV_X1 port map( A => OP2(22), ZN => n181);
   U391 : INV_X1 port map( A => OP2(23), ZN => n182);
   U392 : INV_X1 port map( A => OP2(24), ZN => n183);
   U393 : INV_X1 port map( A => OP2(25), ZN => n184);
   U394 : INV_X1 port map( A => OP2(26), ZN => n185);
   U395 : INV_X1 port map( A => OP2(27), ZN => n186);
   U396 : INV_X1 port map( A => OP2(28), ZN => n187);
   U397 : INV_X1 port map( A => OP2(29), ZN => n188);
   U398 : INV_X1 port map( A => OP2(30), ZN => n190);
   U399 : INV_X1 port map( A => OP2(31), ZN => n191);
   U400 : BUF_X1 port map( A => n82, Z => n37);
   U401 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => OPSel_0_port);
   U402 : OAI22_X1 port map( A1 => n103, A2 => n192, B1 => n104, B2 => n69, ZN 
                           => LOGIC_RES_3_port);
   U403 : OAI22_X1 port map( A1 => n101, A2 => n193, B1 => n102, B2 => n70, ZN 
                           => LOGIC_RES_4_port);
   U404 : OAI22_X1 port map( A1 => n93, A2 => n197, B1 => n94, B2 => n74, ZN =>
                           LOGIC_RES_8_port);
   U405 : OAI22_X1 port map( A1 => n131, A2 => n178, B1 => n132, B2 => n55, ZN 
                           => LOGIC_RES_1_port);
   U406 : OAI22_X1 port map( A1 => n109, A2 => n189, B1 => n110, B2 => n66, ZN 
                           => LOGIC_RES_2_port);
   U407 : OAI22_X1 port map( A1 => n147, A2 => n86, B1 => n148, B2 => n47, ZN 
                           => LOGIC_RES_12_port);
   U408 : OAI22_X1 port map( A1 => n139, A2 => n174, B1 => n140, B2 => n51, ZN 
                           => LOGIC_RES_16_port);
   U409 : OAI22_X1 port map( A1 => n129, A2 => n179, B1 => n130, B2 => n56, ZN 
                           => LOGIC_RES_20_port);
   U410 : OAI22_X1 port map( A1 => n121, A2 => n183, B1 => n122, B2 => n60, ZN 
                           => LOGIC_RES_24_port);
   U411 : OAI22_X1 port map( A1 => n113, A2 => n187, B1 => n114, B2 => n64, ZN 
                           => LOGIC_RES_28_port);
   U412 : INV_X1 port map( A => OP1(16), ZN => n51);
   U413 : INV_X1 port map( A => OP1(17), ZN => n52);
   U414 : INV_X1 port map( A => OP1(18), ZN => n53);
   U415 : INV_X1 port map( A => OP1(19), ZN => n54);
   U416 : INV_X1 port map( A => OP1(20), ZN => n56);
   U417 : INV_X1 port map( A => OP1(21), ZN => n57);
   U418 : INV_X1 port map( A => OP1(22), ZN => n58);
   U419 : INV_X1 port map( A => OP1(23), ZN => n59);
   U420 : INV_X1 port map( A => OP1(24), ZN => n60);
   U421 : INV_X1 port map( A => OP1(25), ZN => n61);
   U422 : INV_X1 port map( A => OP1(26), ZN => n62);
   U423 : INV_X1 port map( A => OP1(27), ZN => n63);
   U424 : INV_X1 port map( A => OP1(28), ZN => n64);
   U425 : INV_X1 port map( A => OP1(29), ZN => n65);
   U426 : INV_X1 port map( A => OP1(30), ZN => n67);
   U433 : INV_X1 port map( A => OP1(31), ZN => n68);
   U437 : NAND2_X1 port map( A1 => n157, A2 => n204, ZN => LOGIC_ARITH);
   U438 : INV_X1 port map( A => LEFT_RIGHT, ZN => n204);
   U439 : INV_X1 port map( A => n84, ZN => n205);
   U440 : INV_X1 port map( A => n87, ZN => n203);
   U441 : INV_X1 port map( A => n80, ZN => n202);
   U442 : NOR3_X1 port map( A1 => n209, A2 => ALU_OPC(1), A3 => n207, ZN => 
                           n162);
   U443 : NOR3_X1 port map( A1 => ALU_OPC(1), A2 => ALU_OPC(0), A3 => 
                           ALU_OPC(2), ZN => n80);
   U444 : NAND4_X1 port map( A1 => ALU_OPC(0), A2 => ALU_OPC(3), A3 => n209, A4
                           => n206, ZN => n88);
   U445 : NAND4_X1 port map( A1 => ALU_OPC(3), A2 => ALU_OPC(1), A3 => 
                           ALU_OPC(2), A4 => n201, ZN => n89);
   U446 : INV_X1 port map( A => ALU_OPC(3), ZN => n208);
   U447 : NAND2_X1 port map( A1 => n158, A2 => n35, ZN => LEFT_RIGHT);
   U448 : NOR3_X1 port map( A1 => ALU_OPC(3), A2 => ALU_OPC(0), A3 => 
                           ALU_OPC(2), ZN => n156);
   U449 : NAND4_X1 port map( A1 => ALU_OPC(3), A2 => ALU_OPC(1), A3 => n161, A4
                           => n209, ZN => n157);
   U450 : NOR2_X1 port map( A1 => ALU_OPC(0), A2 => ALU_OPC(2), ZN => n161);
   U451 : INV_X1 port map( A => ALU_OPC(2), ZN => n207);
   U452 : INV_X1 port map( A => ALU_OPC(1), ZN => n206);
   U453 : OAI211_X1 port map( C1 => n166, C2 => n167, A => n206, B => 
                           ALU_OPC(0), ZN => n87);
   U454 : NOR2_X1 port map( A1 => ALU_OPC(2), A2 => n208, ZN => n167);
   U455 : NOR3_X1 port map( A1 => n207, A2 => ALU_OPC(3), A3 => ALU_OPC(4), ZN 
                           => n166);
   U456 : AND3_X1 port map( A1 => ALU_OPC(3), A2 => ALU_OPC(4), A3 => n155, ZN 
                           => n92);
   U457 : NOR3_X1 port map( A1 => n207, A2 => ALU_OPC(0), A3 => ALU_OPC(1), ZN 
                           => n155);
   U458 : INV_X1 port map( A => ALU_OPC(0), ZN => n201);
   U459 : INV_X1 port map( A => ALU_OPC(4), ZN => n209);
   U460 : OAI21_X1 port map( B1 => n78, B2 => n206, A => n79, ZN => 
                           select_zero_sig);
   U461 : AOI21_X1 port map( B1 => ALU_OPC(2), B2 => n208, A => ALU_OPC(0), ZN 
                           => n78);
   U462 : NAND2_X1 port map( A1 => n165, A2 => n89, ZN => OPSel_1_port);
   U463 : NAND4_X1 port map( A1 => ALU_OPC(0), A2 => n208, A3 => n207, A4 => 
                           n206, ZN => n165);
   U464 : NAND2_X1 port map( A1 => n80, A2 => n169, ZN => n159);
   U465 : XNOR2_X1 port map( A => n208, B => ALU_OPC(4), ZN => n169);
   U466 : AND4_X1 port map( A1 => n164, A2 => n88, A3 => n87, A4 => n200, ZN =>
                           n83);
   U467 : INV_X1 port map( A => OPSel_1_port, ZN => n200);
   U468 : OR4_X1 port map( A1 => n208, A2 => n207, A3 => ALU_OPC(1), A4 => 
                           ALU_OPC(0), ZN => n3);
   U469 : AND2_X1 port map( A1 => n160, A2 => n157, ZN => n81);
   U470 : NAND4_X1 port map( A1 => ALU_OPC(4), A2 => ALU_OPC(1), A3 => n207, A4
                           => n201, ZN => n160);
   U471 : NOR3_X1 port map( A1 => ALU_OPC(3), A2 => ALU_OPC(0), A3 => 
                           ALU_OPC(1), ZN => n163);
   U472 : CLKBUF_X1 port map( A => n205, Z => n12);
   U473 : CLKBUF_X1 port map( A => n92, Z => n24);
   U474 : CLKBUF_X1 port map( A => n83, Z => n34);
   U475 : CLKBUF_X1 port map( A => n81, Z => n43);
   COMP_RES_1_port <= '0';
   COMP_RES_2_port <= '0';
   COMP_RES_3_port <= '0';
   COMP_RES_4_port <= '0';
   COMP_RES_5_port <= '0';
   COMP_RES_6_port <= '0';
   COMP_RES_7_port <= '0';
   COMP_RES_8_port <= '0';
   COMP_RES_9_port <= '0';
   COMP_RES_10_port <= '0';
   COMP_RES_11_port <= '0';
   COMP_RES_12_port <= '0';
   COMP_RES_13_port <= '0';
   COMP_RES_14_port <= '0';
   COMP_RES_15_port <= '0';
   COMP_RES_16_port <= '0';
   COMP_RES_17_port <= '0';
   COMP_RES_18_port <= '0';
   COMP_RES_19_port <= '0';
   COMP_RES_20_port <= '0';
   COMP_RES_21_port <= '0';
   COMP_RES_22_port <= '0';
   COMP_RES_23_port <= '0';
   COMP_RES_24_port <= '0';
   COMP_RES_25_port <= '0';
   COMP_RES_26_port <= '0';
   COMP_RES_27_port <= '0';
   COMP_RES_28_port <= '0';
   COMP_RES_29_port <= '0';
   COMP_RES_30_port <= '0';
   COMP_RES_31_port <= '0';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux41_NBIT32_0 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto 0)
         );

end mux41_NBIT32_0;

architecture SYN_bhv of mux41_NBIT32_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n1, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n6, Z => n72);
   U2 : BUF_X1 port map( A => n6, Z => n73);
   U3 : BUF_X1 port map( A => n4, Z => n78);
   U4 : BUF_X1 port map( A => n4, Z => n79);
   U5 : BUF_X1 port map( A => n7, Z => n1);
   U6 : BUF_X1 port map( A => n7, Z => n70);
   U7 : BUF_X1 port map( A => n5, Z => n75);
   U8 : BUF_X1 port map( A => n5, Z => n76);
   U9 : BUF_X1 port map( A => n6, Z => n74);
   U10 : BUF_X1 port map( A => n4, Z => n80);
   U11 : BUF_X1 port map( A => n7, Z => n71);
   U12 : BUF_X1 port map( A => n5, Z => n77);
   U13 : NOR2_X1 port map( A1 => n81, A2 => S(1), ZN => n6);
   U14 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n7);
   U15 : AND2_X1 port map( A1 => S(1), A2 => S(0), ZN => n4);
   U16 : AND2_X1 port map( A1 => S(1), A2 => n81, ZN => n5);
   U17 : INV_X1 port map( A => S(0), ZN => n81);
   U18 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => Z(0));
   U19 : AOI22_X1 port map( A1 => B(0), A2 => n72, B1 => A(0), B2 => n1, ZN => 
                           n68);
   U20 : AOI22_X1 port map( A1 => D(0), A2 => n78, B1 => C(0), B2 => n75, ZN =>
                           n69);
   U21 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => Z(20));
   U22 : AOI22_X1 port map( A1 => B(20), A2 => n73, B1 => A(20), B2 => n70, ZN 
                           => n44);
   U23 : AOI22_X1 port map( A1 => D(20), A2 => n79, B1 => C(20), B2 => n76, ZN 
                           => n45);
   U24 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => Z(17));
   U25 : AOI22_X1 port map( A1 => B(17), A2 => n72, B1 => A(17), B2 => n1, ZN 
                           => n52);
   U26 : AOI22_X1 port map( A1 => D(17), A2 => n78, B1 => C(17), B2 => n75, ZN 
                           => n53);
   U27 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => Z(13));
   U28 : AOI22_X1 port map( A1 => B(13), A2 => n72, B1 => A(13), B2 => n1, ZN 
                           => n60);
   U29 : AOI22_X1 port map( A1 => D(13), A2 => n78, B1 => C(13), B2 => n75, ZN 
                           => n61);
   U30 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => Z(6));
   U31 : AOI22_X1 port map( A1 => B(6), A2 => n74, B1 => A(6), B2 => n71, ZN =>
                           n12);
   U32 : AOI22_X1 port map( A1 => D(6), A2 => n80, B1 => C(6), B2 => n77, ZN =>
                           n13);
   U33 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => Z(31));
   U34 : AOI22_X1 port map( A1 => B(31), A2 => n74, B1 => A(31), B2 => n71, ZN 
                           => n20);
   U35 : AOI22_X1 port map( A1 => D(31), A2 => n80, B1 => C(31), B2 => n77, ZN 
                           => n21);
   U36 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => Z(28));
   U37 : AOI22_X1 port map( A1 => B(28), A2 => n73, B1 => A(28), B2 => n70, ZN 
                           => n28);
   U38 : AOI22_X1 port map( A1 => D(28), A2 => n79, B1 => C(28), B2 => n76, ZN 
                           => n29);
   U39 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => Z(24));
   U40 : AOI22_X1 port map( A1 => B(24), A2 => n73, B1 => A(24), B2 => n70, ZN 
                           => n36);
   U41 : AOI22_X1 port map( A1 => D(24), A2 => n79, B1 => C(24), B2 => n76, ZN 
                           => n37);
   U42 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => Z(21));
   U43 : AOI22_X1 port map( A1 => B(21), A2 => n73, B1 => A(21), B2 => n70, ZN 
                           => n42);
   U44 : AOI22_X1 port map( A1 => D(21), A2 => n79, B1 => C(21), B2 => n76, ZN 
                           => n43);
   U45 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => Z(18));
   U46 : AOI22_X1 port map( A1 => B(18), A2 => n72, B1 => A(18), B2 => n1, ZN 
                           => n50);
   U47 : AOI22_X1 port map( A1 => D(18), A2 => n78, B1 => C(18), B2 => n75, ZN 
                           => n51);
   U48 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => Z(14));
   U49 : AOI22_X1 port map( A1 => B(14), A2 => n72, B1 => A(14), B2 => n1, ZN 
                           => n58);
   U50 : AOI22_X1 port map( A1 => D(14), A2 => n78, B1 => C(14), B2 => n75, ZN 
                           => n59);
   U51 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => Z(10));
   U52 : AOI22_X1 port map( A1 => B(10), A2 => n72, B1 => A(10), B2 => n1, ZN 
                           => n66);
   U53 : AOI22_X1 port map( A1 => D(10), A2 => n78, B1 => C(10), B2 => n75, ZN 
                           => n67);
   U54 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => Z(7));
   U55 : AOI22_X1 port map( A1 => B(7), A2 => n74, B1 => A(7), B2 => n71, ZN =>
                           n10);
   U56 : AOI22_X1 port map( A1 => D(7), A2 => n80, B1 => C(7), B2 => n77, ZN =>
                           n11);
   U57 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => Z(29));
   U58 : AOI22_X1 port map( A1 => B(29), A2 => n73, B1 => A(29), B2 => n70, ZN 
                           => n26);
   U59 : AOI22_X1 port map( A1 => D(29), A2 => n79, B1 => C(29), B2 => n76, ZN 
                           => n27);
   U60 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => Z(25));
   U61 : AOI22_X1 port map( A1 => B(25), A2 => n73, B1 => A(25), B2 => n70, ZN 
                           => n34);
   U62 : AOI22_X1 port map( A1 => D(25), A2 => n79, B1 => C(25), B2 => n76, ZN 
                           => n35);
   U63 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => Z(3));
   U64 : AOI22_X1 port map( A1 => B(3), A2 => n74, B1 => A(3), B2 => n71, ZN =>
                           n18);
   U65 : AOI22_X1 port map( A1 => D(3), A2 => n80, B1 => C(3), B2 => n77, ZN =>
                           n19);
   U66 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => Z(22));
   U67 : AOI22_X1 port map( A1 => B(22), A2 => n73, B1 => A(22), B2 => n70, ZN 
                           => n40);
   U68 : AOI22_X1 port map( A1 => D(22), A2 => n79, B1 => C(22), B2 => n76, ZN 
                           => n41);
   U69 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => Z(19));
   U70 : AOI22_X1 port map( A1 => B(19), A2 => n72, B1 => A(19), B2 => n1, ZN 
                           => n48);
   U71 : AOI22_X1 port map( A1 => D(19), A2 => n78, B1 => C(19), B2 => n75, ZN 
                           => n49);
   U72 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => Z(15));
   U73 : AOI22_X1 port map( A1 => B(15), A2 => n72, B1 => A(15), B2 => n1, ZN 
                           => n56);
   U74 : AOI22_X1 port map( A1 => D(15), A2 => n78, B1 => C(15), B2 => n75, ZN 
                           => n57);
   U75 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => Z(11));
   U76 : AOI22_X1 port map( A1 => B(11), A2 => n72, B1 => A(11), B2 => n1, ZN 
                           => n64);
   U77 : AOI22_X1 port map( A1 => D(11), A2 => n78, B1 => C(11), B2 => n75, ZN 
                           => n65);
   U78 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => Z(8));
   U79 : AOI22_X1 port map( A1 => B(8), A2 => n74, B1 => A(8), B2 => n71, ZN =>
                           n8);
   U80 : AOI22_X1 port map( A1 => D(8), A2 => n80, B1 => C(8), B2 => n77, ZN =>
                           n9);
   U81 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => Z(4));
   U82 : AOI22_X1 port map( A1 => B(4), A2 => n74, B1 => A(4), B2 => n71, ZN =>
                           n16);
   U83 : AOI22_X1 port map( A1 => D(4), A2 => n80, B1 => C(4), B2 => n77, ZN =>
                           n17);
   U84 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => Z(2));
   U85 : AOI22_X1 port map( A1 => B(2), A2 => n73, B1 => A(2), B2 => n70, ZN =>
                           n24);
   U86 : AOI22_X1 port map( A1 => D(2), A2 => n79, B1 => C(2), B2 => n76, ZN =>
                           n25);
   U87 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => Z(26));
   U88 : AOI22_X1 port map( A1 => B(26), A2 => n73, B1 => A(26), B2 => n70, ZN 
                           => n32);
   U89 : AOI22_X1 port map( A1 => D(26), A2 => n79, B1 => C(26), B2 => n76, ZN 
                           => n33);
   U90 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => Z(23));
   U91 : AOI22_X1 port map( A1 => B(23), A2 => n73, B1 => A(23), B2 => n70, ZN 
                           => n38);
   U92 : AOI22_X1 port map( A1 => D(23), A2 => n79, B1 => C(23), B2 => n76, ZN 
                           => n39);
   U93 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => Z(16));
   U94 : AOI22_X1 port map( A1 => B(16), A2 => n72, B1 => A(16), B2 => n1, ZN 
                           => n54);
   U95 : AOI22_X1 port map( A1 => D(16), A2 => n78, B1 => C(16), B2 => n75, ZN 
                           => n55);
   U96 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => Z(12));
   U97 : AOI22_X1 port map( A1 => B(12), A2 => n72, B1 => A(12), B2 => n1, ZN 
                           => n62);
   U98 : AOI22_X1 port map( A1 => D(12), A2 => n78, B1 => C(12), B2 => n75, ZN 
                           => n63);
   U99 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Z(9));
   U100 : AOI22_X1 port map( A1 => B(9), A2 => n74, B1 => A(9), B2 => n71, ZN 
                           => n2);
   U101 : AOI22_X1 port map( A1 => D(9), A2 => n80, B1 => C(9), B2 => n77, ZN 
                           => n3);
   U102 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => Z(5));
   U103 : AOI22_X1 port map( A1 => B(5), A2 => n74, B1 => A(5), B2 => n71, ZN 
                           => n14);
   U104 : AOI22_X1 port map( A1 => D(5), A2 => n80, B1 => C(5), B2 => n77, ZN 
                           => n15);
   U105 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => Z(30));
   U106 : AOI22_X1 port map( A1 => B(30), A2 => n73, B1 => A(30), B2 => n70, ZN
                           => n22);
   U107 : AOI22_X1 port map( A1 => D(30), A2 => n79, B1 => C(30), B2 => n76, ZN
                           => n23);
   U108 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => Z(27));
   U109 : AOI22_X1 port map( A1 => B(27), A2 => n73, B1 => A(27), B2 => n70, ZN
                           => n30);
   U110 : AOI22_X1 port map( A1 => D(27), A2 => n79, B1 => C(27), B2 => n76, ZN
                           => n31);
   U111 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => Z(1));
   U112 : AOI22_X1 port map( A1 => B(1), A2 => n72, B1 => A(1), B2 => n1, ZN =>
                           n46);
   U113 : AOI22_X1 port map( A1 => D(1), A2 => n78, B1 => C(1), B2 => n75, ZN 
                           => n47);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity FWD_Unit is

   port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB : in 
         std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;  
         FWDA, FWDB : out std_logic_vector (1 downto 0));

end FWD_Unit;

architecture SYN_bhv of FWD_Unit is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42 : std_logic;

begin
   
   U3 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => FWDB(1));
   U4 : AOI21_X1 port map( B1 => n3, B2 => n4, A => n5, ZN => n1);
   U5 : INV_X1 port map( A => n6, ZN => n3);
   U6 : NOR2_X1 port map( A1 => n2, A2 => n7, ZN => FWDB(0));
   U7 : MUX2_X1 port map( A => n6, B => n8, S => n5, Z => n7);
   U8 : AND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => n5);
   U9 : NOR2_X1 port map( A1 => n13, A2 => n14, ZN => n12);
   U10 : XOR2_X1 port map( A => ADD_WR_MEM(4), B => ADD_RS2(4), Z => n14);
   U11 : XOR2_X1 port map( A => ADD_WR_MEM(3), B => ADD_RS2(3), Z => n13);
   U12 : XNOR2_X1 port map( A => ADD_RS2(1), B => ADD_WR_MEM(1), ZN => n11);
   U13 : XNOR2_X1 port map( A => ADD_RS2(2), B => ADD_WR_MEM(2), ZN => n10);
   U14 : XNOR2_X1 port map( A => ADD_RS2(0), B => ADD_WR_MEM(0), ZN => n9);
   U15 : NAND4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           n6);
   U16 : NOR2_X1 port map( A1 => n19, A2 => n20, ZN => n18);
   U17 : XOR2_X1 port map( A => ADD_WR_WB(3), B => ADD_RS2(3), Z => n20);
   U18 : XOR2_X1 port map( A => ADD_WR_WB(2), B => ADD_RS2(2), Z => n19);
   U19 : XNOR2_X1 port map( A => ADD_RS2(4), B => ADD_WR_WB(4), ZN => n17);
   U20 : XNOR2_X1 port map( A => ADD_RS2(1), B => ADD_WR_WB(1), ZN => n16);
   U21 : XNOR2_X1 port map( A => ADD_RS2(0), B => ADD_WR_WB(0), ZN => n15);
   U22 : NOR2_X1 port map( A1 => n21, A2 => n2, ZN => FWDA(1));
   U23 : AOI21_X1 port map( B1 => n22, B2 => n4, A => n23, ZN => n21);
   U24 : OAI21_X1 port map( B1 => n24, B2 => n25, A => RF_WE_WB, ZN => n4);
   U25 : OR2_X1 port map( A1 => ADD_WR_WB(0), A2 => ADD_WR_WB(1), ZN => n25);
   U26 : OR3_X1 port map( A1 => ADD_WR_WB(3), A2 => ADD_WR_WB(4), A3 => 
                           ADD_WR_WB(2), ZN => n24);
   U27 : INV_X1 port map( A => n26, ZN => n22);
   U28 : NOR2_X1 port map( A1 => n2, A2 => n27, ZN => FWDA(0));
   U29 : MUX2_X1 port map( A => n26, B => n8, S => n23, Z => n27);
   U30 : AND4_X1 port map( A1 => n28, A2 => n29, A3 => n30, A4 => n31, ZN => 
                           n23);
   U31 : NOR2_X1 port map( A1 => n32, A2 => n33, ZN => n31);
   U32 : XOR2_X1 port map( A => ADD_WR_MEM(4), B => ADD_RS1(4), Z => n33);
   U33 : XOR2_X1 port map( A => ADD_WR_MEM(3), B => ADD_RS1(3), Z => n32);
   U34 : XNOR2_X1 port map( A => ADD_RS1(1), B => ADD_WR_MEM(1), ZN => n30);
   U35 : XNOR2_X1 port map( A => ADD_RS1(2), B => ADD_WR_MEM(2), ZN => n29);
   U36 : XNOR2_X1 port map( A => ADD_RS1(0), B => ADD_WR_MEM(0), ZN => n28);
   U37 : INV_X1 port map( A => n34, ZN => n8);
   U38 : OAI21_X1 port map( B1 => n35, B2 => n36, A => RF_WE_MEM, ZN => n34);
   U39 : OR2_X1 port map( A1 => ADD_WR_MEM(0), A2 => ADD_WR_MEM(1), ZN => n36);
   U40 : OR3_X1 port map( A1 => ADD_WR_MEM(3), A2 => ADD_WR_MEM(4), A3 => 
                           ADD_WR_MEM(2), ZN => n35);
   U41 : NAND4_X1 port map( A1 => n37, A2 => n38, A3 => n39, A4 => n40, ZN => 
                           n26);
   U42 : NOR2_X1 port map( A1 => n41, A2 => n42, ZN => n40);
   U43 : XOR2_X1 port map( A => ADD_WR_WB(3), B => ADD_RS1(3), Z => n42);
   U44 : XOR2_X1 port map( A => ADD_WR_WB(2), B => ADD_RS1(2), Z => n41);
   U45 : XNOR2_X1 port map( A => ADD_RS1(4), B => ADD_WR_WB(4), ZN => n39);
   U46 : XNOR2_X1 port map( A => ADD_RS1(1), B => ADD_WR_WB(1), ZN => n38);
   U47 : XNOR2_X1 port map( A => ADD_RS1(0), B => ADD_WR_WB(0), ZN => n37);
   U48 : INV_X1 port map( A => RST, ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N2 is

   port( DIN : in std_logic_vector (1 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (1 downto 0));

end regn_N2;

architecture SYN_bhv of regn_N2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   DOUT_reg_1_inst : DFFR_X1 port map( D => n6, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n4);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n5, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n3);
   U2 : OAI21_X1 port map( B1 => n3, B2 => EN, A => n1, ZN => n5);
   U3 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n1);
   U4 : OAI21_X1 port map( B1 => n4, B2 => EN, A => n2, ZN => n6);
   U5 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Branch_Cond_Unit_NBIT32 is

   port( RST : in std_logic;  A : in std_logic_vector (31 downto 0);  ALU_OPC :
         in std_logic_vector (0 to 4);  JUMP_TYPE : in std_logic_vector (1 
         downto 0);  PC_SEL : out std_logic_vector (1 downto 0);  ZERO : out 
         std_logic);

end Branch_Cond_Unit_NBIT32;

architecture SYN_bhv of Branch_Cond_Unit_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n1, n2 : std_logic;

begin
   
   U24 : NAND3_X1 port map( A1 => ALU_OPC(2), A2 => n7, A3 => ALU_OPC(1), ZN =>
                           n9);
   U25 : NAND3_X1 port map( A1 => ALU_OPC(1), A2 => ALU_OPC(2), A3 => n20, ZN 
                           => n7);
   U3 : NOR4_X1 port map( A1 => A(23), A2 => A(22), A3 => A(21), A4 => A(20), 
                           ZN => n15);
   U4 : NOR4_X1 port map( A1 => A(9), A2 => A(8), A3 => A(7), A4 => A(6), ZN =>
                           n19);
   U5 : NOR4_X1 port map( A1 => A(1), A2 => A(19), A3 => A(18), A4 => A(17), ZN
                           => n14);
   U6 : NOR4_X1 port map( A1 => A(5), A2 => A(4), A3 => A(3), A4 => A(31), ZN 
                           => n18);
   U7 : NOR4_X1 port map( A1 => A(16), A2 => A(15), A3 => A(14), A4 => A(13), 
                           ZN => n13);
   U8 : NOR4_X1 port map( A1 => A(30), A2 => A(2), A3 => A(29), A4 => A(28), ZN
                           => n17);
   U9 : NOR4_X1 port map( A1 => A(12), A2 => A(11), A3 => A(10), A4 => A(0), ZN
                           => n12);
   U10 : NOR2_X1 port map( A1 => n10, A2 => n11, ZN => n8);
   U11 : NAND4_X1 port map( A1 => n16, A2 => n17, A3 => n18, A4 => n19, ZN => 
                           n10);
   U12 : NAND4_X1 port map( A1 => n12, A2 => n13, A3 => n14, A4 => n15, ZN => 
                           n11);
   U13 : NOR4_X1 port map( A1 => A(27), A2 => A(26), A3 => A(25), A4 => A(24), 
                           ZN => n16);
   U14 : NOR3_X1 port map( A1 => ALU_OPC(4), A2 => ALU_OPC(0), A3 => ALU_OPC(3)
                           , ZN => n20);
   U15 : OAI211_X1 port map( C1 => n5, C2 => n6, A => JUMP_TYPE(0), B => RST, 
                           ZN => n4);
   U16 : NOR2_X1 port map( A1 => n7, A2 => n1, ZN => n6);
   U17 : NOR4_X1 port map( A1 => n9, A2 => n8, A3 => ALU_OPC(0), A4 => 
                           ALU_OPC(3), ZN => n5);
   U18 : INV_X1 port map( A => n8, ZN => n1);
   U19 : NAND2_X1 port map( A1 => JUMP_TYPE(1), A2 => RST, ZN => n3);
   U20 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => ZERO);
   U21 : OAI22_X1 port map( A1 => JUMP_TYPE(0), A2 => n3, B1 => JUMP_TYPE(1), 
                           B2 => n4, ZN => PC_SEL(0));
   U22 : NOR2_X1 port map( A1 => n2, A2 => n3, ZN => PC_SEL(1));
   U23 : INV_X1 port map( A => JUMP_TYPE(0), ZN => n2);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity register_file_NBIT_ADD5_NBIT_DATA32 is

   port( CLK, RST, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RS1, 
         ADD_RS2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_NBIT_ADD5_NBIT_DATA32;

architecture SYN_bhv of register_file_NBIT_ADD5_NBIT_DATA32 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
      n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
      n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n517, n518, n519, 
      n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n613, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n644, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, 
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n864, n865, n866, n867, n868, n933, n934, n935, 
      n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, 
      n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, 
      n960, n961, n962, n963, n964, n2506, n2507, n2508, n2509, n2510, n2511, 
      n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, 
      n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, 
      n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, 
      n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, 
      n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, 
      n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, 
      n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, 
      n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, 
      n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, 
      n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, 
      n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, 
      n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, 
      n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, 
      n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, 
      n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, 
      n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, 
      n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, 
      n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, 
      n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, 
      n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, 
      n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, 
      n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, 
      n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, 
      n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, 
      n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, 
      n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, 
      n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, 
      n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, 
      n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, 
      n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, 
      n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, 
      n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, 
      n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, 
      n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, 
      n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, 
      n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, 
      n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, 
      n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, 
      n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, 
      n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, 
      n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, 
      n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, 
      n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, 
      n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, 
      n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, 
      n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, 
      n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, 
      n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, 
      n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, 
      n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, 
      n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, 
      n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, 
      n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, 
      n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, 
      n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, 
      n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, 
      n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, 
      n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, 
      n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, 
      n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, 
      n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, 
      n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, 
      n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, 
      n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, 
      n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, 
      n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, 
      n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, 
      n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, 
      n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, 
      n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, 
      n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, 
      n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, 
      n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, 
      n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, 
      n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, 
      n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, 
      n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, 
      n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, 
      n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, 
      n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, 
      n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, 
      n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, 
      n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, 
      n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, 
      n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, 
      n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, 
      n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, 
      n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, 
      n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, 
      n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, 
      n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, 
      n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, 
      n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, 
      n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, 
      n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, 
      n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, 
      n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, 
      n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, 
      n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, 
      n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, 
      n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, 
      n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, 
      n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, 
      n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, 
      n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n293, n294, n295, n296, n297, n298, n299, 
      n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, 
      n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, 
      n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, 
      n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
      n348, n349, n350, n351, n352, n353, n354, n355, n356, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, 
      n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
      n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, 
      n508, n509, n510, n511, n512, n513, n514, n515, n516, n549, n550, n551, 
      n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, 
      n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, 
      n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, 
      n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
      n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, 
      n612, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, 
      n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, 
      n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
      n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
      n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
      n836, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n965, n966, n967, n968, n969, n970, n971, 
      n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, 
      n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, 
      n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, 
      n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, 
      n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, 
      n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, 
      n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
      n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, 
      n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, 
      n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
      n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, 
      n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, 
      n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, 
      n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, 
      n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, 
      n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, 
      n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, 
      n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, 
      n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
      n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, 
      n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
      n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, 
      n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, 
      n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, 
      n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, 
      n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, 
      n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, 
      n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, 
      n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, 
      n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, 
      n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
      n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, 
      n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, 
      n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, 
      n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, 
      n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, 
      n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, 
      n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
      n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, 
      n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, 
      n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
      n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, 
      n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, 
      n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
      n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, 
      n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, 
      n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
      n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, 
      n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n3562, 
      n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, 
      n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, 
      n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, 
      n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, 
      n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, 
      n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, 
      n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, 
      n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, 
      n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, 
      n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, 
      n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, 
      n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, 
      n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, 
      n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, 
      n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, 
      n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, 
      n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, 
      n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, 
      n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, 
      n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, 
      n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, 
      n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, 
      n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, 
      n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, 
      n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, 
      n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, 
      n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, 
      n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, 
      n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, 
      n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, 
      n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, 
      n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, 
      n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, 
      n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, 
      n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, 
      n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, 
      n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, 
      n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, 
      n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, 
      n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, 
      n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, 
      n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, 
      n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, 
      n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, 
      n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, 
      n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, 
      n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, 
      n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, 
      n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, 
      n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, 
      n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, 
      n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, 
      n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, 
      n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, 
      n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, 
      n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, 
      n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, 
      n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, 
      n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, 
      n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, 
      n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, 
      n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, 
      n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, 
      n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, 
      n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, 
      n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, 
      n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, 
      n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, 
      n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, 
      n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, 
      n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, 
      n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, 
      n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, 
      n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, 
      n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, 
      n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, 
      n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, 
      n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, 
      n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, 
      n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, 
      n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, 
      n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, 
      n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, 
      n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, 
      n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, 
      n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, 
      n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, 
      n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, 
      n4443, n4444, n4445, n4446, n_1198, n_1199, n_1200, n_1201, n_1202, 
      n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, 
      n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, 
      n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, 
      n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, 
      n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, 
      n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, 
      n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, 
      n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, 
      n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, 
      n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, 
      n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, 
      n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, 
      n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, 
      n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, 
      n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, 
      n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, 
      n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, 
      n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, 
      n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, 
      n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, 
      n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, 
      n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, 
      n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, 
      n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, 
      n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, 
      n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, 
      n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, 
      n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, 
      n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, 
      n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, 
      n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, 
      n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, 
      n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, 
      n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, 
      n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, 
      n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, 
      n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, 
      n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, 
      n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, 
      n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, 
      n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, 
      n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, 
      n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, 
      n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, 
      n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, 
      n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, 
      n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, 
      n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, 
      n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, 
      n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, 
      n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, 
      n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, 
      n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, 
      n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, 
      n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, 
      n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, 
      n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, 
      n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, 
      n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, 
      n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, 
      n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, 
      n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, 
      n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, 
      n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, 
      n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, 
      n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, 
      n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, 
      n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, 
      n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, 
      n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, 
      n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, 
      n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, 
      n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, 
      n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, 
      n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, 
      n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, 
      n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, 
      n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, 
      n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, 
      n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, 
      n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, 
      n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, 
      n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, 
      n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, 
      n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965 : std_logic;

begin
   
   REGISTERS_reg_8_23_inst : DFFR_X1 port map( D => n3329, CK => CLK, RN => 
                           n665, Q => n_1198, QN => n237);
   REGISTERS_reg_8_22_inst : DFFR_X1 port map( D => n3328, CK => CLK, RN => 
                           n665, Q => n_1199, QN => n238);
   REGISTERS_reg_8_21_inst : DFFR_X1 port map( D => n3327, CK => CLK, RN => 
                           n665, Q => n_1200, QN => n239);
   REGISTERS_reg_8_20_inst : DFFR_X1 port map( D => n3326, CK => CLK, RN => 
                           n665, Q => n_1201, QN => n240);
   REGISTERS_reg_8_19_inst : DFFR_X1 port map( D => n3325, CK => CLK, RN => 
                           n665, Q => n_1202, QN => n241);
   REGISTERS_reg_8_18_inst : DFFR_X1 port map( D => n3324, CK => CLK, RN => 
                           n664, Q => n_1203, QN => n242);
   REGISTERS_reg_8_17_inst : DFFR_X1 port map( D => n3323, CK => CLK, RN => 
                           n664, Q => n_1204, QN => n243);
   REGISTERS_reg_8_16_inst : DFFR_X1 port map( D => n3322, CK => CLK, RN => 
                           n664, Q => n_1205, QN => n244);
   REGISTERS_reg_8_15_inst : DFFR_X1 port map( D => n3321, CK => CLK, RN => 
                           n664, Q => n_1206, QN => n245);
   REGISTERS_reg_8_14_inst : DFFR_X1 port map( D => n3320, CK => CLK, RN => 
                           n664, Q => n_1207, QN => n246);
   REGISTERS_reg_8_13_inst : DFFR_X1 port map( D => n3319, CK => CLK, RN => 
                           n664, Q => n_1208, QN => n247);
   REGISTERS_reg_8_12_inst : DFFR_X1 port map( D => n3318, CK => CLK, RN => 
                           n664, Q => n_1209, QN => n248);
   REGISTERS_reg_8_11_inst : DFFR_X1 port map( D => n3317, CK => CLK, RN => 
                           n664, Q => n_1210, QN => n249);
   REGISTERS_reg_8_10_inst : DFFR_X1 port map( D => n3316, CK => CLK, RN => 
                           n664, Q => n_1211, QN => n250);
   REGISTERS_reg_8_9_inst : DFFR_X1 port map( D => n3315, CK => CLK, RN => n664
                           , Q => n_1212, QN => n251);
   REGISTERS_reg_8_8_inst : DFFR_X1 port map( D => n3314, CK => CLK, RN => n664
                           , Q => n_1213, QN => n252);
   REGISTERS_reg_8_7_inst : DFFR_X1 port map( D => n3313, CK => CLK, RN => n669
                           , Q => n_1214, QN => n253);
   REGISTERS_reg_8_6_inst : DFFR_X1 port map( D => n3312, CK => CLK, RN => n611
                           , Q => n_1215, QN => n254);
   REGISTERS_reg_8_5_inst : DFFR_X1 port map( D => n3311, CK => CLK, RN => n611
                           , Q => n_1216, QN => n255);
   REGISTERS_reg_8_4_inst : DFFR_X1 port map( D => n3310, CK => CLK, RN => n611
                           , Q => n_1217, QN => n256);
   REGISTERS_reg_8_3_inst : DFFR_X1 port map( D => n3309, CK => CLK, RN => n611
                           , Q => n_1218, QN => n257);
   REGISTERS_reg_8_2_inst : DFFR_X1 port map( D => n3308, CK => CLK, RN => n611
                           , Q => n_1219, QN => n258);
   REGISTERS_reg_8_1_inst : DFFR_X1 port map( D => n3307, CK => CLK, RN => n610
                           , Q => n_1220, QN => n259);
   REGISTERS_reg_8_0_inst : DFFR_X1 port map( D => n3306, CK => CLK, RN => n610
                           , Q => n_1221, QN => n260);
   REGISTERS_reg_9_23_inst : DFFR_X1 port map( D => n3297, CK => CLK, RN => 
                           n610, Q => n_1222, QN => n269);
   REGISTERS_reg_9_22_inst : DFFR_X1 port map( D => n3296, CK => CLK, RN => 
                           n610, Q => n_1223, QN => n270);
   REGISTERS_reg_9_21_inst : DFFR_X1 port map( D => n3295, CK => CLK, RN => 
                           n609, Q => n_1224, QN => n271);
   REGISTERS_reg_9_20_inst : DFFR_X1 port map( D => n3294, CK => CLK, RN => 
                           n609, Q => n_1225, QN => n272);
   REGISTERS_reg_9_19_inst : DFFR_X1 port map( D => n3293, CK => CLK, RN => 
                           n609, Q => n_1226, QN => n273);
   REGISTERS_reg_9_18_inst : DFFR_X1 port map( D => n3292, CK => CLK, RN => 
                           n609, Q => n_1227, QN => n274);
   REGISTERS_reg_9_17_inst : DFFR_X1 port map( D => n3291, CK => CLK, RN => 
                           n609, Q => n_1228, QN => n275);
   REGISTERS_reg_9_16_inst : DFFR_X1 port map( D => n3290, CK => CLK, RN => 
                           n609, Q => n_1229, QN => n276);
   REGISTERS_reg_9_15_inst : DFFR_X1 port map( D => n3289, CK => CLK, RN => 
                           n609, Q => n_1230, QN => n277);
   REGISTERS_reg_9_14_inst : DFFR_X1 port map( D => n3288, CK => CLK, RN => 
                           n609, Q => n_1231, QN => n278);
   REGISTERS_reg_9_13_inst : DFFR_X1 port map( D => n3287, CK => CLK, RN => 
                           n609, Q => n_1232, QN => n279);
   REGISTERS_reg_9_12_inst : DFFR_X1 port map( D => n3286, CK => CLK, RN => 
                           n609, Q => n_1233, QN => n280);
   REGISTERS_reg_9_11_inst : DFFR_X1 port map( D => n3285, CK => CLK, RN => 
                           n609, Q => n_1234, QN => n281);
   REGISTERS_reg_9_10_inst : DFFR_X1 port map( D => n3284, CK => CLK, RN => 
                           n609, Q => n_1235, QN => n282);
   REGISTERS_reg_9_9_inst : DFFR_X1 port map( D => n3283, CK => CLK, RN => n608
                           , Q => n_1236, QN => n283);
   REGISTERS_reg_9_8_inst : DFFR_X1 port map( D => n3282, CK => CLK, RN => n608
                           , Q => n_1237, QN => n284);
   REGISTERS_reg_9_7_inst : DFFR_X1 port map( D => n3281, CK => CLK, RN => n608
                           , Q => n_1238, QN => n285);
   REGISTERS_reg_9_6_inst : DFFR_X1 port map( D => n3280, CK => CLK, RN => n608
                           , Q => n_1239, QN => n286);
   REGISTERS_reg_9_5_inst : DFFR_X1 port map( D => n3279, CK => CLK, RN => n608
                           , Q => n_1240, QN => n287);
   REGISTERS_reg_9_4_inst : DFFR_X1 port map( D => n3278, CK => CLK, RN => n608
                           , Q => n_1241, QN => n288);
   REGISTERS_reg_9_3_inst : DFFR_X1 port map( D => n3277, CK => CLK, RN => n608
                           , Q => n_1242, QN => n289);
   REGISTERS_reg_9_2_inst : DFFR_X1 port map( D => n3276, CK => CLK, RN => n608
                           , Q => n_1243, QN => n290);
   REGISTERS_reg_9_1_inst : DFFR_X1 port map( D => n3275, CK => CLK, RN => n608
                           , Q => n_1244, QN => n291);
   REGISTERS_reg_9_0_inst : DFFR_X1 port map( D => n3274, CK => CLK, RN => n608
                           , Q => n_1245, QN => n292);
   REGISTERS_reg_12_14_inst : DFFR_X1 port map( D => n3192, CK => CLK, RN => 
                           n601, Q => n_1246, QN => n374);
   REGISTERS_reg_12_13_inst : DFFR_X1 port map( D => n3191, CK => CLK, RN => 
                           n601, Q => n_1247, QN => n375);
   REGISTERS_reg_12_12_inst : DFFR_X1 port map( D => n3190, CK => CLK, RN => 
                           n601, Q => n_1248, QN => n376);
   REGISTERS_reg_12_11_inst : DFFR_X1 port map( D => n3189, CK => CLK, RN => 
                           n606, Q => n_1249, QN => n377);
   REGISTERS_reg_12_10_inst : DFFR_X1 port map( D => n3188, CK => CLK, RN => 
                           n653, Q => n_1250, QN => n378);
   REGISTERS_reg_12_9_inst : DFFR_X1 port map( D => n3187, CK => CLK, RN => 
                           n653, Q => n_1251, QN => n379);
   REGISTERS_reg_12_8_inst : DFFR_X1 port map( D => n3186, CK => CLK, RN => 
                           n653, Q => n_1252, QN => n380);
   REGISTERS_reg_12_7_inst : DFFR_X1 port map( D => n3185, CK => CLK, RN => 
                           n653, Q => n_1253, QN => n381);
   REGISTERS_reg_12_6_inst : DFFR_X1 port map( D => n3184, CK => CLK, RN => 
                           n653, Q => n_1254, QN => n382);
   REGISTERS_reg_12_5_inst : DFFR_X1 port map( D => n3183, CK => CLK, RN => 
                           n653, Q => n_1255, QN => n383);
   REGISTERS_reg_12_4_inst : DFFR_X1 port map( D => n3182, CK => CLK, RN => 
                           n653, Q => n_1256, QN => n384);
   REGISTERS_reg_12_3_inst : DFFR_X1 port map( D => n3181, CK => CLK, RN => 
                           n653, Q => n_1257, QN => n385);
   REGISTERS_reg_12_2_inst : DFFR_X1 port map( D => n3180, CK => CLK, RN => 
                           n652, Q => n_1258, QN => n386);
   REGISTERS_reg_12_1_inst : DFFR_X1 port map( D => n3179, CK => CLK, RN => 
                           n652, Q => n_1259, QN => n387);
   REGISTERS_reg_12_0_inst : DFFR_X1 port map( D => n3178, CK => CLK, RN => 
                           n652, Q => n_1260, QN => n388);
   REGISTERS_reg_17_23_inst : DFFR_X1 port map( D => n3041, CK => CLK, RN => 
                           n703, Q => n_1261, QN => n525);
   REGISTERS_reg_17_22_inst : DFFR_X1 port map( D => n3040, CK => CLK, RN => 
                           n703, Q => n_1262, QN => n526);
   REGISTERS_reg_17_21_inst : DFFR_X1 port map( D => n3039, CK => CLK, RN => 
                           n703, Q => n_1263, QN => n527);
   REGISTERS_reg_17_20_inst : DFFR_X1 port map( D => n3038, CK => CLK, RN => 
                           n703, Q => n_1264, QN => n528);
   REGISTERS_reg_17_19_inst : DFFR_X1 port map( D => n3037, CK => CLK, RN => 
                           n703, Q => n_1265, QN => n529);
   REGISTERS_reg_17_18_inst : DFFR_X1 port map( D => n3036, CK => CLK, RN => 
                           n703, Q => n_1266, QN => n530);
   REGISTERS_reg_17_17_inst : DFFR_X1 port map( D => n3035, CK => CLK, RN => 
                           n702, Q => n_1267, QN => n531);
   REGISTERS_reg_17_16_inst : DFFR_X1 port map( D => n3034, CK => CLK, RN => 
                           n702, Q => n_1268, QN => n532);
   REGISTERS_reg_17_15_inst : DFFR_X1 port map( D => n3033, CK => CLK, RN => 
                           n702, Q => n_1269, QN => n533);
   REGISTERS_reg_17_14_inst : DFFR_X1 port map( D => n3032, CK => CLK, RN => 
                           n702, Q => n_1270, QN => n534);
   REGISTERS_reg_17_13_inst : DFFR_X1 port map( D => n3031, CK => CLK, RN => 
                           n702, Q => n_1271, QN => n535);
   REGISTERS_reg_17_12_inst : DFFR_X1 port map( D => n3030, CK => CLK, RN => 
                           n702, Q => n_1272, QN => n536);
   REGISTERS_reg_17_11_inst : DFFR_X1 port map( D => n3029, CK => CLK, RN => 
                           n702, Q => n_1273, QN => n537);
   REGISTERS_reg_17_10_inst : DFFR_X1 port map( D => n3028, CK => CLK, RN => 
                           n702, Q => n_1274, QN => n538);
   REGISTERS_reg_17_9_inst : DFFR_X1 port map( D => n3027, CK => CLK, RN => 
                           n702, Q => n_1275, QN => n539);
   REGISTERS_reg_17_8_inst : DFFR_X1 port map( D => n3026, CK => CLK, RN => 
                           n702, Q => n_1276, QN => n540);
   REGISTERS_reg_17_7_inst : DFFR_X1 port map( D => n3025, CK => CLK, RN => 
                           n702, Q => n_1277, QN => n541);
   REGISTERS_reg_17_6_inst : DFFR_X1 port map( D => n3024, CK => CLK, RN => 
                           n702, Q => n_1278, QN => n542);
   REGISTERS_reg_17_5_inst : DFFR_X1 port map( D => n3023, CK => CLK, RN => 
                           n701, Q => n_1279, QN => n543);
   REGISTERS_reg_17_4_inst : DFFR_X1 port map( D => n3022, CK => CLK, RN => 
                           n701, Q => n_1280, QN => n544);
   REGISTERS_reg_17_3_inst : DFFR_X1 port map( D => n3021, CK => CLK, RN => 
                           n701, Q => n_1281, QN => n545);
   REGISTERS_reg_17_2_inst : DFFR_X1 port map( D => n3020, CK => CLK, RN => 
                           n701, Q => n_1282, QN => n546);
   REGISTERS_reg_17_1_inst : DFFR_X1 port map( D => n3019, CK => CLK, RN => 
                           n701, Q => n_1283, QN => n547);
   REGISTERS_reg_17_0_inst : DFFR_X1 port map( D => n3018, CK => CLK, RN => 
                           n701, Q => n_1284, QN => n548);
   REGISTERS_reg_20_23_inst : DFFR_X1 port map( D => n2945, CK => CLK, RN => 
                           n695, Q => n_1285, QN => n621);
   REGISTERS_reg_20_22_inst : DFFR_X1 port map( D => n2944, CK => CLK, RN => 
                           n695, Q => n_1286, QN => n622);
   REGISTERS_reg_20_21_inst : DFFR_X1 port map( D => n2943, CK => CLK, RN => 
                           n695, Q => n_1287, QN => n623);
   REGISTERS_reg_20_20_inst : DFFR_X1 port map( D => n2942, CK => CLK, RN => 
                           n695, Q => n_1288, QN => n624);
   REGISTERS_reg_20_19_inst : DFFR_X1 port map( D => n2941, CK => CLK, RN => 
                           n700, Q => n_1289, QN => n625);
   REGISTERS_reg_20_18_inst : DFFR_X1 port map( D => n2940, CK => CLK, RN => 
                           n715, Q => n_1290, QN => n626);
   REGISTERS_reg_20_17_inst : DFFR_X1 port map( D => n2939, CK => CLK, RN => 
                           n715, Q => n_1291, QN => n627);
   REGISTERS_reg_20_16_inst : DFFR_X1 port map( D => n2938, CK => CLK, RN => 
                           n715, Q => n_1292, QN => n628);
   REGISTERS_reg_20_15_inst : DFFR_X1 port map( D => n2937, CK => CLK, RN => 
                           n715, Q => n_1293, QN => n629);
   REGISTERS_reg_20_14_inst : DFFR_X1 port map( D => n2936, CK => CLK, RN => 
                           n715, Q => n_1294, QN => n630);
   REGISTERS_reg_20_13_inst : DFFR_X1 port map( D => n2935, CK => CLK, RN => 
                           n715, Q => n_1295, QN => n631);
   REGISTERS_reg_20_12_inst : DFFR_X1 port map( D => n2934, CK => CLK, RN => 
                           n715, Q => n_1296, QN => n632);
   REGISTERS_reg_20_11_inst : DFFR_X1 port map( D => n2933, CK => CLK, RN => 
                           n715, Q => n_1297, QN => n633);
   REGISTERS_reg_20_10_inst : DFFR_X1 port map( D => n2932, CK => CLK, RN => 
                           n714, Q => n_1298, QN => n634);
   REGISTERS_reg_20_9_inst : DFFR_X1 port map( D => n2931, CK => CLK, RN => 
                           n714, Q => n_1299, QN => n635);
   REGISTERS_reg_20_8_inst : DFFR_X1 port map( D => n2930, CK => CLK, RN => 
                           n714, Q => n_1300, QN => n636);
   REGISTERS_reg_20_7_inst : DFFR_X1 port map( D => n2929, CK => CLK, RN => 
                           n714, Q => n_1301, QN => n637);
   REGISTERS_reg_20_6_inst : DFFR_X1 port map( D => n2928, CK => CLK, RN => 
                           n714, Q => n_1302, QN => n638);
   REGISTERS_reg_20_5_inst : DFFR_X1 port map( D => n2927, CK => CLK, RN => 
                           n714, Q => n_1303, QN => n639);
   REGISTERS_reg_20_4_inst : DFFR_X1 port map( D => n2926, CK => CLK, RN => 
                           n714, Q => n_1304, QN => n640);
   REGISTERS_reg_20_3_inst : DFFR_X1 port map( D => n2925, CK => CLK, RN => 
                           n714, Q => n_1305, QN => n641);
   REGISTERS_reg_20_2_inst : DFFR_X1 port map( D => n2924, CK => CLK, RN => 
                           n714, Q => n_1306, QN => n642);
   REGISTERS_reg_20_1_inst : DFFR_X1 port map( D => n2923, CK => CLK, RN => 
                           n714, Q => n_1307, QN => n643);
   REGISTERS_reg_20_0_inst : DFFR_X1 port map( D => n2922, CK => CLK, RN => 
                           n714, Q => n_1308, QN => n644);
   REGISTERS_reg_24_3_inst : DFFR_X1 port map( D => n2797, CK => CLK, RN => 
                           n683, Q => n4034, QN => n_1309);
   REGISTERS_reg_24_2_inst : DFFR_X1 port map( D => n2796, CK => CLK, RN => 
                           n682, Q => n4033, QN => n_1310);
   REGISTERS_reg_24_1_inst : DFFR_X1 port map( D => n2795, CK => CLK, RN => 
                           n682, Q => n4032, QN => n_1311);
   REGISTERS_reg_24_0_inst : DFFR_X1 port map( D => n2794, CK => CLK, RN => 
                           n682, Q => n4031, QN => n_1312);
   REGISTERS_reg_27_23_inst : DFFR_X1 port map( D => n2721, CK => CLK, RN => 
                           n676, Q => n_1313, QN => n845);
   REGISTERS_reg_27_22_inst : DFFR_X1 port map( D => n2720, CK => CLK, RN => 
                           n676, Q => n_1314, QN => n846);
   REGISTERS_reg_27_21_inst : DFFR_X1 port map( D => n2719, CK => CLK, RN => 
                           n676, Q => n_1315, QN => n847);
   REGISTERS_reg_27_20_inst : DFFR_X1 port map( D => n2718, CK => CLK, RN => 
                           n676, Q => n_1316, QN => n848);
   REGISTERS_reg_27_19_inst : DFFR_X1 port map( D => n2717, CK => CLK, RN => 
                           n676, Q => n_1317, QN => n849);
   REGISTERS_reg_27_18_inst : DFFR_X1 port map( D => n2716, CK => CLK, RN => 
                           n676, Q => n_1318, QN => n850);
   REGISTERS_reg_27_17_inst : DFFR_X1 port map( D => n2715, CK => CLK, RN => 
                           n676, Q => n_1319, QN => n851);
   REGISTERS_reg_27_16_inst : DFFR_X1 port map( D => n2714, CK => CLK, RN => 
                           n676, Q => n_1320, QN => n852);
   REGISTERS_reg_27_15_inst : DFFR_X1 port map( D => n2713, CK => CLK, RN => 
                           n675, Q => n_1321, QN => n853);
   REGISTERS_reg_27_14_inst : DFFR_X1 port map( D => n2712, CK => CLK, RN => 
                           n675, Q => n_1322, QN => n854);
   REGISTERS_reg_27_13_inst : DFFR_X1 port map( D => n2711, CK => CLK, RN => 
                           n675, Q => n_1323, QN => n855);
   REGISTERS_reg_27_12_inst : DFFR_X1 port map( D => n2710, CK => CLK, RN => 
                           n675, Q => n_1324, QN => n856);
   REGISTERS_reg_27_11_inst : DFFR_X1 port map( D => n2709, CK => CLK, RN => 
                           n675, Q => n_1325, QN => n857);
   REGISTERS_reg_27_10_inst : DFFR_X1 port map( D => n2708, CK => CLK, RN => 
                           n675, Q => n_1326, QN => n858);
   REGISTERS_reg_27_9_inst : DFFR_X1 port map( D => n2707, CK => CLK, RN => 
                           n675, Q => n_1327, QN => n859);
   REGISTERS_reg_27_8_inst : DFFR_X1 port map( D => n2706, CK => CLK, RN => 
                           n675, Q => n_1328, QN => n860);
   REGISTERS_reg_27_7_inst : DFFR_X1 port map( D => n2705, CK => CLK, RN => 
                           n675, Q => n_1329, QN => n861);
   REGISTERS_reg_27_6_inst : DFFR_X1 port map( D => n2704, CK => CLK, RN => 
                           n675, Q => n_1330, QN => n862);
   REGISTERS_reg_27_5_inst : DFFR_X1 port map( D => n2703, CK => CLK, RN => 
                           n675, Q => n_1331, QN => n863);
   REGISTERS_reg_27_4_inst : DFFR_X1 port map( D => n2702, CK => CLK, RN => 
                           n675, Q => n_1332, QN => n864);
   REGISTERS_reg_27_3_inst : DFFR_X1 port map( D => n2701, CK => CLK, RN => 
                           n674, Q => n_1333, QN => n865);
   REGISTERS_reg_27_2_inst : DFFR_X1 port map( D => n2700, CK => CLK, RN => 
                           n674, Q => n_1334, QN => n866);
   REGISTERS_reg_27_1_inst : DFFR_X1 port map( D => n2699, CK => CLK, RN => 
                           n674, Q => n_1335, QN => n867);
   REGISTERS_reg_27_0_inst : DFFR_X1 port map( D => n2698, CK => CLK, RN => 
                           n674, Q => n_1336, QN => n868);
   REGISTERS_reg_30_23_inst : DFFR_X1 port map( D => n2625, CK => CLK, RN => 
                           n689, Q => n_1337, QN => n941);
   REGISTERS_reg_30_22_inst : DFFR_X1 port map( D => n2624, CK => CLK, RN => 
                           n689, Q => n_1338, QN => n942);
   REGISTERS_reg_30_21_inst : DFFR_X1 port map( D => n2623, CK => CLK, RN => 
                           n689, Q => n_1339, QN => n943);
   REGISTERS_reg_30_20_inst : DFFR_X1 port map( D => n2622, CK => CLK, RN => 
                           n689, Q => n_1340, QN => n944);
   REGISTERS_reg_30_19_inst : DFFR_X1 port map( D => n2621, CK => CLK, RN => 
                           n688, Q => n_1341, QN => n945);
   REGISTERS_reg_30_18_inst : DFFR_X1 port map( D => n2620, CK => CLK, RN => 
                           n688, Q => n_1342, QN => n946);
   REGISTERS_reg_30_17_inst : DFFR_X1 port map( D => n2619, CK => CLK, RN => 
                           n688, Q => n_1343, QN => n947);
   REGISTERS_reg_30_16_inst : DFFR_X1 port map( D => n2618, CK => CLK, RN => 
                           n688, Q => n_1344, QN => n948);
   REGISTERS_reg_30_15_inst : DFFR_X1 port map( D => n2617, CK => CLK, RN => 
                           n688, Q => n_1345, QN => n949);
   REGISTERS_reg_30_14_inst : DFFR_X1 port map( D => n2616, CK => CLK, RN => 
                           n688, Q => n_1346, QN => n950);
   REGISTERS_reg_30_13_inst : DFFR_X1 port map( D => n2615, CK => CLK, RN => 
                           n688, Q => n_1347, QN => n951);
   REGISTERS_reg_30_12_inst : DFFR_X1 port map( D => n2614, CK => CLK, RN => 
                           n688, Q => n_1348, QN => n952);
   REGISTERS_reg_30_11_inst : DFFR_X1 port map( D => n2613, CK => CLK, RN => 
                           n688, Q => n_1349, QN => n953);
   REGISTERS_reg_30_10_inst : DFFR_X1 port map( D => n2612, CK => CLK, RN => 
                           n688, Q => n_1350, QN => n954);
   REGISTERS_reg_30_9_inst : DFFR_X1 port map( D => n2611, CK => CLK, RN => 
                           n688, Q => n_1351, QN => n955);
   REGISTERS_reg_30_8_inst : DFFR_X1 port map( D => n2610, CK => CLK, RN => 
                           n688, Q => n_1352, QN => n956);
   REGISTERS_reg_30_7_inst : DFFR_X1 port map( D => n2609, CK => CLK, RN => 
                           n687, Q => n_1353, QN => n957);
   REGISTERS_reg_30_6_inst : DFFR_X1 port map( D => n2608, CK => CLK, RN => 
                           n687, Q => n_1354, QN => n958);
   REGISTERS_reg_30_5_inst : DFFR_X1 port map( D => n2607, CK => CLK, RN => 
                           n687, Q => n_1355, QN => n959);
   REGISTERS_reg_30_4_inst : DFFR_X1 port map( D => n2606, CK => CLK, RN => 
                           n687, Q => n_1356, QN => n960);
   REGISTERS_reg_30_3_inst : DFFR_X1 port map( D => n2605, CK => CLK, RN => 
                           n687, Q => n_1357, QN => n961);
   REGISTERS_reg_30_2_inst : DFFR_X1 port map( D => n2604, CK => CLK, RN => 
                           n687, Q => n_1358, QN => n962);
   REGISTERS_reg_30_1_inst : DFFR_X1 port map( D => n2603, CK => CLK, RN => 
                           n687, Q => n_1359, QN => n963);
   REGISTERS_reg_30_0_inst : DFFR_X1 port map( D => n2602, CK => CLK, RN => 
                           n687, Q => n_1360, QN => n964);
   REGISTERS_reg_5_31_inst : DFFR_X1 port map( D => n3433, CK => CLK, RN => RST
                           , Q => n803, QN => n_1361);
   REGISTERS_reg_5_30_inst : DFFR_X1 port map( D => n3432, CK => CLK, RN => 
                           n674, Q => n805, QN => n_1362);
   REGISTERS_reg_5_29_inst : DFFR_X1 port map( D => n3431, CK => CLK, RN => 
                           n673, Q => n806, QN => n_1363);
   REGISTERS_reg_5_28_inst : DFFR_X1 port map( D => n3430, CK => CLK, RN => 
                           n673, Q => n807, QN => n_1364);
   REGISTERS_reg_5_27_inst : DFFR_X1 port map( D => n3429, CK => CLK, RN => 
                           n673, Q => n808, QN => n_1365);
   REGISTERS_reg_5_26_inst : DFFR_X1 port map( D => n3428, CK => CLK, RN => 
                           n673, Q => n809, QN => n_1366);
   REGISTERS_reg_5_25_inst : DFFR_X1 port map( D => n3427, CK => CLK, RN => 
                           n673, Q => n810, QN => n_1367);
   REGISTERS_reg_5_24_inst : DFFR_X1 port map( D => n3426, CK => CLK, RN => 
                           n673, Q => n811, QN => n_1368);
   REGISTERS_reg_4_31_inst : DFFR_X1 port map( D => n3465, CK => CLK, RN => 
                           n656, Q => n769, QN => n_1369);
   REGISTERS_reg_4_30_inst : DFFR_X1 port map( D => n3464, CK => CLK, RN => 
                           n656, Q => n771, QN => n_1370);
   REGISTERS_reg_4_29_inst : DFFR_X1 port map( D => n3463, CK => CLK, RN => 
                           n655, Q => n772, QN => n_1371);
   REGISTERS_reg_4_28_inst : DFFR_X1 port map( D => n3462, CK => CLK, RN => 
                           n655, Q => n773, QN => n_1372);
   REGISTERS_reg_4_27_inst : DFFR_X1 port map( D => n3461, CK => CLK, RN => 
                           n655, Q => n774, QN => n_1373);
   REGISTERS_reg_4_26_inst : DFFR_X1 port map( D => n3460, CK => CLK, RN => 
                           n655, Q => n775, QN => n_1374);
   REGISTERS_reg_4_25_inst : DFFR_X1 port map( D => n3459, CK => CLK, RN => 
                           n655, Q => n776, QN => n_1375);
   REGISTERS_reg_4_24_inst : DFFR_X1 port map( D => n3458, CK => CLK, RN => 
                           n655, Q => n777, QN => n_1376);
   REGISTERS_reg_1_31_inst : DFFR_X1 port map( D => n3561, CK => CLK, RN => 
                           n674, Q => n730, QN => n_1377);
   REGISTERS_reg_1_30_inst : DFFR_X1 port map( D => n3560, CK => CLK, RN => 
                           n601, Q => n732, QN => n_1378);
   REGISTERS_reg_1_29_inst : DFFR_X1 port map( D => n3559, CK => CLK, RN => 
                           n664, Q => n733, QN => n_1379);
   REGISTERS_reg_1_28_inst : DFFR_X1 port map( D => n3558, CK => CLK, RN => 
                           n663, Q => n734, QN => n_1380);
   REGISTERS_reg_1_27_inst : DFFR_X1 port map( D => n3557, CK => CLK, RN => 
                           n663, Q => n735, QN => n_1381);
   REGISTERS_reg_1_26_inst : DFFR_X1 port map( D => n3556, CK => CLK, RN => 
                           n663, Q => n736, QN => n_1382);
   REGISTERS_reg_1_25_inst : DFFR_X1 port map( D => n3555, CK => CLK, RN => 
                           n663, Q => n737, QN => n_1383);
   REGISTERS_reg_1_24_inst : DFFR_X1 port map( D => n3554, CK => CLK, RN => 
                           n663, Q => n738, QN => n_1384);
   REGISTERS_reg_21_31_inst : DFFR_X1 port map( D => n2921, CK => CLK, RN => 
                           n714, Q => n1148, QN => n_1385);
   REGISTERS_reg_21_30_inst : DFFR_X1 port map( D => n2920, CK => CLK, RN => 
                           n713, Q => n1150, QN => n_1386);
   REGISTERS_reg_21_29_inst : DFFR_X1 port map( D => n2919, CK => CLK, RN => 
                           n713, Q => n1151, QN => n_1387);
   REGISTERS_reg_21_28_inst : DFFR_X1 port map( D => n2918, CK => CLK, RN => 
                           n713, Q => n1152, QN => n_1388);
   REGISTERS_reg_21_27_inst : DFFR_X1 port map( D => n2917, CK => CLK, RN => 
                           n713, Q => n1153, QN => n_1389);
   REGISTERS_reg_21_26_inst : DFFR_X1 port map( D => n2916, CK => CLK, RN => 
                           n713, Q => n1154, QN => n_1390);
   REGISTERS_reg_21_25_inst : DFFR_X1 port map( D => n2915, CK => CLK, RN => 
                           n713, Q => n1155, QN => n_1391);
   REGISTERS_reg_21_24_inst : DFFR_X1 port map( D => n2914, CK => CLK, RN => 
                           n713, Q => n1156, QN => n_1392);
   REGISTERS_reg_16_31_inst : DFFR_X1 port map( D => n3081, CK => CLK, RN => 
                           n612, Q => n1046, QN => n_1393);
   REGISTERS_reg_16_30_inst : DFFR_X1 port map( D => n3080, CK => CLK, RN => 
                           n612, Q => n1048, QN => n_1394);
   REGISTERS_reg_16_29_inst : DFFR_X1 port map( D => n3079, CK => CLK, RN => 
                           n612, Q => n1049, QN => n_1395);
   REGISTERS_reg_16_28_inst : DFFR_X1 port map( D => n3078, CK => CLK, RN => 
                           n612, Q => n1050, QN => n_1396);
   REGISTERS_reg_16_27_inst : DFFR_X1 port map( D => n3077, CK => CLK, RN => 
                           n612, Q => n1051, QN => n_1397);
   REGISTERS_reg_16_26_inst : DFFR_X1 port map( D => n3076, CK => CLK, RN => 
                           n612, Q => n1052, QN => n_1398);
   REGISTERS_reg_16_25_inst : DFFR_X1 port map( D => n3075, CK => CLK, RN => 
                           n612, Q => n1053, QN => n_1399);
   REGISTERS_reg_16_24_inst : DFFR_X1 port map( D => n3074, CK => CLK, RN => 
                           n612, Q => n1054, QN => n_1400);
   REGISTERS_reg_31_31_inst : DFFR_X1 port map( D => n2601, CK => CLK, RN => 
                           n687, Q => n1289, QN => n_1401);
   REGISTERS_reg_31_30_inst : DFFR_X1 port map( D => n2600, CK => CLK, RN => 
                           n687, Q => n1291, QN => n_1402);
   REGISTERS_reg_31_29_inst : DFFR_X1 port map( D => n2599, CK => CLK, RN => 
                           n687, Q => n1292, QN => n_1403);
   REGISTERS_reg_31_28_inst : DFFR_X1 port map( D => n2598, CK => CLK, RN => 
                           n687, Q => n1293, QN => n_1404);
   REGISTERS_reg_31_27_inst : DFFR_X1 port map( D => n2597, CK => CLK, RN => 
                           n686, Q => n1294, QN => n_1405);
   REGISTERS_reg_31_26_inst : DFFR_X1 port map( D => n2596, CK => CLK, RN => 
                           n686, Q => n1295, QN => n_1406);
   REGISTERS_reg_31_25_inst : DFFR_X1 port map( D => n2595, CK => CLK, RN => 
                           n686, Q => n1296, QN => n_1407);
   REGISTERS_reg_31_24_inst : DFFR_X1 port map( D => n2594, CK => CLK, RN => 
                           n686, Q => n1297, QN => n_1408);
   REGISTERS_reg_26_31_inst : DFFR_X1 port map( D => n2761, CK => CLK, RN => 
                           n680, Q => n1187, QN => n_1409);
   REGISTERS_reg_26_30_inst : DFFR_X1 port map( D => n2760, CK => CLK, RN => 
                           n679, Q => n1189, QN => n_1410);
   REGISTERS_reg_26_29_inst : DFFR_X1 port map( D => n2759, CK => CLK, RN => 
                           n679, Q => n1190, QN => n_1411);
   REGISTERS_reg_26_28_inst : DFFR_X1 port map( D => n2758, CK => CLK, RN => 
                           n679, Q => n1191, QN => n_1412);
   REGISTERS_reg_26_27_inst : DFFR_X1 port map( D => n2757, CK => CLK, RN => 
                           n679, Q => n1192, QN => n_1413);
   REGISTERS_reg_26_26_inst : DFFR_X1 port map( D => n2756, CK => CLK, RN => 
                           n679, Q => n1193, QN => n_1414);
   REGISTERS_reg_26_25_inst : DFFR_X1 port map( D => n2755, CK => CLK, RN => 
                           n679, Q => n1194, QN => n_1415);
   REGISTERS_reg_26_24_inst : DFFR_X1 port map( D => n2754, CK => CLK, RN => 
                           n679, Q => n1195, QN => n_1416);
   REGISTERS_reg_5_23_inst : DFFR_X1 port map( D => n3425, CK => CLK, RN => 
                           n673, Q => n812, QN => n_1417);
   REGISTERS_reg_5_22_inst : DFFR_X1 port map( D => n3424, CK => CLK, RN => 
                           n673, Q => n813, QN => n_1418);
   REGISTERS_reg_5_21_inst : DFFR_X1 port map( D => n3423, CK => CLK, RN => 
                           n673, Q => n814, QN => n_1419);
   REGISTERS_reg_5_20_inst : DFFR_X1 port map( D => n3422, CK => CLK, RN => 
                           n673, Q => n815, QN => n_1420);
   REGISTERS_reg_5_19_inst : DFFR_X1 port map( D => n3421, CK => CLK, RN => 
                           n673, Q => n816, QN => n_1421);
   REGISTERS_reg_5_18_inst : DFFR_X1 port map( D => n3420, CK => CLK, RN => 
                           n673, Q => n817, QN => n_1422);
   REGISTERS_reg_5_17_inst : DFFR_X1 port map( D => n3419, CK => CLK, RN => 
                           n672, Q => n818, QN => n_1423);
   REGISTERS_reg_5_16_inst : DFFR_X1 port map( D => n3418, CK => CLK, RN => 
                           n672, Q => n819, QN => n_1424);
   REGISTERS_reg_5_15_inst : DFFR_X1 port map( D => n3417, CK => CLK, RN => 
                           n672, Q => n820, QN => n_1425);
   REGISTERS_reg_5_14_inst : DFFR_X1 port map( D => n3416, CK => CLK, RN => 
                           n672, Q => n821, QN => n_1426);
   REGISTERS_reg_5_13_inst : DFFR_X1 port map( D => n3415, CK => CLK, RN => 
                           n672, Q => n822, QN => n_1427);
   REGISTERS_reg_5_12_inst : DFFR_X1 port map( D => n3414, CK => CLK, RN => 
                           n672, Q => n823, QN => n_1428);
   REGISTERS_reg_5_11_inst : DFFR_X1 port map( D => n3413, CK => CLK, RN => 
                           n672, Q => n824, QN => n_1429);
   REGISTERS_reg_5_10_inst : DFFR_X1 port map( D => n3412, CK => CLK, RN => 
                           n672, Q => n825, QN => n_1430);
   REGISTERS_reg_5_9_inst : DFFR_X1 port map( D => n3411, CK => CLK, RN => n672
                           , Q => n826, QN => n_1431);
   REGISTERS_reg_5_8_inst : DFFR_X1 port map( D => n3410, CK => CLK, RN => n672
                           , Q => n827, QN => n_1432);
   REGISTERS_reg_5_7_inst : DFFR_X1 port map( D => n3409, CK => CLK, RN => n672
                           , Q => n828, QN => n_1433);
   REGISTERS_reg_5_6_inst : DFFR_X1 port map( D => n3408, CK => CLK, RN => n672
                           , Q => n829, QN => n_1434);
   REGISTERS_reg_5_5_inst : DFFR_X1 port map( D => n3407, CK => CLK, RN => n671
                           , Q => n830, QN => n_1435);
   REGISTERS_reg_5_4_inst : DFFR_X1 port map( D => n3406, CK => CLK, RN => n671
                           , Q => n831, QN => n_1436);
   REGISTERS_reg_5_3_inst : DFFR_X1 port map( D => n3405, CK => CLK, RN => n671
                           , Q => n832, QN => n_1437);
   REGISTERS_reg_5_2_inst : DFFR_X1 port map( D => n3404, CK => CLK, RN => n671
                           , Q => n833, QN => n_1438);
   REGISTERS_reg_5_1_inst : DFFR_X1 port map( D => n3403, CK => CLK, RN => n671
                           , Q => n834, QN => n_1439);
   REGISTERS_reg_5_0_inst : DFFR_X1 port map( D => n3402, CK => CLK, RN => n671
                           , Q => n835, QN => n_1440);
   REGISTERS_reg_4_23_inst : DFFR_X1 port map( D => n3457, CK => CLK, RN => 
                           n655, Q => n778, QN => n_1441);
   REGISTERS_reg_4_22_inst : DFFR_X1 port map( D => n3456, CK => CLK, RN => 
                           n655, Q => n779, QN => n_1442);
   REGISTERS_reg_4_21_inst : DFFR_X1 port map( D => n3455, CK => CLK, RN => 
                           n655, Q => n780, QN => n_1443);
   REGISTERS_reg_4_20_inst : DFFR_X1 port map( D => n3454, CK => CLK, RN => 
                           n655, Q => n781, QN => n_1444);
   REGISTERS_reg_4_19_inst : DFFR_X1 port map( D => n3453, CK => CLK, RN => 
                           n655, Q => n782, QN => n_1445);
   REGISTERS_reg_4_18_inst : DFFR_X1 port map( D => n3452, CK => CLK, RN => 
                           n655, Q => n783, QN => n_1446);
   REGISTERS_reg_4_17_inst : DFFR_X1 port map( D => n3451, CK => CLK, RN => 
                           n654, Q => n784, QN => n_1447);
   REGISTERS_reg_4_16_inst : DFFR_X1 port map( D => n3450, CK => CLK, RN => 
                           n654, Q => n785, QN => n_1448);
   REGISTERS_reg_4_15_inst : DFFR_X1 port map( D => n3449, CK => CLK, RN => 
                           n654, Q => n786, QN => n_1449);
   REGISTERS_reg_4_14_inst : DFFR_X1 port map( D => n3448, CK => CLK, RN => 
                           n654, Q => n787, QN => n_1450);
   REGISTERS_reg_4_13_inst : DFFR_X1 port map( D => n3447, CK => CLK, RN => 
                           n654, Q => n788, QN => n_1451);
   REGISTERS_reg_4_12_inst : DFFR_X1 port map( D => n3446, CK => CLK, RN => 
                           n654, Q => n789, QN => n_1452);
   REGISTERS_reg_4_11_inst : DFFR_X1 port map( D => n3445, CK => CLK, RN => 
                           n654, Q => n790, QN => n_1453);
   REGISTERS_reg_4_10_inst : DFFR_X1 port map( D => n3444, CK => CLK, RN => 
                           n654, Q => n791, QN => n_1454);
   REGISTERS_reg_4_9_inst : DFFR_X1 port map( D => n3443, CK => CLK, RN => n654
                           , Q => n792, QN => n_1455);
   REGISTERS_reg_4_8_inst : DFFR_X1 port map( D => n3442, CK => CLK, RN => n654
                           , Q => n793, QN => n_1456);
   REGISTERS_reg_4_7_inst : DFFR_X1 port map( D => n3441, CK => CLK, RN => n654
                           , Q => n794, QN => n_1457);
   REGISTERS_reg_4_6_inst : DFFR_X1 port map( D => n3440, CK => CLK, RN => n654
                           , Q => n795, QN => n_1458);
   REGISTERS_reg_4_5_inst : DFFR_X1 port map( D => n3439, CK => CLK, RN => n653
                           , Q => n796, QN => n_1459);
   REGISTERS_reg_4_4_inst : DFFR_X1 port map( D => n3438, CK => CLK, RN => n653
                           , Q => n797, QN => n_1460);
   REGISTERS_reg_4_3_inst : DFFR_X1 port map( D => n3437, CK => CLK, RN => n653
                           , Q => n798, QN => n_1461);
   REGISTERS_reg_4_2_inst : DFFR_X1 port map( D => n3436, CK => CLK, RN => n658
                           , Q => n799, QN => n_1462);
   REGISTERS_reg_4_1_inst : DFFR_X1 port map( D => n3435, CK => CLK, RN => n674
                           , Q => n800, QN => n_1463);
   REGISTERS_reg_4_0_inst : DFFR_X1 port map( D => n3434, CK => CLK, RN => n674
                           , Q => n801, QN => n_1464);
   REGISTERS_reg_1_23_inst : DFFR_X1 port map( D => n3553, CK => CLK, RN => 
                           n663, Q => n739, QN => n_1465);
   REGISTERS_reg_1_22_inst : DFFR_X1 port map( D => n3552, CK => CLK, RN => 
                           n663, Q => n740, QN => n_1466);
   REGISTERS_reg_1_21_inst : DFFR_X1 port map( D => n3551, CK => CLK, RN => 
                           n663, Q => n741, QN => n_1467);
   REGISTERS_reg_1_20_inst : DFFR_X1 port map( D => n3550, CK => CLK, RN => 
                           n663, Q => n742, QN => n_1468);
   REGISTERS_reg_1_19_inst : DFFR_X1 port map( D => n3549, CK => CLK, RN => 
                           n663, Q => n743, QN => n_1469);
   REGISTERS_reg_1_18_inst : DFFR_X1 port map( D => n3548, CK => CLK, RN => 
                           n663, Q => n744, QN => n_1470);
   REGISTERS_reg_1_17_inst : DFFR_X1 port map( D => n3547, CK => CLK, RN => 
                           n663, Q => n745, QN => n_1471);
   REGISTERS_reg_1_16_inst : DFFR_X1 port map( D => n3546, CK => CLK, RN => 
                           n662, Q => n746, QN => n_1472);
   REGISTERS_reg_1_15_inst : DFFR_X1 port map( D => n3545, CK => CLK, RN => 
                           n662, Q => n747, QN => n_1473);
   REGISTERS_reg_1_14_inst : DFFR_X1 port map( D => n3544, CK => CLK, RN => 
                           n662, Q => n748, QN => n_1474);
   REGISTERS_reg_1_13_inst : DFFR_X1 port map( D => n3543, CK => CLK, RN => 
                           n662, Q => n749, QN => n_1475);
   REGISTERS_reg_1_12_inst : DFFR_X1 port map( D => n3542, CK => CLK, RN => 
                           n662, Q => n750, QN => n_1476);
   REGISTERS_reg_1_11_inst : DFFR_X1 port map( D => n3541, CK => CLK, RN => 
                           n662, Q => n751, QN => n_1477);
   REGISTERS_reg_1_10_inst : DFFR_X1 port map( D => n3540, CK => CLK, RN => 
                           n662, Q => n752, QN => n_1478);
   REGISTERS_reg_1_9_inst : DFFR_X1 port map( D => n3539, CK => CLK, RN => n662
                           , Q => n753, QN => n_1479);
   REGISTERS_reg_1_8_inst : DFFR_X1 port map( D => n3538, CK => CLK, RN => n662
                           , Q => n754, QN => n_1480);
   REGISTERS_reg_1_7_inst : DFFR_X1 port map( D => n3537, CK => CLK, RN => n662
                           , Q => n755, QN => n_1481);
   REGISTERS_reg_1_6_inst : DFFR_X1 port map( D => n3536, CK => CLK, RN => n662
                           , Q => n756, QN => n_1482);
   REGISTERS_reg_1_5_inst : DFFR_X1 port map( D => n3535, CK => CLK, RN => n662
                           , Q => n757, QN => n_1483);
   REGISTERS_reg_1_4_inst : DFFR_X1 port map( D => n3534, CK => CLK, RN => n661
                           , Q => n758, QN => n_1484);
   REGISTERS_reg_1_3_inst : DFFR_X1 port map( D => n3533, CK => CLK, RN => n661
                           , Q => n759, QN => n_1485);
   REGISTERS_reg_1_2_inst : DFFR_X1 port map( D => n3532, CK => CLK, RN => n661
                           , Q => n760, QN => n_1486);
   REGISTERS_reg_1_1_inst : DFFR_X1 port map( D => n3531, CK => CLK, RN => n661
                           , Q => n761, QN => n_1487);
   REGISTERS_reg_1_0_inst : DFFR_X1 port map( D => n3530, CK => CLK, RN => n661
                           , Q => n762, QN => n_1488);
   REGISTERS_reg_13_31_inst : DFFR_X1 port map( D => n3177, CK => CLK, RN => 
                           n652, Q => n_1489, QN => n389);
   REGISTERS_reg_13_30_inst : DFFR_X1 port map( D => n3176, CK => CLK, RN => 
                           n652, Q => n_1490, QN => n390);
   REGISTERS_reg_13_29_inst : DFFR_X1 port map( D => n3175, CK => CLK, RN => 
                           n652, Q => n_1491, QN => n391);
   REGISTERS_reg_13_28_inst : DFFR_X1 port map( D => n3174, CK => CLK, RN => 
                           n652, Q => n_1492, QN => n392);
   REGISTERS_reg_13_27_inst : DFFR_X1 port map( D => n3173, CK => CLK, RN => 
                           n652, Q => n_1493, QN => n393);
   REGISTERS_reg_13_26_inst : DFFR_X1 port map( D => n3172, CK => CLK, RN => 
                           n652, Q => n_1494, QN => n394);
   REGISTERS_reg_13_25_inst : DFFR_X1 port map( D => n3171, CK => CLK, RN => 
                           n652, Q => n_1495, QN => n395);
   REGISTERS_reg_13_24_inst : DFFR_X1 port map( D => n3170, CK => CLK, RN => 
                           n652, Q => n_1496, QN => n396);
   REGISTERS_reg_12_31_inst : DFFR_X1 port map( D => n3209, CK => CLK, RN => 
                           n602, Q => n_1497, QN => n357);
   REGISTERS_reg_12_30_inst : DFFR_X1 port map( D => n3208, CK => CLK, RN => 
                           n602, Q => n_1498, QN => n358);
   REGISTERS_reg_12_29_inst : DFFR_X1 port map( D => n3207, CK => CLK, RN => 
                           n602, Q => n_1499, QN => n359);
   REGISTERS_reg_12_28_inst : DFFR_X1 port map( D => n3206, CK => CLK, RN => 
                           n602, Q => n_1500, QN => n360);
   REGISTERS_reg_12_27_inst : DFFR_X1 port map( D => n3205, CK => CLK, RN => 
                           n602, Q => n_1501, QN => n361);
   REGISTERS_reg_12_26_inst : DFFR_X1 port map( D => n3204, CK => CLK, RN => 
                           n602, Q => n_1502, QN => n362);
   REGISTERS_reg_12_25_inst : DFFR_X1 port map( D => n3203, CK => CLK, RN => 
                           n602, Q => n_1503, QN => n363);
   REGISTERS_reg_12_24_inst : DFFR_X1 port map( D => n3202, CK => CLK, RN => 
                           n602, Q => n_1504, QN => n364);
   REGISTERS_reg_20_31_inst : DFFR_X1 port map( D => n2953, CK => CLK, RN => 
                           n696, Q => n_1505, QN => n613);
   REGISTERS_reg_20_30_inst : DFFR_X1 port map( D => n2952, CK => CLK, RN => 
                           n695, Q => n_1506, QN => n614);
   REGISTERS_reg_20_29_inst : DFFR_X1 port map( D => n2951, CK => CLK, RN => 
                           n695, Q => n_1507, QN => n615);
   REGISTERS_reg_20_28_inst : DFFR_X1 port map( D => n2950, CK => CLK, RN => 
                           n695, Q => n_1508, QN => n616);
   REGISTERS_reg_20_27_inst : DFFR_X1 port map( D => n2949, CK => CLK, RN => 
                           n695, Q => n_1509, QN => n617);
   REGISTERS_reg_20_26_inst : DFFR_X1 port map( D => n2948, CK => CLK, RN => 
                           n695, Q => n_1510, QN => n618);
   REGISTERS_reg_20_25_inst : DFFR_X1 port map( D => n2947, CK => CLK, RN => 
                           n695, Q => n_1511, QN => n619);
   REGISTERS_reg_20_24_inst : DFFR_X1 port map( D => n2946, CK => CLK, RN => 
                           n695, Q => n_1512, QN => n620);
   REGISTERS_reg_9_31_inst : DFFR_X1 port map( D => n3305, CK => CLK, RN => 
                           n610, Q => n_1513, QN => n261);
   REGISTERS_reg_9_30_inst : DFFR_X1 port map( D => n3304, CK => CLK, RN => 
                           n610, Q => n_1514, QN => n262);
   REGISTERS_reg_9_29_inst : DFFR_X1 port map( D => n3303, CK => CLK, RN => 
                           n610, Q => n_1515, QN => n263);
   REGISTERS_reg_9_28_inst : DFFR_X1 port map( D => n3302, CK => CLK, RN => 
                           n610, Q => n_1516, QN => n264);
   REGISTERS_reg_9_27_inst : DFFR_X1 port map( D => n3301, CK => CLK, RN => 
                           n610, Q => n_1517, QN => n265);
   REGISTERS_reg_9_26_inst : DFFR_X1 port map( D => n3300, CK => CLK, RN => 
                           n610, Q => n_1518, QN => n266);
   REGISTERS_reg_9_25_inst : DFFR_X1 port map( D => n3299, CK => CLK, RN => 
                           n610, Q => n_1519, QN => n267);
   REGISTERS_reg_9_24_inst : DFFR_X1 port map( D => n3298, CK => CLK, RN => 
                           n610, Q => n_1520, QN => n268);
   REGISTERS_reg_17_31_inst : DFFR_X1 port map( D => n3049, CK => CLK, RN => 
                           n704, Q => n_1521, QN => n517);
   REGISTERS_reg_17_30_inst : DFFR_X1 port map( D => n3048, CK => CLK, RN => 
                           n704, Q => n_1522, QN => n518);
   REGISTERS_reg_17_29_inst : DFFR_X1 port map( D => n3047, CK => CLK, RN => 
                           n703, Q => n_1523, QN => n519);
   REGISTERS_reg_17_28_inst : DFFR_X1 port map( D => n3046, CK => CLK, RN => 
                           n703, Q => n_1524, QN => n520);
   REGISTERS_reg_17_27_inst : DFFR_X1 port map( D => n3045, CK => CLK, RN => 
                           n703, Q => n_1525, QN => n521);
   REGISTERS_reg_17_26_inst : DFFR_X1 port map( D => n3044, CK => CLK, RN => 
                           n703, Q => n_1526, QN => n522);
   REGISTERS_reg_17_25_inst : DFFR_X1 port map( D => n3043, CK => CLK, RN => 
                           n703, Q => n_1527, QN => n523);
   REGISTERS_reg_17_24_inst : DFFR_X1 port map( D => n3042, CK => CLK, RN => 
                           n703, Q => n_1528, QN => n524);
   REGISTERS_reg_8_31_inst : DFFR_X1 port map( D => n3337, CK => CLK, RN => 
                           n666, Q => n_1529, QN => n229);
   REGISTERS_reg_8_30_inst : DFFR_X1 port map( D => n3336, CK => CLK, RN => 
                           n665, Q => n_1530, QN => n230);
   REGISTERS_reg_8_29_inst : DFFR_X1 port map( D => n3335, CK => CLK, RN => 
                           n665, Q => n_1531, QN => n231);
   REGISTERS_reg_8_28_inst : DFFR_X1 port map( D => n3334, CK => CLK, RN => 
                           n665, Q => n_1532, QN => n232);
   REGISTERS_reg_8_27_inst : DFFR_X1 port map( D => n3333, CK => CLK, RN => 
                           n665, Q => n_1533, QN => n233);
   REGISTERS_reg_8_26_inst : DFFR_X1 port map( D => n3332, CK => CLK, RN => 
                           n665, Q => n_1534, QN => n234);
   REGISTERS_reg_8_25_inst : DFFR_X1 port map( D => n3331, CK => CLK, RN => 
                           n665, Q => n_1535, QN => n235);
   REGISTERS_reg_8_24_inst : DFFR_X1 port map( D => n3330, CK => CLK, RN => 
                           n665, Q => n_1536, QN => n236);
   REGISTERS_reg_30_31_inst : DFFR_X1 port map( D => n2633, CK => CLK, RN => 
                           n690, Q => n_1537, QN => n933);
   REGISTERS_reg_30_30_inst : DFFR_X1 port map( D => n2632, CK => CLK, RN => 
                           n689, Q => n_1538, QN => n934);
   REGISTERS_reg_30_29_inst : DFFR_X1 port map( D => n2631, CK => CLK, RN => 
                           n689, Q => n_1539, QN => n935);
   REGISTERS_reg_30_28_inst : DFFR_X1 port map( D => n2630, CK => CLK, RN => 
                           n689, Q => n_1540, QN => n936);
   REGISTERS_reg_30_27_inst : DFFR_X1 port map( D => n2629, CK => CLK, RN => 
                           n689, Q => n_1541, QN => n937);
   REGISTERS_reg_30_26_inst : DFFR_X1 port map( D => n2628, CK => CLK, RN => 
                           n689, Q => n_1542, QN => n938);
   REGISTERS_reg_30_25_inst : DFFR_X1 port map( D => n2627, CK => CLK, RN => 
                           n689, Q => n_1543, QN => n939);
   REGISTERS_reg_30_24_inst : DFFR_X1 port map( D => n2626, CK => CLK, RN => 
                           n689, Q => n_1544, QN => n940);
   REGISTERS_reg_27_31_inst : DFFR_X1 port map( D => n2729, CK => CLK, RN => 
                           n677, Q => n_1545, QN => n837);
   REGISTERS_reg_27_30_inst : DFFR_X1 port map( D => n2728, CK => CLK, RN => 
                           n677, Q => n_1546, QN => n838);
   REGISTERS_reg_27_29_inst : DFFR_X1 port map( D => n2727, CK => CLK, RN => 
                           n677, Q => n_1547, QN => n839);
   REGISTERS_reg_27_28_inst : DFFR_X1 port map( D => n2726, CK => CLK, RN => 
                           n677, Q => n_1548, QN => n840);
   REGISTERS_reg_27_27_inst : DFFR_X1 port map( D => n2725, CK => CLK, RN => 
                           n676, Q => n_1549, QN => n841);
   REGISTERS_reg_27_26_inst : DFFR_X1 port map( D => n2724, CK => CLK, RN => 
                           n676, Q => n_1550, QN => n842);
   REGISTERS_reg_27_25_inst : DFFR_X1 port map( D => n2723, CK => CLK, RN => 
                           n676, Q => n_1551, QN => n843);
   REGISTERS_reg_27_24_inst : DFFR_X1 port map( D => n2722, CK => CLK, RN => 
                           n676, Q => n_1552, QN => n844);
   REGISTERS_reg_21_23_inst : DFFR_X1 port map( D => n2913, CK => CLK, RN => 
                           n713, Q => n1157, QN => n_1553);
   REGISTERS_reg_21_22_inst : DFFR_X1 port map( D => n2912, CK => CLK, RN => 
                           n713, Q => n1158, QN => n_1554);
   REGISTERS_reg_21_21_inst : DFFR_X1 port map( D => n2911, CK => CLK, RN => 
                           n713, Q => n1159, QN => n_1555);
   REGISTERS_reg_21_20_inst : DFFR_X1 port map( D => n2910, CK => CLK, RN => 
                           n713, Q => n1160, QN => n_1556);
   REGISTERS_reg_21_19_inst : DFFR_X1 port map( D => n2909, CK => CLK, RN => 
                           n713, Q => n1161, QN => n_1557);
   REGISTERS_reg_21_18_inst : DFFR_X1 port map( D => n2908, CK => CLK, RN => 
                           n712, Q => n1162, QN => n_1558);
   REGISTERS_reg_21_17_inst : DFFR_X1 port map( D => n2907, CK => CLK, RN => 
                           n712, Q => n1163, QN => n_1559);
   REGISTERS_reg_21_16_inst : DFFR_X1 port map( D => n2906, CK => CLK, RN => 
                           n712, Q => n1164, QN => n_1560);
   REGISTERS_reg_21_15_inst : DFFR_X1 port map( D => n2905, CK => CLK, RN => 
                           n712, Q => n1165, QN => n_1561);
   REGISTERS_reg_21_14_inst : DFFR_X1 port map( D => n2904, CK => CLK, RN => 
                           n712, Q => n1166, QN => n_1562);
   REGISTERS_reg_21_13_inst : DFFR_X1 port map( D => n2903, CK => CLK, RN => 
                           n712, Q => n1167, QN => n_1563);
   REGISTERS_reg_21_12_inst : DFFR_X1 port map( D => n2902, CK => CLK, RN => 
                           n712, Q => n1168, QN => n_1564);
   REGISTERS_reg_21_11_inst : DFFR_X1 port map( D => n2901, CK => CLK, RN => 
                           n712, Q => n1169, QN => n_1565);
   REGISTERS_reg_21_10_inst : DFFR_X1 port map( D => n2900, CK => CLK, RN => 
                           n712, Q => n1170, QN => n_1566);
   REGISTERS_reg_21_9_inst : DFFR_X1 port map( D => n2899, CK => CLK, RN => 
                           n712, Q => n1171, QN => n_1567);
   REGISTERS_reg_21_8_inst : DFFR_X1 port map( D => n2898, CK => CLK, RN => 
                           n712, Q => n1172, QN => n_1568);
   REGISTERS_reg_21_7_inst : DFFR_X1 port map( D => n2897, CK => CLK, RN => 
                           n712, Q => n1173, QN => n_1569);
   REGISTERS_reg_21_6_inst : DFFR_X1 port map( D => n2896, CK => CLK, RN => 
                           n711, Q => n1174, QN => n_1570);
   REGISTERS_reg_21_5_inst : DFFR_X1 port map( D => n2895, CK => CLK, RN => 
                           n711, Q => n1175, QN => n_1571);
   REGISTERS_reg_21_4_inst : DFFR_X1 port map( D => n2894, CK => CLK, RN => 
                           n711, Q => n1176, QN => n_1572);
   REGISTERS_reg_21_3_inst : DFFR_X1 port map( D => n2893, CK => CLK, RN => 
                           n711, Q => n1177, QN => n_1573);
   REGISTERS_reg_21_2_inst : DFFR_X1 port map( D => n2892, CK => CLK, RN => 
                           n711, Q => n1178, QN => n_1574);
   REGISTERS_reg_21_1_inst : DFFR_X1 port map( D => n2891, CK => CLK, RN => 
                           n711, Q => n1179, QN => n_1575);
   REGISTERS_reg_21_0_inst : DFFR_X1 port map( D => n2890, CK => CLK, RN => 
                           n711, Q => n1180, QN => n_1576);
   REGISTERS_reg_16_23_inst : DFFR_X1 port map( D => n3073, CK => CLK, RN => 
                           n611, Q => n1055, QN => n_1577);
   REGISTERS_reg_16_22_inst : DFFR_X1 port map( D => n3072, CK => CLK, RN => 
                           n611, Q => n1056, QN => n_1578);
   REGISTERS_reg_16_21_inst : DFFR_X1 port map( D => n3071, CK => CLK, RN => 
                           n611, Q => n1057, QN => n_1579);
   REGISTERS_reg_16_20_inst : DFFR_X1 port map( D => n3070, CK => CLK, RN => 
                           n611, Q => n1058, QN => n_1580);
   REGISTERS_reg_16_19_inst : DFFR_X1 port map( D => n3069, CK => CLK, RN => 
                           n611, Q => n1059, QN => n_1581);
   REGISTERS_reg_16_18_inst : DFFR_X1 port map( D => n3068, CK => CLK, RN => 
                           n611, Q => n1060, QN => n_1582);
   REGISTERS_reg_16_17_inst : DFFR_X1 port map( D => n3067, CK => CLK, RN => 
                           n611, Q => n1061, QN => n_1583);
   REGISTERS_reg_16_16_inst : DFFR_X1 port map( D => n3066, CK => CLK, RN => 
                           n648, Q => n1062, QN => n_1584);
   REGISTERS_reg_16_15_inst : DFFR_X1 port map( D => n3065, CK => CLK, RN => 
                           n653, Q => n1063, QN => n_1585);
   REGISTERS_reg_16_14_inst : DFFR_X1 port map( D => n3064, CK => CLK, RN => 
                           n705, Q => n1064, QN => n_1586);
   REGISTERS_reg_16_13_inst : DFFR_X1 port map( D => n3063, CK => CLK, RN => 
                           n705, Q => n1065, QN => n_1587);
   REGISTERS_reg_16_12_inst : DFFR_X1 port map( D => n3062, CK => CLK, RN => 
                           n705, Q => n1066, QN => n_1588);
   REGISTERS_reg_16_11_inst : DFFR_X1 port map( D => n3061, CK => CLK, RN => 
                           n705, Q => n1067, QN => n_1589);
   REGISTERS_reg_16_10_inst : DFFR_X1 port map( D => n3060, CK => CLK, RN => 
                           n705, Q => n1068, QN => n_1590);
   REGISTERS_reg_16_9_inst : DFFR_X1 port map( D => n3059, CK => CLK, RN => 
                           n704, Q => n1069, QN => n_1591);
   REGISTERS_reg_16_8_inst : DFFR_X1 port map( D => n3058, CK => CLK, RN => 
                           n704, Q => n1070, QN => n_1592);
   REGISTERS_reg_16_7_inst : DFFR_X1 port map( D => n3057, CK => CLK, RN => 
                           n704, Q => n1071, QN => n_1593);
   REGISTERS_reg_16_6_inst : DFFR_X1 port map( D => n3056, CK => CLK, RN => 
                           n704, Q => n1072, QN => n_1594);
   REGISTERS_reg_16_5_inst : DFFR_X1 port map( D => n3055, CK => CLK, RN => 
                           n704, Q => n1073, QN => n_1595);
   REGISTERS_reg_16_4_inst : DFFR_X1 port map( D => n3054, CK => CLK, RN => 
                           n704, Q => n1074, QN => n_1596);
   REGISTERS_reg_16_3_inst : DFFR_X1 port map( D => n3053, CK => CLK, RN => 
                           n704, Q => n1075, QN => n_1597);
   REGISTERS_reg_16_2_inst : DFFR_X1 port map( D => n3052, CK => CLK, RN => 
                           n704, Q => n1076, QN => n_1598);
   REGISTERS_reg_16_1_inst : DFFR_X1 port map( D => n3051, CK => CLK, RN => 
                           n704, Q => n1077, QN => n_1599);
   REGISTERS_reg_16_0_inst : DFFR_X1 port map( D => n3050, CK => CLK, RN => 
                           n704, Q => n1078, QN => n_1600);
   REGISTERS_reg_31_23_inst : DFFR_X1 port map( D => n2593, CK => CLK, RN => 
                           n686, Q => n1298, QN => n_1601);
   REGISTERS_reg_31_22_inst : DFFR_X1 port map( D => n2592, CK => CLK, RN => 
                           n686, Q => n1299, QN => n_1602);
   REGISTERS_reg_31_21_inst : DFFR_X1 port map( D => n2591, CK => CLK, RN => 
                           n686, Q => n1300, QN => n_1603);
   REGISTERS_reg_31_20_inst : DFFR_X1 port map( D => n2590, CK => CLK, RN => 
                           n686, Q => n1301, QN => n_1604);
   REGISTERS_reg_31_19_inst : DFFR_X1 port map( D => n2589, CK => CLK, RN => 
                           n686, Q => n1302, QN => n_1605);
   REGISTERS_reg_31_18_inst : DFFR_X1 port map( D => n2588, CK => CLK, RN => 
                           n686, Q => n1303, QN => n_1606);
   REGISTERS_reg_31_17_inst : DFFR_X1 port map( D => n2587, CK => CLK, RN => 
                           n686, Q => n1304, QN => n_1607);
   REGISTERS_reg_31_16_inst : DFFR_X1 port map( D => n2586, CK => CLK, RN => 
                           n686, Q => n1305, QN => n_1608);
   REGISTERS_reg_31_15_inst : DFFR_X1 port map( D => n2585, CK => CLK, RN => 
                           n685, Q => n1306, QN => n_1609);
   REGISTERS_reg_31_14_inst : DFFR_X1 port map( D => n2584, CK => CLK, RN => 
                           n685, Q => n1307, QN => n_1610);
   REGISTERS_reg_31_13_inst : DFFR_X1 port map( D => n2583, CK => CLK, RN => 
                           n685, Q => n1308, QN => n_1611);
   REGISTERS_reg_31_12_inst : DFFR_X1 port map( D => n2582, CK => CLK, RN => 
                           n685, Q => n1309, QN => n_1612);
   REGISTERS_reg_31_11_inst : DFFR_X1 port map( D => n2581, CK => CLK, RN => 
                           n685, Q => n1310, QN => n_1613);
   REGISTERS_reg_31_10_inst : DFFR_X1 port map( D => n2580, CK => CLK, RN => 
                           n685, Q => n1311, QN => n_1614);
   REGISTERS_reg_31_9_inst : DFFR_X1 port map( D => n2579, CK => CLK, RN => 
                           n685, Q => n1312, QN => n_1615);
   REGISTERS_reg_31_8_inst : DFFR_X1 port map( D => n2578, CK => CLK, RN => 
                           n685, Q => n1313, QN => n_1616);
   REGISTERS_reg_31_7_inst : DFFR_X1 port map( D => n2577, CK => CLK, RN => 
                           n685, Q => n1314, QN => n_1617);
   REGISTERS_reg_31_6_inst : DFFR_X1 port map( D => n2576, CK => CLK, RN => 
                           n685, Q => n1315, QN => n_1618);
   REGISTERS_reg_31_5_inst : DFFR_X1 port map( D => n2575, CK => CLK, RN => 
                           n685, Q => n1316, QN => n_1619);
   REGISTERS_reg_31_4_inst : DFFR_X1 port map( D => n2574, CK => CLK, RN => 
                           n685, Q => n1317, QN => n_1620);
   REGISTERS_reg_31_3_inst : DFFR_X1 port map( D => n2573, CK => CLK, RN => 
                           n684, Q => n1318, QN => n_1621);
   REGISTERS_reg_31_2_inst : DFFR_X1 port map( D => n2572, CK => CLK, RN => 
                           n684, Q => n1319, QN => n_1622);
   REGISTERS_reg_31_1_inst : DFFR_X1 port map( D => n2571, CK => CLK, RN => 
                           n684, Q => n1320, QN => n_1623);
   REGISTERS_reg_31_0_inst : DFFR_X1 port map( D => n2570, CK => CLK, RN => 
                           n689, Q => n1321, QN => n_1624);
   REGISTERS_reg_26_23_inst : DFFR_X1 port map( D => n2753, CK => CLK, RN => 
                           n679, Q => n1196, QN => n_1625);
   REGISTERS_reg_26_22_inst : DFFR_X1 port map( D => n2752, CK => CLK, RN => 
                           n679, Q => n1197, QN => n_1626);
   REGISTERS_reg_26_21_inst : DFFR_X1 port map( D => n2751, CK => CLK, RN => 
                           n679, Q => n1198, QN => n_1627);
   REGISTERS_reg_26_20_inst : DFFR_X1 port map( D => n2750, CK => CLK, RN => 
                           n679, Q => n1199, QN => n_1628);
   REGISTERS_reg_26_19_inst : DFFR_X1 port map( D => n2749, CK => CLK, RN => 
                           n678, Q => n1200, QN => n_1629);
   REGISTERS_reg_26_18_inst : DFFR_X1 port map( D => n2748, CK => CLK, RN => 
                           n678, Q => n1201, QN => n_1630);
   REGISTERS_reg_26_17_inst : DFFR_X1 port map( D => n2747, CK => CLK, RN => 
                           n678, Q => n1202, QN => n_1631);
   REGISTERS_reg_26_16_inst : DFFR_X1 port map( D => n2746, CK => CLK, RN => 
                           n678, Q => n1203, QN => n_1632);
   REGISTERS_reg_26_15_inst : DFFR_X1 port map( D => n2745, CK => CLK, RN => 
                           n678, Q => n1204, QN => n_1633);
   REGISTERS_reg_26_14_inst : DFFR_X1 port map( D => n2744, CK => CLK, RN => 
                           n678, Q => n1205, QN => n_1634);
   REGISTERS_reg_26_13_inst : DFFR_X1 port map( D => n2743, CK => CLK, RN => 
                           n678, Q => n1206, QN => n_1635);
   REGISTERS_reg_26_12_inst : DFFR_X1 port map( D => n2742, CK => CLK, RN => 
                           n678, Q => n1207, QN => n_1636);
   REGISTERS_reg_26_11_inst : DFFR_X1 port map( D => n2741, CK => CLK, RN => 
                           n678, Q => n1208, QN => n_1637);
   REGISTERS_reg_26_10_inst : DFFR_X1 port map( D => n2740, CK => CLK, RN => 
                           n678, Q => n1209, QN => n_1638);
   REGISTERS_reg_26_9_inst : DFFR_X1 port map( D => n2739, CK => CLK, RN => 
                           n678, Q => n1210, QN => n_1639);
   REGISTERS_reg_26_8_inst : DFFR_X1 port map( D => n2738, CK => CLK, RN => 
                           n678, Q => n1211, QN => n_1640);
   REGISTERS_reg_26_7_inst : DFFR_X1 port map( D => n2737, CK => CLK, RN => 
                           n677, Q => n1212, QN => n_1641);
   REGISTERS_reg_26_6_inst : DFFR_X1 port map( D => n2736, CK => CLK, RN => 
                           n677, Q => n1213, QN => n_1642);
   REGISTERS_reg_26_5_inst : DFFR_X1 port map( D => n2735, CK => CLK, RN => 
                           n677, Q => n1214, QN => n_1643);
   REGISTERS_reg_26_4_inst : DFFR_X1 port map( D => n2734, CK => CLK, RN => 
                           n677, Q => n1215, QN => n_1644);
   REGISTERS_reg_26_3_inst : DFFR_X1 port map( D => n2733, CK => CLK, RN => 
                           n677, Q => n1216, QN => n_1645);
   REGISTERS_reg_26_2_inst : DFFR_X1 port map( D => n2732, CK => CLK, RN => 
                           n677, Q => n1217, QN => n_1646);
   REGISTERS_reg_26_1_inst : DFFR_X1 port map( D => n2731, CK => CLK, RN => 
                           n677, Q => n1218, QN => n_1647);
   REGISTERS_reg_26_0_inst : DFFR_X1 port map( D => n2730, CK => CLK, RN => 
                           n677, Q => n1219, QN => n_1648);
   REGISTERS_reg_13_23_inst : DFFR_X1 port map( D => n3169, CK => CLK, RN => 
                           n652, Q => n_1649, QN => n397);
   REGISTERS_reg_13_22_inst : DFFR_X1 port map( D => n3168, CK => CLK, RN => 
                           n651, Q => n_1650, QN => n398);
   REGISTERS_reg_13_21_inst : DFFR_X1 port map( D => n3167, CK => CLK, RN => 
                           n651, Q => n_1651, QN => n399);
   REGISTERS_reg_13_20_inst : DFFR_X1 port map( D => n3166, CK => CLK, RN => 
                           n651, Q => n_1652, QN => n400);
   REGISTERS_reg_13_19_inst : DFFR_X1 port map( D => n3165, CK => CLK, RN => 
                           n651, Q => n_1653, QN => n401);
   REGISTERS_reg_13_18_inst : DFFR_X1 port map( D => n3164, CK => CLK, RN => 
                           n651, Q => n_1654, QN => n402);
   REGISTERS_reg_13_17_inst : DFFR_X1 port map( D => n3163, CK => CLK, RN => 
                           n651, Q => n_1655, QN => n403);
   REGISTERS_reg_13_16_inst : DFFR_X1 port map( D => n3162, CK => CLK, RN => 
                           n651, Q => n_1656, QN => n404);
   REGISTERS_reg_13_15_inst : DFFR_X1 port map( D => n3161, CK => CLK, RN => 
                           n651, Q => n_1657, QN => n405);
   REGISTERS_reg_13_14_inst : DFFR_X1 port map( D => n3160, CK => CLK, RN => 
                           n651, Q => n_1658, QN => n406);
   REGISTERS_reg_13_13_inst : DFFR_X1 port map( D => n3159, CK => CLK, RN => 
                           n651, Q => n_1659, QN => n407);
   REGISTERS_reg_13_12_inst : DFFR_X1 port map( D => n3158, CK => CLK, RN => 
                           n651, Q => n_1660, QN => n408);
   REGISTERS_reg_13_11_inst : DFFR_X1 port map( D => n3157, CK => CLK, RN => 
                           n651, Q => n_1661, QN => n409);
   REGISTERS_reg_13_10_inst : DFFR_X1 port map( D => n3156, CK => CLK, RN => 
                           n650, Q => n_1662, QN => n410);
   REGISTERS_reg_13_9_inst : DFFR_X1 port map( D => n3155, CK => CLK, RN => 
                           n650, Q => n_1663, QN => n411);
   REGISTERS_reg_13_8_inst : DFFR_X1 port map( D => n3154, CK => CLK, RN => 
                           n650, Q => n_1664, QN => n412);
   REGISTERS_reg_13_7_inst : DFFR_X1 port map( D => n3153, CK => CLK, RN => 
                           n650, Q => n_1665, QN => n413);
   REGISTERS_reg_13_6_inst : DFFR_X1 port map( D => n3152, CK => CLK, RN => 
                           n650, Q => n_1666, QN => n414);
   REGISTERS_reg_13_5_inst : DFFR_X1 port map( D => n3151, CK => CLK, RN => 
                           n650, Q => n_1667, QN => n415);
   REGISTERS_reg_13_4_inst : DFFR_X1 port map( D => n3150, CK => CLK, RN => 
                           n650, Q => n_1668, QN => n416);
   REGISTERS_reg_13_3_inst : DFFR_X1 port map( D => n3149, CK => CLK, RN => 
                           n650, Q => n_1669, QN => n417);
   REGISTERS_reg_13_2_inst : DFFR_X1 port map( D => n3148, CK => CLK, RN => 
                           n650, Q => n_1670, QN => n418);
   REGISTERS_reg_13_1_inst : DFFR_X1 port map( D => n3147, CK => CLK, RN => 
                           n650, Q => n_1671, QN => n419);
   REGISTERS_reg_13_0_inst : DFFR_X1 port map( D => n3146, CK => CLK, RN => 
                           n650, Q => n_1672, QN => n420);
   REGISTERS_reg_12_23_inst : DFFR_X1 port map( D => n3201, CK => CLK, RN => 
                           n602, Q => n_1673, QN => n365);
   REGISTERS_reg_12_22_inst : DFFR_X1 port map( D => n3200, CK => CLK, RN => 
                           n601, Q => n_1674, QN => n366);
   REGISTERS_reg_12_21_inst : DFFR_X1 port map( D => n3199, CK => CLK, RN => 
                           n601, Q => n_1675, QN => n367);
   REGISTERS_reg_12_20_inst : DFFR_X1 port map( D => n3198, CK => CLK, RN => 
                           n601, Q => n_1676, QN => n368);
   REGISTERS_reg_12_19_inst : DFFR_X1 port map( D => n3197, CK => CLK, RN => 
                           n601, Q => n_1677, QN => n369);
   REGISTERS_reg_12_18_inst : DFFR_X1 port map( D => n3196, CK => CLK, RN => 
                           n601, Q => n_1678, QN => n370);
   REGISTERS_reg_12_17_inst : DFFR_X1 port map( D => n3195, CK => CLK, RN => 
                           n601, Q => n_1679, QN => n371);
   REGISTERS_reg_12_16_inst : DFFR_X1 port map( D => n3194, CK => CLK, RN => 
                           n601, Q => n_1680, QN => n372);
   REGISTERS_reg_12_15_inst : DFFR_X1 port map( D => n3193, CK => CLK, RN => 
                           n601, Q => n_1681, QN => n373);
   REGISTERS_reg_7_31_inst : DFFR_X1 port map( D => n3369, CK => CLK, RN => 
                           n668, Q => n4350, QN => n1374);
   REGISTERS_reg_7_30_inst : DFFR_X1 port map( D => n3368, CK => CLK, RN => 
                           n668, Q => n4349, QN => n1404);
   REGISTERS_reg_7_29_inst : DFFR_X1 port map( D => n3367, CK => CLK, RN => 
                           n668, Q => n4348, QN => n1429);
   REGISTERS_reg_7_28_inst : DFFR_X1 port map( D => n3366, CK => CLK, RN => 
                           n668, Q => n4347, QN => n1454);
   REGISTERS_reg_7_27_inst : DFFR_X1 port map( D => n3365, CK => CLK, RN => 
                           n668, Q => n4346, QN => n1479);
   REGISTERS_reg_7_26_inst : DFFR_X1 port map( D => n3364, CK => CLK, RN => 
                           n668, Q => n4345, QN => n1504);
   REGISTERS_reg_7_25_inst : DFFR_X1 port map( D => n3363, CK => CLK, RN => 
                           n668, Q => n4344, QN => n1529);
   REGISTERS_reg_7_24_inst : DFFR_X1 port map( D => n3362, CK => CLK, RN => 
                           n668, Q => n4343, QN => n1554);
   REGISTERS_reg_6_31_inst : DFFR_X1 port map( D => n3401, CK => CLK, RN => 
                           n671, Q => n4382, QN => n1372);
   REGISTERS_reg_6_30_inst : DFFR_X1 port map( D => n3400, CK => CLK, RN => 
                           n671, Q => n4381, QN => n1403);
   REGISTERS_reg_6_29_inst : DFFR_X1 port map( D => n3399, CK => CLK, RN => 
                           n671, Q => n4380, QN => n1428);
   REGISTERS_reg_6_28_inst : DFFR_X1 port map( D => n3398, CK => CLK, RN => 
                           n671, Q => n4379, QN => n1453);
   REGISTERS_reg_6_27_inst : DFFR_X1 port map( D => n3397, CK => CLK, RN => 
                           n671, Q => n4378, QN => n1478);
   REGISTERS_reg_6_26_inst : DFFR_X1 port map( D => n3396, CK => CLK, RN => 
                           n671, Q => n4377, QN => n1503);
   REGISTERS_reg_6_25_inst : DFFR_X1 port map( D => n3395, CK => CLK, RN => 
                           n670, Q => n4376, QN => n1528);
   REGISTERS_reg_6_24_inst : DFFR_X1 port map( D => n3394, CK => CLK, RN => 
                           n670, Q => n4375, QN => n1553);
   REGISTERS_reg_3_31_inst : DFFR_X1 port map( D => n3497, CK => CLK, RN => 
                           n658, Q => n4414, QN => n1381);
   REGISTERS_reg_3_30_inst : DFFR_X1 port map( D => n3496, CK => CLK, RN => 
                           n658, Q => n4413, QN => n1407);
   REGISTERS_reg_3_29_inst : DFFR_X1 port map( D => n3495, CK => CLK, RN => 
                           n658, Q => n4412, QN => n1432);
   REGISTERS_reg_3_28_inst : DFFR_X1 port map( D => n3494, CK => CLK, RN => 
                           n658, Q => n4411, QN => n1457);
   REGISTERS_reg_3_27_inst : DFFR_X1 port map( D => n3493, CK => CLK, RN => 
                           n658, Q => n4410, QN => n1482);
   REGISTERS_reg_3_26_inst : DFFR_X1 port map( D => n3492, CK => CLK, RN => 
                           n658, Q => n4409, QN => n1507);
   REGISTERS_reg_3_25_inst : DFFR_X1 port map( D => n3491, CK => CLK, RN => 
                           n658, Q => n4408, QN => n1532);
   REGISTERS_reg_3_24_inst : DFFR_X1 port map( D => n3490, CK => CLK, RN => 
                           n658, Q => n4407, QN => n1557);
   REGISTERS_reg_2_31_inst : DFFR_X1 port map( D => n3529, CK => CLK, RN => 
                           n661, Q => n4446, QN => n1379);
   REGISTERS_reg_2_30_inst : DFFR_X1 port map( D => n3528, CK => CLK, RN => 
                           n661, Q => n4445, QN => n1406);
   REGISTERS_reg_2_29_inst : DFFR_X1 port map( D => n3527, CK => CLK, RN => 
                           n661, Q => n4444, QN => n1431);
   REGISTERS_reg_2_28_inst : DFFR_X1 port map( D => n3526, CK => CLK, RN => 
                           n661, Q => n4443, QN => n1456);
   REGISTERS_reg_2_27_inst : DFFR_X1 port map( D => n3525, CK => CLK, RN => 
                           n661, Q => n4442, QN => n1481);
   REGISTERS_reg_2_26_inst : DFFR_X1 port map( D => n3524, CK => CLK, RN => 
                           n661, Q => n4441, QN => n1506);
   REGISTERS_reg_2_25_inst : DFFR_X1 port map( D => n3523, CK => CLK, RN => 
                           n661, Q => n4440, QN => n1531);
   REGISTERS_reg_2_24_inst : DFFR_X1 port map( D => n3522, CK => CLK, RN => 
                           n660, Q => n4439, QN => n1556);
   REGISTERS_reg_15_31_inst : DFFR_X1 port map( D => n3113, CK => CLK, RN => 
                           n647, Q => n4222, QN => n_1682);
   REGISTERS_reg_15_30_inst : DFFR_X1 port map( D => n3112, CK => CLK, RN => 
                           n647, Q => n4221, QN => n_1683);
   REGISTERS_reg_15_29_inst : DFFR_X1 port map( D => n3111, CK => CLK, RN => 
                           n647, Q => n4220, QN => n_1684);
   REGISTERS_reg_15_28_inst : DFFR_X1 port map( D => n3110, CK => CLK, RN => 
                           n647, Q => n4219, QN => n_1685);
   REGISTERS_reg_15_27_inst : DFFR_X1 port map( D => n3109, CK => CLK, RN => 
                           n646, Q => n4218, QN => n_1686);
   REGISTERS_reg_15_26_inst : DFFR_X1 port map( D => n3108, CK => CLK, RN => 
                           n646, Q => n4217, QN => n_1687);
   REGISTERS_reg_15_25_inst : DFFR_X1 port map( D => n3107, CK => CLK, RN => 
                           n646, Q => n4216, QN => n_1688);
   REGISTERS_reg_15_24_inst : DFFR_X1 port map( D => n3106, CK => CLK, RN => 
                           n646, Q => n4215, QN => n_1689);
   REGISTERS_reg_14_31_inst : DFFR_X1 port map( D => n3145, CK => CLK, RN => 
                           n650, Q => n4254, QN => n_1690);
   REGISTERS_reg_14_30_inst : DFFR_X1 port map( D => n3144, CK => CLK, RN => 
                           n649, Q => n4253, QN => n_1691);
   REGISTERS_reg_14_29_inst : DFFR_X1 port map( D => n3143, CK => CLK, RN => 
                           n649, Q => n4252, QN => n_1692);
   REGISTERS_reg_14_28_inst : DFFR_X1 port map( D => n3142, CK => CLK, RN => 
                           n649, Q => n4251, QN => n_1693);
   REGISTERS_reg_14_27_inst : DFFR_X1 port map( D => n3141, CK => CLK, RN => 
                           n649, Q => n4250, QN => n_1694);
   REGISTERS_reg_14_26_inst : DFFR_X1 port map( D => n3140, CK => CLK, RN => 
                           n649, Q => n4249, QN => n_1695);
   REGISTERS_reg_14_25_inst : DFFR_X1 port map( D => n3139, CK => CLK, RN => 
                           n649, Q => n4248, QN => n_1696);
   REGISTERS_reg_14_24_inst : DFFR_X1 port map( D => n3138, CK => CLK, RN => 
                           n649, Q => n4247, QN => n_1697);
   REGISTERS_reg_23_31_inst : DFFR_X1 port map( D => n2857, CK => CLK, RN => 
                           n708, Q => n4094, QN => n1333);
   REGISTERS_reg_23_30_inst : DFFR_X1 port map( D => n2856, CK => CLK, RN => 
                           n708, Q => n4093, QN => n1388);
   REGISTERS_reg_23_29_inst : DFFR_X1 port map( D => n2855, CK => CLK, RN => 
                           n708, Q => n4092, QN => n1413);
   REGISTERS_reg_23_28_inst : DFFR_X1 port map( D => n2854, CK => CLK, RN => 
                           n708, Q => n4091, QN => n1438);
   REGISTERS_reg_23_27_inst : DFFR_X1 port map( D => n2853, CK => CLK, RN => 
                           n708, Q => n4090, QN => n1463);
   REGISTERS_reg_23_26_inst : DFFR_X1 port map( D => n2852, CK => CLK, RN => 
                           n708, Q => n4089, QN => n1488);
   REGISTERS_reg_23_25_inst : DFFR_X1 port map( D => n2851, CK => CLK, RN => 
                           n708, Q => n4088, QN => n1513);
   REGISTERS_reg_23_24_inst : DFFR_X1 port map( D => n2850, CK => CLK, RN => 
                           n708, Q => n4087, QN => n1538);
   REGISTERS_reg_22_31_inst : DFFR_X1 port map( D => n2889, CK => CLK, RN => 
                           n711, Q => n4126, QN => n1351);
   REGISTERS_reg_22_30_inst : DFFR_X1 port map( D => n2888, CK => CLK, RN => 
                           n711, Q => n4125, QN => n1395);
   REGISTERS_reg_22_29_inst : DFFR_X1 port map( D => n2887, CK => CLK, RN => 
                           n711, Q => n4124, QN => n1420);
   REGISTERS_reg_22_28_inst : DFFR_X1 port map( D => n2886, CK => CLK, RN => 
                           n711, Q => n4123, QN => n1445);
   REGISTERS_reg_22_27_inst : DFFR_X1 port map( D => n2885, CK => CLK, RN => 
                           n711, Q => n4122, QN => n1470);
   REGISTERS_reg_22_26_inst : DFFR_X1 port map( D => n2884, CK => CLK, RN => 
                           n710, Q => n4121, QN => n1495);
   REGISTERS_reg_22_25_inst : DFFR_X1 port map( D => n2883, CK => CLK, RN => 
                           n710, Q => n4120, QN => n1520);
   REGISTERS_reg_22_24_inst : DFFR_X1 port map( D => n2882, CK => CLK, RN => 
                           n710, Q => n4119, QN => n1545);
   REGISTERS_reg_11_31_inst : DFFR_X1 port map( D => n3241, CK => CLK, RN => 
                           n605, Q => n4286, QN => n_1698);
   REGISTERS_reg_11_30_inst : DFFR_X1 port map( D => n3240, CK => CLK, RN => 
                           n605, Q => n4285, QN => n_1699);
   REGISTERS_reg_11_29_inst : DFFR_X1 port map( D => n3239, CK => CLK, RN => 
                           n605, Q => n4284, QN => n_1700);
   REGISTERS_reg_11_28_inst : DFFR_X1 port map( D => n3238, CK => CLK, RN => 
                           n605, Q => n4283, QN => n_1701);
   REGISTERS_reg_11_27_inst : DFFR_X1 port map( D => n3237, CK => CLK, RN => 
                           n605, Q => n4282, QN => n_1702);
   REGISTERS_reg_11_26_inst : DFFR_X1 port map( D => n3236, CK => CLK, RN => 
                           n604, Q => n4281, QN => n_1703);
   REGISTERS_reg_11_25_inst : DFFR_X1 port map( D => n3235, CK => CLK, RN => 
                           n604, Q => n4280, QN => n_1704);
   REGISTERS_reg_11_24_inst : DFFR_X1 port map( D => n3234, CK => CLK, RN => 
                           n604, Q => n4279, QN => n_1705);
   REGISTERS_reg_10_31_inst : DFFR_X1 port map( D => n3273, CK => CLK, RN => 
                           n608, Q => n4318, QN => n_1706);
   REGISTERS_reg_10_30_inst : DFFR_X1 port map( D => n3272, CK => CLK, RN => 
                           n608, Q => n4317, QN => n_1707);
   REGISTERS_reg_10_29_inst : DFFR_X1 port map( D => n3271, CK => CLK, RN => 
                           n607, Q => n4316, QN => n_1708);
   REGISTERS_reg_10_28_inst : DFFR_X1 port map( D => n3270, CK => CLK, RN => 
                           n607, Q => n4315, QN => n_1709);
   REGISTERS_reg_10_27_inst : DFFR_X1 port map( D => n3269, CK => CLK, RN => 
                           n607, Q => n4314, QN => n_1710);
   REGISTERS_reg_10_26_inst : DFFR_X1 port map( D => n3268, CK => CLK, RN => 
                           n607, Q => n4313, QN => n_1711);
   REGISTERS_reg_10_25_inst : DFFR_X1 port map( D => n3267, CK => CLK, RN => 
                           n607, Q => n4312, QN => n_1712);
   REGISTERS_reg_10_24_inst : DFFR_X1 port map( D => n3266, CK => CLK, RN => 
                           n607, Q => n4311, QN => n_1713);
   REGISTERS_reg_19_31_inst : DFFR_X1 port map( D => n2985, CK => CLK, RN => 
                           n698, Q => n4158, QN => n_1714);
   REGISTERS_reg_19_30_inst : DFFR_X1 port map( D => n2984, CK => CLK, RN => 
                           n698, Q => n4157, QN => n_1715);
   REGISTERS_reg_19_29_inst : DFFR_X1 port map( D => n2983, CK => CLK, RN => 
                           n698, Q => n4156, QN => n_1716);
   REGISTERS_reg_19_28_inst : DFFR_X1 port map( D => n2982, CK => CLK, RN => 
                           n698, Q => n4155, QN => n_1717);
   REGISTERS_reg_19_27_inst : DFFR_X1 port map( D => n2981, CK => CLK, RN => 
                           n698, Q => n4154, QN => n_1718);
   REGISTERS_reg_19_26_inst : DFFR_X1 port map( D => n2980, CK => CLK, RN => 
                           n698, Q => n4153, QN => n_1719);
   REGISTERS_reg_19_25_inst : DFFR_X1 port map( D => n2979, CK => CLK, RN => 
                           n698, Q => n4152, QN => n_1720);
   REGISTERS_reg_19_24_inst : DFFR_X1 port map( D => n2978, CK => CLK, RN => 
                           n698, Q => n4151, QN => n_1721);
   REGISTERS_reg_18_31_inst : DFFR_X1 port map( D => n3017, CK => CLK, RN => 
                           n701, Q => n4190, QN => n_1722);
   REGISTERS_reg_18_30_inst : DFFR_X1 port map( D => n3016, CK => CLK, RN => 
                           n701, Q => n4189, QN => n_1723);
   REGISTERS_reg_18_29_inst : DFFR_X1 port map( D => n3015, CK => CLK, RN => 
                           n701, Q => n4188, QN => n_1724);
   REGISTERS_reg_18_28_inst : DFFR_X1 port map( D => n3014, CK => CLK, RN => 
                           n701, Q => n4187, QN => n_1725);
   REGISTERS_reg_18_27_inst : DFFR_X1 port map( D => n3013, CK => CLK, RN => 
                           n701, Q => n4186, QN => n_1726);
   REGISTERS_reg_18_26_inst : DFFR_X1 port map( D => n3012, CK => CLK, RN => 
                           n701, Q => n4185, QN => n_1727);
   REGISTERS_reg_18_25_inst : DFFR_X1 port map( D => n3011, CK => CLK, RN => 
                           n700, Q => n4184, QN => n_1728);
   REGISTERS_reg_18_24_inst : DFFR_X1 port map( D => n3010, CK => CLK, RN => 
                           n700, Q => n4183, QN => n_1729);
   REGISTERS_reg_29_31_inst : DFFR_X1 port map( D => n2665, CK => CLK, RN => 
                           n692, Q => n3966, QN => n_1730);
   REGISTERS_reg_29_30_inst : DFFR_X1 port map( D => n2664, CK => CLK, RN => 
                           n692, Q => n3965, QN => n_1731);
   REGISTERS_reg_29_29_inst : DFFR_X1 port map( D => n2663, CK => CLK, RN => 
                           n692, Q => n3964, QN => n_1732);
   REGISTERS_reg_29_28_inst : DFFR_X1 port map( D => n2662, CK => CLK, RN => 
                           n692, Q => n3963, QN => n_1733);
   REGISTERS_reg_29_27_inst : DFFR_X1 port map( D => n2661, CK => CLK, RN => 
                           n692, Q => n3962, QN => n_1734);
   REGISTERS_reg_29_26_inst : DFFR_X1 port map( D => n2660, CK => CLK, RN => 
                           n692, Q => n3961, QN => n_1735);
   REGISTERS_reg_29_25_inst : DFFR_X1 port map( D => n2659, CK => CLK, RN => 
                           n692, Q => n3960, QN => n_1736);
   REGISTERS_reg_29_24_inst : DFFR_X1 port map( D => n2658, CK => CLK, RN => 
                           n692, Q => n3959, QN => n_1737);
   REGISTERS_reg_28_31_inst : DFFR_X1 port map( D => n2697, CK => CLK, RN => 
                           n674, Q => n3998, QN => n1338);
   REGISTERS_reg_28_30_inst : DFFR_X1 port map( D => n2696, CK => CLK, RN => 
                           n674, Q => n3997, QN => n1390);
   REGISTERS_reg_28_29_inst : DFFR_X1 port map( D => n2695, CK => CLK, RN => 
                           n674, Q => n3996, QN => n1415);
   REGISTERS_reg_28_28_inst : DFFR_X1 port map( D => n2694, CK => CLK, RN => 
                           n679, Q => n3995, QN => n1440);
   REGISTERS_reg_28_27_inst : DFFR_X1 port map( D => n2693, CK => CLK, RN => 
                           n694, Q => n3994, QN => n1465);
   REGISTERS_reg_28_26_inst : DFFR_X1 port map( D => n2692, CK => CLK, RN => 
                           n695, Q => n3993, QN => n1490);
   REGISTERS_reg_28_25_inst : DFFR_X1 port map( D => n2691, CK => CLK, RN => 
                           n694, Q => n3992, QN => n1515);
   REGISTERS_reg_28_24_inst : DFFR_X1 port map( D => n2690, CK => CLK, RN => 
                           n694, Q => n3991, QN => n1540);
   REGISTERS_reg_25_31_inst : DFFR_X1 port map( D => n2793, CK => CLK, RN => 
                           n682, Q => n4030, QN => n_1738);
   REGISTERS_reg_25_30_inst : DFFR_X1 port map( D => n2792, CK => CLK, RN => 
                           n682, Q => n4029, QN => n_1739);
   REGISTERS_reg_25_29_inst : DFFR_X1 port map( D => n2791, CK => CLK, RN => 
                           n682, Q => n4028, QN => n_1740);
   REGISTERS_reg_25_28_inst : DFFR_X1 port map( D => n2790, CK => CLK, RN => 
                           n682, Q => n4027, QN => n_1741);
   REGISTERS_reg_25_27_inst : DFFR_X1 port map( D => n2789, CK => CLK, RN => 
                           n682, Q => n4026, QN => n_1742);
   REGISTERS_reg_25_26_inst : DFFR_X1 port map( D => n2788, CK => CLK, RN => 
                           n682, Q => n4025, QN => n_1743);
   REGISTERS_reg_25_25_inst : DFFR_X1 port map( D => n2787, CK => CLK, RN => 
                           n682, Q => n4024, QN => n_1744);
   REGISTERS_reg_25_24_inst : DFFR_X1 port map( D => n2786, CK => CLK, RN => 
                           n682, Q => n4023, QN => n_1745);
   REGISTERS_reg_24_31_inst : DFFR_X1 port map( D => n2825, CK => CLK, RN => 
                           n705, Q => n4062, QN => n_1746);
   REGISTERS_reg_24_30_inst : DFFR_X1 port map( D => n2824, CK => CLK, RN => 
                           n705, Q => n4061, QN => n_1747);
   REGISTERS_reg_24_29_inst : DFFR_X1 port map( D => n2823, CK => CLK, RN => 
                           n705, Q => n4060, QN => n_1748);
   REGISTERS_reg_24_28_inst : DFFR_X1 port map( D => n2822, CK => CLK, RN => 
                           n705, Q => n4059, QN => n_1749);
   REGISTERS_reg_24_27_inst : DFFR_X1 port map( D => n2821, CK => CLK, RN => 
                           n705, Q => n4058, QN => n_1750);
   REGISTERS_reg_24_26_inst : DFFR_X1 port map( D => n2820, CK => CLK, RN => 
                           n705, Q => n4057, QN => n_1751);
   REGISTERS_reg_24_25_inst : DFFR_X1 port map( D => n2819, CK => CLK, RN => 
                           n705, Q => n4056, QN => n_1752);
   REGISTERS_reg_24_24_inst : DFFR_X1 port map( D => n2818, CK => CLK, RN => 
                           n710, Q => n4055, QN => n_1753);
   REGISTERS_reg_7_23_inst : DFFR_X1 port map( D => n3361, CK => CLK, RN => 
                           n668, Q => n4342, QN => n1579);
   REGISTERS_reg_7_22_inst : DFFR_X1 port map( D => n3360, CK => CLK, RN => 
                           n667, Q => n4341, QN => n1604);
   REGISTERS_reg_7_21_inst : DFFR_X1 port map( D => n3359, CK => CLK, RN => 
                           n667, Q => n4340, QN => n1629);
   REGISTERS_reg_7_20_inst : DFFR_X1 port map( D => n3358, CK => CLK, RN => 
                           n667, Q => n4339, QN => n1654);
   REGISTERS_reg_7_19_inst : DFFR_X1 port map( D => n3357, CK => CLK, RN => 
                           n667, Q => n4338, QN => n1679);
   REGISTERS_reg_7_18_inst : DFFR_X1 port map( D => n3356, CK => CLK, RN => 
                           n667, Q => n4337, QN => n1704);
   REGISTERS_reg_7_17_inst : DFFR_X1 port map( D => n3355, CK => CLK, RN => 
                           n667, Q => n4336, QN => n1729);
   REGISTERS_reg_7_16_inst : DFFR_X1 port map( D => n3354, CK => CLK, RN => 
                           n667, Q => n4335, QN => n1754);
   REGISTERS_reg_7_15_inst : DFFR_X1 port map( D => n3353, CK => CLK, RN => 
                           n667, Q => n4334, QN => n1779);
   REGISTERS_reg_7_14_inst : DFFR_X1 port map( D => n3352, CK => CLK, RN => 
                           n667, Q => n4333, QN => n1804);
   REGISTERS_reg_7_13_inst : DFFR_X1 port map( D => n3351, CK => CLK, RN => 
                           n667, Q => n4332, QN => n1829);
   REGISTERS_reg_7_12_inst : DFFR_X1 port map( D => n3350, CK => CLK, RN => 
                           n667, Q => n4331, QN => n1854);
   REGISTERS_reg_7_11_inst : DFFR_X1 port map( D => n3349, CK => CLK, RN => 
                           n667, Q => n4330, QN => n1879);
   REGISTERS_reg_7_10_inst : DFFR_X1 port map( D => n3348, CK => CLK, RN => 
                           n666, Q => n4329, QN => n1904);
   REGISTERS_reg_7_9_inst : DFFR_X1 port map( D => n3347, CK => CLK, RN => n666
                           , Q => n4328, QN => n1929);
   REGISTERS_reg_7_8_inst : DFFR_X1 port map( D => n3346, CK => CLK, RN => n666
                           , Q => n4327, QN => n1954);
   REGISTERS_reg_7_7_inst : DFFR_X1 port map( D => n3345, CK => CLK, RN => n666
                           , Q => n4326, QN => n1979);
   REGISTERS_reg_7_6_inst : DFFR_X1 port map( D => n3344, CK => CLK, RN => n666
                           , Q => n4325, QN => n2004);
   REGISTERS_reg_7_5_inst : DFFR_X1 port map( D => n3343, CK => CLK, RN => n666
                           , Q => n4324, QN => n2029);
   REGISTERS_reg_7_4_inst : DFFR_X1 port map( D => n3342, CK => CLK, RN => n666
                           , Q => n4323, QN => n2054);
   REGISTERS_reg_7_3_inst : DFFR_X1 port map( D => n3341, CK => CLK, RN => n666
                           , Q => n4322, QN => n2079);
   REGISTERS_reg_7_2_inst : DFFR_X1 port map( D => n3340, CK => CLK, RN => n666
                           , Q => n4321, QN => n2104);
   REGISTERS_reg_7_1_inst : DFFR_X1 port map( D => n3339, CK => CLK, RN => n666
                           , Q => n4320, QN => n2129);
   REGISTERS_reg_7_0_inst : DFFR_X1 port map( D => n3338, CK => CLK, RN => n666
                           , Q => n4319, QN => n2167);
   REGISTERS_reg_6_23_inst : DFFR_X1 port map( D => n3393, CK => CLK, RN => 
                           n670, Q => n4374, QN => n1578);
   REGISTERS_reg_6_22_inst : DFFR_X1 port map( D => n3392, CK => CLK, RN => 
                           n670, Q => n4373, QN => n1603);
   REGISTERS_reg_6_21_inst : DFFR_X1 port map( D => n3391, CK => CLK, RN => 
                           n670, Q => n4372, QN => n1628);
   REGISTERS_reg_6_20_inst : DFFR_X1 port map( D => n3390, CK => CLK, RN => 
                           n670, Q => n4371, QN => n1653);
   REGISTERS_reg_6_19_inst : DFFR_X1 port map( D => n3389, CK => CLK, RN => 
                           n670, Q => n4370, QN => n1678);
   REGISTERS_reg_6_18_inst : DFFR_X1 port map( D => n3388, CK => CLK, RN => 
                           n670, Q => n4369, QN => n1703);
   REGISTERS_reg_6_17_inst : DFFR_X1 port map( D => n3387, CK => CLK, RN => 
                           n670, Q => n4368, QN => n1728);
   REGISTERS_reg_6_16_inst : DFFR_X1 port map( D => n3386, CK => CLK, RN => 
                           n670, Q => n4367, QN => n1753);
   REGISTERS_reg_6_15_inst : DFFR_X1 port map( D => n3385, CK => CLK, RN => 
                           n670, Q => n4366, QN => n1778);
   REGISTERS_reg_6_14_inst : DFFR_X1 port map( D => n3384, CK => CLK, RN => 
                           n670, Q => n4365, QN => n1803);
   REGISTERS_reg_6_13_inst : DFFR_X1 port map( D => n3383, CK => CLK, RN => 
                           n669, Q => n4364, QN => n1828);
   REGISTERS_reg_6_12_inst : DFFR_X1 port map( D => n3382, CK => CLK, RN => 
                           n669, Q => n4363, QN => n1853);
   REGISTERS_reg_6_11_inst : DFFR_X1 port map( D => n3381, CK => CLK, RN => 
                           n669, Q => n4362, QN => n1878);
   REGISTERS_reg_6_10_inst : DFFR_X1 port map( D => n3380, CK => CLK, RN => 
                           n669, Q => n4361, QN => n1903);
   REGISTERS_reg_6_9_inst : DFFR_X1 port map( D => n3379, CK => CLK, RN => n669
                           , Q => n4360, QN => n1928);
   REGISTERS_reg_6_8_inst : DFFR_X1 port map( D => n3378, CK => CLK, RN => n669
                           , Q => n4359, QN => n1953);
   REGISTERS_reg_6_7_inst : DFFR_X1 port map( D => n3377, CK => CLK, RN => n669
                           , Q => n4358, QN => n1978);
   REGISTERS_reg_6_6_inst : DFFR_X1 port map( D => n3376, CK => CLK, RN => n669
                           , Q => n4357, QN => n2003);
   REGISTERS_reg_6_5_inst : DFFR_X1 port map( D => n3375, CK => CLK, RN => n669
                           , Q => n4356, QN => n2028);
   REGISTERS_reg_6_4_inst : DFFR_X1 port map( D => n3374, CK => CLK, RN => n669
                           , Q => n4355, QN => n2053);
   REGISTERS_reg_6_3_inst : DFFR_X1 port map( D => n3373, CK => CLK, RN => n669
                           , Q => n4354, QN => n2078);
   REGISTERS_reg_6_2_inst : DFFR_X1 port map( D => n3372, CK => CLK, RN => n668
                           , Q => n4353, QN => n2103);
   REGISTERS_reg_6_1_inst : DFFR_X1 port map( D => n3371, CK => CLK, RN => n668
                           , Q => n4352, QN => n2128);
   REGISTERS_reg_6_0_inst : DFFR_X1 port map( D => n3370, CK => CLK, RN => n668
                           , Q => n4351, QN => n2166);
   REGISTERS_reg_3_23_inst : DFFR_X1 port map( D => n3489, CK => CLK, RN => 
                           n658, Q => n4406, QN => n1582);
   REGISTERS_reg_3_22_inst : DFFR_X1 port map( D => n3488, CK => CLK, RN => 
                           n658, Q => n4405, QN => n1607);
   REGISTERS_reg_3_21_inst : DFFR_X1 port map( D => n3487, CK => CLK, RN => 
                           n657, Q => n4404, QN => n1632);
   REGISTERS_reg_3_20_inst : DFFR_X1 port map( D => n3486, CK => CLK, RN => 
                           n657, Q => n4403, QN => n1657);
   REGISTERS_reg_3_19_inst : DFFR_X1 port map( D => n3485, CK => CLK, RN => 
                           n657, Q => n4402, QN => n1682);
   REGISTERS_reg_3_18_inst : DFFR_X1 port map( D => n3484, CK => CLK, RN => 
                           n657, Q => n4401, QN => n1707);
   REGISTERS_reg_3_17_inst : DFFR_X1 port map( D => n3483, CK => CLK, RN => 
                           n657, Q => n4400, QN => n1732);
   REGISTERS_reg_3_16_inst : DFFR_X1 port map( D => n3482, CK => CLK, RN => 
                           n657, Q => n4399, QN => n1757);
   REGISTERS_reg_3_15_inst : DFFR_X1 port map( D => n3481, CK => CLK, RN => 
                           n657, Q => n4398, QN => n1782);
   REGISTERS_reg_3_14_inst : DFFR_X1 port map( D => n3480, CK => CLK, RN => 
                           n657, Q => n4397, QN => n1807);
   REGISTERS_reg_3_13_inst : DFFR_X1 port map( D => n3479, CK => CLK, RN => 
                           n657, Q => n4396, QN => n1832);
   REGISTERS_reg_3_12_inst : DFFR_X1 port map( D => n3478, CK => CLK, RN => 
                           n657, Q => n4395, QN => n1857);
   REGISTERS_reg_3_11_inst : DFFR_X1 port map( D => n3477, CK => CLK, RN => 
                           n657, Q => n4394, QN => n1882);
   REGISTERS_reg_3_10_inst : DFFR_X1 port map( D => n3476, CK => CLK, RN => 
                           n657, Q => n4393, QN => n1907);
   REGISTERS_reg_3_9_inst : DFFR_X1 port map( D => n3475, CK => CLK, RN => n656
                           , Q => n4392, QN => n1932);
   REGISTERS_reg_3_8_inst : DFFR_X1 port map( D => n3474, CK => CLK, RN => n656
                           , Q => n4391, QN => n1957);
   REGISTERS_reg_3_7_inst : DFFR_X1 port map( D => n3473, CK => CLK, RN => n656
                           , Q => n4390, QN => n1982);
   REGISTERS_reg_3_6_inst : DFFR_X1 port map( D => n3472, CK => CLK, RN => n656
                           , Q => n4389, QN => n2007);
   REGISTERS_reg_3_5_inst : DFFR_X1 port map( D => n3471, CK => CLK, RN => n656
                           , Q => n4388, QN => n2032);
   REGISTERS_reg_3_4_inst : DFFR_X1 port map( D => n3470, CK => CLK, RN => n656
                           , Q => n4387, QN => n2057);
   REGISTERS_reg_3_3_inst : DFFR_X1 port map( D => n3469, CK => CLK, RN => n656
                           , Q => n4386, QN => n2082);
   REGISTERS_reg_3_2_inst : DFFR_X1 port map( D => n3468, CK => CLK, RN => n656
                           , Q => n4385, QN => n2107);
   REGISTERS_reg_3_1_inst : DFFR_X1 port map( D => n3467, CK => CLK, RN => n656
                           , Q => n4384, QN => n2132);
   REGISTERS_reg_3_0_inst : DFFR_X1 port map( D => n3466, CK => CLK, RN => n656
                           , Q => n4383, QN => n2172);
   REGISTERS_reg_2_23_inst : DFFR_X1 port map( D => n3521, CK => CLK, RN => 
                           n660, Q => n4438, QN => n1581);
   REGISTERS_reg_2_22_inst : DFFR_X1 port map( D => n3520, CK => CLK, RN => 
                           n660, Q => n4437, QN => n1606);
   REGISTERS_reg_2_21_inst : DFFR_X1 port map( D => n3519, CK => CLK, RN => 
                           n660, Q => n4436, QN => n1631);
   REGISTERS_reg_2_20_inst : DFFR_X1 port map( D => n3518, CK => CLK, RN => 
                           n660, Q => n4435, QN => n1656);
   REGISTERS_reg_2_19_inst : DFFR_X1 port map( D => n3517, CK => CLK, RN => 
                           n660, Q => n4434, QN => n1681);
   REGISTERS_reg_2_18_inst : DFFR_X1 port map( D => n3516, CK => CLK, RN => 
                           n660, Q => n4433, QN => n1706);
   REGISTERS_reg_2_17_inst : DFFR_X1 port map( D => n3515, CK => CLK, RN => 
                           n660, Q => n4432, QN => n1731);
   REGISTERS_reg_2_16_inst : DFFR_X1 port map( D => n3514, CK => CLK, RN => 
                           n660, Q => n4431, QN => n1756);
   REGISTERS_reg_2_15_inst : DFFR_X1 port map( D => n3513, CK => CLK, RN => 
                           n660, Q => n4430, QN => n1781);
   REGISTERS_reg_2_14_inst : DFFR_X1 port map( D => n3512, CK => CLK, RN => 
                           n660, Q => n4429, QN => n1806);
   REGISTERS_reg_2_13_inst : DFFR_X1 port map( D => n3511, CK => CLK, RN => 
                           n660, Q => n4428, QN => n1831);
   REGISTERS_reg_2_12_inst : DFFR_X1 port map( D => n3510, CK => CLK, RN => 
                           n659, Q => n4427, QN => n1856);
   REGISTERS_reg_2_11_inst : DFFR_X1 port map( D => n3509, CK => CLK, RN => 
                           n659, Q => n4426, QN => n1881);
   REGISTERS_reg_2_10_inst : DFFR_X1 port map( D => n3508, CK => CLK, RN => 
                           n659, Q => n4425, QN => n1906);
   REGISTERS_reg_2_9_inst : DFFR_X1 port map( D => n3507, CK => CLK, RN => n659
                           , Q => n4424, QN => n1931);
   REGISTERS_reg_2_8_inst : DFFR_X1 port map( D => n3506, CK => CLK, RN => n659
                           , Q => n4423, QN => n1956);
   REGISTERS_reg_2_7_inst : DFFR_X1 port map( D => n3505, CK => CLK, RN => n659
                           , Q => n4422, QN => n1981);
   REGISTERS_reg_2_6_inst : DFFR_X1 port map( D => n3504, CK => CLK, RN => n659
                           , Q => n4421, QN => n2006);
   REGISTERS_reg_2_5_inst : DFFR_X1 port map( D => n3503, CK => CLK, RN => n659
                           , Q => n4420, QN => n2031);
   REGISTERS_reg_2_4_inst : DFFR_X1 port map( D => n3502, CK => CLK, RN => n659
                           , Q => n4419, QN => n2056);
   REGISTERS_reg_2_3_inst : DFFR_X1 port map( D => n3501, CK => CLK, RN => n659
                           , Q => n4418, QN => n2081);
   REGISTERS_reg_2_2_inst : DFFR_X1 port map( D => n3500, CK => CLK, RN => n659
                           , Q => n4417, QN => n2106);
   REGISTERS_reg_2_1_inst : DFFR_X1 port map( D => n3499, CK => CLK, RN => n659
                           , Q => n4416, QN => n2131);
   REGISTERS_reg_2_0_inst : DFFR_X1 port map( D => n3498, CK => CLK, RN => n658
                           , Q => n4415, QN => n2171);
   REGISTERS_reg_15_23_inst : DFFR_X1 port map( D => n3105, CK => CLK, RN => 
                           n646, Q => n4214, QN => n_1754);
   REGISTERS_reg_15_22_inst : DFFR_X1 port map( D => n3104, CK => CLK, RN => 
                           n646, Q => n4213, QN => n_1755);
   REGISTERS_reg_15_21_inst : DFFR_X1 port map( D => n3103, CK => CLK, RN => 
                           n646, Q => n4212, QN => n_1756);
   REGISTERS_reg_15_20_inst : DFFR_X1 port map( D => n3102, CK => CLK, RN => 
                           n646, Q => n4211, QN => n_1757);
   REGISTERS_reg_15_19_inst : DFFR_X1 port map( D => n3101, CK => CLK, RN => 
                           n646, Q => n4210, QN => n_1758);
   REGISTERS_reg_15_18_inst : DFFR_X1 port map( D => n3100, CK => CLK, RN => 
                           n646, Q => n4209, QN => n_1759);
   REGISTERS_reg_15_17_inst : DFFR_X1 port map( D => n3099, CK => CLK, RN => 
                           n646, Q => n4208, QN => n_1760);
   REGISTERS_reg_15_16_inst : DFFR_X1 port map( D => n3098, CK => CLK, RN => 
                           n646, Q => n4207, QN => n_1761);
   REGISTERS_reg_15_15_inst : DFFR_X1 port map( D => n3097, CK => CLK, RN => 
                           n645, Q => n4206, QN => n_1762);
   REGISTERS_reg_15_14_inst : DFFR_X1 port map( D => n3096, CK => CLK, RN => 
                           n645, Q => n4205, QN => n_1763);
   REGISTERS_reg_15_13_inst : DFFR_X1 port map( D => n3095, CK => CLK, RN => 
                           n645, Q => n4204, QN => n_1764);
   REGISTERS_reg_15_12_inst : DFFR_X1 port map( D => n3094, CK => CLK, RN => 
                           n645, Q => n4203, QN => n_1765);
   REGISTERS_reg_15_11_inst : DFFR_X1 port map( D => n3093, CK => CLK, RN => 
                           n645, Q => n4202, QN => n_1766);
   REGISTERS_reg_15_10_inst : DFFR_X1 port map( D => n3092, CK => CLK, RN => 
                           n645, Q => n4201, QN => n_1767);
   REGISTERS_reg_15_9_inst : DFFR_X1 port map( D => n3091, CK => CLK, RN => 
                           n645, Q => n4200, QN => n_1768);
   REGISTERS_reg_15_8_inst : DFFR_X1 port map( D => n3090, CK => CLK, RN => 
                           n645, Q => n4199, QN => n_1769);
   REGISTERS_reg_15_7_inst : DFFR_X1 port map( D => n3089, CK => CLK, RN => 
                           n645, Q => n4198, QN => n_1770);
   REGISTERS_reg_15_6_inst : DFFR_X1 port map( D => n3088, CK => CLK, RN => 
                           n645, Q => n4197, QN => n_1771);
   REGISTERS_reg_15_5_inst : DFFR_X1 port map( D => n3087, CK => CLK, RN => 
                           n645, Q => n4196, QN => n_1772);
   REGISTERS_reg_15_4_inst : DFFR_X1 port map( D => n3086, CK => CLK, RN => 
                           n645, Q => n4195, QN => n_1773);
   REGISTERS_reg_15_3_inst : DFFR_X1 port map( D => n3085, CK => CLK, RN => 
                           n612, Q => n4194, QN => n_1774);
   REGISTERS_reg_15_2_inst : DFFR_X1 port map( D => n3084, CK => CLK, RN => 
                           n612, Q => n4193, QN => n_1775);
   REGISTERS_reg_15_1_inst : DFFR_X1 port map( D => n3083, CK => CLK, RN => 
                           n612, Q => n4192, QN => n_1776);
   REGISTERS_reg_15_0_inst : DFFR_X1 port map( D => n3082, CK => CLK, RN => 
                           n612, Q => n4191, QN => n_1777);
   REGISTERS_reg_14_23_inst : DFFR_X1 port map( D => n3137, CK => CLK, RN => 
                           n649, Q => n4246, QN => n_1778);
   REGISTERS_reg_14_22_inst : DFFR_X1 port map( D => n3136, CK => CLK, RN => 
                           n649, Q => n4245, QN => n_1779);
   REGISTERS_reg_14_21_inst : DFFR_X1 port map( D => n3135, CK => CLK, RN => 
                           n649, Q => n4244, QN => n_1780);
   REGISTERS_reg_14_20_inst : DFFR_X1 port map( D => n3134, CK => CLK, RN => 
                           n649, Q => n4243, QN => n_1781);
   REGISTERS_reg_14_19_inst : DFFR_X1 port map( D => n3133, CK => CLK, RN => 
                           n649, Q => n4242, QN => n_1782);
   REGISTERS_reg_14_18_inst : DFFR_X1 port map( D => n3132, CK => CLK, RN => 
                           n648, Q => n4241, QN => n_1783);
   REGISTERS_reg_14_17_inst : DFFR_X1 port map( D => n3131, CK => CLK, RN => 
                           n648, Q => n4240, QN => n_1784);
   REGISTERS_reg_14_16_inst : DFFR_X1 port map( D => n3130, CK => CLK, RN => 
                           n648, Q => n4239, QN => n_1785);
   REGISTERS_reg_14_15_inst : DFFR_X1 port map( D => n3129, CK => CLK, RN => 
                           n648, Q => n4238, QN => n_1786);
   REGISTERS_reg_14_14_inst : DFFR_X1 port map( D => n3128, CK => CLK, RN => 
                           n648, Q => n4237, QN => n_1787);
   REGISTERS_reg_14_13_inst : DFFR_X1 port map( D => n3127, CK => CLK, RN => 
                           n648, Q => n4236, QN => n_1788);
   REGISTERS_reg_14_12_inst : DFFR_X1 port map( D => n3126, CK => CLK, RN => 
                           n648, Q => n4235, QN => n_1789);
   REGISTERS_reg_14_11_inst : DFFR_X1 port map( D => n3125, CK => CLK, RN => 
                           n648, Q => n4234, QN => n_1790);
   REGISTERS_reg_14_10_inst : DFFR_X1 port map( D => n3124, CK => CLK, RN => 
                           n648, Q => n4233, QN => n_1791);
   REGISTERS_reg_14_9_inst : DFFR_X1 port map( D => n3123, CK => CLK, RN => 
                           n648, Q => n4232, QN => n_1792);
   REGISTERS_reg_14_8_inst : DFFR_X1 port map( D => n3122, CK => CLK, RN => 
                           n648, Q => n4231, QN => n_1793);
   REGISTERS_reg_14_7_inst : DFFR_X1 port map( D => n3121, CK => CLK, RN => 
                           n647, Q => n4230, QN => n_1794);
   REGISTERS_reg_14_6_inst : DFFR_X1 port map( D => n3120, CK => CLK, RN => 
                           n647, Q => n4229, QN => n_1795);
   REGISTERS_reg_14_5_inst : DFFR_X1 port map( D => n3119, CK => CLK, RN => 
                           n647, Q => n4228, QN => n_1796);
   REGISTERS_reg_14_4_inst : DFFR_X1 port map( D => n3118, CK => CLK, RN => 
                           n647, Q => n4227, QN => n_1797);
   REGISTERS_reg_14_3_inst : DFFR_X1 port map( D => n3117, CK => CLK, RN => 
                           n647, Q => n4226, QN => n_1798);
   REGISTERS_reg_14_2_inst : DFFR_X1 port map( D => n3116, CK => CLK, RN => 
                           n647, Q => n4225, QN => n_1799);
   REGISTERS_reg_14_1_inst : DFFR_X1 port map( D => n3115, CK => CLK, RN => 
                           n647, Q => n4224, QN => n_1800);
   REGISTERS_reg_14_0_inst : DFFR_X1 port map( D => n3114, CK => CLK, RN => 
                           n647, Q => n4223, QN => n_1801);
   REGISTERS_reg_23_23_inst : DFFR_X1 port map( D => n2849, CK => CLK, RN => 
                           n707, Q => n4086, QN => n1563);
   REGISTERS_reg_23_22_inst : DFFR_X1 port map( D => n2848, CK => CLK, RN => 
                           n707, Q => n4085, QN => n1588);
   REGISTERS_reg_23_21_inst : DFFR_X1 port map( D => n2847, CK => CLK, RN => 
                           n707, Q => n4084, QN => n1613);
   REGISTERS_reg_23_20_inst : DFFR_X1 port map( D => n2846, CK => CLK, RN => 
                           n707, Q => n4083, QN => n1638);
   REGISTERS_reg_23_19_inst : DFFR_X1 port map( D => n2845, CK => CLK, RN => 
                           n707, Q => n4082, QN => n1663);
   REGISTERS_reg_23_18_inst : DFFR_X1 port map( D => n2844, CK => CLK, RN => 
                           n707, Q => n4081, QN => n1688);
   REGISTERS_reg_23_17_inst : DFFR_X1 port map( D => n2843, CK => CLK, RN => 
                           n707, Q => n4080, QN => n1713);
   REGISTERS_reg_23_16_inst : DFFR_X1 port map( D => n2842, CK => CLK, RN => 
                           n707, Q => n4079, QN => n1738);
   REGISTERS_reg_23_15_inst : DFFR_X1 port map( D => n2841, CK => CLK, RN => 
                           n707, Q => n4078, QN => n1763);
   REGISTERS_reg_23_14_inst : DFFR_X1 port map( D => n2840, CK => CLK, RN => 
                           n707, Q => n4077, QN => n1788);
   REGISTERS_reg_23_13_inst : DFFR_X1 port map( D => n2839, CK => CLK, RN => 
                           n707, Q => n4076, QN => n1813);
   REGISTERS_reg_23_12_inst : DFFR_X1 port map( D => n2838, CK => CLK, RN => 
                           n707, Q => n4075, QN => n1838);
   REGISTERS_reg_23_11_inst : DFFR_X1 port map( D => n2837, CK => CLK, RN => 
                           n706, Q => n4074, QN => n1863);
   REGISTERS_reg_23_10_inst : DFFR_X1 port map( D => n2836, CK => CLK, RN => 
                           n706, Q => n4073, QN => n1888);
   REGISTERS_reg_23_9_inst : DFFR_X1 port map( D => n2835, CK => CLK, RN => 
                           n706, Q => n4072, QN => n1913);
   REGISTERS_reg_23_8_inst : DFFR_X1 port map( D => n2834, CK => CLK, RN => 
                           n706, Q => n4071, QN => n1938);
   REGISTERS_reg_23_7_inst : DFFR_X1 port map( D => n2833, CK => CLK, RN => 
                           n706, Q => n4070, QN => n1963);
   REGISTERS_reg_23_6_inst : DFFR_X1 port map( D => n2832, CK => CLK, RN => 
                           n706, Q => n4069, QN => n1988);
   REGISTERS_reg_23_5_inst : DFFR_X1 port map( D => n2831, CK => CLK, RN => 
                           n706, Q => n4068, QN => n2013);
   REGISTERS_reg_23_4_inst : DFFR_X1 port map( D => n2830, CK => CLK, RN => 
                           n706, Q => n4067, QN => n2038);
   REGISTERS_reg_23_3_inst : DFFR_X1 port map( D => n2829, CK => CLK, RN => 
                           n706, Q => n4066, QN => n2063);
   REGISTERS_reg_23_2_inst : DFFR_X1 port map( D => n2828, CK => CLK, RN => 
                           n706, Q => n4065, QN => n2088);
   REGISTERS_reg_23_1_inst : DFFR_X1 port map( D => n2827, CK => CLK, RN => 
                           n706, Q => n4064, QN => n2113);
   REGISTERS_reg_23_0_inst : DFFR_X1 port map( D => n2826, CK => CLK, RN => 
                           n706, Q => n4063, QN => n2139);
   REGISTERS_reg_22_23_inst : DFFR_X1 port map( D => n2881, CK => CLK, RN => 
                           n710, Q => n4118, QN => n1570);
   REGISTERS_reg_22_22_inst : DFFR_X1 port map( D => n2880, CK => CLK, RN => 
                           n710, Q => n4117, QN => n1595);
   REGISTERS_reg_22_21_inst : DFFR_X1 port map( D => n2879, CK => CLK, RN => 
                           n710, Q => n4116, QN => n1620);
   REGISTERS_reg_22_20_inst : DFFR_X1 port map( D => n2878, CK => CLK, RN => 
                           n710, Q => n4115, QN => n1645);
   REGISTERS_reg_22_19_inst : DFFR_X1 port map( D => n2877, CK => CLK, RN => 
                           n710, Q => n4114, QN => n1670);
   REGISTERS_reg_22_18_inst : DFFR_X1 port map( D => n2876, CK => CLK, RN => 
                           n710, Q => n4113, QN => n1695);
   REGISTERS_reg_22_17_inst : DFFR_X1 port map( D => n2875, CK => CLK, RN => 
                           n710, Q => n4112, QN => n1720);
   REGISTERS_reg_22_16_inst : DFFR_X1 port map( D => n2874, CK => CLK, RN => 
                           n710, Q => n4111, QN => n1745);
   REGISTERS_reg_22_15_inst : DFFR_X1 port map( D => n2873, CK => CLK, RN => 
                           n709, Q => n4110, QN => n1770);
   REGISTERS_reg_22_14_inst : DFFR_X1 port map( D => n2872, CK => CLK, RN => 
                           n709, Q => n4109, QN => n1795);
   REGISTERS_reg_22_13_inst : DFFR_X1 port map( D => n2871, CK => CLK, RN => 
                           n709, Q => n4108, QN => n1820);
   REGISTERS_reg_22_12_inst : DFFR_X1 port map( D => n2870, CK => CLK, RN => 
                           n709, Q => n4107, QN => n1845);
   REGISTERS_reg_22_11_inst : DFFR_X1 port map( D => n2869, CK => CLK, RN => 
                           n709, Q => n4106, QN => n1870);
   REGISTERS_reg_22_10_inst : DFFR_X1 port map( D => n2868, CK => CLK, RN => 
                           n709, Q => n4105, QN => n1895);
   REGISTERS_reg_22_9_inst : DFFR_X1 port map( D => n2867, CK => CLK, RN => 
                           n709, Q => n4104, QN => n1920);
   REGISTERS_reg_22_8_inst : DFFR_X1 port map( D => n2866, CK => CLK, RN => 
                           n709, Q => n4103, QN => n1945);
   REGISTERS_reg_22_7_inst : DFFR_X1 port map( D => n2865, CK => CLK, RN => 
                           n709, Q => n4102, QN => n1970);
   REGISTERS_reg_22_6_inst : DFFR_X1 port map( D => n2864, CK => CLK, RN => 
                           n709, Q => n4101, QN => n1995);
   REGISTERS_reg_22_5_inst : DFFR_X1 port map( D => n2863, CK => CLK, RN => 
                           n709, Q => n4100, QN => n2020);
   REGISTERS_reg_22_4_inst : DFFR_X1 port map( D => n2862, CK => CLK, RN => 
                           n709, Q => n4099, QN => n2045);
   REGISTERS_reg_22_3_inst : DFFR_X1 port map( D => n2861, CK => CLK, RN => 
                           n708, Q => n4098, QN => n2070);
   REGISTERS_reg_22_2_inst : DFFR_X1 port map( D => n2860, CK => CLK, RN => 
                           n708, Q => n4097, QN => n2095);
   REGISTERS_reg_22_1_inst : DFFR_X1 port map( D => n2859, CK => CLK, RN => 
                           n708, Q => n4096, QN => n2120);
   REGISTERS_reg_22_0_inst : DFFR_X1 port map( D => n2858, CK => CLK, RN => 
                           n708, Q => n4095, QN => n2155);
   REGISTERS_reg_11_23_inst : DFFR_X1 port map( D => n3233, CK => CLK, RN => 
                           n604, Q => n4278, QN => n_1802);
   REGISTERS_reg_11_22_inst : DFFR_X1 port map( D => n3232, CK => CLK, RN => 
                           n604, Q => n4277, QN => n_1803);
   REGISTERS_reg_11_21_inst : DFFR_X1 port map( D => n3231, CK => CLK, RN => 
                           n604, Q => n4276, QN => n_1804);
   REGISTERS_reg_11_20_inst : DFFR_X1 port map( D => n3230, CK => CLK, RN => 
                           n604, Q => n4275, QN => n_1805);
   REGISTERS_reg_11_19_inst : DFFR_X1 port map( D => n3229, CK => CLK, RN => 
                           n604, Q => n4274, QN => n_1806);
   REGISTERS_reg_11_18_inst : DFFR_X1 port map( D => n3228, CK => CLK, RN => 
                           n604, Q => n4273, QN => n_1807);
   REGISTERS_reg_11_17_inst : DFFR_X1 port map( D => n3227, CK => CLK, RN => 
                           n604, Q => n4272, QN => n_1808);
   REGISTERS_reg_11_16_inst : DFFR_X1 port map( D => n3226, CK => CLK, RN => 
                           n604, Q => n4271, QN => n_1809);
   REGISTERS_reg_11_15_inst : DFFR_X1 port map( D => n3225, CK => CLK, RN => 
                           n604, Q => n4270, QN => n_1810);
   REGISTERS_reg_11_14_inst : DFFR_X1 port map( D => n3224, CK => CLK, RN => 
                           n603, Q => n4269, QN => n_1811);
   REGISTERS_reg_11_13_inst : DFFR_X1 port map( D => n3223, CK => CLK, RN => 
                           n603, Q => n4268, QN => n_1812);
   REGISTERS_reg_11_12_inst : DFFR_X1 port map( D => n3222, CK => CLK, RN => 
                           n603, Q => n4267, QN => n_1813);
   REGISTERS_reg_11_11_inst : DFFR_X1 port map( D => n3221, CK => CLK, RN => 
                           n603, Q => n4266, QN => n_1814);
   REGISTERS_reg_11_10_inst : DFFR_X1 port map( D => n3220, CK => CLK, RN => 
                           n603, Q => n4265, QN => n_1815);
   REGISTERS_reg_11_9_inst : DFFR_X1 port map( D => n3219, CK => CLK, RN => 
                           n603, Q => n4264, QN => n_1816);
   REGISTERS_reg_11_8_inst : DFFR_X1 port map( D => n3218, CK => CLK, RN => 
                           n603, Q => n4263, QN => n_1817);
   REGISTERS_reg_11_7_inst : DFFR_X1 port map( D => n3217, CK => CLK, RN => 
                           n603, Q => n4262, QN => n_1818);
   REGISTERS_reg_11_6_inst : DFFR_X1 port map( D => n3216, CK => CLK, RN => 
                           n603, Q => n4261, QN => n_1819);
   REGISTERS_reg_11_5_inst : DFFR_X1 port map( D => n3215, CK => CLK, RN => 
                           n603, Q => n4260, QN => n_1820);
   REGISTERS_reg_11_4_inst : DFFR_X1 port map( D => n3214, CK => CLK, RN => 
                           n603, Q => n4259, QN => n_1821);
   REGISTERS_reg_11_3_inst : DFFR_X1 port map( D => n3213, CK => CLK, RN => 
                           n603, Q => n4258, QN => n_1822);
   REGISTERS_reg_11_2_inst : DFFR_X1 port map( D => n3212, CK => CLK, RN => 
                           n602, Q => n4257, QN => n_1823);
   REGISTERS_reg_11_1_inst : DFFR_X1 port map( D => n3211, CK => CLK, RN => 
                           n602, Q => n4256, QN => n_1824);
   REGISTERS_reg_11_0_inst : DFFR_X1 port map( D => n3210, CK => CLK, RN => 
                           n602, Q => n4255, QN => n_1825);
   REGISTERS_reg_10_23_inst : DFFR_X1 port map( D => n3265, CK => CLK, RN => 
                           n607, Q => n4310, QN => n_1826);
   REGISTERS_reg_10_22_inst : DFFR_X1 port map( D => n3264, CK => CLK, RN => 
                           n607, Q => n4309, QN => n_1827);
   REGISTERS_reg_10_21_inst : DFFR_X1 port map( D => n3263, CK => CLK, RN => 
                           n607, Q => n4308, QN => n_1828);
   REGISTERS_reg_10_20_inst : DFFR_X1 port map( D => n3262, CK => CLK, RN => 
                           n607, Q => n4307, QN => n_1829);
   REGISTERS_reg_10_19_inst : DFFR_X1 port map( D => n3261, CK => CLK, RN => 
                           n607, Q => n4306, QN => n_1830);
   REGISTERS_reg_10_18_inst : DFFR_X1 port map( D => n3260, CK => CLK, RN => 
                           n607, Q => n4305, QN => n_1831);
   REGISTERS_reg_10_17_inst : DFFR_X1 port map( D => n3259, CK => CLK, RN => 
                           n606, Q => n4304, QN => n_1832);
   REGISTERS_reg_10_16_inst : DFFR_X1 port map( D => n3258, CK => CLK, RN => 
                           n606, Q => n4303, QN => n_1833);
   REGISTERS_reg_10_15_inst : DFFR_X1 port map( D => n3257, CK => CLK, RN => 
                           n606, Q => n4302, QN => n_1834);
   REGISTERS_reg_10_14_inst : DFFR_X1 port map( D => n3256, CK => CLK, RN => 
                           n606, Q => n4301, QN => n_1835);
   REGISTERS_reg_10_13_inst : DFFR_X1 port map( D => n3255, CK => CLK, RN => 
                           n606, Q => n4300, QN => n_1836);
   REGISTERS_reg_10_12_inst : DFFR_X1 port map( D => n3254, CK => CLK, RN => 
                           n606, Q => n4299, QN => n_1837);
   REGISTERS_reg_10_11_inst : DFFR_X1 port map( D => n3253, CK => CLK, RN => 
                           n606, Q => n4298, QN => n_1838);
   REGISTERS_reg_10_10_inst : DFFR_X1 port map( D => n3252, CK => CLK, RN => 
                           n606, Q => n4297, QN => n_1839);
   REGISTERS_reg_10_9_inst : DFFR_X1 port map( D => n3251, CK => CLK, RN => 
                           n606, Q => n4296, QN => n_1840);
   REGISTERS_reg_10_8_inst : DFFR_X1 port map( D => n3250, CK => CLK, RN => 
                           n606, Q => n4295, QN => n_1841);
   REGISTERS_reg_10_7_inst : DFFR_X1 port map( D => n3249, CK => CLK, RN => 
                           n606, Q => n4294, QN => n_1842);
   REGISTERS_reg_10_6_inst : DFFR_X1 port map( D => n3248, CK => CLK, RN => 
                           n605, Q => n4293, QN => n_1843);
   REGISTERS_reg_10_5_inst : DFFR_X1 port map( D => n3247, CK => CLK, RN => 
                           n605, Q => n4292, QN => n_1844);
   REGISTERS_reg_10_4_inst : DFFR_X1 port map( D => n3246, CK => CLK, RN => 
                           n605, Q => n4291, QN => n_1845);
   REGISTERS_reg_10_3_inst : DFFR_X1 port map( D => n3245, CK => CLK, RN => 
                           n605, Q => n4290, QN => n_1846);
   REGISTERS_reg_10_2_inst : DFFR_X1 port map( D => n3244, CK => CLK, RN => 
                           n605, Q => n4289, QN => n_1847);
   REGISTERS_reg_10_1_inst : DFFR_X1 port map( D => n3243, CK => CLK, RN => 
                           n605, Q => n4288, QN => n_1848);
   REGISTERS_reg_10_0_inst : DFFR_X1 port map( D => n3242, CK => CLK, RN => 
                           n605, Q => n4287, QN => n_1849);
   REGISTERS_reg_19_23_inst : DFFR_X1 port map( D => n2977, CK => CLK, RN => 
                           n698, Q => n4150, QN => n_1850);
   REGISTERS_reg_19_22_inst : DFFR_X1 port map( D => n2976, CK => CLK, RN => 
                           n697, Q => n4149, QN => n_1851);
   REGISTERS_reg_19_21_inst : DFFR_X1 port map( D => n2975, CK => CLK, RN => 
                           n697, Q => n4148, QN => n_1852);
   REGISTERS_reg_19_20_inst : DFFR_X1 port map( D => n2974, CK => CLK, RN => 
                           n697, Q => n4147, QN => n_1853);
   REGISTERS_reg_19_19_inst : DFFR_X1 port map( D => n2973, CK => CLK, RN => 
                           n697, Q => n4146, QN => n_1854);
   REGISTERS_reg_19_18_inst : DFFR_X1 port map( D => n2972, CK => CLK, RN => 
                           n697, Q => n4145, QN => n_1855);
   REGISTERS_reg_19_17_inst : DFFR_X1 port map( D => n2971, CK => CLK, RN => 
                           n697, Q => n4144, QN => n_1856);
   REGISTERS_reg_19_16_inst : DFFR_X1 port map( D => n2970, CK => CLK, RN => 
                           n697, Q => n4143, QN => n_1857);
   REGISTERS_reg_19_15_inst : DFFR_X1 port map( D => n2969, CK => CLK, RN => 
                           n697, Q => n4142, QN => n_1858);
   REGISTERS_reg_19_14_inst : DFFR_X1 port map( D => n2968, CK => CLK, RN => 
                           n697, Q => n4141, QN => n_1859);
   REGISTERS_reg_19_13_inst : DFFR_X1 port map( D => n2967, CK => CLK, RN => 
                           n697, Q => n4140, QN => n_1860);
   REGISTERS_reg_19_12_inst : DFFR_X1 port map( D => n2966, CK => CLK, RN => 
                           n697, Q => n4139, QN => n_1861);
   REGISTERS_reg_19_11_inst : DFFR_X1 port map( D => n2965, CK => CLK, RN => 
                           n697, Q => n4138, QN => n_1862);
   REGISTERS_reg_19_10_inst : DFFR_X1 port map( D => n2964, CK => CLK, RN => 
                           n696, Q => n4137, QN => n_1863);
   REGISTERS_reg_19_9_inst : DFFR_X1 port map( D => n2963, CK => CLK, RN => 
                           n696, Q => n4136, QN => n_1864);
   REGISTERS_reg_19_8_inst : DFFR_X1 port map( D => n2962, CK => CLK, RN => 
                           n696, Q => n4135, QN => n_1865);
   REGISTERS_reg_19_7_inst : DFFR_X1 port map( D => n2961, CK => CLK, RN => 
                           n696, Q => n4134, QN => n_1866);
   REGISTERS_reg_19_6_inst : DFFR_X1 port map( D => n2960, CK => CLK, RN => 
                           n696, Q => n4133, QN => n_1867);
   REGISTERS_reg_19_5_inst : DFFR_X1 port map( D => n2959, CK => CLK, RN => 
                           n696, Q => n4132, QN => n_1868);
   REGISTERS_reg_19_4_inst : DFFR_X1 port map( D => n2958, CK => CLK, RN => 
                           n696, Q => n4131, QN => n_1869);
   REGISTERS_reg_19_3_inst : DFFR_X1 port map( D => n2957, CK => CLK, RN => 
                           n696, Q => n4130, QN => n_1870);
   REGISTERS_reg_19_2_inst : DFFR_X1 port map( D => n2956, CK => CLK, RN => 
                           n696, Q => n4129, QN => n_1871);
   REGISTERS_reg_19_1_inst : DFFR_X1 port map( D => n2955, CK => CLK, RN => 
                           n696, Q => n4128, QN => n_1872);
   REGISTERS_reg_19_0_inst : DFFR_X1 port map( D => n2954, CK => CLK, RN => 
                           n696, Q => n4127, QN => n_1873);
   REGISTERS_reg_18_23_inst : DFFR_X1 port map( D => n3009, CK => CLK, RN => 
                           n700, Q => n4182, QN => n_1874);
   REGISTERS_reg_18_22_inst : DFFR_X1 port map( D => n3008, CK => CLK, RN => 
                           n700, Q => n4181, QN => n_1875);
   REGISTERS_reg_18_21_inst : DFFR_X1 port map( D => n3007, CK => CLK, RN => 
                           n700, Q => n4180, QN => n_1876);
   REGISTERS_reg_18_20_inst : DFFR_X1 port map( D => n3006, CK => CLK, RN => 
                           n700, Q => n4179, QN => n_1877);
   REGISTERS_reg_18_19_inst : DFFR_X1 port map( D => n3005, CK => CLK, RN => 
                           n700, Q => n4178, QN => n_1878);
   REGISTERS_reg_18_18_inst : DFFR_X1 port map( D => n3004, CK => CLK, RN => 
                           n700, Q => n4177, QN => n_1879);
   REGISTERS_reg_18_17_inst : DFFR_X1 port map( D => n3003, CK => CLK, RN => 
                           n700, Q => n4176, QN => n_1880);
   REGISTERS_reg_18_16_inst : DFFR_X1 port map( D => n3002, CK => CLK, RN => 
                           n700, Q => n4175, QN => n_1881);
   REGISTERS_reg_18_15_inst : DFFR_X1 port map( D => n3001, CK => CLK, RN => 
                           n700, Q => n4174, QN => n_1882);
   REGISTERS_reg_18_14_inst : DFFR_X1 port map( D => n3000, CK => CLK, RN => 
                           n699, Q => n4173, QN => n_1883);
   REGISTERS_reg_18_13_inst : DFFR_X1 port map( D => n2999, CK => CLK, RN => 
                           n699, Q => n4172, QN => n_1884);
   REGISTERS_reg_18_12_inst : DFFR_X1 port map( D => n2998, CK => CLK, RN => 
                           n699, Q => n4171, QN => n_1885);
   REGISTERS_reg_18_11_inst : DFFR_X1 port map( D => n2997, CK => CLK, RN => 
                           n699, Q => n4170, QN => n_1886);
   REGISTERS_reg_18_10_inst : DFFR_X1 port map( D => n2996, CK => CLK, RN => 
                           n699, Q => n4169, QN => n_1887);
   REGISTERS_reg_18_9_inst : DFFR_X1 port map( D => n2995, CK => CLK, RN => 
                           n699, Q => n4168, QN => n_1888);
   REGISTERS_reg_18_8_inst : DFFR_X1 port map( D => n2994, CK => CLK, RN => 
                           n699, Q => n4167, QN => n_1889);
   REGISTERS_reg_18_7_inst : DFFR_X1 port map( D => n2993, CK => CLK, RN => 
                           n699, Q => n4166, QN => n_1890);
   REGISTERS_reg_18_6_inst : DFFR_X1 port map( D => n2992, CK => CLK, RN => 
                           n699, Q => n4165, QN => n_1891);
   REGISTERS_reg_18_5_inst : DFFR_X1 port map( D => n2991, CK => CLK, RN => 
                           n699, Q => n4164, QN => n_1892);
   REGISTERS_reg_18_4_inst : DFFR_X1 port map( D => n2990, CK => CLK, RN => 
                           n699, Q => n4163, QN => n_1893);
   REGISTERS_reg_18_3_inst : DFFR_X1 port map( D => n2989, CK => CLK, RN => 
                           n699, Q => n4162, QN => n_1894);
   REGISTERS_reg_18_2_inst : DFFR_X1 port map( D => n2988, CK => CLK, RN => 
                           n698, Q => n4161, QN => n_1895);
   REGISTERS_reg_18_1_inst : DFFR_X1 port map( D => n2987, CK => CLK, RN => 
                           n698, Q => n4160, QN => n_1896);
   REGISTERS_reg_18_0_inst : DFFR_X1 port map( D => n2986, CK => CLK, RN => 
                           n698, Q => n4159, QN => n_1897);
   REGISTERS_reg_29_23_inst : DFFR_X1 port map( D => n2657, CK => CLK, RN => 
                           n692, Q => n3958, QN => n_1898);
   REGISTERS_reg_29_22_inst : DFFR_X1 port map( D => n2656, CK => CLK, RN => 
                           n691, Q => n3957, QN => n_1899);
   REGISTERS_reg_29_21_inst : DFFR_X1 port map( D => n2655, CK => CLK, RN => 
                           n691, Q => n3956, QN => n_1900);
   REGISTERS_reg_29_20_inst : DFFR_X1 port map( D => n2654, CK => CLK, RN => 
                           n691, Q => n3955, QN => n_1901);
   REGISTERS_reg_29_19_inst : DFFR_X1 port map( D => n2653, CK => CLK, RN => 
                           n691, Q => n3954, QN => n_1902);
   REGISTERS_reg_29_18_inst : DFFR_X1 port map( D => n2652, CK => CLK, RN => 
                           n691, Q => n3953, QN => n_1903);
   REGISTERS_reg_29_17_inst : DFFR_X1 port map( D => n2651, CK => CLK, RN => 
                           n691, Q => n3952, QN => n_1904);
   REGISTERS_reg_29_16_inst : DFFR_X1 port map( D => n2650, CK => CLK, RN => 
                           n691, Q => n3951, QN => n_1905);
   REGISTERS_reg_29_15_inst : DFFR_X1 port map( D => n2649, CK => CLK, RN => 
                           n691, Q => n3950, QN => n_1906);
   REGISTERS_reg_29_14_inst : DFFR_X1 port map( D => n2648, CK => CLK, RN => 
                           n691, Q => n3949, QN => n_1907);
   REGISTERS_reg_29_13_inst : DFFR_X1 port map( D => n2647, CK => CLK, RN => 
                           n691, Q => n3948, QN => n_1908);
   REGISTERS_reg_29_12_inst : DFFR_X1 port map( D => n2646, CK => CLK, RN => 
                           n691, Q => n3947, QN => n_1909);
   REGISTERS_reg_29_11_inst : DFFR_X1 port map( D => n2645, CK => CLK, RN => 
                           n691, Q => n3946, QN => n_1910);
   REGISTERS_reg_29_10_inst : DFFR_X1 port map( D => n2644, CK => CLK, RN => 
                           n690, Q => n3945, QN => n_1911);
   REGISTERS_reg_29_9_inst : DFFR_X1 port map( D => n2643, CK => CLK, RN => 
                           n690, Q => n3944, QN => n_1912);
   REGISTERS_reg_29_8_inst : DFFR_X1 port map( D => n2642, CK => CLK, RN => 
                           n690, Q => n3943, QN => n_1913);
   REGISTERS_reg_29_7_inst : DFFR_X1 port map( D => n2641, CK => CLK, RN => 
                           n690, Q => n3942, QN => n_1914);
   REGISTERS_reg_29_6_inst : DFFR_X1 port map( D => n2640, CK => CLK, RN => 
                           n690, Q => n3941, QN => n_1915);
   REGISTERS_reg_29_5_inst : DFFR_X1 port map( D => n2639, CK => CLK, RN => 
                           n690, Q => n3940, QN => n_1916);
   REGISTERS_reg_29_4_inst : DFFR_X1 port map( D => n2638, CK => CLK, RN => 
                           n690, Q => n3939, QN => n_1917);
   REGISTERS_reg_29_3_inst : DFFR_X1 port map( D => n2637, CK => CLK, RN => 
                           n690, Q => n3938, QN => n_1918);
   REGISTERS_reg_29_2_inst : DFFR_X1 port map( D => n2636, CK => CLK, RN => 
                           n690, Q => n3937, QN => n_1919);
   REGISTERS_reg_29_1_inst : DFFR_X1 port map( D => n2635, CK => CLK, RN => 
                           n690, Q => n3936, QN => n_1920);
   REGISTERS_reg_29_0_inst : DFFR_X1 port map( D => n2634, CK => CLK, RN => 
                           n690, Q => n3935, QN => n_1921);
   REGISTERS_reg_28_23_inst : DFFR_X1 port map( D => n2689, CK => CLK, RN => 
                           n694, Q => n3990, QN => n1565);
   REGISTERS_reg_28_22_inst : DFFR_X1 port map( D => n2688, CK => CLK, RN => 
                           n694, Q => n3989, QN => n1590);
   REGISTERS_reg_28_21_inst : DFFR_X1 port map( D => n2687, CK => CLK, RN => 
                           n694, Q => n3988, QN => n1615);
   REGISTERS_reg_28_20_inst : DFFR_X1 port map( D => n2686, CK => CLK, RN => 
                           n694, Q => n3987, QN => n1640);
   REGISTERS_reg_28_19_inst : DFFR_X1 port map( D => n2685, CK => CLK, RN => 
                           n694, Q => n3986, QN => n1665);
   REGISTERS_reg_28_18_inst : DFFR_X1 port map( D => n2684, CK => CLK, RN => 
                           n694, Q => n3985, QN => n1690);
   REGISTERS_reg_28_17_inst : DFFR_X1 port map( D => n2683, CK => CLK, RN => 
                           n694, Q => n3984, QN => n1715);
   REGISTERS_reg_28_16_inst : DFFR_X1 port map( D => n2682, CK => CLK, RN => 
                           n694, Q => n3983, QN => n1740);
   REGISTERS_reg_28_15_inst : DFFR_X1 port map( D => n2681, CK => CLK, RN => 
                           n694, Q => n3982, QN => n1765);
   REGISTERS_reg_28_14_inst : DFFR_X1 port map( D => n2680, CK => CLK, RN => 
                           n693, Q => n3981, QN => n1790);
   REGISTERS_reg_28_13_inst : DFFR_X1 port map( D => n2679, CK => CLK, RN => 
                           n693, Q => n3980, QN => n1815);
   REGISTERS_reg_28_12_inst : DFFR_X1 port map( D => n2678, CK => CLK, RN => 
                           n693, Q => n3979, QN => n1840);
   REGISTERS_reg_28_11_inst : DFFR_X1 port map( D => n2677, CK => CLK, RN => 
                           n693, Q => n3978, QN => n1865);
   REGISTERS_reg_28_10_inst : DFFR_X1 port map( D => n2676, CK => CLK, RN => 
                           n693, Q => n3977, QN => n1890);
   REGISTERS_reg_28_9_inst : DFFR_X1 port map( D => n2675, CK => CLK, RN => 
                           n693, Q => n3976, QN => n1915);
   REGISTERS_reg_28_8_inst : DFFR_X1 port map( D => n2674, CK => CLK, RN => 
                           n693, Q => n3975, QN => n1940);
   REGISTERS_reg_28_7_inst : DFFR_X1 port map( D => n2673, CK => CLK, RN => 
                           n693, Q => n3974, QN => n1965);
   REGISTERS_reg_28_6_inst : DFFR_X1 port map( D => n2672, CK => CLK, RN => 
                           n693, Q => n3973, QN => n1990);
   REGISTERS_reg_28_5_inst : DFFR_X1 port map( D => n2671, CK => CLK, RN => 
                           n693, Q => n3972, QN => n2015);
   REGISTERS_reg_28_4_inst : DFFR_X1 port map( D => n2670, CK => CLK, RN => 
                           n693, Q => n3971, QN => n2040);
   REGISTERS_reg_28_3_inst : DFFR_X1 port map( D => n2669, CK => CLK, RN => 
                           n693, Q => n3970, QN => n2065);
   REGISTERS_reg_28_2_inst : DFFR_X1 port map( D => n2668, CK => CLK, RN => 
                           n692, Q => n3969, QN => n2090);
   REGISTERS_reg_28_1_inst : DFFR_X1 port map( D => n2667, CK => CLK, RN => 
                           n692, Q => n3968, QN => n2115);
   REGISTERS_reg_28_0_inst : DFFR_X1 port map( D => n2666, CK => CLK, RN => 
                           n692, Q => n3967, QN => n2147);
   REGISTERS_reg_25_23_inst : DFFR_X1 port map( D => n2785, CK => CLK, RN => 
                           n682, Q => n4022, QN => n_1922);
   REGISTERS_reg_25_22_inst : DFFR_X1 port map( D => n2784, CK => CLK, RN => 
                           n681, Q => n4021, QN => n_1923);
   REGISTERS_reg_25_21_inst : DFFR_X1 port map( D => n2783, CK => CLK, RN => 
                           n681, Q => n4020, QN => n_1924);
   REGISTERS_reg_25_20_inst : DFFR_X1 port map( D => n2782, CK => CLK, RN => 
                           n681, Q => n4019, QN => n_1925);
   REGISTERS_reg_25_19_inst : DFFR_X1 port map( D => n2781, CK => CLK, RN => 
                           n681, Q => n4018, QN => n_1926);
   REGISTERS_reg_25_18_inst : DFFR_X1 port map( D => n2780, CK => CLK, RN => 
                           n681, Q => n4017, QN => n_1927);
   REGISTERS_reg_25_17_inst : DFFR_X1 port map( D => n2779, CK => CLK, RN => 
                           n681, Q => n4016, QN => n_1928);
   REGISTERS_reg_25_16_inst : DFFR_X1 port map( D => n2778, CK => CLK, RN => 
                           n681, Q => n4015, QN => n_1929);
   REGISTERS_reg_25_15_inst : DFFR_X1 port map( D => n2777, CK => CLK, RN => 
                           n681, Q => n4014, QN => n_1930);
   REGISTERS_reg_25_14_inst : DFFR_X1 port map( D => n2776, CK => CLK, RN => 
                           n681, Q => n4013, QN => n_1931);
   REGISTERS_reg_25_13_inst : DFFR_X1 port map( D => n2775, CK => CLK, RN => 
                           n681, Q => n4012, QN => n_1932);
   REGISTERS_reg_25_12_inst : DFFR_X1 port map( D => n2774, CK => CLK, RN => 
                           n681, Q => n4011, QN => n_1933);
   REGISTERS_reg_25_11_inst : DFFR_X1 port map( D => n2773, CK => CLK, RN => 
                           n681, Q => n4010, QN => n_1934);
   REGISTERS_reg_25_10_inst : DFFR_X1 port map( D => n2772, CK => CLK, RN => 
                           n680, Q => n4009, QN => n_1935);
   REGISTERS_reg_25_9_inst : DFFR_X1 port map( D => n2771, CK => CLK, RN => 
                           n680, Q => n4008, QN => n_1936);
   REGISTERS_reg_25_8_inst : DFFR_X1 port map( D => n2770, CK => CLK, RN => 
                           n680, Q => n4007, QN => n_1937);
   REGISTERS_reg_25_7_inst : DFFR_X1 port map( D => n2769, CK => CLK, RN => 
                           n680, Q => n4006, QN => n_1938);
   REGISTERS_reg_25_6_inst : DFFR_X1 port map( D => n2768, CK => CLK, RN => 
                           n680, Q => n4005, QN => n_1939);
   REGISTERS_reg_25_5_inst : DFFR_X1 port map( D => n2767, CK => CLK, RN => 
                           n680, Q => n4004, QN => n_1940);
   REGISTERS_reg_25_4_inst : DFFR_X1 port map( D => n2766, CK => CLK, RN => 
                           n680, Q => n4003, QN => n_1941);
   REGISTERS_reg_25_3_inst : DFFR_X1 port map( D => n2765, CK => CLK, RN => 
                           n680, Q => n4002, QN => n_1942);
   REGISTERS_reg_25_2_inst : DFFR_X1 port map( D => n2764, CK => CLK, RN => 
                           n680, Q => n4001, QN => n_1943);
   REGISTERS_reg_25_1_inst : DFFR_X1 port map( D => n2763, CK => CLK, RN => 
                           n680, Q => n4000, QN => n_1944);
   REGISTERS_reg_25_0_inst : DFFR_X1 port map( D => n2762, CK => CLK, RN => 
                           n680, Q => n3999, QN => n_1945);
   REGISTERS_reg_24_23_inst : DFFR_X1 port map( D => n2817, CK => CLK, RN => 
                           n684, Q => n4054, QN => n_1946);
   REGISTERS_reg_24_22_inst : DFFR_X1 port map( D => n2816, CK => CLK, RN => 
                           n684, Q => n4053, QN => n_1947);
   REGISTERS_reg_24_21_inst : DFFR_X1 port map( D => n2815, CK => CLK, RN => 
                           n684, Q => n4052, QN => n_1948);
   REGISTERS_reg_24_20_inst : DFFR_X1 port map( D => n2814, CK => CLK, RN => 
                           n684, Q => n4051, QN => n_1949);
   REGISTERS_reg_24_19_inst : DFFR_X1 port map( D => n2813, CK => CLK, RN => 
                           n684, Q => n4050, QN => n_1950);
   REGISTERS_reg_24_18_inst : DFFR_X1 port map( D => n2812, CK => CLK, RN => 
                           n684, Q => n4049, QN => n_1951);
   REGISTERS_reg_24_17_inst : DFFR_X1 port map( D => n2811, CK => CLK, RN => 
                           n684, Q => n4048, QN => n_1952);
   REGISTERS_reg_24_16_inst : DFFR_X1 port map( D => n2810, CK => CLK, RN => 
                           n684, Q => n4047, QN => n_1953);
   REGISTERS_reg_24_15_inst : DFFR_X1 port map( D => n2809, CK => CLK, RN => 
                           n684, Q => n4046, QN => n_1954);
   REGISTERS_reg_24_14_inst : DFFR_X1 port map( D => n2808, CK => CLK, RN => 
                           n683, Q => n4045, QN => n_1955);
   REGISTERS_reg_24_13_inst : DFFR_X1 port map( D => n2807, CK => CLK, RN => 
                           n683, Q => n4044, QN => n_1956);
   REGISTERS_reg_24_12_inst : DFFR_X1 port map( D => n2806, CK => CLK, RN => 
                           n683, Q => n4043, QN => n_1957);
   REGISTERS_reg_24_11_inst : DFFR_X1 port map( D => n2805, CK => CLK, RN => 
                           n683, Q => n4042, QN => n_1958);
   REGISTERS_reg_24_10_inst : DFFR_X1 port map( D => n2804, CK => CLK, RN => 
                           n683, Q => n4041, QN => n_1959);
   REGISTERS_reg_24_9_inst : DFFR_X1 port map( D => n2803, CK => CLK, RN => 
                           n683, Q => n4040, QN => n_1960);
   REGISTERS_reg_24_8_inst : DFFR_X1 port map( D => n2802, CK => CLK, RN => 
                           n683, Q => n4039, QN => n_1961);
   REGISTERS_reg_24_7_inst : DFFR_X1 port map( D => n2801, CK => CLK, RN => 
                           n683, Q => n4038, QN => n_1962);
   REGISTERS_reg_24_6_inst : DFFR_X1 port map( D => n2800, CK => CLK, RN => 
                           n683, Q => n4037, QN => n_1963);
   REGISTERS_reg_24_5_inst : DFFR_X1 port map( D => n2799, CK => CLK, RN => 
                           n683, Q => n4036, QN => n_1964);
   REGISTERS_reg_24_4_inst : DFFR_X1 port map( D => n2798, CK => CLK, RN => 
                           n683, Q => n4035, QN => n_1965);
   OUT1_reg_8_inst : DFF_X1 port map( D => n2514, CK => CLK, Q => OUT1(8), QN 
                           => n3879);
   OUT1_reg_2_inst : DFF_X1 port map( D => n2508, CK => CLK, Q => OUT1(2), QN 
                           => n3873);
   OUT1_reg_13_inst : DFF_X1 port map( D => n2519, CK => CLK, Q => OUT1(13), QN
                           => n3884);
   OUT1_reg_12_inst : DFF_X1 port map( D => n2518, CK => CLK, Q => OUT1(12), QN
                           => n3883);
   OUT1_reg_9_inst : DFF_X1 port map( D => n2515, CK => CLK, Q => OUT1(9), QN 
                           => n3880);
   OUT1_reg_4_inst : DFF_X1 port map( D => n2510, CK => CLK, Q => OUT1(4), QN 
                           => n3875);
   OUT1_reg_3_inst : DFF_X1 port map( D => n2509, CK => CLK, Q => OUT1(3), QN 
                           => n3874);
   OUT1_reg_1_inst : DFF_X1 port map( D => n2507, CK => CLK, Q => OUT1(1), QN 
                           => n3872);
   OUT1_reg_17_inst : DFF_X1 port map( D => n2523, CK => CLK, Q => OUT1(17), QN
                           => n3888);
   OUT1_reg_16_inst : DFF_X1 port map( D => n2522, CK => CLK, Q => OUT1(16), QN
                           => n3887);
   OUT1_reg_15_inst : DFF_X1 port map( D => n2521, CK => CLK, Q => OUT1(15), QN
                           => n3886);
   OUT1_reg_14_inst : DFF_X1 port map( D => n2520, CK => CLK, Q => OUT1(14), QN
                           => n3885);
   OUT2_reg_10_inst : DFF_X1 port map( D => n2548, CK => CLK, Q => OUT2(10), QN
                           => n3913);
   OUT2_reg_8_inst : DFF_X1 port map( D => n2546, CK => CLK, Q => OUT2(8), QN 
                           => n3911);
   OUT2_reg_6_inst : DFF_X1 port map( D => n2544, CK => CLK, Q => OUT2(6), QN 
                           => n3909);
   OUT2_reg_4_inst : DFF_X1 port map( D => n2542, CK => CLK, Q => OUT2(4), QN 
                           => n3907);
   OUT2_reg_22_inst : DFF_X1 port map( D => n2560, CK => CLK, Q => OUT2(22), QN
                           => n3925);
   OUT2_reg_20_inst : DFF_X1 port map( D => n2558, CK => CLK, Q => OUT2(20), QN
                           => n3923);
   OUT2_reg_18_inst : DFF_X1 port map( D => n2556, CK => CLK, Q => OUT2(18), QN
                           => n3921);
   OUT2_reg_16_inst : DFF_X1 port map( D => n2554, CK => CLK, Q => OUT2(16), QN
                           => n3919);
   OUT2_reg_14_inst : DFF_X1 port map( D => n2552, CK => CLK, Q => OUT2(14), QN
                           => n3917);
   OUT2_reg_12_inst : DFF_X1 port map( D => n2550, CK => CLK, Q => OUT2(12), QN
                           => n3915);
   OUT1_reg_0_inst : DFF_X1 port map( D => n2506, CK => CLK, Q => OUT1(0), QN 
                           => n3871);
   OUT1_reg_31_inst : DFF_X1 port map( D => n2537, CK => CLK, Q => OUT1(31), QN
                           => n3902);
   OUT1_reg_30_inst : DFF_X1 port map( D => n2536, CK => CLK, Q => OUT1(30), QN
                           => n3901);
   OUT1_reg_29_inst : DFF_X1 port map( D => n2535, CK => CLK, Q => OUT1(29), QN
                           => n3900);
   OUT1_reg_28_inst : DFF_X1 port map( D => n2534, CK => CLK, Q => OUT1(28), QN
                           => n3899);
   OUT1_reg_27_inst : DFF_X1 port map( D => n2533, CK => CLK, Q => OUT1(27), QN
                           => n3898);
   OUT1_reg_26_inst : DFF_X1 port map( D => n2532, CK => CLK, Q => OUT1(26), QN
                           => n3897);
   OUT1_reg_25_inst : DFF_X1 port map( D => n2531, CK => CLK, Q => OUT1(25), QN
                           => n3896);
   OUT1_reg_24_inst : DFF_X1 port map( D => n2530, CK => CLK, Q => OUT1(24), QN
                           => n3895);
   OUT1_reg_6_inst : DFF_X1 port map( D => n2512, CK => CLK, Q => OUT1(6), QN 
                           => n3877);
   OUT1_reg_5_inst : DFF_X1 port map( D => n2511, CK => CLK, Q => OUT1(5), QN 
                           => n3876);
   OUT2_reg_0_inst : DFF_X1 port map( D => n2538, CK => CLK, Q => OUT2(0), QN 
                           => n3903);
   OUT2_reg_1_inst : DFF_X1 port map( D => n2539, CK => CLK, Q => OUT2(1), QN 
                           => n3904);
   OUT2_reg_2_inst : DFF_X1 port map( D => n2540, CK => CLK, Q => OUT2(2), QN 
                           => n3905);
   OUT1_reg_23_inst : DFF_X1 port map( D => n2529, CK => CLK, Q => OUT1(23), QN
                           => n3894);
   OUT1_reg_22_inst : DFF_X1 port map( D => n2528, CK => CLK, Q => OUT1(22), QN
                           => n3893);
   OUT1_reg_21_inst : DFF_X1 port map( D => n2527, CK => CLK, Q => OUT1(21), QN
                           => n3892);
   OUT1_reg_20_inst : DFF_X1 port map( D => n2526, CK => CLK, Q => OUT1(20), QN
                           => n3891);
   OUT1_reg_19_inst : DFF_X1 port map( D => n2525, CK => CLK, Q => OUT1(19), QN
                           => n3890);
   OUT1_reg_18_inst : DFF_X1 port map( D => n2524, CK => CLK, Q => OUT1(18), QN
                           => n3889);
   OUT1_reg_11_inst : DFF_X1 port map( D => n2517, CK => CLK, Q => OUT1(11), QN
                           => n3882);
   OUT1_reg_10_inst : DFF_X1 port map( D => n2516, CK => CLK, Q => OUT1(10), QN
                           => n3881);
   OUT1_reg_7_inst : DFF_X1 port map( D => n2513, CK => CLK, Q => OUT1(7), QN 
                           => n3878);
   OUT2_reg_19_inst : DFF_X1 port map( D => n2557, CK => CLK, Q => OUT2(19), QN
                           => n3922);
   OUT2_reg_17_inst : DFF_X1 port map( D => n2555, CK => CLK, Q => OUT2(17), QN
                           => n3920);
   OUT2_reg_15_inst : DFF_X1 port map( D => n2553, CK => CLK, Q => OUT2(15), QN
                           => n3918);
   OUT2_reg_23_inst : DFF_X1 port map( D => n2561, CK => CLK, Q => OUT2(23), QN
                           => n3926);
   OUT2_reg_21_inst : DFF_X1 port map( D => n2559, CK => CLK, Q => OUT2(21), QN
                           => n3924);
   OUT2_reg_13_inst : DFF_X1 port map( D => n2551, CK => CLK, Q => OUT2(13), QN
                           => n3916);
   OUT2_reg_9_inst : DFF_X1 port map( D => n2547, CK => CLK, Q => OUT2(9), QN 
                           => n3912);
   OUT2_reg_7_inst : DFF_X1 port map( D => n2545, CK => CLK, Q => OUT2(7), QN 
                           => n3910);
   OUT2_reg_5_inst : DFF_X1 port map( D => n2543, CK => CLK, Q => OUT2(5), QN 
                           => n3908);
   OUT2_reg_31_inst : DFF_X1 port map( D => n2569, CK => CLK, Q => OUT2(31), QN
                           => n3934);
   OUT2_reg_30_inst : DFF_X1 port map( D => n2568, CK => CLK, Q => OUT2(30), QN
                           => n3933);
   OUT2_reg_29_inst : DFF_X1 port map( D => n2567, CK => CLK, Q => OUT2(29), QN
                           => n3932);
   OUT2_reg_28_inst : DFF_X1 port map( D => n2566, CK => CLK, Q => OUT2(28), QN
                           => n3931);
   OUT2_reg_27_inst : DFF_X1 port map( D => n2565, CK => CLK, Q => OUT2(27), QN
                           => n3930);
   OUT2_reg_26_inst : DFF_X1 port map( D => n2564, CK => CLK, Q => OUT2(26), QN
                           => n3929);
   OUT2_reg_25_inst : DFF_X1 port map( D => n2563, CK => CLK, Q => OUT2(25), QN
                           => n3928);
   OUT2_reg_24_inst : DFF_X1 port map( D => n2562, CK => CLK, Q => OUT2(24), QN
                           => n3927);
   OUT2_reg_11_inst : DFF_X1 port map( D => n2549, CK => CLK, Q => OUT2(11), QN
                           => n3914);
   OUT2_reg_3_inst : DFF_X2 port map( D => n2541, CK => CLK, Q => OUT2(3), QN 
                           => n3906);
   U2 : CLKBUF_X1 port map( A => ADD_RS2(0), Z => n1);
   U3 : NOR3_X1 port map( A1 => ADD_RS1(0), A2 => ADD_RS1(3), A3 => n56, ZN => 
                           n2);
   U4 : CLKBUF_X1 port map( A => n3858, Z => n3);
   U5 : BUF_X2 port map( A => n1354, Z => n323);
   U6 : BUF_X2 port map( A => n1353, Z => n320);
   U7 : BUF_X2 port map( A => n1347, Z => n309);
   U8 : BUF_X2 port map( A => n1354, Z => n322);
   U9 : BUF_X2 port map( A => n1353, Z => n319);
   U10 : BUF_X2 port map( A => n1350, Z => n315);
   U11 : BUF_X2 port map( A => n1352, Z => n318);
   U12 : BUF_X2 port map( A => n1343, Z => n302);
   U13 : BUF_X2 port map( A => n1343, Z => n301);
   U14 : OAI211_X1 port map( C1 => n535, C2 => n305, A => n1817, B => n1818, ZN
                           => n1810);
   U15 : OAI211_X1 port map( C1 => n547, C2 => n304, A => n2117, B => n2118, ZN
                           => n2110);
   U16 : BUF_X1 port map( A => n2195, Z => n457);
   U17 : CLKBUF_X1 port map( A => ADD_RS2(1), Z => n4);
   U18 : BUF_X2 port map( A => n1367, Z => n342);
   U19 : BUF_X2 port map( A => n1367, Z => n33);
   U20 : BUF_X2 port map( A => n1367, Z => n34);
   U21 : BUF_X2 port map( A => n1367, Z => n341);
   U22 : BUF_X2 port map( A => n1367, Z => n340);
   U23 : CLKBUF_X3 port map( A => n1382, Z => n5);
   U24 : BUF_X2 port map( A => n1369, Z => n346);
   U25 : BUF_X2 port map( A => n1369, Z => n347);
   U26 : CLKBUF_X3 port map( A => n1375, Z => n356);
   U27 : OR2_X1 port map( A1 => n1812, A2 => n1811, ZN => n6);
   U28 : OR2_X1 port map( A1 => n2470, A2 => n2471, ZN => n7);
   U29 : OR2_X1 port map( A1 => n2489, A2 => n2488, ZN => n8);
   U30 : OR2_X1 port map( A1 => n3725, A2 => n3724, ZN => n9);
   U31 : OR2_X1 port map( A1 => n3563, A2 => n3562, ZN => n10);
   U32 : OR2_X1 port map( A1 => n3743, A2 => n3742, ZN => n11);
   U33 : OR2_X1 port map( A1 => n3581, A2 => n3580, ZN => n12);
   U34 : OR2_X1 port map( A1 => n2061, A2 => n2062, ZN => n13);
   U35 : OR2_X1 port map( A1 => n3599, A2 => n3598, ZN => n14);
   U36 : OR2_X1 port map( A1 => n2111, A2 => n2112, ZN => n15);
   U37 : OR2_X1 port map( A1 => n3617, A2 => n3616, ZN => n16);
   U38 : OR2_X1 port map( A1 => n2137, A2 => n2138, ZN => n17);
   U39 : CLKBUF_X1 port map( A => n2162, Z => n19);
   U40 : CLKBUF_X3 port map( A => n1350, Z => n313);
   U41 : BUF_X2 port map( A => n1347, Z => n307);
   U42 : CLKBUF_X3 port map( A => n1350, Z => n314);
   U43 : BUF_X2 port map( A => n2206, Z => n477);
   U44 : CLKBUF_X3 port map( A => n2206, Z => n476);
   U45 : CLKBUF_X3 port map( A => n2206, Z => n478);
   U46 : CLKBUF_X1 port map( A => n2143, Z => n18);
   U47 : BUF_X2 port map( A => n1370, Z => n349);
   U48 : AND2_X2 port map( A1 => ADD_RS2(1), A2 => n2173, ZN => n2142);
   U49 : BUF_X1 port map( A => ADD_RS2(3), Z => n80);
   U50 : CLKBUF_X3 port map( A => n1363, Z => n20);
   U51 : CLKBUF_X3 port map( A => n1363, Z => n21);
   U52 : CLKBUF_X3 port map( A => n1382, Z => n22);
   U53 : CLKBUF_X3 port map( A => n1382, Z => n23);
   U54 : CLKBUF_X3 port map( A => n2222, Z => n24);
   U55 : CLKBUF_X3 port map( A => n2222, Z => n25);
   U56 : CLKBUF_X1 port map( A => n2149, Z => n78);
   U57 : CLKBUF_X1 port map( A => n2156, Z => n26);
   U58 : NOR3_X1 port map( A1 => n2469, A2 => n2468, A3 => n7, ZN => n2467);
   U59 : BUF_X1 port map( A => n2205, Z => n27);
   U60 : BUF_X1 port map( A => n2205, Z => n28);
   U61 : BUF_X1 port map( A => n1337, Z => n29);
   U62 : BUF_X1 port map( A => n1337, Z => n30);
   U63 : NOR3_X1 port map( A1 => n2487, A2 => n2486, A3 => n8, ZN => n2485);
   U64 : NOR3_X1 port map( A1 => n3723, A2 => n3722, A3 => n9, ZN => n3721);
   U65 : NOR3_X1 port map( A1 => n2505, A2 => n2504, A3 => n10, ZN => n2503);
   U66 : NOR3_X1 port map( A1 => n3741, A2 => n3740, A3 => n11, ZN => n3739);
   U67 : NOR3_X1 port map( A1 => n3579, A2 => n3578, A3 => n12, ZN => n3577);
   U68 : BUF_X1 port map( A => n1362, Z => n31);
   U69 : BUF_X1 port map( A => n1362, Z => n32);
   U70 : NOR3_X1 port map( A1 => n1809, A2 => n1810, A3 => n6, ZN => n1808);
   U71 : CLKBUF_X3 port map( A => n1368, Z => n344);
   U72 : CLKBUF_X2 port map( A => n1368, Z => n345);
   U73 : CLKBUF_X3 port map( A => n1368, Z => n343);
   U74 : NOR3_X1 port map( A1 => n2059, A2 => n2060, A3 => n13, ZN => n2058);
   U75 : CLKBUF_X3 port map( A => n1380, Z => n428);
   U76 : NOR3_X1 port map( A1 => n3596, A2 => n3597, A3 => n14, ZN => n3595);
   U77 : CLKBUF_X3 port map( A => n2216, Z => n492);
   U78 : NOR3_X1 port map( A1 => n2109, A2 => n2110, A3 => n15, ZN => n2108);
   U79 : NOR3_X1 port map( A1 => n3614, A2 => n3615, A3 => n16, ZN => n3613);
   U80 : CLKBUF_X3 port map( A => n2217, Z => n496);
   U81 : CLKBUF_X3 port map( A => n2217, Z => n495);
   U82 : NOR3_X1 port map( A1 => n2135, A2 => n2136, A3 => n17, ZN => n2133);
   U83 : CLKBUF_X3 port map( A => n1380, Z => n429);
   U84 : BUF_X1 port map( A => n2163, Z => n35);
   U85 : CLKBUF_X1 port map( A => n3854, Z => n36);
   U86 : BUF_X2 port map( A => n1377, Z => n425);
   U87 : BUF_X2 port map( A => n1339, Z => n228);
   U88 : BUF_X1 port map( A => n1339, Z => n293);
   U89 : BUF_X1 port map( A => n1377, Z => n427);
   U90 : BUF_X1 port map( A => n716, Z => n715);
   U91 : BUF_X1 port map( A => n1347, Z => n308);
   U92 : BUF_X2 port map( A => n1336, Z => n222);
   U93 : BUF_X2 port map( A => n1336, Z => n223);
   U94 : BUF_X2 port map( A => n1360, Z => n329);
   U95 : BUF_X2 port map( A => n1348, Z => n310);
   U96 : BUF_X2 port map( A => n1348, Z => n311);
   U97 : BUF_X2 port map( A => n1365, Z => n337);
   U98 : BUF_X2 port map( A => n1365, Z => n338);
   U99 : BUF_X2 port map( A => n1352, Z => n316);
   U100 : BUF_X2 port map( A => n1375, Z => n355);
   U101 : BUF_X2 port map( A => n1352, Z => n317);
   U102 : BUF_X2 port map( A => n1332, Z => n216);
   U103 : BUF_X2 port map( A => n1332, Z => n217);
   U104 : BUF_X2 port map( A => n1373, Z => n352);
   U105 : BUF_X2 port map( A => n1373, Z => n353);
   U106 : BUF_X2 port map( A => n1334, Z => n219);
   U107 : BUF_X2 port map( A => n1340, Z => n295);
   U108 : BUF_X2 port map( A => n1334, Z => n220);
   U109 : BUF_X2 port map( A => n1340, Z => n296);
   U110 : BUF_X2 port map( A => n1337, Z => n225);
   U111 : BUF_X1 port map( A => n1337, Z => n226);
   U112 : BUF_X2 port map( A => n1359, Z => n326);
   U113 : BUF_X2 port map( A => n1364, Z => n334);
   U114 : BUF_X2 port map( A => n1364, Z => n335);
   U115 : BUF_X2 port map( A => n1344, Z => n304);
   U116 : BUF_X2 port map( A => n1344, Z => n305);
   U117 : BUF_X1 port map( A => n1362, Z => n333);
   U118 : BUF_X1 port map( A => n1362, Z => n332);
   U119 : BUF_X2 port map( A => n1376, Z => n422);
   U120 : BUF_X2 port map( A => n1376, Z => n423);
   U121 : BUF_X1 port map( A => n1362, Z => n331);
   U122 : BUF_X2 port map( A => n1353, Z => n321);
   U123 : BUF_X2 port map( A => n1342, Z => n300);
   U124 : BUF_X1 port map( A => n1336, Z => n224);
   U125 : BUF_X2 port map( A => n1360, Z => n330);
   U126 : BUF_X2 port map( A => n1348, Z => n312);
   U127 : BUF_X2 port map( A => n1365, Z => n339);
   U128 : BUF_X2 port map( A => n1375, Z => n421);
   U129 : BUF_X1 port map( A => n1332, Z => n218);
   U130 : BUF_X2 port map( A => n1373, Z => n354);
   U131 : BUF_X1 port map( A => n1340, Z => n297);
   U132 : BUF_X1 port map( A => n1334, Z => n221);
   U133 : BUF_X2 port map( A => n1380, Z => n430);
   U134 : BUF_X2 port map( A => n1354, Z => n324);
   U135 : BUF_X1 port map( A => n1343, Z => n303);
   U136 : BUF_X1 port map( A => n1337, Z => n227);
   U137 : BUF_X1 port map( A => n1359, Z => n327);
   U138 : BUF_X1 port map( A => n1364, Z => n336);
   U139 : BUF_X1 port map( A => n1369, Z => n348);
   U140 : BUF_X1 port map( A => n1344, Z => n306);
   U141 : BUF_X1 port map( A => n594, Z => n716);
   U142 : BUF_X1 port map( A => n595, Z => n720);
   U143 : BUF_X1 port map( A => n595, Z => n721);
   U144 : BUF_X1 port map( A => n595, Z => n719);
   U145 : BUF_X1 port map( A => n594, Z => n718);
   U146 : BUF_X1 port map( A => n594, Z => n717);
   U147 : BUF_X1 port map( A => n597, Z => n727);
   U148 : BUF_X1 port map( A => n596, Z => n723);
   U149 : BUF_X1 port map( A => n597, Z => n726);
   U150 : BUF_X1 port map( A => n597, Z => n725);
   U151 : BUF_X1 port map( A => n596, Z => n724);
   U152 : BUF_X1 port map( A => n596, Z => n722);
   U153 : BUF_X1 port map( A => n598, Z => n728);
   U154 : BUF_X1 port map( A => n598, Z => n729);
   U155 : BUF_X2 port map( A => n2192, Z => n446);
   U156 : BUF_X2 port map( A => n2192, Z => n447);
   U157 : BUF_X2 port map( A => n2207, Z => n479);
   U158 : BUF_X2 port map( A => n2197, Z => n458);
   U159 : BUF_X2 port map( A => n2207, Z => n480);
   U160 : BUF_X2 port map( A => n2197, Z => n459);
   U161 : BUF_X2 port map( A => n2203, Z => n471);
   U162 : BUF_X2 port map( A => n2224, Z => n510);
   U163 : BUF_X2 port map( A => n2229, Z => n554);
   U164 : BUF_X2 port map( A => n2214, Z => n488);
   U165 : BUF_X2 port map( A => n2214, Z => n489);
   U166 : BUF_X2 port map( A => n2219, Z => n500);
   U167 : BUF_X2 port map( A => n2219, Z => n501);
   U168 : BUF_X2 port map( A => n2217, Z => n494);
   U169 : BUF_X2 port map( A => n2232, Z => n559);
   U170 : BUF_X2 port map( A => n2232, Z => n560);
   U171 : BUF_X2 port map( A => n2189, Z => n440);
   U172 : BUF_X2 port map( A => n2189, Z => n441);
   U173 : BUF_X2 port map( A => n2194, Z => n452);
   U174 : BUF_X2 port map( A => n2194, Z => n453);
   U175 : BUF_X2 port map( A => n2231, Z => n556);
   U176 : BUF_X2 port map( A => n2231, Z => n557);
   U177 : BUF_X2 port map( A => n2221, Z => n503);
   U178 : BUF_X2 port map( A => n2216, Z => n491);
   U179 : BUF_X2 port map( A => n2226, Z => n512);
   U180 : BUF_X2 port map( A => n2221, Z => n504);
   U181 : BUF_X2 port map( A => n2226, Z => n513);
   U182 : BUF_X1 port map( A => n2205, Z => n473);
   U183 : BUF_X1 port map( A => n2205, Z => n474);
   U184 : BUF_X2 port map( A => n2190, Z => n443);
   U185 : BUF_X2 port map( A => n2195, Z => n455);
   U186 : BUF_X2 port map( A => n2190, Z => n444);
   U187 : BUF_X2 port map( A => n2195, Z => n456);
   U188 : BUF_X2 port map( A => n2208, Z => n482);
   U189 : BUF_X2 port map( A => n2198, Z => n461);
   U190 : BUF_X2 port map( A => n2208, Z => n483);
   U191 : BUF_X2 port map( A => n2193, Z => n450);
   U192 : BUF_X2 port map( A => n2198, Z => n462);
   U193 : BUF_X1 port map( A => n2193, Z => n449);
   U194 : BUF_X2 port map( A => n2202, Z => n468);
   U195 : BUF_X2 port map( A => n2228, Z => n551);
   U196 : BUF_X2 port map( A => n2223, Z => n507);
   U197 : BUF_X2 port map( A => n2218, Z => n497);
   U198 : BUF_X2 port map( A => n2213, Z => n485);
   U199 : BUF_X2 port map( A => n2213, Z => n486);
   U200 : BUF_X2 port map( A => n2218, Z => n498);
   U201 : BUF_X2 port map( A => n2199, Z => n464);
   U202 : BUF_X2 port map( A => n2199, Z => n465);
   U203 : BUF_X2 port map( A => n2227, Z => n516);
   U204 : BUF_X2 port map( A => n2227, Z => n549);
   U205 : BUF_X1 port map( A => n2192, Z => n448);
   U206 : BUF_X1 port map( A => n2197, Z => n460);
   U207 : BUF_X1 port map( A => n2207, Z => n481);
   U208 : BUF_X1 port map( A => n2203, Z => n472);
   U209 : BUF_X1 port map( A => n2224, Z => n511);
   U210 : BUF_X1 port map( A => n2229, Z => n555);
   U211 : BUF_X1 port map( A => n2214, Z => n490);
   U212 : BUF_X1 port map( A => n2219, Z => n502);
   U213 : BUF_X1 port map( A => n2189, Z => n442);
   U214 : BUF_X2 port map( A => n2194, Z => n454);
   U215 : BUF_X2 port map( A => n2231, Z => n558);
   U216 : BUF_X2 port map( A => n2226, Z => n514);
   U217 : BUF_X2 port map( A => n2221, Z => n505);
   U218 : BUF_X2 port map( A => n2216, Z => n493);
   U219 : BUF_X2 port map( A => n2205, Z => n475);
   U220 : BUF_X2 port map( A => n2190, Z => n445);
   U221 : BUF_X1 port map( A => n2202, Z => n469);
   U222 : BUF_X1 port map( A => n2228, Z => n552);
   U223 : BUF_X1 port map( A => n2193, Z => n451);
   U224 : BUF_X1 port map( A => n2208, Z => n484);
   U225 : BUF_X1 port map( A => n2198, Z => n463);
   U226 : BUF_X1 port map( A => n2223, Z => n508);
   U227 : BUF_X1 port map( A => n2218, Z => n499);
   U228 : BUF_X1 port map( A => n2213, Z => n487);
   U229 : BUF_X1 port map( A => n2199, Z => n466);
   U230 : BUF_X1 port map( A => n599, Z => n597);
   U231 : BUF_X1 port map( A => n599, Z => n596);
   U232 : BUF_X1 port map( A => n600, Z => n595);
   U233 : BUF_X1 port map( A => n600, Z => n594);
   U234 : BUF_X1 port map( A => n599, Z => n598);
   U235 : BUF_X1 port map( A => n1257, Z => n201);
   U236 : BUF_X1 port map( A => n1257, Z => n202);
   U237 : BUF_X1 port map( A => n1222, Z => n192);
   U238 : BUF_X1 port map( A => n1222, Z => n193);
   U239 : BUF_X1 port map( A => n1116, Z => n171);
   U240 : BUF_X1 port map( A => n1116, Z => n172);
   U241 : BUF_X1 port map( A => n1081, Z => n162);
   U242 : BUF_X1 port map( A => n1081, Z => n163);
   U243 : BUF_X1 port map( A => n1012, Z => n150);
   U244 : BUF_X1 port map( A => n1012, Z => n151);
   U245 : BUF_X1 port map( A => n979, Z => n147);
   U246 : BUF_X1 port map( A => n979, Z => n148);
   U247 : BUF_X1 port map( A => n912, Z => n138);
   U248 : BUF_X1 port map( A => n912, Z => n139);
   U249 : BUF_X1 port map( A => n877, Z => n135);
   U250 : BUF_X1 port map( A => n877, Z => n136);
   U251 : BUF_X1 port map( A => n1290, Z => n204);
   U252 : BUF_X1 port map( A => n1290, Z => n205);
   U253 : BUF_X1 port map( A => n1255, Z => n198);
   U254 : BUF_X1 port map( A => n1255, Z => n199);
   U255 : BUF_X1 port map( A => n1254, Z => n195);
   U256 : BUF_X1 port map( A => n1254, Z => n196);
   U257 : BUF_X1 port map( A => n1188, Z => n189);
   U258 : BUF_X1 port map( A => n1188, Z => n190);
   U259 : BUF_X1 port map( A => n1185, Z => n186);
   U260 : BUF_X1 port map( A => n1185, Z => n187);
   U261 : BUF_X1 port map( A => n1183, Z => n183);
   U262 : BUF_X1 port map( A => n1183, Z => n184);
   U263 : BUF_X1 port map( A => n1182, Z => n180);
   U264 : BUF_X1 port map( A => n1182, Z => n181);
   U265 : BUF_X1 port map( A => n1181, Z => n177);
   U266 : BUF_X1 port map( A => n1181, Z => n178);
   U267 : BUF_X1 port map( A => n1149, Z => n174);
   U268 : BUF_X1 port map( A => n1149, Z => n175);
   U269 : BUF_X1 port map( A => n1114, Z => n168);
   U270 : BUF_X1 port map( A => n1114, Z => n169);
   U271 : BUF_X1 port map( A => n1113, Z => n165);
   U272 : BUF_X1 port map( A => n1113, Z => n166);
   U273 : BUF_X1 port map( A => n1047, Z => n159);
   U274 : BUF_X1 port map( A => n1047, Z => n160);
   U275 : BUF_X1 port map( A => n1045, Z => n156);
   U276 : BUF_X1 port map( A => n1045, Z => n157);
   U277 : BUF_X1 port map( A => n1044, Z => n153);
   U278 : BUF_X1 port map( A => n1044, Z => n154);
   U279 : BUF_X1 port map( A => n977, Z => n144);
   U280 : BUF_X1 port map( A => n977, Z => n145);
   U281 : BUF_X1 port map( A => n976, Z => n141);
   U282 : BUF_X1 port map( A => n976, Z => n142);
   U283 : BUF_X1 port map( A => n871, Z => n132);
   U284 : BUF_X1 port map( A => n871, Z => n133);
   U285 : BUF_X1 port map( A => n869, Z => n129);
   U286 : BUF_X1 port map( A => n869, Z => n130);
   U287 : BUF_X1 port map( A => n804, Z => n126);
   U288 : BUF_X1 port map( A => n804, Z => n127);
   U289 : BUF_X1 port map( A => n770, Z => n123);
   U290 : BUF_X1 port map( A => n770, Z => n124);
   U291 : BUF_X1 port map( A => n767, Z => n120);
   U292 : BUF_X1 port map( A => n767, Z => n121);
   U293 : BUF_X1 port map( A => n765, Z => n117);
   U294 : BUF_X1 port map( A => n765, Z => n118);
   U295 : BUF_X1 port map( A => n731, Z => n114);
   U296 : BUF_X1 port map( A => n731, Z => n115);
   U297 : BUF_X2 port map( A => n2183, Z => n434);
   U298 : BUF_X2 port map( A => n2183, Z => n435);
   U299 : BUF_X2 port map( A => n1324, Z => n207);
   U300 : BUF_X2 port map( A => n1324, Z => n208);
   U301 : BUF_X2 port map( A => n2181, Z => n431);
   U302 : BUF_X2 port map( A => n2181, Z => n432);
   U303 : BUF_X1 port map( A => n1257, Z => n203);
   U304 : BUF_X1 port map( A => n1222, Z => n194);
   U305 : BUF_X1 port map( A => n1116, Z => n173);
   U306 : BUF_X1 port map( A => n1081, Z => n164);
   U307 : BUF_X1 port map( A => n1012, Z => n152);
   U308 : BUF_X1 port map( A => n979, Z => n149);
   U309 : BUF_X1 port map( A => n912, Z => n140);
   U310 : BUF_X1 port map( A => n877, Z => n137);
   U311 : BUF_X1 port map( A => n1290, Z => n206);
   U312 : BUF_X1 port map( A => n1255, Z => n200);
   U313 : BUF_X1 port map( A => n1254, Z => n197);
   U314 : BUF_X1 port map( A => n1188, Z => n191);
   U315 : BUF_X1 port map( A => n1185, Z => n188);
   U316 : BUF_X1 port map( A => n1183, Z => n185);
   U317 : BUF_X1 port map( A => n1182, Z => n182);
   U318 : BUF_X1 port map( A => n1181, Z => n179);
   U319 : BUF_X1 port map( A => n1149, Z => n176);
   U320 : BUF_X1 port map( A => n1114, Z => n170);
   U321 : BUF_X1 port map( A => n1113, Z => n167);
   U322 : BUF_X1 port map( A => n1047, Z => n161);
   U323 : BUF_X1 port map( A => n767, Z => n122);
   U324 : BUF_X1 port map( A => n765, Z => n119);
   U325 : BUF_X1 port map( A => n731, Z => n116);
   U326 : BUF_X1 port map( A => n1045, Z => n158);
   U327 : BUF_X1 port map( A => n1044, Z => n155);
   U328 : BUF_X1 port map( A => n977, Z => n146);
   U329 : BUF_X1 port map( A => n976, Z => n143);
   U330 : BUF_X1 port map( A => n871, Z => n134);
   U331 : BUF_X1 port map( A => n869, Z => n131);
   U332 : BUF_X1 port map( A => n804, Z => n128);
   U333 : BUF_X1 port map( A => n770, Z => n125);
   U334 : BUF_X1 port map( A => n2183, Z => n436);
   U335 : BUF_X1 port map( A => n1326, Z => n212);
   U336 : BUF_X1 port map( A => n2181, Z => n433);
   U337 : BUF_X1 port map( A => n1324, Z => n209);
   U338 : BUF_X1 port map( A => RST, Z => n599);
   U339 : BUF_X1 port map( A => RST, Z => n600);
   U340 : BUF_X1 port map( A => n2184, Z => n437);
   U341 : BUF_X1 port map( A => n1327, Z => n213);
   U342 : BUF_X1 port map( A => n2184, Z => n438);
   U343 : BUF_X1 port map( A => n1327, Z => n214);
   U344 : BUF_X1 port map( A => n2184, Z => n439);
   U345 : BUF_X1 port map( A => n1327, Z => n215);
   U346 : INV_X1 port map( A => DATAIN(2), ZN => n564);
   U347 : INV_X1 port map( A => DATAIN(4), ZN => n566);
   U348 : INV_X1 port map( A => DATAIN(5), ZN => n567);
   U349 : INV_X1 port map( A => DATAIN(6), ZN => n568);
   U350 : INV_X1 port map( A => DATAIN(7), ZN => n569);
   U351 : INV_X1 port map( A => DATAIN(8), ZN => n570);
   U352 : INV_X1 port map( A => DATAIN(10), ZN => n572);
   U353 : INV_X1 port map( A => DATAIN(11), ZN => n573);
   U354 : INV_X1 port map( A => DATAIN(12), ZN => n574);
   U355 : INV_X1 port map( A => DATAIN(13), ZN => n575);
   U356 : INV_X1 port map( A => DATAIN(14), ZN => n576);
   U357 : INV_X1 port map( A => DATAIN(15), ZN => n577);
   U358 : INV_X1 port map( A => DATAIN(16), ZN => n578);
   U359 : INV_X1 port map( A => DATAIN(17), ZN => n579);
   U360 : INV_X1 port map( A => DATAIN(18), ZN => n580);
   U361 : INV_X1 port map( A => DATAIN(19), ZN => n581);
   U362 : INV_X1 port map( A => DATAIN(20), ZN => n582);
   U363 : INV_X1 port map( A => DATAIN(21), ZN => n583);
   U364 : INV_X1 port map( A => DATAIN(22), ZN => n584);
   U365 : INV_X1 port map( A => DATAIN(23), ZN => n585);
   U366 : INV_X1 port map( A => DATAIN(24), ZN => n586);
   U367 : INV_X1 port map( A => DATAIN(25), ZN => n587);
   U368 : INV_X1 port map( A => DATAIN(26), ZN => n588);
   U369 : INV_X1 port map( A => DATAIN(27), ZN => n589);
   U370 : INV_X1 port map( A => DATAIN(28), ZN => n590);
   U371 : INV_X1 port map( A => DATAIN(29), ZN => n591);
   U372 : INV_X1 port map( A => DATAIN(30), ZN => n592);
   U373 : INV_X1 port map( A => DATAIN(31), ZN => n593);
   U374 : INV_X1 port map( A => DATAIN(0), ZN => n562);
   U375 : INV_X1 port map( A => DATAIN(1), ZN => n563);
   U376 : INV_X1 port map( A => DATAIN(3), ZN => n565);
   U377 : INV_X1 port map( A => DATAIN(9), ZN => n571);
   U378 : OR2_X1 port map( A1 => n3815, A2 => n3814, ZN => n37);
   U379 : OR2_X1 port map( A1 => n3797, A2 => n3796, ZN => n38);
   U380 : OR2_X1 port map( A1 => n3779, A2 => n3778, ZN => n39);
   U381 : OR2_X1 port map( A1 => n2037, A2 => n2036, ZN => n40);
   U382 : OR2_X1 port map( A1 => n1987, A2 => n1986, ZN => n41);
   U383 : OR2_X1 port map( A1 => n1937, A2 => n1936, ZN => n42);
   U384 : OR2_X1 port map( A1 => n1887, A2 => n1886, ZN => n43);
   U385 : OR2_X1 port map( A1 => n1837, A2 => n1836, ZN => n44);
   U386 : OR2_X1 port map( A1 => n1787, A2 => n1786, ZN => n45);
   U387 : OR2_X1 port map( A1 => n1737, A2 => n1736, ZN => n46);
   U388 : OR2_X1 port map( A1 => n1687, A2 => n1686, ZN => n47);
   U389 : OR2_X1 port map( A1 => n1637, A2 => n1636, ZN => n48);
   U390 : OR2_X1 port map( A1 => n1587, A2 => n1586, ZN => n49);
   U391 : OR2_X1 port map( A1 => n2087, A2 => n2086, ZN => n50);
   U392 : OR2_X1 port map( A1 => n3761, A2 => n3760, ZN => n51);
   U393 : OR2_X1 port map( A1 => n3689, A2 => n3688, ZN => n52);
   U394 : OR2_X1 port map( A1 => n3671, A2 => n3670, ZN => n53);
   U395 : CLKBUF_X1 port map( A => n2168, Z => n79);
   U396 : AND3_X1 port map( A1 => ADD_RS1(0), A2 => n56, A3 => ADD_RS1(3), ZN 
                           => n3855);
   U397 : BUF_X1 port map( A => n2141, Z => n54);
   U398 : INV_X1 port map( A => ADD_RS1(4), ZN => n55);
   U399 : INV_X1 port map( A => ADD_RS1(4), ZN => n56);
   U400 : CLKBUF_X1 port map( A => ADD_RS1(2), Z => n57);
   U401 : CLKBUF_X1 port map( A => n2, Z => n58);
   U402 : NAND2_X1 port map( A1 => n424, A2 => n739, ZN => n59);
   U403 : NAND2_X1 port map( A1 => n426, A2 => n3958, ZN => n60);
   U404 : INV_X1 port map( A => n1580, ZN => n61);
   U405 : AND3_X1 port map( A1 => n59, A2 => n60, A3 => n61, ZN => n1571);
   U406 : NAND2_X1 port map( A1 => n424, A2 => n741, ZN => n62);
   U407 : NAND2_X1 port map( A1 => n426, A2 => n3956, ZN => n63);
   U408 : INV_X1 port map( A => n1630, ZN => n64);
   U409 : AND3_X1 port map( A1 => n62, A2 => n63, A3 => n64, ZN => n1621);
   U410 : NAND2_X1 port map( A1 => n424, A2 => n743, ZN => n65);
   U411 : NAND2_X1 port map( A1 => n426, A2 => n3954, ZN => n66);
   U412 : INV_X1 port map( A => n1680, ZN => n67);
   U413 : AND3_X1 port map( A1 => n65, A2 => n66, A3 => n67, ZN => n1671);
   U414 : NAND2_X1 port map( A1 => n424, A2 => n745, ZN => n68);
   U415 : NAND2_X1 port map( A1 => n426, A2 => n3952, ZN => n69);
   U416 : INV_X1 port map( A => n1730, ZN => n70);
   U417 : AND3_X1 port map( A1 => n68, A2 => n69, A3 => n70, ZN => n1721);
   U418 : NAND2_X1 port map( A1 => n424, A2 => n747, ZN => n71);
   U419 : NAND2_X1 port map( A1 => n426, A2 => n3950, ZN => n72);
   U420 : INV_X1 port map( A => n1780, ZN => n73);
   U421 : AND3_X1 port map( A1 => n71, A2 => n72, A3 => n73, ZN => n1771);
   U422 : NAND2_X1 port map( A1 => n424, A2 => n749, ZN => n74);
   U423 : NAND2_X1 port map( A1 => n426, A2 => n3948, ZN => n75);
   U424 : INV_X1 port map( A => n1830, ZN => n76);
   U425 : AND3_X1 port map( A1 => n74, A2 => n75, A3 => n76, ZN => n1821);
   U426 : BUF_X2 port map( A => n1376, Z => n424);
   U427 : BUF_X2 port map( A => n1377, Z => n426);
   U428 : CLKBUF_X1 port map( A => n1339, Z => n294);
   U429 : CLKBUF_X1 port map( A => n2149, Z => n85);
   U430 : INV_X1 port map( A => ADD_RS2(0), ZN => n77);
   U431 : BUF_X1 port map( A => n1370, Z => n350);
   U432 : BUF_X1 port map( A => n1370, Z => n351);
   U433 : AND2_X1 port map( A1 => n325, A2 => n4194, ZN => n81);
   U434 : AND2_X1 port map( A1 => n328, A2 => n4226, ZN => n82);
   U435 : NOR3_X1 port map( A1 => n81, A2 => n82, A3 => n2075, ZN => n2074);
   U436 : BUF_X2 port map( A => n1359, Z => n325);
   U437 : BUF_X2 port map( A => n1360, Z => n328);
   U438 : INV_X1 port map( A => ADD_RS1(0), ZN => n83);
   U439 : INV_X1 port map( A => ADD_RS1(0), ZN => n84);
   U440 : CLKBUF_X2 port map( A => n2232, Z => n561);
   U441 : CLKBUF_X2 port map( A => n2227, Z => n515);
   U442 : AND2_X1 port map( A1 => ADD_RS2(2), A2 => ADD_RS2(1), ZN => n2145);
   U443 : NOR3_X1 port map( A1 => n77, A2 => ADD_RS2(4), A3 => ADD_RS2(3), ZN 
                           => n2168);
   U444 : INV_X1 port map( A => ADD_RS2(4), ZN => n86);
   U445 : NOR3_X1 port map( A1 => n1584, A2 => n1585, A3 => n49, ZN => n1583);
   U446 : NOR3_X1 port map( A1 => n1634, A2 => n1635, A3 => n48, ZN => n1633);
   U447 : NOR3_X1 port map( A1 => n1684, A2 => n1685, A3 => n47, ZN => n1683);
   U448 : NOR3_X1 port map( A1 => n1734, A2 => n1735, A3 => n46, ZN => n1733);
   U449 : NOR3_X1 port map( A1 => n1784, A2 => n1785, A3 => n45, ZN => n1783);
   U450 : NOR3_X1 port map( A1 => n1834, A2 => n1835, A3 => n44, ZN => n1833);
   U451 : NOR3_X1 port map( A1 => n1884, A2 => n1885, A3 => n43, ZN => n1883);
   U452 : NOR3_X1 port map( A1 => n1934, A2 => n1935, A3 => n42, ZN => n1933);
   U453 : NOR3_X1 port map( A1 => n1984, A2 => n1985, A3 => n41, ZN => n1983);
   U454 : NOR3_X1 port map( A1 => n2034, A2 => n2035, A3 => n40, ZN => n2033);
   U455 : AND2_X1 port map( A1 => n346, A2 => n799, ZN => n87);
   U456 : AND2_X1 port map( A1 => n349, A2 => n833, ZN => n88);
   U457 : NOR3_X1 port map( A1 => n87, A2 => n88, A3 => n2102, ZN => n2097);
   U458 : NOR3_X1 port map( A1 => n2085, A2 => n2084, A3 => n50, ZN => n2083);
   U459 : AND2_X1 port map( A1 => n346, A2 => n800, ZN => n89);
   U460 : AND2_X1 port map( A1 => n349, A2 => n834, ZN => n90);
   U461 : NOR3_X1 port map( A1 => n89, A2 => n90, A3 => n2127, ZN => n2122);
   U462 : AND2_X1 port map( A1 => n550, A2 => n762, ZN => n91);
   U463 : AND2_X1 port map( A1 => n553, A2 => n3935, ZN => n92);
   U464 : NOR3_X1 port map( A1 => n91, A2 => n92, A3 => n3860, ZN => n3849);
   U465 : BUF_X2 port map( A => n2228, Z => n550);
   U466 : BUF_X2 port map( A => n2229, Z => n553);
   U467 : AND2_X1 port map( A1 => n346, A2 => n801, ZN => n93);
   U468 : AND2_X1 port map( A1 => n349, A2 => n835, ZN => n94);
   U469 : NOR3_X1 port map( A1 => n93, A2 => n94, A3 => n2165, ZN => n2158);
   U470 : AND2_X1 port map( A1 => n506, A2 => n790, ZN => n95);
   U471 : AND2_X1 port map( A1 => n509, A2 => n824, ZN => n96);
   U472 : NOR3_X1 port map( A1 => n95, A2 => n96, A3 => n3647, ZN => n3642);
   U473 : AND2_X1 port map( A1 => n506, A2 => n791, ZN => n97);
   U474 : AND2_X1 port map( A1 => n509, A2 => n825, ZN => n98);
   U475 : NOR3_X1 port map( A1 => n97, A2 => n98, A3 => n3665, ZN => n3660);
   U476 : NOR3_X1 port map( A1 => n3668, A2 => n3669, A3 => n53, ZN => n3667);
   U477 : AND2_X1 port map( A1 => n506, A2 => n793, ZN => n99);
   U478 : AND2_X1 port map( A1 => n509, A2 => n827, ZN => n100);
   U479 : NOR3_X1 port map( A1 => n99, A2 => n100, A3 => n3701, ZN => n3696);
   U480 : NOR3_X1 port map( A1 => n3686, A2 => n3687, A3 => n52, ZN => n3685);
   U481 : AND2_X1 port map( A1 => n506, A2 => n794, ZN => n101);
   U482 : AND2_X1 port map( A1 => n509, A2 => n828, ZN => n102);
   U483 : NOR3_X1 port map( A1 => n101, A2 => n102, A3 => n3719, ZN => n3714);
   U484 : AND2_X1 port map( A1 => n506, A2 => n795, ZN => n103);
   U485 : AND2_X1 port map( A1 => n509, A2 => n829, ZN => n104);
   U486 : NOR3_X1 port map( A1 => n103, A2 => n104, A3 => n3737, ZN => n3732);
   U487 : AND2_X1 port map( A1 => n506, A2 => n796, ZN => n105);
   U488 : AND2_X1 port map( A1 => n509, A2 => n830, ZN => n106);
   U489 : NOR3_X1 port map( A1 => n105, A2 => n106, A3 => n3755, ZN => n3750);
   U490 : NOR3_X1 port map( A1 => n3758, A2 => n3759, A3 => n51, ZN => n3757);
   U491 : AND2_X2 port map( A1 => ADD_RS1(2), A2 => ADD_RS1(1), ZN => n3840);
   U492 : NOR3_X1 port map( A1 => n3776, A2 => n3777, A3 => n39, ZN => n3775);
   U493 : AND2_X1 port map( A1 => n506, A2 => n799, ZN => n107);
   U494 : AND2_X1 port map( A1 => n509, A2 => n833, ZN => n108);
   U495 : NOR3_X1 port map( A1 => n107, A2 => n108, A3 => n3809, ZN => n3804);
   U496 : NOR3_X1 port map( A1 => n3794, A2 => n3795, A3 => n38, ZN => n3793);
   U497 : NOR3_X1 port map( A1 => n3812, A2 => n3813, A3 => n37, ZN => n3811);
   U498 : AND2_X1 port map( A1 => n506, A2 => n801, ZN => n109);
   U499 : AND2_X1 port map( A1 => n509, A2 => n835, ZN => n110);
   U500 : NOR3_X1 port map( A1 => n109, A2 => n110, A3 => n3857, ZN => n3850);
   U501 : BUF_X2 port map( A => n2223, Z => n506);
   U502 : BUF_X2 port map( A => n2224, Z => n509);
   U503 : AND2_X1 port map( A1 => n467, A2 => n1180, ZN => n111);
   U504 : AND2_X1 port map( A1 => n470, A2 => n4127, ZN => n112);
   U505 : NOR3_X1 port map( A1 => n111, A2 => n112, A3 => n3847, ZN => n3846);
   U506 : NOR2_X1 port map( A1 => n3861, A2 => ADD_RS1(1), ZN => n113);
   U507 : BUF_X2 port map( A => n2202, Z => n467);
   U508 : BUF_X2 port map( A => n2203, Z => n470);
   U509 : CLKBUF_X3 port map( A => n1326, Z => n210);
   U510 : CLKBUF_X3 port map( A => n1326, Z => n211);
   U511 : CLKBUF_X3 port map( A => n1342, Z => n298);
   U512 : CLKBUF_X3 port map( A => n1342, Z => n299);
   U513 : CLKBUF_X1 port map( A => n729, Z => n601);
   U514 : CLKBUF_X1 port map( A => n729, Z => n602);
   U515 : CLKBUF_X1 port map( A => n729, Z => n603);
   U516 : CLKBUF_X1 port map( A => n729, Z => n604);
   U517 : CLKBUF_X1 port map( A => n729, Z => n605);
   U518 : CLKBUF_X1 port map( A => n728, Z => n606);
   U519 : CLKBUF_X1 port map( A => n728, Z => n607);
   U520 : CLKBUF_X1 port map( A => n728, Z => n608);
   U521 : CLKBUF_X1 port map( A => n728, Z => n609);
   U522 : CLKBUF_X1 port map( A => n728, Z => n610);
   U523 : CLKBUF_X1 port map( A => n728, Z => n611);
   U524 : CLKBUF_X1 port map( A => n727, Z => n612);
   U525 : CLKBUF_X1 port map( A => n727, Z => n645);
   U526 : CLKBUF_X1 port map( A => n727, Z => n646);
   U527 : CLKBUF_X1 port map( A => n727, Z => n647);
   U528 : CLKBUF_X1 port map( A => n727, Z => n648);
   U529 : CLKBUF_X1 port map( A => n727, Z => n649);
   U530 : CLKBUF_X1 port map( A => n726, Z => n650);
   U531 : CLKBUF_X1 port map( A => n726, Z => n651);
   U532 : CLKBUF_X1 port map( A => n726, Z => n652);
   U533 : CLKBUF_X1 port map( A => n726, Z => n653);
   U534 : CLKBUF_X1 port map( A => n726, Z => n654);
   U535 : CLKBUF_X1 port map( A => n726, Z => n655);
   U536 : CLKBUF_X1 port map( A => n725, Z => n656);
   U537 : CLKBUF_X1 port map( A => n725, Z => n657);
   U538 : CLKBUF_X1 port map( A => n725, Z => n658);
   U539 : CLKBUF_X1 port map( A => n725, Z => n659);
   U540 : CLKBUF_X1 port map( A => n725, Z => n660);
   U541 : CLKBUF_X1 port map( A => n725, Z => n661);
   U542 : CLKBUF_X1 port map( A => n724, Z => n662);
   U543 : CLKBUF_X1 port map( A => n724, Z => n663);
   U544 : CLKBUF_X1 port map( A => n724, Z => n664);
   U545 : CLKBUF_X1 port map( A => n724, Z => n665);
   U546 : CLKBUF_X1 port map( A => n724, Z => n666);
   U547 : CLKBUF_X1 port map( A => n724, Z => n667);
   U548 : CLKBUF_X1 port map( A => n723, Z => n668);
   U549 : CLKBUF_X1 port map( A => n723, Z => n669);
   U550 : CLKBUF_X1 port map( A => n723, Z => n670);
   U551 : CLKBUF_X1 port map( A => n723, Z => n671);
   U552 : CLKBUF_X1 port map( A => n723, Z => n672);
   U553 : CLKBUF_X1 port map( A => n723, Z => n673);
   U554 : CLKBUF_X1 port map( A => n722, Z => n674);
   U555 : CLKBUF_X1 port map( A => n722, Z => n675);
   U556 : CLKBUF_X1 port map( A => n722, Z => n676);
   U557 : CLKBUF_X1 port map( A => n722, Z => n677);
   U558 : CLKBUF_X1 port map( A => n722, Z => n678);
   U559 : CLKBUF_X1 port map( A => n722, Z => n679);
   U560 : CLKBUF_X1 port map( A => n721, Z => n680);
   U561 : CLKBUF_X1 port map( A => n721, Z => n681);
   U562 : CLKBUF_X1 port map( A => n721, Z => n682);
   U563 : CLKBUF_X1 port map( A => n721, Z => n683);
   U564 : CLKBUF_X1 port map( A => n721, Z => n684);
   U565 : CLKBUF_X1 port map( A => n721, Z => n685);
   U566 : CLKBUF_X1 port map( A => n720, Z => n686);
   U567 : CLKBUF_X1 port map( A => n720, Z => n687);
   U568 : CLKBUF_X1 port map( A => n720, Z => n688);
   U569 : CLKBUF_X1 port map( A => n720, Z => n689);
   U570 : CLKBUF_X1 port map( A => n720, Z => n690);
   U571 : CLKBUF_X1 port map( A => n720, Z => n691);
   U572 : CLKBUF_X1 port map( A => n719, Z => n692);
   U573 : CLKBUF_X1 port map( A => n719, Z => n693);
   U574 : CLKBUF_X1 port map( A => n719, Z => n694);
   U575 : CLKBUF_X1 port map( A => n719, Z => n695);
   U576 : CLKBUF_X1 port map( A => n719, Z => n696);
   U577 : CLKBUF_X1 port map( A => n719, Z => n697);
   U578 : CLKBUF_X1 port map( A => n718, Z => n698);
   U579 : CLKBUF_X1 port map( A => n718, Z => n699);
   U580 : CLKBUF_X1 port map( A => n718, Z => n700);
   U581 : CLKBUF_X1 port map( A => n718, Z => n701);
   U582 : CLKBUF_X1 port map( A => n718, Z => n702);
   U583 : CLKBUF_X1 port map( A => n718, Z => n703);
   U584 : CLKBUF_X1 port map( A => n717, Z => n704);
   U585 : CLKBUF_X1 port map( A => n717, Z => n705);
   U586 : CLKBUF_X1 port map( A => n717, Z => n706);
   U587 : CLKBUF_X1 port map( A => n717, Z => n707);
   U588 : CLKBUF_X1 port map( A => n717, Z => n708);
   U589 : CLKBUF_X1 port map( A => n717, Z => n709);
   U590 : CLKBUF_X1 port map( A => n716, Z => n710);
   U591 : CLKBUF_X1 port map( A => n716, Z => n711);
   U592 : CLKBUF_X1 port map( A => n716, Z => n712);
   U593 : CLKBUF_X1 port map( A => n716, Z => n713);
   U594 : CLKBUF_X1 port map( A => n716, Z => n714);
   U595 : MUX2_X1 port map( A => n730, B => DATAIN(31), S => n116, Z => n3561);
   U596 : MUX2_X1 port map( A => n732, B => DATAIN(30), S => n116, Z => n3560);
   U597 : MUX2_X1 port map( A => n733, B => DATAIN(29), S => n116, Z => n3559);
   U598 : MUX2_X1 port map( A => n734, B => DATAIN(28), S => n116, Z => n3558);
   U599 : MUX2_X1 port map( A => n735, B => DATAIN(27), S => n116, Z => n3557);
   U600 : MUX2_X1 port map( A => n736, B => DATAIN(26), S => n116, Z => n3556);
   U601 : MUX2_X1 port map( A => n737, B => DATAIN(25), S => n116, Z => n3555);
   U602 : MUX2_X1 port map( A => n738, B => DATAIN(24), S => n116, Z => n3554);
   U603 : MUX2_X1 port map( A => n739, B => DATAIN(23), S => n115, Z => n3553);
   U604 : MUX2_X1 port map( A => n740, B => DATAIN(22), S => n115, Z => n3552);
   U605 : MUX2_X1 port map( A => n741, B => DATAIN(21), S => n115, Z => n3551);
   U606 : MUX2_X1 port map( A => n742, B => DATAIN(20), S => n115, Z => n3550);
   U607 : MUX2_X1 port map( A => n743, B => DATAIN(19), S => n115, Z => n3549);
   U608 : MUX2_X1 port map( A => n744, B => DATAIN(18), S => n115, Z => n3548);
   U609 : MUX2_X1 port map( A => n745, B => DATAIN(17), S => n115, Z => n3547);
   U610 : MUX2_X1 port map( A => n746, B => DATAIN(16), S => n115, Z => n3546);
   U611 : MUX2_X1 port map( A => n747, B => DATAIN(15), S => n115, Z => n3545);
   U612 : MUX2_X1 port map( A => n748, B => DATAIN(14), S => n115, Z => n3544);
   U613 : MUX2_X1 port map( A => n749, B => DATAIN(13), S => n115, Z => n3543);
   U614 : MUX2_X1 port map( A => n750, B => DATAIN(12), S => n115, Z => n3542);
   U615 : MUX2_X1 port map( A => n751, B => DATAIN(11), S => n114, Z => n3541);
   U616 : MUX2_X1 port map( A => n752, B => DATAIN(10), S => n114, Z => n3540);
   U617 : MUX2_X1 port map( A => n753, B => DATAIN(9), S => n114, Z => n3539);
   U618 : MUX2_X1 port map( A => n754, B => DATAIN(8), S => n114, Z => n3538);
   U619 : MUX2_X1 port map( A => n755, B => DATAIN(7), S => n114, Z => n3537);
   U620 : MUX2_X1 port map( A => n756, B => DATAIN(6), S => n114, Z => n3536);
   U621 : MUX2_X1 port map( A => n757, B => DATAIN(5), S => n114, Z => n3535);
   U622 : MUX2_X1 port map( A => n758, B => DATAIN(4), S => n114, Z => n3534);
   U623 : MUX2_X1 port map( A => n759, B => DATAIN(3), S => n114, Z => n3533);
   U624 : MUX2_X1 port map( A => n760, B => DATAIN(2), S => n114, Z => n3532);
   U625 : MUX2_X1 port map( A => n761, B => DATAIN(1), S => n114, Z => n3531);
   U626 : MUX2_X1 port map( A => n762, B => DATAIN(0), S => n114, Z => n3530);
   U627 : AND2_X1 port map( A1 => n763, A2 => n764, ZN => n731);
   U628 : MUX2_X1 port map( A => n4446, B => DATAIN(31), S => n119, Z => n3529)
                           ;
   U629 : MUX2_X1 port map( A => n4445, B => DATAIN(30), S => n119, Z => n3528)
                           ;
   U630 : MUX2_X1 port map( A => n4444, B => DATAIN(29), S => n119, Z => n3527)
                           ;
   U631 : MUX2_X1 port map( A => n4443, B => DATAIN(28), S => n119, Z => n3526)
                           ;
   U632 : MUX2_X1 port map( A => n4442, B => DATAIN(27), S => n119, Z => n3525)
                           ;
   U633 : MUX2_X1 port map( A => n4441, B => DATAIN(26), S => n119, Z => n3524)
                           ;
   U634 : MUX2_X1 port map( A => n4440, B => DATAIN(25), S => n119, Z => n3523)
                           ;
   U635 : MUX2_X1 port map( A => n4439, B => DATAIN(24), S => n119, Z => n3522)
                           ;
   U636 : MUX2_X1 port map( A => n4438, B => DATAIN(23), S => n118, Z => n3521)
                           ;
   U637 : MUX2_X1 port map( A => n4437, B => DATAIN(22), S => n118, Z => n3520)
                           ;
   U638 : MUX2_X1 port map( A => n4436, B => DATAIN(21), S => n118, Z => n3519)
                           ;
   U639 : MUX2_X1 port map( A => n4435, B => DATAIN(20), S => n118, Z => n3518)
                           ;
   U640 : MUX2_X1 port map( A => n4434, B => DATAIN(19), S => n118, Z => n3517)
                           ;
   U641 : MUX2_X1 port map( A => n4433, B => DATAIN(18), S => n118, Z => n3516)
                           ;
   U642 : MUX2_X1 port map( A => n4432, B => DATAIN(17), S => n118, Z => n3515)
                           ;
   U643 : MUX2_X1 port map( A => n4431, B => DATAIN(16), S => n118, Z => n3514)
                           ;
   U644 : MUX2_X1 port map( A => n4430, B => DATAIN(15), S => n118, Z => n3513)
                           ;
   U645 : MUX2_X1 port map( A => n4429, B => DATAIN(14), S => n118, Z => n3512)
                           ;
   U646 : MUX2_X1 port map( A => n4428, B => DATAIN(13), S => n118, Z => n3511)
                           ;
   U647 : MUX2_X1 port map( A => n4427, B => DATAIN(12), S => n118, Z => n3510)
                           ;
   U648 : MUX2_X1 port map( A => n4426, B => DATAIN(11), S => n117, Z => n3509)
                           ;
   U649 : MUX2_X1 port map( A => n4425, B => DATAIN(10), S => n117, Z => n3508)
                           ;
   U650 : MUX2_X1 port map( A => n4424, B => DATAIN(9), S => n117, Z => n3507);
   U651 : MUX2_X1 port map( A => n4423, B => DATAIN(8), S => n117, Z => n3506);
   U652 : MUX2_X1 port map( A => n4422, B => DATAIN(7), S => n117, Z => n3505);
   U653 : MUX2_X1 port map( A => n4421, B => DATAIN(6), S => n117, Z => n3504);
   U654 : MUX2_X1 port map( A => n4420, B => DATAIN(5), S => n117, Z => n3503);
   U655 : MUX2_X1 port map( A => n4419, B => DATAIN(4), S => n117, Z => n3502);
   U656 : MUX2_X1 port map( A => n4418, B => DATAIN(3), S => n117, Z => n3501);
   U657 : MUX2_X1 port map( A => n4417, B => DATAIN(2), S => n117, Z => n3500);
   U658 : MUX2_X1 port map( A => n4416, B => DATAIN(1), S => n117, Z => n3499);
   U659 : MUX2_X1 port map( A => n4415, B => DATAIN(0), S => n117, Z => n3498);
   U660 : AND2_X1 port map( A1 => n766, A2 => n764, ZN => n765);
   U661 : MUX2_X1 port map( A => n4414, B => DATAIN(31), S => n122, Z => n3497)
                           ;
   U662 : MUX2_X1 port map( A => n4413, B => DATAIN(30), S => n122, Z => n3496)
                           ;
   U663 : MUX2_X1 port map( A => n4412, B => DATAIN(29), S => n122, Z => n3495)
                           ;
   U664 : MUX2_X1 port map( A => n4411, B => DATAIN(28), S => n122, Z => n3494)
                           ;
   U665 : MUX2_X1 port map( A => n4410, B => DATAIN(27), S => n122, Z => n3493)
                           ;
   U666 : MUX2_X1 port map( A => n4409, B => DATAIN(26), S => n122, Z => n3492)
                           ;
   U667 : MUX2_X1 port map( A => n4408, B => DATAIN(25), S => n122, Z => n3491)
                           ;
   U668 : MUX2_X1 port map( A => n4407, B => DATAIN(24), S => n122, Z => n3490)
                           ;
   U669 : MUX2_X1 port map( A => n4406, B => DATAIN(23), S => n121, Z => n3489)
                           ;
   U670 : MUX2_X1 port map( A => n4405, B => DATAIN(22), S => n121, Z => n3488)
                           ;
   U671 : MUX2_X1 port map( A => n4404, B => DATAIN(21), S => n121, Z => n3487)
                           ;
   U672 : MUX2_X1 port map( A => n4403, B => DATAIN(20), S => n121, Z => n3486)
                           ;
   U673 : MUX2_X1 port map( A => n4402, B => DATAIN(19), S => n121, Z => n3485)
                           ;
   U674 : MUX2_X1 port map( A => n4401, B => DATAIN(18), S => n121, Z => n3484)
                           ;
   U675 : MUX2_X1 port map( A => n4400, B => DATAIN(17), S => n121, Z => n3483)
                           ;
   U676 : MUX2_X1 port map( A => n4399, B => DATAIN(16), S => n121, Z => n3482)
                           ;
   U677 : MUX2_X1 port map( A => n4398, B => DATAIN(15), S => n121, Z => n3481)
                           ;
   U678 : MUX2_X1 port map( A => n4397, B => DATAIN(14), S => n121, Z => n3480)
                           ;
   U679 : MUX2_X1 port map( A => n4396, B => DATAIN(13), S => n121, Z => n3479)
                           ;
   U680 : MUX2_X1 port map( A => n4395, B => DATAIN(12), S => n121, Z => n3478)
                           ;
   U681 : MUX2_X1 port map( A => n4394, B => DATAIN(11), S => n120, Z => n3477)
                           ;
   U682 : MUX2_X1 port map( A => n4393, B => DATAIN(10), S => n120, Z => n3476)
                           ;
   U683 : MUX2_X1 port map( A => n4392, B => DATAIN(9), S => n120, Z => n3475);
   U684 : MUX2_X1 port map( A => n4391, B => DATAIN(8), S => n120, Z => n3474);
   U685 : MUX2_X1 port map( A => n4390, B => DATAIN(7), S => n120, Z => n3473);
   U686 : MUX2_X1 port map( A => n4389, B => DATAIN(6), S => n120, Z => n3472);
   U687 : MUX2_X1 port map( A => n4388, B => DATAIN(5), S => n120, Z => n3471);
   U688 : MUX2_X1 port map( A => n4387, B => DATAIN(4), S => n120, Z => n3470);
   U689 : MUX2_X1 port map( A => n4386, B => DATAIN(3), S => n120, Z => n3469);
   U690 : MUX2_X1 port map( A => n4385, B => DATAIN(2), S => n120, Z => n3468);
   U691 : MUX2_X1 port map( A => n4384, B => DATAIN(1), S => n120, Z => n3467);
   U692 : MUX2_X1 port map( A => n4383, B => DATAIN(0), S => n120, Z => n3466);
   U693 : AND2_X1 port map( A1 => n768, A2 => n764, ZN => n767);
   U694 : MUX2_X1 port map( A => n769, B => DATAIN(31), S => n125, Z => n3465);
   U695 : MUX2_X1 port map( A => n771, B => DATAIN(30), S => n125, Z => n3464);
   U696 : MUX2_X1 port map( A => n772, B => DATAIN(29), S => n125, Z => n3463);
   U697 : MUX2_X1 port map( A => n773, B => DATAIN(28), S => n125, Z => n3462);
   U698 : MUX2_X1 port map( A => n774, B => DATAIN(27), S => n125, Z => n3461);
   U699 : MUX2_X1 port map( A => n775, B => DATAIN(26), S => n125, Z => n3460);
   U700 : MUX2_X1 port map( A => n776, B => DATAIN(25), S => n125, Z => n3459);
   U701 : MUX2_X1 port map( A => n777, B => DATAIN(24), S => n125, Z => n3458);
   U702 : MUX2_X1 port map( A => n778, B => DATAIN(23), S => n124, Z => n3457);
   U703 : MUX2_X1 port map( A => n779, B => DATAIN(22), S => n124, Z => n3456);
   U704 : MUX2_X1 port map( A => n780, B => DATAIN(21), S => n124, Z => n3455);
   U705 : MUX2_X1 port map( A => n781, B => DATAIN(20), S => n124, Z => n3454);
   U706 : MUX2_X1 port map( A => n782, B => DATAIN(19), S => n124, Z => n3453);
   U707 : MUX2_X1 port map( A => n783, B => DATAIN(18), S => n124, Z => n3452);
   U708 : MUX2_X1 port map( A => n784, B => DATAIN(17), S => n124, Z => n3451);
   U709 : MUX2_X1 port map( A => n785, B => DATAIN(16), S => n124, Z => n3450);
   U710 : MUX2_X1 port map( A => n786, B => DATAIN(15), S => n124, Z => n3449);
   U711 : MUX2_X1 port map( A => n787, B => DATAIN(14), S => n124, Z => n3448);
   U712 : MUX2_X1 port map( A => n788, B => DATAIN(13), S => n124, Z => n3447);
   U713 : MUX2_X1 port map( A => n789, B => DATAIN(12), S => n124, Z => n3446);
   U714 : MUX2_X1 port map( A => n790, B => DATAIN(11), S => n123, Z => n3445);
   U715 : MUX2_X1 port map( A => n791, B => DATAIN(10), S => n123, Z => n3444);
   U716 : MUX2_X1 port map( A => n792, B => DATAIN(9), S => n123, Z => n3443);
   U717 : MUX2_X1 port map( A => n793, B => DATAIN(8), S => n123, Z => n3442);
   U718 : MUX2_X1 port map( A => n794, B => DATAIN(7), S => n123, Z => n3441);
   U719 : MUX2_X1 port map( A => n795, B => DATAIN(6), S => n123, Z => n3440);
   U720 : MUX2_X1 port map( A => n796, B => DATAIN(5), S => n123, Z => n3439);
   U721 : MUX2_X1 port map( A => n797, B => DATAIN(4), S => n123, Z => n3438);
   U722 : MUX2_X1 port map( A => n798, B => DATAIN(3), S => n123, Z => n3437);
   U723 : MUX2_X1 port map( A => n799, B => DATAIN(2), S => n123, Z => n3436);
   U724 : MUX2_X1 port map( A => n800, B => DATAIN(1), S => n123, Z => n3435);
   U725 : MUX2_X1 port map( A => n801, B => DATAIN(0), S => n123, Z => n3434);
   U726 : AND2_X1 port map( A1 => n802, A2 => n764, ZN => n770);
   U727 : MUX2_X1 port map( A => n803, B => DATAIN(31), S => n128, Z => n3433);
   U728 : MUX2_X1 port map( A => n805, B => DATAIN(30), S => n128, Z => n3432);
   U729 : MUX2_X1 port map( A => n806, B => DATAIN(29), S => n128, Z => n3431);
   U730 : MUX2_X1 port map( A => n807, B => DATAIN(28), S => n128, Z => n3430);
   U731 : MUX2_X1 port map( A => n808, B => DATAIN(27), S => n128, Z => n3429);
   U732 : MUX2_X1 port map( A => n809, B => DATAIN(26), S => n128, Z => n3428);
   U733 : MUX2_X1 port map( A => n810, B => DATAIN(25), S => n128, Z => n3427);
   U734 : MUX2_X1 port map( A => n811, B => DATAIN(24), S => n128, Z => n3426);
   U735 : MUX2_X1 port map( A => n812, B => DATAIN(23), S => n127, Z => n3425);
   U736 : MUX2_X1 port map( A => n813, B => DATAIN(22), S => n127, Z => n3424);
   U737 : MUX2_X1 port map( A => n814, B => DATAIN(21), S => n127, Z => n3423);
   U738 : MUX2_X1 port map( A => n815, B => DATAIN(20), S => n127, Z => n3422);
   U739 : MUX2_X1 port map( A => n816, B => DATAIN(19), S => n127, Z => n3421);
   U740 : MUX2_X1 port map( A => n817, B => DATAIN(18), S => n127, Z => n3420);
   U741 : MUX2_X1 port map( A => n818, B => DATAIN(17), S => n127, Z => n3419);
   U742 : MUX2_X1 port map( A => n819, B => DATAIN(16), S => n127, Z => n3418);
   U743 : MUX2_X1 port map( A => n820, B => DATAIN(15), S => n127, Z => n3417);
   U744 : MUX2_X1 port map( A => n821, B => DATAIN(14), S => n127, Z => n3416);
   U745 : MUX2_X1 port map( A => n822, B => DATAIN(13), S => n127, Z => n3415);
   U746 : MUX2_X1 port map( A => n823, B => DATAIN(12), S => n127, Z => n3414);
   U747 : MUX2_X1 port map( A => n824, B => DATAIN(11), S => n126, Z => n3413);
   U748 : MUX2_X1 port map( A => n825, B => DATAIN(10), S => n126, Z => n3412);
   U749 : MUX2_X1 port map( A => n826, B => DATAIN(9), S => n126, Z => n3411);
   U750 : MUX2_X1 port map( A => n827, B => DATAIN(8), S => n126, Z => n3410);
   U751 : MUX2_X1 port map( A => n828, B => DATAIN(7), S => n126, Z => n3409);
   U752 : MUX2_X1 port map( A => n829, B => DATAIN(6), S => n126, Z => n3408);
   U753 : MUX2_X1 port map( A => n830, B => DATAIN(5), S => n126, Z => n3407);
   U754 : MUX2_X1 port map( A => n831, B => DATAIN(4), S => n126, Z => n3406);
   U755 : MUX2_X1 port map( A => n832, B => DATAIN(3), S => n126, Z => n3405);
   U756 : MUX2_X1 port map( A => n833, B => DATAIN(2), S => n126, Z => n3404);
   U757 : MUX2_X1 port map( A => n834, B => DATAIN(1), S => n126, Z => n3403);
   U758 : MUX2_X1 port map( A => n835, B => DATAIN(0), S => n126, Z => n3402);
   U759 : AND2_X1 port map( A1 => n836, A2 => n764, ZN => n804);
   U760 : MUX2_X1 port map( A => n4382, B => DATAIN(31), S => n131, Z => n3401)
                           ;
   U761 : MUX2_X1 port map( A => n4381, B => DATAIN(30), S => n131, Z => n3400)
                           ;
   U762 : MUX2_X1 port map( A => n4380, B => DATAIN(29), S => n131, Z => n3399)
                           ;
   U763 : MUX2_X1 port map( A => n4379, B => DATAIN(28), S => n131, Z => n3398)
                           ;
   U764 : MUX2_X1 port map( A => n4378, B => DATAIN(27), S => n131, Z => n3397)
                           ;
   U765 : MUX2_X1 port map( A => n4377, B => DATAIN(26), S => n131, Z => n3396)
                           ;
   U766 : MUX2_X1 port map( A => n4376, B => DATAIN(25), S => n131, Z => n3395)
                           ;
   U767 : MUX2_X1 port map( A => n4375, B => DATAIN(24), S => n131, Z => n3394)
                           ;
   U768 : MUX2_X1 port map( A => n4374, B => DATAIN(23), S => n130, Z => n3393)
                           ;
   U769 : MUX2_X1 port map( A => n4373, B => DATAIN(22), S => n130, Z => n3392)
                           ;
   U770 : MUX2_X1 port map( A => n4372, B => DATAIN(21), S => n130, Z => n3391)
                           ;
   U771 : MUX2_X1 port map( A => n4371, B => DATAIN(20), S => n130, Z => n3390)
                           ;
   U772 : MUX2_X1 port map( A => n4370, B => DATAIN(19), S => n130, Z => n3389)
                           ;
   U773 : MUX2_X1 port map( A => n4369, B => DATAIN(18), S => n130, Z => n3388)
                           ;
   U774 : MUX2_X1 port map( A => n4368, B => DATAIN(17), S => n130, Z => n3387)
                           ;
   U775 : MUX2_X1 port map( A => n4367, B => DATAIN(16), S => n130, Z => n3386)
                           ;
   U776 : MUX2_X1 port map( A => n4366, B => DATAIN(15), S => n130, Z => n3385)
                           ;
   U777 : MUX2_X1 port map( A => n4365, B => DATAIN(14), S => n130, Z => n3384)
                           ;
   U778 : MUX2_X1 port map( A => n4364, B => DATAIN(13), S => n130, Z => n3383)
                           ;
   U779 : MUX2_X1 port map( A => n4363, B => DATAIN(12), S => n130, Z => n3382)
                           ;
   U780 : MUX2_X1 port map( A => n4362, B => DATAIN(11), S => n129, Z => n3381)
                           ;
   U781 : MUX2_X1 port map( A => n4361, B => DATAIN(10), S => n129, Z => n3380)
                           ;
   U782 : MUX2_X1 port map( A => n4360, B => DATAIN(9), S => n129, Z => n3379);
   U783 : MUX2_X1 port map( A => n4359, B => DATAIN(8), S => n129, Z => n3378);
   U784 : MUX2_X1 port map( A => n4358, B => DATAIN(7), S => n129, Z => n3377);
   U785 : MUX2_X1 port map( A => n4357, B => DATAIN(6), S => n129, Z => n3376);
   U786 : MUX2_X1 port map( A => n4356, B => DATAIN(5), S => n129, Z => n3375);
   U787 : MUX2_X1 port map( A => n4355, B => DATAIN(4), S => n129, Z => n3374);
   U788 : MUX2_X1 port map( A => n4354, B => DATAIN(3), S => n129, Z => n3373);
   U789 : MUX2_X1 port map( A => n4353, B => DATAIN(2), S => n129, Z => n3372);
   U790 : MUX2_X1 port map( A => n4352, B => DATAIN(1), S => n129, Z => n3371);
   U791 : MUX2_X1 port map( A => n4351, B => DATAIN(0), S => n129, Z => n3370);
   U792 : AND2_X1 port map( A1 => n870, A2 => n764, ZN => n869);
   U793 : MUX2_X1 port map( A => n4350, B => DATAIN(31), S => n134, Z => n3369)
                           ;
   U794 : MUX2_X1 port map( A => n4349, B => DATAIN(30), S => n134, Z => n3368)
                           ;
   U795 : MUX2_X1 port map( A => n4348, B => DATAIN(29), S => n134, Z => n3367)
                           ;
   U796 : MUX2_X1 port map( A => n4347, B => DATAIN(28), S => n134, Z => n3366)
                           ;
   U797 : MUX2_X1 port map( A => n4346, B => DATAIN(27), S => n134, Z => n3365)
                           ;
   U798 : MUX2_X1 port map( A => n4345, B => DATAIN(26), S => n134, Z => n3364)
                           ;
   U799 : MUX2_X1 port map( A => n4344, B => DATAIN(25), S => n134, Z => n3363)
                           ;
   U800 : MUX2_X1 port map( A => n4343, B => DATAIN(24), S => n134, Z => n3362)
                           ;
   U801 : MUX2_X1 port map( A => n4342, B => DATAIN(23), S => n133, Z => n3361)
                           ;
   U802 : MUX2_X1 port map( A => n4341, B => DATAIN(22), S => n133, Z => n3360)
                           ;
   U803 : MUX2_X1 port map( A => n4340, B => DATAIN(21), S => n133, Z => n3359)
                           ;
   U804 : MUX2_X1 port map( A => n4339, B => DATAIN(20), S => n133, Z => n3358)
                           ;
   U805 : MUX2_X1 port map( A => n4338, B => DATAIN(19), S => n133, Z => n3357)
                           ;
   U806 : MUX2_X1 port map( A => n4337, B => DATAIN(18), S => n133, Z => n3356)
                           ;
   U807 : MUX2_X1 port map( A => n4336, B => DATAIN(17), S => n133, Z => n3355)
                           ;
   U808 : MUX2_X1 port map( A => n4335, B => DATAIN(16), S => n133, Z => n3354)
                           ;
   U809 : MUX2_X1 port map( A => n4334, B => DATAIN(15), S => n133, Z => n3353)
                           ;
   U810 : MUX2_X1 port map( A => n4333, B => DATAIN(14), S => n133, Z => n3352)
                           ;
   U811 : MUX2_X1 port map( A => n4332, B => DATAIN(13), S => n133, Z => n3351)
                           ;
   U812 : MUX2_X1 port map( A => n4331, B => DATAIN(12), S => n133, Z => n3350)
                           ;
   U813 : MUX2_X1 port map( A => n4330, B => DATAIN(11), S => n132, Z => n3349)
                           ;
   U814 : MUX2_X1 port map( A => n4329, B => DATAIN(10), S => n132, Z => n3348)
                           ;
   U815 : MUX2_X1 port map( A => n4328, B => DATAIN(9), S => n132, Z => n3347);
   U816 : MUX2_X1 port map( A => n4327, B => DATAIN(8), S => n132, Z => n3346);
   U817 : MUX2_X1 port map( A => n4326, B => DATAIN(7), S => n132, Z => n3345);
   U818 : MUX2_X1 port map( A => n4325, B => DATAIN(6), S => n132, Z => n3344);
   U819 : MUX2_X1 port map( A => n4324, B => DATAIN(5), S => n132, Z => n3343);
   U820 : MUX2_X1 port map( A => n4323, B => DATAIN(4), S => n132, Z => n3342);
   U821 : MUX2_X1 port map( A => n4322, B => DATAIN(3), S => n132, Z => n3341);
   U822 : MUX2_X1 port map( A => n4321, B => DATAIN(2), S => n132, Z => n3340);
   U823 : MUX2_X1 port map( A => n4320, B => DATAIN(1), S => n132, Z => n3339);
   U824 : MUX2_X1 port map( A => n4319, B => DATAIN(0), S => n132, Z => n3338);
   U825 : AND2_X1 port map( A1 => n872, A2 => n764, ZN => n871);
   U826 : AND3_X1 port map( A1 => n873, A2 => n874, A3 => n875, ZN => n764);
   U827 : INV_X1 port map( A => n876, ZN => n3337);
   U828 : MUX2_X1 port map( A => n229, B => n593, S => n137, Z => n876);
   U829 : INV_X1 port map( A => n878, ZN => n3336);
   U830 : MUX2_X1 port map( A => n230, B => n592, S => n137, Z => n878);
   U831 : INV_X1 port map( A => n879, ZN => n3335);
   U832 : MUX2_X1 port map( A => n231, B => n591, S => n137, Z => n879);
   U833 : INV_X1 port map( A => n880, ZN => n3334);
   U834 : MUX2_X1 port map( A => n232, B => n590, S => n137, Z => n880);
   U835 : INV_X1 port map( A => n881, ZN => n3333);
   U836 : MUX2_X1 port map( A => n233, B => n589, S => n137, Z => n881);
   U837 : INV_X1 port map( A => n882, ZN => n3332);
   U838 : MUX2_X1 port map( A => n234, B => n588, S => n137, Z => n882);
   U839 : INV_X1 port map( A => n883, ZN => n3331);
   U840 : MUX2_X1 port map( A => n235, B => n587, S => n137, Z => n883);
   U841 : INV_X1 port map( A => n884, ZN => n3330);
   U842 : MUX2_X1 port map( A => n236, B => n586, S => n137, Z => n884);
   U843 : INV_X1 port map( A => n885, ZN => n3329);
   U844 : MUX2_X1 port map( A => n237, B => n585, S => n136, Z => n885);
   U845 : INV_X1 port map( A => n886, ZN => n3328);
   U846 : MUX2_X1 port map( A => n238, B => n584, S => n136, Z => n886);
   U847 : INV_X1 port map( A => n887, ZN => n3327);
   U848 : MUX2_X1 port map( A => n239, B => n583, S => n136, Z => n887);
   U849 : INV_X1 port map( A => n888, ZN => n3326);
   U850 : MUX2_X1 port map( A => n240, B => n582, S => n136, Z => n888);
   U851 : INV_X1 port map( A => n889, ZN => n3325);
   U852 : MUX2_X1 port map( A => n241, B => n581, S => n136, Z => n889);
   U853 : INV_X1 port map( A => n890, ZN => n3324);
   U854 : MUX2_X1 port map( A => n242, B => n580, S => n136, Z => n890);
   U855 : INV_X1 port map( A => n891, ZN => n3323);
   U856 : MUX2_X1 port map( A => n243, B => n579, S => n136, Z => n891);
   U857 : INV_X1 port map( A => n892, ZN => n3322);
   U858 : MUX2_X1 port map( A => n244, B => n578, S => n136, Z => n892);
   U859 : INV_X1 port map( A => n893, ZN => n3321);
   U860 : MUX2_X1 port map( A => n245, B => n577, S => n136, Z => n893);
   U861 : INV_X1 port map( A => n894, ZN => n3320);
   U862 : MUX2_X1 port map( A => n246, B => n576, S => n136, Z => n894);
   U863 : INV_X1 port map( A => n895, ZN => n3319);
   U864 : MUX2_X1 port map( A => n247, B => n575, S => n136, Z => n895);
   U865 : INV_X1 port map( A => n896, ZN => n3318);
   U866 : MUX2_X1 port map( A => n248, B => n574, S => n136, Z => n896);
   U867 : INV_X1 port map( A => n897, ZN => n3317);
   U868 : MUX2_X1 port map( A => n249, B => n573, S => n135, Z => n897);
   U869 : INV_X1 port map( A => n898, ZN => n3316);
   U870 : MUX2_X1 port map( A => n250, B => n572, S => n135, Z => n898);
   U871 : INV_X1 port map( A => n899, ZN => n3315);
   U872 : MUX2_X1 port map( A => n251, B => n571, S => n135, Z => n899);
   U873 : INV_X1 port map( A => n900, ZN => n3314);
   U874 : MUX2_X1 port map( A => n252, B => n570, S => n135, Z => n900);
   U875 : INV_X1 port map( A => n901, ZN => n3313);
   U876 : MUX2_X1 port map( A => n253, B => n569, S => n135, Z => n901);
   U877 : INV_X1 port map( A => n902, ZN => n3312);
   U878 : MUX2_X1 port map( A => n254, B => n568, S => n135, Z => n902);
   U879 : INV_X1 port map( A => n903, ZN => n3311);
   U880 : MUX2_X1 port map( A => n255, B => n567, S => n135, Z => n903);
   U881 : INV_X1 port map( A => n904, ZN => n3310);
   U882 : MUX2_X1 port map( A => n256, B => n566, S => n135, Z => n904);
   U883 : INV_X1 port map( A => n905, ZN => n3309);
   U884 : MUX2_X1 port map( A => n257, B => n565, S => n135, Z => n905);
   U885 : INV_X1 port map( A => n906, ZN => n3308);
   U886 : MUX2_X1 port map( A => n258, B => n564, S => n135, Z => n906);
   U887 : INV_X1 port map( A => n907, ZN => n3307);
   U888 : MUX2_X1 port map( A => n259, B => n563, S => n135, Z => n907);
   U889 : INV_X1 port map( A => n908, ZN => n3306);
   U890 : MUX2_X1 port map( A => n260, B => n562, S => n135, Z => n908);
   U891 : AND2_X1 port map( A1 => n909, A2 => n910, ZN => n877);
   U892 : INV_X1 port map( A => n911, ZN => n3305);
   U893 : MUX2_X1 port map( A => n261, B => n593, S => n140, Z => n911);
   U894 : INV_X1 port map( A => n913, ZN => n3304);
   U895 : MUX2_X1 port map( A => n262, B => n592, S => n140, Z => n913);
   U896 : INV_X1 port map( A => n914, ZN => n3303);
   U897 : MUX2_X1 port map( A => n263, B => n591, S => n140, Z => n914);
   U898 : INV_X1 port map( A => n915, ZN => n3302);
   U899 : MUX2_X1 port map( A => n264, B => n590, S => n140, Z => n915);
   U900 : INV_X1 port map( A => n916, ZN => n3301);
   U901 : MUX2_X1 port map( A => n265, B => n589, S => n140, Z => n916);
   U902 : INV_X1 port map( A => n917, ZN => n3300);
   U903 : MUX2_X1 port map( A => n266, B => n588, S => n140, Z => n917);
   U904 : INV_X1 port map( A => n918, ZN => n3299);
   U905 : MUX2_X1 port map( A => n267, B => n587, S => n140, Z => n918);
   U906 : INV_X1 port map( A => n919, ZN => n3298);
   U907 : MUX2_X1 port map( A => n268, B => n586, S => n140, Z => n919);
   U908 : INV_X1 port map( A => n920, ZN => n3297);
   U909 : MUX2_X1 port map( A => n269, B => n585, S => n139, Z => n920);
   U910 : INV_X1 port map( A => n921, ZN => n3296);
   U911 : MUX2_X1 port map( A => n270, B => n584, S => n139, Z => n921);
   U912 : INV_X1 port map( A => n922, ZN => n3295);
   U913 : MUX2_X1 port map( A => n271, B => n583, S => n139, Z => n922);
   U914 : INV_X1 port map( A => n923, ZN => n3294);
   U915 : MUX2_X1 port map( A => n272, B => n582, S => n139, Z => n923);
   U916 : INV_X1 port map( A => n924, ZN => n3293);
   U917 : MUX2_X1 port map( A => n273, B => n581, S => n139, Z => n924);
   U918 : INV_X1 port map( A => n925, ZN => n3292);
   U919 : MUX2_X1 port map( A => n274, B => n580, S => n139, Z => n925);
   U920 : INV_X1 port map( A => n926, ZN => n3291);
   U921 : MUX2_X1 port map( A => n275, B => n579, S => n139, Z => n926);
   U922 : INV_X1 port map( A => n927, ZN => n3290);
   U923 : MUX2_X1 port map( A => n276, B => n578, S => n139, Z => n927);
   U924 : INV_X1 port map( A => n928, ZN => n3289);
   U925 : MUX2_X1 port map( A => n277, B => n577, S => n139, Z => n928);
   U926 : INV_X1 port map( A => n929, ZN => n3288);
   U927 : MUX2_X1 port map( A => n278, B => n576, S => n139, Z => n929);
   U928 : INV_X1 port map( A => n930, ZN => n3287);
   U929 : MUX2_X1 port map( A => n279, B => n575, S => n139, Z => n930);
   U930 : INV_X1 port map( A => n931, ZN => n3286);
   U931 : MUX2_X1 port map( A => n280, B => n574, S => n139, Z => n931);
   U932 : INV_X1 port map( A => n932, ZN => n3285);
   U933 : MUX2_X1 port map( A => n281, B => n573, S => n138, Z => n932);
   U934 : INV_X1 port map( A => n965, ZN => n3284);
   U935 : MUX2_X1 port map( A => n282, B => n572, S => n138, Z => n965);
   U936 : INV_X1 port map( A => n966, ZN => n3283);
   U937 : MUX2_X1 port map( A => n283, B => n571, S => n138, Z => n966);
   U938 : INV_X1 port map( A => n967, ZN => n3282);
   U939 : MUX2_X1 port map( A => n284, B => n570, S => n138, Z => n967);
   U940 : INV_X1 port map( A => n968, ZN => n3281);
   U941 : MUX2_X1 port map( A => n285, B => n569, S => n138, Z => n968);
   U942 : INV_X1 port map( A => n969, ZN => n3280);
   U943 : MUX2_X1 port map( A => n286, B => n568, S => n138, Z => n969);
   U944 : INV_X1 port map( A => n970, ZN => n3279);
   U945 : MUX2_X1 port map( A => n287, B => n567, S => n138, Z => n970);
   U946 : INV_X1 port map( A => n971, ZN => n3278);
   U947 : MUX2_X1 port map( A => n288, B => n566, S => n138, Z => n971);
   U948 : INV_X1 port map( A => n972, ZN => n3277);
   U949 : MUX2_X1 port map( A => n289, B => n565, S => n138, Z => n972);
   U950 : INV_X1 port map( A => n973, ZN => n3276);
   U951 : MUX2_X1 port map( A => n290, B => n564, S => n138, Z => n973);
   U952 : INV_X1 port map( A => n974, ZN => n3275);
   U953 : MUX2_X1 port map( A => n291, B => n563, S => n138, Z => n974);
   U954 : INV_X1 port map( A => n975, ZN => n3274);
   U955 : MUX2_X1 port map( A => n292, B => n562, S => n138, Z => n975);
   U956 : AND2_X1 port map( A1 => n909, A2 => n763, ZN => n912);
   U957 : MUX2_X1 port map( A => n4318, B => DATAIN(31), S => n143, Z => n3273)
                           ;
   U958 : MUX2_X1 port map( A => n4317, B => DATAIN(30), S => n143, Z => n3272)
                           ;
   U959 : MUX2_X1 port map( A => n4316, B => DATAIN(29), S => n143, Z => n3271)
                           ;
   U960 : MUX2_X1 port map( A => n4315, B => DATAIN(28), S => n143, Z => n3270)
                           ;
   U961 : MUX2_X1 port map( A => n4314, B => DATAIN(27), S => n143, Z => n3269)
                           ;
   U962 : MUX2_X1 port map( A => n4313, B => DATAIN(26), S => n143, Z => n3268)
                           ;
   U963 : MUX2_X1 port map( A => n4312, B => DATAIN(25), S => n143, Z => n3267)
                           ;
   U964 : MUX2_X1 port map( A => n4311, B => DATAIN(24), S => n143, Z => n3266)
                           ;
   U965 : MUX2_X1 port map( A => n4310, B => DATAIN(23), S => n142, Z => n3265)
                           ;
   U966 : MUX2_X1 port map( A => n4309, B => DATAIN(22), S => n142, Z => n3264)
                           ;
   U967 : MUX2_X1 port map( A => n4308, B => DATAIN(21), S => n142, Z => n3263)
                           ;
   U968 : MUX2_X1 port map( A => n4307, B => DATAIN(20), S => n142, Z => n3262)
                           ;
   U969 : MUX2_X1 port map( A => n4306, B => DATAIN(19), S => n142, Z => n3261)
                           ;
   U970 : MUX2_X1 port map( A => n4305, B => DATAIN(18), S => n142, Z => n3260)
                           ;
   U971 : MUX2_X1 port map( A => n4304, B => DATAIN(17), S => n142, Z => n3259)
                           ;
   U972 : MUX2_X1 port map( A => n4303, B => DATAIN(16), S => n142, Z => n3258)
                           ;
   U973 : MUX2_X1 port map( A => n4302, B => DATAIN(15), S => n142, Z => n3257)
                           ;
   U974 : MUX2_X1 port map( A => n4301, B => DATAIN(14), S => n142, Z => n3256)
                           ;
   U975 : MUX2_X1 port map( A => n4300, B => DATAIN(13), S => n142, Z => n3255)
                           ;
   U976 : MUX2_X1 port map( A => n4299, B => DATAIN(12), S => n142, Z => n3254)
                           ;
   U977 : MUX2_X1 port map( A => n4298, B => DATAIN(11), S => n141, Z => n3253)
                           ;
   U978 : MUX2_X1 port map( A => n4297, B => DATAIN(10), S => n141, Z => n3252)
                           ;
   U979 : MUX2_X1 port map( A => n4296, B => DATAIN(9), S => n141, Z => n3251);
   U980 : MUX2_X1 port map( A => n4295, B => DATAIN(8), S => n141, Z => n3250);
   U981 : MUX2_X1 port map( A => n4294, B => DATAIN(7), S => n141, Z => n3249);
   U982 : MUX2_X1 port map( A => n4293, B => DATAIN(6), S => n141, Z => n3248);
   U983 : MUX2_X1 port map( A => n4292, B => DATAIN(5), S => n141, Z => n3247);
   U984 : MUX2_X1 port map( A => n4291, B => DATAIN(4), S => n141, Z => n3246);
   U985 : MUX2_X1 port map( A => n4290, B => DATAIN(3), S => n141, Z => n3245);
   U986 : MUX2_X1 port map( A => n4289, B => DATAIN(2), S => n141, Z => n3244);
   U987 : MUX2_X1 port map( A => n4288, B => DATAIN(1), S => n141, Z => n3243);
   U988 : MUX2_X1 port map( A => n4287, B => DATAIN(0), S => n141, Z => n3242);
   U989 : AND2_X1 port map( A1 => n909, A2 => n766, ZN => n976);
   U990 : MUX2_X1 port map( A => n4286, B => DATAIN(31), S => n146, Z => n3241)
                           ;
   U991 : MUX2_X1 port map( A => n4285, B => DATAIN(30), S => n146, Z => n3240)
                           ;
   U992 : MUX2_X1 port map( A => n4284, B => DATAIN(29), S => n146, Z => n3239)
                           ;
   U993 : MUX2_X1 port map( A => n4283, B => DATAIN(28), S => n146, Z => n3238)
                           ;
   U994 : MUX2_X1 port map( A => n4282, B => DATAIN(27), S => n146, Z => n3237)
                           ;
   U995 : MUX2_X1 port map( A => n4281, B => DATAIN(26), S => n146, Z => n3236)
                           ;
   U996 : MUX2_X1 port map( A => n4280, B => DATAIN(25), S => n146, Z => n3235)
                           ;
   U997 : MUX2_X1 port map( A => n4279, B => DATAIN(24), S => n146, Z => n3234)
                           ;
   U998 : MUX2_X1 port map( A => n4278, B => DATAIN(23), S => n145, Z => n3233)
                           ;
   U999 : MUX2_X1 port map( A => n4277, B => DATAIN(22), S => n145, Z => n3232)
                           ;
   U1000 : MUX2_X1 port map( A => n4276, B => DATAIN(21), S => n145, Z => n3231
                           );
   U1001 : MUX2_X1 port map( A => n4275, B => DATAIN(20), S => n145, Z => n3230
                           );
   U1002 : MUX2_X1 port map( A => n4274, B => DATAIN(19), S => n145, Z => n3229
                           );
   U1003 : MUX2_X1 port map( A => n4273, B => DATAIN(18), S => n145, Z => n3228
                           );
   U1004 : MUX2_X1 port map( A => n4272, B => DATAIN(17), S => n145, Z => n3227
                           );
   U1005 : MUX2_X1 port map( A => n4271, B => DATAIN(16), S => n145, Z => n3226
                           );
   U1006 : MUX2_X1 port map( A => n4270, B => DATAIN(15), S => n145, Z => n3225
                           );
   U1007 : MUX2_X1 port map( A => n4269, B => DATAIN(14), S => n145, Z => n3224
                           );
   U1008 : MUX2_X1 port map( A => n4268, B => DATAIN(13), S => n145, Z => n3223
                           );
   U1009 : MUX2_X1 port map( A => n4267, B => DATAIN(12), S => n145, Z => n3222
                           );
   U1010 : MUX2_X1 port map( A => n4266, B => DATAIN(11), S => n144, Z => n3221
                           );
   U1011 : MUX2_X1 port map( A => n4265, B => DATAIN(10), S => n144, Z => n3220
                           );
   U1012 : MUX2_X1 port map( A => n4264, B => DATAIN(9), S => n144, Z => n3219)
                           ;
   U1013 : MUX2_X1 port map( A => n4263, B => DATAIN(8), S => n144, Z => n3218)
                           ;
   U1014 : MUX2_X1 port map( A => n4262, B => DATAIN(7), S => n144, Z => n3217)
                           ;
   U1015 : MUX2_X1 port map( A => n4261, B => DATAIN(6), S => n144, Z => n3216)
                           ;
   U1016 : MUX2_X1 port map( A => n4260, B => DATAIN(5), S => n144, Z => n3215)
                           ;
   U1017 : MUX2_X1 port map( A => n4259, B => DATAIN(4), S => n144, Z => n3214)
                           ;
   U1018 : MUX2_X1 port map( A => n4258, B => DATAIN(3), S => n144, Z => n3213)
                           ;
   U1019 : MUX2_X1 port map( A => n4257, B => DATAIN(2), S => n144, Z => n3212)
                           ;
   U1020 : MUX2_X1 port map( A => n4256, B => DATAIN(1), S => n144, Z => n3211)
                           ;
   U1021 : MUX2_X1 port map( A => n4255, B => DATAIN(0), S => n144, Z => n3210)
                           ;
   U1022 : AND2_X1 port map( A1 => n909, A2 => n768, ZN => n977);
   U1023 : INV_X1 port map( A => n978, ZN => n3209);
   U1024 : MUX2_X1 port map( A => n357, B => n593, S => n149, Z => n978);
   U1025 : INV_X1 port map( A => n980, ZN => n3208);
   U1026 : MUX2_X1 port map( A => n358, B => n592, S => n149, Z => n980);
   U1027 : INV_X1 port map( A => n981, ZN => n3207);
   U1028 : MUX2_X1 port map( A => n359, B => n591, S => n149, Z => n981);
   U1029 : INV_X1 port map( A => n982, ZN => n3206);
   U1030 : MUX2_X1 port map( A => n360, B => n590, S => n149, Z => n982);
   U1031 : INV_X1 port map( A => n983, ZN => n3205);
   U1032 : MUX2_X1 port map( A => n361, B => n589, S => n149, Z => n983);
   U1033 : INV_X1 port map( A => n984, ZN => n3204);
   U1034 : MUX2_X1 port map( A => n362, B => n588, S => n149, Z => n984);
   U1035 : INV_X1 port map( A => n985, ZN => n3203);
   U1036 : MUX2_X1 port map( A => n363, B => n587, S => n149, Z => n985);
   U1037 : INV_X1 port map( A => n986, ZN => n3202);
   U1038 : MUX2_X1 port map( A => n364, B => n586, S => n149, Z => n986);
   U1039 : INV_X1 port map( A => n987, ZN => n3201);
   U1040 : MUX2_X1 port map( A => n365, B => n585, S => n148, Z => n987);
   U1041 : INV_X1 port map( A => n988, ZN => n3200);
   U1042 : MUX2_X1 port map( A => n366, B => n584, S => n148, Z => n988);
   U1043 : INV_X1 port map( A => n989, ZN => n3199);
   U1044 : MUX2_X1 port map( A => n367, B => n583, S => n148, Z => n989);
   U1045 : INV_X1 port map( A => n990, ZN => n3198);
   U1046 : MUX2_X1 port map( A => n368, B => n582, S => n148, Z => n990);
   U1047 : INV_X1 port map( A => n991, ZN => n3197);
   U1048 : MUX2_X1 port map( A => n369, B => n581, S => n148, Z => n991);
   U1049 : INV_X1 port map( A => n992, ZN => n3196);
   U1050 : MUX2_X1 port map( A => n370, B => n580, S => n148, Z => n992);
   U1051 : INV_X1 port map( A => n993, ZN => n3195);
   U1052 : MUX2_X1 port map( A => n371, B => n579, S => n148, Z => n993);
   U1053 : INV_X1 port map( A => n994, ZN => n3194);
   U1054 : MUX2_X1 port map( A => n372, B => n578, S => n148, Z => n994);
   U1055 : INV_X1 port map( A => n995, ZN => n3193);
   U1056 : MUX2_X1 port map( A => n373, B => n577, S => n148, Z => n995);
   U1057 : INV_X1 port map( A => n996, ZN => n3192);
   U1058 : MUX2_X1 port map( A => n374, B => n576, S => n148, Z => n996);
   U1059 : INV_X1 port map( A => n997, ZN => n3191);
   U1060 : MUX2_X1 port map( A => n375, B => n575, S => n148, Z => n997);
   U1061 : INV_X1 port map( A => n998, ZN => n3190);
   U1062 : MUX2_X1 port map( A => n376, B => n574, S => n148, Z => n998);
   U1063 : INV_X1 port map( A => n999, ZN => n3189);
   U1064 : MUX2_X1 port map( A => n377, B => n573, S => n147, Z => n999);
   U1065 : INV_X1 port map( A => n1000, ZN => n3188);
   U1066 : MUX2_X1 port map( A => n378, B => n572, S => n147, Z => n1000);
   U1067 : INV_X1 port map( A => n1001, ZN => n3187);
   U1068 : MUX2_X1 port map( A => n379, B => n571, S => n147, Z => n1001);
   U1069 : INV_X1 port map( A => n1002, ZN => n3186);
   U1070 : MUX2_X1 port map( A => n380, B => n570, S => n147, Z => n1002);
   U1071 : INV_X1 port map( A => n1003, ZN => n3185);
   U1072 : MUX2_X1 port map( A => n381, B => n569, S => n147, Z => n1003);
   U1073 : INV_X1 port map( A => n1004, ZN => n3184);
   U1074 : MUX2_X1 port map( A => n382, B => n568, S => n147, Z => n1004);
   U1075 : INV_X1 port map( A => n1005, ZN => n3183);
   U1076 : MUX2_X1 port map( A => n383, B => n567, S => n147, Z => n1005);
   U1077 : INV_X1 port map( A => n1006, ZN => n3182);
   U1078 : MUX2_X1 port map( A => n384, B => n566, S => n147, Z => n1006);
   U1079 : INV_X1 port map( A => n1007, ZN => n3181);
   U1080 : MUX2_X1 port map( A => n385, B => n565, S => n147, Z => n1007);
   U1081 : INV_X1 port map( A => n1008, ZN => n3180);
   U1082 : MUX2_X1 port map( A => n386, B => n564, S => n147, Z => n1008);
   U1083 : INV_X1 port map( A => n1009, ZN => n3179);
   U1084 : MUX2_X1 port map( A => n387, B => n563, S => n147, Z => n1009);
   U1085 : INV_X1 port map( A => n1010, ZN => n3178);
   U1086 : MUX2_X1 port map( A => n388, B => n562, S => n147, Z => n1010);
   U1087 : AND2_X1 port map( A1 => n909, A2 => n802, ZN => n979);
   U1088 : INV_X1 port map( A => n1011, ZN => n3177);
   U1089 : MUX2_X1 port map( A => n389, B => n593, S => n152, Z => n1011);
   U1090 : INV_X1 port map( A => n1013, ZN => n3176);
   U1091 : MUX2_X1 port map( A => n390, B => n592, S => n152, Z => n1013);
   U1092 : INV_X1 port map( A => n1014, ZN => n3175);
   U1093 : MUX2_X1 port map( A => n391, B => n591, S => n152, Z => n1014);
   U1094 : INV_X1 port map( A => n1015, ZN => n3174);
   U1095 : MUX2_X1 port map( A => n392, B => n590, S => n152, Z => n1015);
   U1096 : INV_X1 port map( A => n1016, ZN => n3173);
   U1097 : MUX2_X1 port map( A => n393, B => n589, S => n152, Z => n1016);
   U1098 : INV_X1 port map( A => n1017, ZN => n3172);
   U1099 : MUX2_X1 port map( A => n394, B => n588, S => n152, Z => n1017);
   U1100 : INV_X1 port map( A => n1018, ZN => n3171);
   U1101 : MUX2_X1 port map( A => n395, B => n587, S => n152, Z => n1018);
   U1102 : INV_X1 port map( A => n1019, ZN => n3170);
   U1103 : MUX2_X1 port map( A => n396, B => n586, S => n152, Z => n1019);
   U1104 : INV_X1 port map( A => n1020, ZN => n3169);
   U1105 : MUX2_X1 port map( A => n397, B => n585, S => n151, Z => n1020);
   U1106 : INV_X1 port map( A => n1021, ZN => n3168);
   U1107 : MUX2_X1 port map( A => n398, B => n584, S => n151, Z => n1021);
   U1108 : INV_X1 port map( A => n1022, ZN => n3167);
   U1109 : MUX2_X1 port map( A => n399, B => n583, S => n151, Z => n1022);
   U1110 : INV_X1 port map( A => n1023, ZN => n3166);
   U1111 : MUX2_X1 port map( A => n400, B => n582, S => n151, Z => n1023);
   U1112 : INV_X1 port map( A => n1024, ZN => n3165);
   U1113 : MUX2_X1 port map( A => n401, B => n581, S => n151, Z => n1024);
   U1114 : INV_X1 port map( A => n1025, ZN => n3164);
   U1115 : MUX2_X1 port map( A => n402, B => n580, S => n151, Z => n1025);
   U1116 : INV_X1 port map( A => n1026, ZN => n3163);
   U1117 : MUX2_X1 port map( A => n403, B => n579, S => n151, Z => n1026);
   U1118 : INV_X1 port map( A => n1027, ZN => n3162);
   U1119 : MUX2_X1 port map( A => n404, B => n578, S => n151, Z => n1027);
   U1120 : INV_X1 port map( A => n1028, ZN => n3161);
   U1121 : MUX2_X1 port map( A => n405, B => n577, S => n151, Z => n1028);
   U1122 : INV_X1 port map( A => n1029, ZN => n3160);
   U1123 : MUX2_X1 port map( A => n406, B => n576, S => n151, Z => n1029);
   U1124 : INV_X1 port map( A => n1030, ZN => n3159);
   U1125 : MUX2_X1 port map( A => n407, B => n575, S => n151, Z => n1030);
   U1126 : INV_X1 port map( A => n1031, ZN => n3158);
   U1127 : MUX2_X1 port map( A => n408, B => n574, S => n151, Z => n1031);
   U1128 : INV_X1 port map( A => n1032, ZN => n3157);
   U1129 : MUX2_X1 port map( A => n409, B => n573, S => n150, Z => n1032);
   U1130 : INV_X1 port map( A => n1033, ZN => n3156);
   U1131 : MUX2_X1 port map( A => n410, B => n572, S => n150, Z => n1033);
   U1132 : INV_X1 port map( A => n1034, ZN => n3155);
   U1133 : MUX2_X1 port map( A => n411, B => n571, S => n150, Z => n1034);
   U1134 : INV_X1 port map( A => n1035, ZN => n3154);
   U1135 : MUX2_X1 port map( A => n412, B => n570, S => n150, Z => n1035);
   U1136 : INV_X1 port map( A => n1036, ZN => n3153);
   U1137 : MUX2_X1 port map( A => n413, B => n569, S => n150, Z => n1036);
   U1138 : INV_X1 port map( A => n1037, ZN => n3152);
   U1139 : MUX2_X1 port map( A => n414, B => n568, S => n150, Z => n1037);
   U1140 : INV_X1 port map( A => n1038, ZN => n3151);
   U1141 : MUX2_X1 port map( A => n415, B => n567, S => n150, Z => n1038);
   U1142 : INV_X1 port map( A => n1039, ZN => n3150);
   U1143 : MUX2_X1 port map( A => n416, B => n566, S => n150, Z => n1039);
   U1144 : INV_X1 port map( A => n1040, ZN => n3149);
   U1145 : MUX2_X1 port map( A => n417, B => n565, S => n150, Z => n1040);
   U1146 : INV_X1 port map( A => n1041, ZN => n3148);
   U1147 : MUX2_X1 port map( A => n418, B => n564, S => n150, Z => n1041);
   U1148 : INV_X1 port map( A => n1042, ZN => n3147);
   U1149 : MUX2_X1 port map( A => n419, B => n563, S => n150, Z => n1042);
   U1150 : INV_X1 port map( A => n1043, ZN => n3146);
   U1151 : MUX2_X1 port map( A => n420, B => n562, S => n150, Z => n1043);
   U1152 : AND2_X1 port map( A1 => n909, A2 => n836, ZN => n1012);
   U1153 : MUX2_X1 port map( A => n4254, B => DATAIN(31), S => n155, Z => n3145
                           );
   U1154 : MUX2_X1 port map( A => n4253, B => DATAIN(30), S => n155, Z => n3144
                           );
   U1155 : MUX2_X1 port map( A => n4252, B => DATAIN(29), S => n155, Z => n3143
                           );
   U1156 : MUX2_X1 port map( A => n4251, B => DATAIN(28), S => n155, Z => n3142
                           );
   U1157 : MUX2_X1 port map( A => n4250, B => DATAIN(27), S => n155, Z => n3141
                           );
   U1158 : MUX2_X1 port map( A => n4249, B => DATAIN(26), S => n155, Z => n3140
                           );
   U1159 : MUX2_X1 port map( A => n4248, B => DATAIN(25), S => n155, Z => n3139
                           );
   U1160 : MUX2_X1 port map( A => n4247, B => DATAIN(24), S => n155, Z => n3138
                           );
   U1161 : MUX2_X1 port map( A => n4246, B => DATAIN(23), S => n154, Z => n3137
                           );
   U1162 : MUX2_X1 port map( A => n4245, B => DATAIN(22), S => n154, Z => n3136
                           );
   U1163 : MUX2_X1 port map( A => n4244, B => DATAIN(21), S => n154, Z => n3135
                           );
   U1164 : MUX2_X1 port map( A => n4243, B => DATAIN(20), S => n154, Z => n3134
                           );
   U1165 : MUX2_X1 port map( A => n4242, B => DATAIN(19), S => n154, Z => n3133
                           );
   U1166 : MUX2_X1 port map( A => n4241, B => DATAIN(18), S => n154, Z => n3132
                           );
   U1167 : MUX2_X1 port map( A => n4240, B => DATAIN(17), S => n154, Z => n3131
                           );
   U1168 : MUX2_X1 port map( A => n4239, B => DATAIN(16), S => n154, Z => n3130
                           );
   U1169 : MUX2_X1 port map( A => n4238, B => DATAIN(15), S => n154, Z => n3129
                           );
   U1170 : MUX2_X1 port map( A => n4237, B => DATAIN(14), S => n154, Z => n3128
                           );
   U1171 : MUX2_X1 port map( A => n4236, B => DATAIN(13), S => n154, Z => n3127
                           );
   U1172 : MUX2_X1 port map( A => n4235, B => DATAIN(12), S => n154, Z => n3126
                           );
   U1173 : MUX2_X1 port map( A => n4234, B => DATAIN(11), S => n153, Z => n3125
                           );
   U1174 : MUX2_X1 port map( A => n4233, B => DATAIN(10), S => n153, Z => n3124
                           );
   U1175 : MUX2_X1 port map( A => n4232, B => DATAIN(9), S => n153, Z => n3123)
                           ;
   U1176 : MUX2_X1 port map( A => n4231, B => DATAIN(8), S => n153, Z => n3122)
                           ;
   U1177 : MUX2_X1 port map( A => n4230, B => DATAIN(7), S => n153, Z => n3121)
                           ;
   U1178 : MUX2_X1 port map( A => n4229, B => DATAIN(6), S => n153, Z => n3120)
                           ;
   U1179 : MUX2_X1 port map( A => n4228, B => DATAIN(5), S => n153, Z => n3119)
                           ;
   U1180 : MUX2_X1 port map( A => n4227, B => DATAIN(4), S => n153, Z => n3118)
                           ;
   U1181 : MUX2_X1 port map( A => n4226, B => DATAIN(3), S => n153, Z => n3117)
                           ;
   U1182 : MUX2_X1 port map( A => n4225, B => DATAIN(2), S => n153, Z => n3116)
                           ;
   U1183 : MUX2_X1 port map( A => n4224, B => DATAIN(1), S => n153, Z => n3115)
                           ;
   U1184 : MUX2_X1 port map( A => n4223, B => DATAIN(0), S => n153, Z => n3114)
                           ;
   U1185 : AND2_X1 port map( A1 => n909, A2 => n870, ZN => n1044);
   U1186 : MUX2_X1 port map( A => n4222, B => DATAIN(31), S => n158, Z => n3113
                           );
   U1187 : MUX2_X1 port map( A => n4221, B => DATAIN(30), S => n158, Z => n3112
                           );
   U1188 : MUX2_X1 port map( A => n4220, B => DATAIN(29), S => n158, Z => n3111
                           );
   U1189 : MUX2_X1 port map( A => n4219, B => DATAIN(28), S => n158, Z => n3110
                           );
   U1190 : MUX2_X1 port map( A => n4218, B => DATAIN(27), S => n158, Z => n3109
                           );
   U1191 : MUX2_X1 port map( A => n4217, B => DATAIN(26), S => n158, Z => n3108
                           );
   U1192 : MUX2_X1 port map( A => n4216, B => DATAIN(25), S => n158, Z => n3107
                           );
   U1193 : MUX2_X1 port map( A => n4215, B => DATAIN(24), S => n158, Z => n3106
                           );
   U1194 : MUX2_X1 port map( A => n4214, B => DATAIN(23), S => n157, Z => n3105
                           );
   U1195 : MUX2_X1 port map( A => n4213, B => DATAIN(22), S => n157, Z => n3104
                           );
   U1196 : MUX2_X1 port map( A => n4212, B => DATAIN(21), S => n157, Z => n3103
                           );
   U1197 : MUX2_X1 port map( A => n4211, B => DATAIN(20), S => n157, Z => n3102
                           );
   U1198 : MUX2_X1 port map( A => n4210, B => DATAIN(19), S => n157, Z => n3101
                           );
   U1199 : MUX2_X1 port map( A => n4209, B => DATAIN(18), S => n157, Z => n3100
                           );
   U1200 : MUX2_X1 port map( A => n4208, B => DATAIN(17), S => n157, Z => n3099
                           );
   U1201 : MUX2_X1 port map( A => n4207, B => DATAIN(16), S => n157, Z => n3098
                           );
   U1202 : MUX2_X1 port map( A => n4206, B => DATAIN(15), S => n157, Z => n3097
                           );
   U1203 : MUX2_X1 port map( A => n4205, B => DATAIN(14), S => n157, Z => n3096
                           );
   U1204 : MUX2_X1 port map( A => n4204, B => DATAIN(13), S => n157, Z => n3095
                           );
   U1205 : MUX2_X1 port map( A => n4203, B => DATAIN(12), S => n157, Z => n3094
                           );
   U1206 : MUX2_X1 port map( A => n4202, B => DATAIN(11), S => n156, Z => n3093
                           );
   U1207 : MUX2_X1 port map( A => n4201, B => DATAIN(10), S => n156, Z => n3092
                           );
   U1208 : MUX2_X1 port map( A => n4200, B => DATAIN(9), S => n156, Z => n3091)
                           ;
   U1209 : MUX2_X1 port map( A => n4199, B => DATAIN(8), S => n156, Z => n3090)
                           ;
   U1210 : MUX2_X1 port map( A => n4198, B => DATAIN(7), S => n156, Z => n3089)
                           ;
   U1211 : MUX2_X1 port map( A => n4197, B => DATAIN(6), S => n156, Z => n3088)
                           ;
   U1212 : MUX2_X1 port map( A => n4196, B => DATAIN(5), S => n156, Z => n3087)
                           ;
   U1213 : MUX2_X1 port map( A => n4195, B => DATAIN(4), S => n156, Z => n3086)
                           ;
   U1214 : MUX2_X1 port map( A => n4194, B => DATAIN(3), S => n156, Z => n3085)
                           ;
   U1215 : MUX2_X1 port map( A => n4193, B => DATAIN(2), S => n156, Z => n3084)
                           ;
   U1216 : MUX2_X1 port map( A => n4192, B => DATAIN(1), S => n156, Z => n3083)
                           ;
   U1217 : MUX2_X1 port map( A => n4191, B => DATAIN(0), S => n156, Z => n3082)
                           ;
   U1218 : AND2_X1 port map( A1 => n909, A2 => n872, ZN => n1045);
   U1219 : AND3_X1 port map( A1 => n875, A2 => n874, A3 => ADD_WR(3), ZN => 
                           n909);
   U1220 : MUX2_X1 port map( A => n1046, B => DATAIN(31), S => n161, Z => n3081
                           );
   U1221 : MUX2_X1 port map( A => n1048, B => DATAIN(30), S => n161, Z => n3080
                           );
   U1222 : MUX2_X1 port map( A => n1049, B => DATAIN(29), S => n161, Z => n3079
                           );
   U1223 : MUX2_X1 port map( A => n1050, B => DATAIN(28), S => n161, Z => n3078
                           );
   U1224 : MUX2_X1 port map( A => n1051, B => DATAIN(27), S => n161, Z => n3077
                           );
   U1225 : MUX2_X1 port map( A => n1052, B => DATAIN(26), S => n161, Z => n3076
                           );
   U1226 : MUX2_X1 port map( A => n1053, B => DATAIN(25), S => n161, Z => n3075
                           );
   U1227 : MUX2_X1 port map( A => n1054, B => DATAIN(24), S => n161, Z => n3074
                           );
   U1228 : MUX2_X1 port map( A => n1055, B => DATAIN(23), S => n160, Z => n3073
                           );
   U1229 : MUX2_X1 port map( A => n1056, B => DATAIN(22), S => n160, Z => n3072
                           );
   U1230 : MUX2_X1 port map( A => n1057, B => DATAIN(21), S => n160, Z => n3071
                           );
   U1231 : MUX2_X1 port map( A => n1058, B => DATAIN(20), S => n160, Z => n3070
                           );
   U1232 : MUX2_X1 port map( A => n1059, B => DATAIN(19), S => n160, Z => n3069
                           );
   U1233 : MUX2_X1 port map( A => n1060, B => DATAIN(18), S => n160, Z => n3068
                           );
   U1234 : MUX2_X1 port map( A => n1061, B => DATAIN(17), S => n160, Z => n3067
                           );
   U1235 : MUX2_X1 port map( A => n1062, B => DATAIN(16), S => n160, Z => n3066
                           );
   U1236 : MUX2_X1 port map( A => n1063, B => DATAIN(15), S => n160, Z => n3065
                           );
   U1237 : MUX2_X1 port map( A => n1064, B => DATAIN(14), S => n160, Z => n3064
                           );
   U1238 : MUX2_X1 port map( A => n1065, B => DATAIN(13), S => n160, Z => n3063
                           );
   U1239 : MUX2_X1 port map( A => n1066, B => DATAIN(12), S => n160, Z => n3062
                           );
   U1240 : MUX2_X1 port map( A => n1067, B => DATAIN(11), S => n159, Z => n3061
                           );
   U1241 : MUX2_X1 port map( A => n1068, B => DATAIN(10), S => n159, Z => n3060
                           );
   U1242 : MUX2_X1 port map( A => n1069, B => DATAIN(9), S => n159, Z => n3059)
                           ;
   U1243 : MUX2_X1 port map( A => n1070, B => DATAIN(8), S => n159, Z => n3058)
                           ;
   U1244 : MUX2_X1 port map( A => n1071, B => DATAIN(7), S => n159, Z => n3057)
                           ;
   U1245 : MUX2_X1 port map( A => n1072, B => DATAIN(6), S => n159, Z => n3056)
                           ;
   U1246 : MUX2_X1 port map( A => n1073, B => DATAIN(5), S => n159, Z => n3055)
                           ;
   U1247 : MUX2_X1 port map( A => n1074, B => DATAIN(4), S => n159, Z => n3054)
                           ;
   U1248 : MUX2_X1 port map( A => n1075, B => DATAIN(3), S => n159, Z => n3053)
                           ;
   U1249 : MUX2_X1 port map( A => n1076, B => DATAIN(2), S => n159, Z => n3052)
                           ;
   U1250 : MUX2_X1 port map( A => n1077, B => DATAIN(1), S => n159, Z => n3051)
                           ;
   U1251 : MUX2_X1 port map( A => n1078, B => DATAIN(0), S => n159, Z => n3050)
                           ;
   U1252 : AND2_X1 port map( A1 => n1079, A2 => n910, ZN => n1047);
   U1253 : INV_X1 port map( A => n1080, ZN => n3049);
   U1254 : MUX2_X1 port map( A => n517, B => n593, S => n164, Z => n1080);
   U1255 : INV_X1 port map( A => n1082, ZN => n3048);
   U1256 : MUX2_X1 port map( A => n518, B => n592, S => n164, Z => n1082);
   U1257 : INV_X1 port map( A => n1083, ZN => n3047);
   U1258 : MUX2_X1 port map( A => n519, B => n591, S => n164, Z => n1083);
   U1259 : INV_X1 port map( A => n1084, ZN => n3046);
   U1260 : MUX2_X1 port map( A => n520, B => n590, S => n164, Z => n1084);
   U1261 : INV_X1 port map( A => n1085, ZN => n3045);
   U1262 : MUX2_X1 port map( A => n521, B => n589, S => n164, Z => n1085);
   U1263 : INV_X1 port map( A => n1086, ZN => n3044);
   U1264 : MUX2_X1 port map( A => n522, B => n588, S => n164, Z => n1086);
   U1265 : INV_X1 port map( A => n1087, ZN => n3043);
   U1266 : MUX2_X1 port map( A => n523, B => n587, S => n164, Z => n1087);
   U1267 : INV_X1 port map( A => n1088, ZN => n3042);
   U1268 : MUX2_X1 port map( A => n524, B => n586, S => n164, Z => n1088);
   U1269 : INV_X1 port map( A => n1089, ZN => n3041);
   U1270 : MUX2_X1 port map( A => n525, B => n585, S => n163, Z => n1089);
   U1271 : INV_X1 port map( A => n1090, ZN => n3040);
   U1272 : MUX2_X1 port map( A => n526, B => n584, S => n163, Z => n1090);
   U1273 : INV_X1 port map( A => n1091, ZN => n3039);
   U1274 : MUX2_X1 port map( A => n527, B => n583, S => n163, Z => n1091);
   U1275 : INV_X1 port map( A => n1092, ZN => n3038);
   U1276 : MUX2_X1 port map( A => n528, B => n582, S => n163, Z => n1092);
   U1277 : INV_X1 port map( A => n1093, ZN => n3037);
   U1278 : MUX2_X1 port map( A => n529, B => n581, S => n163, Z => n1093);
   U1279 : INV_X1 port map( A => n1094, ZN => n3036);
   U1280 : MUX2_X1 port map( A => n530, B => n580, S => n163, Z => n1094);
   U1281 : INV_X1 port map( A => n1095, ZN => n3035);
   U1282 : MUX2_X1 port map( A => n531, B => n579, S => n163, Z => n1095);
   U1283 : INV_X1 port map( A => n1096, ZN => n3034);
   U1284 : MUX2_X1 port map( A => n532, B => n578, S => n163, Z => n1096);
   U1285 : INV_X1 port map( A => n1097, ZN => n3033);
   U1286 : MUX2_X1 port map( A => n533, B => n577, S => n163, Z => n1097);
   U1287 : INV_X1 port map( A => n1098, ZN => n3032);
   U1288 : MUX2_X1 port map( A => n534, B => n576, S => n163, Z => n1098);
   U1289 : INV_X1 port map( A => n1099, ZN => n3031);
   U1290 : MUX2_X1 port map( A => n535, B => n575, S => n163, Z => n1099);
   U1291 : INV_X1 port map( A => n1100, ZN => n3030);
   U1292 : MUX2_X1 port map( A => n536, B => n574, S => n163, Z => n1100);
   U1293 : INV_X1 port map( A => n1101, ZN => n3029);
   U1294 : MUX2_X1 port map( A => n537, B => n573, S => n162, Z => n1101);
   U1295 : INV_X1 port map( A => n1102, ZN => n3028);
   U1296 : MUX2_X1 port map( A => n538, B => n572, S => n162, Z => n1102);
   U1297 : INV_X1 port map( A => n1103, ZN => n3027);
   U1298 : MUX2_X1 port map( A => n539, B => n571, S => n162, Z => n1103);
   U1299 : INV_X1 port map( A => n1104, ZN => n3026);
   U1300 : MUX2_X1 port map( A => n540, B => n570, S => n162, Z => n1104);
   U1301 : INV_X1 port map( A => n1105, ZN => n3025);
   U1302 : MUX2_X1 port map( A => n541, B => n569, S => n162, Z => n1105);
   U1303 : INV_X1 port map( A => n1106, ZN => n3024);
   U1304 : MUX2_X1 port map( A => n542, B => n568, S => n162, Z => n1106);
   U1305 : INV_X1 port map( A => n1107, ZN => n3023);
   U1306 : MUX2_X1 port map( A => n543, B => n567, S => n162, Z => n1107);
   U1307 : INV_X1 port map( A => n1108, ZN => n3022);
   U1308 : MUX2_X1 port map( A => n544, B => n566, S => n162, Z => n1108);
   U1309 : INV_X1 port map( A => n1109, ZN => n3021);
   U1310 : MUX2_X1 port map( A => n545, B => n565, S => n162, Z => n1109);
   U1311 : INV_X1 port map( A => n1110, ZN => n3020);
   U1312 : MUX2_X1 port map( A => n546, B => n564, S => n162, Z => n1110);
   U1313 : INV_X1 port map( A => n1111, ZN => n3019);
   U1314 : MUX2_X1 port map( A => n547, B => n563, S => n162, Z => n1111);
   U1315 : INV_X1 port map( A => n1112, ZN => n3018);
   U1316 : MUX2_X1 port map( A => n548, B => n562, S => n162, Z => n1112);
   U1317 : AND2_X1 port map( A1 => n1079, A2 => n763, ZN => n1081);
   U1318 : MUX2_X1 port map( A => n4190, B => DATAIN(31), S => n167, Z => n3017
                           );
   U1319 : MUX2_X1 port map( A => n4189, B => DATAIN(30), S => n167, Z => n3016
                           );
   U1320 : MUX2_X1 port map( A => n4188, B => DATAIN(29), S => n167, Z => n3015
                           );
   U1321 : MUX2_X1 port map( A => n4187, B => DATAIN(28), S => n167, Z => n3014
                           );
   U1322 : MUX2_X1 port map( A => n4186, B => DATAIN(27), S => n167, Z => n3013
                           );
   U1323 : MUX2_X1 port map( A => n4185, B => DATAIN(26), S => n167, Z => n3012
                           );
   U1324 : MUX2_X1 port map( A => n4184, B => DATAIN(25), S => n167, Z => n3011
                           );
   U1325 : MUX2_X1 port map( A => n4183, B => DATAIN(24), S => n167, Z => n3010
                           );
   U1326 : MUX2_X1 port map( A => n4182, B => DATAIN(23), S => n166, Z => n3009
                           );
   U1327 : MUX2_X1 port map( A => n4181, B => DATAIN(22), S => n166, Z => n3008
                           );
   U1328 : MUX2_X1 port map( A => n4180, B => DATAIN(21), S => n166, Z => n3007
                           );
   U1329 : MUX2_X1 port map( A => n4179, B => DATAIN(20), S => n166, Z => n3006
                           );
   U1330 : MUX2_X1 port map( A => n4178, B => DATAIN(19), S => n166, Z => n3005
                           );
   U1331 : MUX2_X1 port map( A => n4177, B => DATAIN(18), S => n166, Z => n3004
                           );
   U1332 : MUX2_X1 port map( A => n4176, B => DATAIN(17), S => n166, Z => n3003
                           );
   U1333 : MUX2_X1 port map( A => n4175, B => DATAIN(16), S => n166, Z => n3002
                           );
   U1334 : MUX2_X1 port map( A => n4174, B => DATAIN(15), S => n166, Z => n3001
                           );
   U1335 : MUX2_X1 port map( A => n4173, B => DATAIN(14), S => n166, Z => n3000
                           );
   U1336 : MUX2_X1 port map( A => n4172, B => DATAIN(13), S => n166, Z => n2999
                           );
   U1337 : MUX2_X1 port map( A => n4171, B => DATAIN(12), S => n166, Z => n2998
                           );
   U1338 : MUX2_X1 port map( A => n4170, B => DATAIN(11), S => n165, Z => n2997
                           );
   U1339 : MUX2_X1 port map( A => n4169, B => DATAIN(10), S => n165, Z => n2996
                           );
   U1340 : MUX2_X1 port map( A => n4168, B => DATAIN(9), S => n165, Z => n2995)
                           ;
   U1341 : MUX2_X1 port map( A => n4167, B => DATAIN(8), S => n165, Z => n2994)
                           ;
   U1342 : MUX2_X1 port map( A => n4166, B => DATAIN(7), S => n165, Z => n2993)
                           ;
   U1343 : MUX2_X1 port map( A => n4165, B => DATAIN(6), S => n165, Z => n2992)
                           ;
   U1344 : MUX2_X1 port map( A => n4164, B => DATAIN(5), S => n165, Z => n2991)
                           ;
   U1345 : MUX2_X1 port map( A => n4163, B => DATAIN(4), S => n165, Z => n2990)
                           ;
   U1346 : MUX2_X1 port map( A => n4162, B => DATAIN(3), S => n165, Z => n2989)
                           ;
   U1347 : MUX2_X1 port map( A => n4161, B => DATAIN(2), S => n165, Z => n2988)
                           ;
   U1348 : MUX2_X1 port map( A => n4160, B => DATAIN(1), S => n165, Z => n2987)
                           ;
   U1349 : MUX2_X1 port map( A => n4159, B => DATAIN(0), S => n165, Z => n2986)
                           ;
   U1350 : AND2_X1 port map( A1 => n1079, A2 => n766, ZN => n1113);
   U1351 : MUX2_X1 port map( A => n4158, B => DATAIN(31), S => n170, Z => n2985
                           );
   U1352 : MUX2_X1 port map( A => n4157, B => DATAIN(30), S => n170, Z => n2984
                           );
   U1353 : MUX2_X1 port map( A => n4156, B => DATAIN(29), S => n170, Z => n2983
                           );
   U1354 : MUX2_X1 port map( A => n4155, B => DATAIN(28), S => n170, Z => n2982
                           );
   U1355 : MUX2_X1 port map( A => n4154, B => DATAIN(27), S => n170, Z => n2981
                           );
   U1356 : MUX2_X1 port map( A => n4153, B => DATAIN(26), S => n170, Z => n2980
                           );
   U1357 : MUX2_X1 port map( A => n4152, B => DATAIN(25), S => n170, Z => n2979
                           );
   U1358 : MUX2_X1 port map( A => n4151, B => DATAIN(24), S => n170, Z => n2978
                           );
   U1359 : MUX2_X1 port map( A => n4150, B => DATAIN(23), S => n169, Z => n2977
                           );
   U1360 : MUX2_X1 port map( A => n4149, B => DATAIN(22), S => n169, Z => n2976
                           );
   U1361 : MUX2_X1 port map( A => n4148, B => DATAIN(21), S => n169, Z => n2975
                           );
   U1362 : MUX2_X1 port map( A => n4147, B => DATAIN(20), S => n169, Z => n2974
                           );
   U1363 : MUX2_X1 port map( A => n4146, B => DATAIN(19), S => n169, Z => n2973
                           );
   U1364 : MUX2_X1 port map( A => n4145, B => DATAIN(18), S => n169, Z => n2972
                           );
   U1365 : MUX2_X1 port map( A => n4144, B => DATAIN(17), S => n169, Z => n2971
                           );
   U1366 : MUX2_X1 port map( A => n4143, B => DATAIN(16), S => n169, Z => n2970
                           );
   U1367 : MUX2_X1 port map( A => n4142, B => DATAIN(15), S => n169, Z => n2969
                           );
   U1368 : MUX2_X1 port map( A => n4141, B => DATAIN(14), S => n169, Z => n2968
                           );
   U1369 : MUX2_X1 port map( A => n4140, B => DATAIN(13), S => n169, Z => n2967
                           );
   U1370 : MUX2_X1 port map( A => n4139, B => DATAIN(12), S => n169, Z => n2966
                           );
   U1371 : MUX2_X1 port map( A => n4138, B => DATAIN(11), S => n168, Z => n2965
                           );
   U1372 : MUX2_X1 port map( A => n4137, B => DATAIN(10), S => n168, Z => n2964
                           );
   U1373 : MUX2_X1 port map( A => n4136, B => DATAIN(9), S => n168, Z => n2963)
                           ;
   U1374 : MUX2_X1 port map( A => n4135, B => DATAIN(8), S => n168, Z => n2962)
                           ;
   U1375 : MUX2_X1 port map( A => n4134, B => DATAIN(7), S => n168, Z => n2961)
                           ;
   U1376 : MUX2_X1 port map( A => n4133, B => DATAIN(6), S => n168, Z => n2960)
                           ;
   U1377 : MUX2_X1 port map( A => n4132, B => DATAIN(5), S => n168, Z => n2959)
                           ;
   U1378 : MUX2_X1 port map( A => n4131, B => DATAIN(4), S => n168, Z => n2958)
                           ;
   U1379 : MUX2_X1 port map( A => n4130, B => DATAIN(3), S => n168, Z => n2957)
                           ;
   U1380 : MUX2_X1 port map( A => n4129, B => DATAIN(2), S => n168, Z => n2956)
                           ;
   U1381 : MUX2_X1 port map( A => n4128, B => DATAIN(1), S => n168, Z => n2955)
                           ;
   U1382 : MUX2_X1 port map( A => n4127, B => DATAIN(0), S => n168, Z => n2954)
                           ;
   U1383 : AND2_X1 port map( A1 => n1079, A2 => n768, ZN => n1114);
   U1384 : INV_X1 port map( A => n1115, ZN => n2953);
   U1385 : MUX2_X1 port map( A => n613, B => n593, S => n173, Z => n1115);
   U1386 : INV_X1 port map( A => n1117, ZN => n2952);
   U1387 : MUX2_X1 port map( A => n614, B => n592, S => n173, Z => n1117);
   U1388 : INV_X1 port map( A => n1118, ZN => n2951);
   U1389 : MUX2_X1 port map( A => n615, B => n591, S => n173, Z => n1118);
   U1390 : INV_X1 port map( A => n1119, ZN => n2950);
   U1391 : MUX2_X1 port map( A => n616, B => n590, S => n173, Z => n1119);
   U1392 : INV_X1 port map( A => n1120, ZN => n2949);
   U1393 : MUX2_X1 port map( A => n617, B => n589, S => n173, Z => n1120);
   U1394 : INV_X1 port map( A => n1121, ZN => n2948);
   U1395 : MUX2_X1 port map( A => n618, B => n588, S => n173, Z => n1121);
   U1396 : INV_X1 port map( A => n1122, ZN => n2947);
   U1397 : MUX2_X1 port map( A => n619, B => n587, S => n173, Z => n1122);
   U1398 : INV_X1 port map( A => n1123, ZN => n2946);
   U1399 : MUX2_X1 port map( A => n620, B => n586, S => n173, Z => n1123);
   U1400 : INV_X1 port map( A => n1124, ZN => n2945);
   U1401 : MUX2_X1 port map( A => n621, B => n585, S => n172, Z => n1124);
   U1402 : INV_X1 port map( A => n1125, ZN => n2944);
   U1403 : MUX2_X1 port map( A => n622, B => n584, S => n172, Z => n1125);
   U1404 : INV_X1 port map( A => n1126, ZN => n2943);
   U1405 : MUX2_X1 port map( A => n623, B => n583, S => n172, Z => n1126);
   U1406 : INV_X1 port map( A => n1127, ZN => n2942);
   U1407 : MUX2_X1 port map( A => n624, B => n582, S => n172, Z => n1127);
   U1408 : INV_X1 port map( A => n1128, ZN => n2941);
   U1409 : MUX2_X1 port map( A => n625, B => n581, S => n172, Z => n1128);
   U1410 : INV_X1 port map( A => n1129, ZN => n2940);
   U1411 : MUX2_X1 port map( A => n626, B => n580, S => n172, Z => n1129);
   U1412 : INV_X1 port map( A => n1130, ZN => n2939);
   U1413 : MUX2_X1 port map( A => n627, B => n579, S => n172, Z => n1130);
   U1414 : INV_X1 port map( A => n1131, ZN => n2938);
   U1415 : MUX2_X1 port map( A => n628, B => n578, S => n172, Z => n1131);
   U1416 : INV_X1 port map( A => n1132, ZN => n2937);
   U1417 : MUX2_X1 port map( A => n629, B => n577, S => n172, Z => n1132);
   U1418 : INV_X1 port map( A => n1133, ZN => n2936);
   U1419 : MUX2_X1 port map( A => n630, B => n576, S => n172, Z => n1133);
   U1420 : INV_X1 port map( A => n1134, ZN => n2935);
   U1421 : MUX2_X1 port map( A => n631, B => n575, S => n172, Z => n1134);
   U1422 : INV_X1 port map( A => n1135, ZN => n2934);
   U1423 : MUX2_X1 port map( A => n632, B => n574, S => n172, Z => n1135);
   U1424 : INV_X1 port map( A => n1136, ZN => n2933);
   U1425 : MUX2_X1 port map( A => n633, B => n573, S => n171, Z => n1136);
   U1426 : INV_X1 port map( A => n1137, ZN => n2932);
   U1427 : MUX2_X1 port map( A => n634, B => n572, S => n171, Z => n1137);
   U1428 : INV_X1 port map( A => n1138, ZN => n2931);
   U1429 : MUX2_X1 port map( A => n635, B => n571, S => n171, Z => n1138);
   U1430 : INV_X1 port map( A => n1139, ZN => n2930);
   U1431 : MUX2_X1 port map( A => n636, B => n570, S => n171, Z => n1139);
   U1432 : INV_X1 port map( A => n1140, ZN => n2929);
   U1433 : MUX2_X1 port map( A => n637, B => n569, S => n171, Z => n1140);
   U1434 : INV_X1 port map( A => n1141, ZN => n2928);
   U1435 : MUX2_X1 port map( A => n638, B => n568, S => n171, Z => n1141);
   U1436 : INV_X1 port map( A => n1142, ZN => n2927);
   U1437 : MUX2_X1 port map( A => n639, B => n567, S => n171, Z => n1142);
   U1438 : INV_X1 port map( A => n1143, ZN => n2926);
   U1439 : MUX2_X1 port map( A => n640, B => n566, S => n171, Z => n1143);
   U1440 : INV_X1 port map( A => n1144, ZN => n2925);
   U1441 : MUX2_X1 port map( A => n641, B => n565, S => n171, Z => n1144);
   U1442 : INV_X1 port map( A => n1145, ZN => n2924);
   U1443 : MUX2_X1 port map( A => n642, B => n564, S => n171, Z => n1145);
   U1444 : INV_X1 port map( A => n1146, ZN => n2923);
   U1445 : MUX2_X1 port map( A => n643, B => n563, S => n171, Z => n1146);
   U1446 : INV_X1 port map( A => n1147, ZN => n2922);
   U1447 : MUX2_X1 port map( A => n644, B => n562, S => n171, Z => n1147);
   U1448 : AND2_X1 port map( A1 => n1079, A2 => n802, ZN => n1116);
   U1449 : MUX2_X1 port map( A => n1148, B => DATAIN(31), S => n176, Z => n2921
                           );
   U1450 : MUX2_X1 port map( A => n1150, B => DATAIN(30), S => n176, Z => n2920
                           );
   U1451 : MUX2_X1 port map( A => n1151, B => DATAIN(29), S => n176, Z => n2919
                           );
   U1452 : MUX2_X1 port map( A => n1152, B => DATAIN(28), S => n176, Z => n2918
                           );
   U1453 : MUX2_X1 port map( A => n1153, B => DATAIN(27), S => n176, Z => n2917
                           );
   U1454 : MUX2_X1 port map( A => n1154, B => DATAIN(26), S => n176, Z => n2916
                           );
   U1455 : MUX2_X1 port map( A => n1155, B => DATAIN(25), S => n176, Z => n2915
                           );
   U1456 : MUX2_X1 port map( A => n1156, B => DATAIN(24), S => n176, Z => n2914
                           );
   U1457 : MUX2_X1 port map( A => n1157, B => DATAIN(23), S => n175, Z => n2913
                           );
   U1458 : MUX2_X1 port map( A => n1158, B => DATAIN(22), S => n175, Z => n2912
                           );
   U1459 : MUX2_X1 port map( A => n1159, B => DATAIN(21), S => n175, Z => n2911
                           );
   U1460 : MUX2_X1 port map( A => n1160, B => DATAIN(20), S => n175, Z => n2910
                           );
   U1461 : MUX2_X1 port map( A => n1161, B => DATAIN(19), S => n175, Z => n2909
                           );
   U1462 : MUX2_X1 port map( A => n1162, B => DATAIN(18), S => n175, Z => n2908
                           );
   U1463 : MUX2_X1 port map( A => n1163, B => DATAIN(17), S => n175, Z => n2907
                           );
   U1464 : MUX2_X1 port map( A => n1164, B => DATAIN(16), S => n175, Z => n2906
                           );
   U1465 : MUX2_X1 port map( A => n1165, B => DATAIN(15), S => n175, Z => n2905
                           );
   U1466 : MUX2_X1 port map( A => n1166, B => DATAIN(14), S => n175, Z => n2904
                           );
   U1467 : MUX2_X1 port map( A => n1167, B => DATAIN(13), S => n175, Z => n2903
                           );
   U1468 : MUX2_X1 port map( A => n1168, B => DATAIN(12), S => n175, Z => n2902
                           );
   U1469 : MUX2_X1 port map( A => n1169, B => DATAIN(11), S => n174, Z => n2901
                           );
   U1470 : MUX2_X1 port map( A => n1170, B => DATAIN(10), S => n174, Z => n2900
                           );
   U1471 : MUX2_X1 port map( A => n1171, B => DATAIN(9), S => n174, Z => n2899)
                           ;
   U1472 : MUX2_X1 port map( A => n1172, B => DATAIN(8), S => n174, Z => n2898)
                           ;
   U1473 : MUX2_X1 port map( A => n1173, B => DATAIN(7), S => n174, Z => n2897)
                           ;
   U1474 : MUX2_X1 port map( A => n1174, B => DATAIN(6), S => n174, Z => n2896)
                           ;
   U1475 : MUX2_X1 port map( A => n1175, B => DATAIN(5), S => n174, Z => n2895)
                           ;
   U1476 : MUX2_X1 port map( A => n1176, B => DATAIN(4), S => n174, Z => n2894)
                           ;
   U1477 : MUX2_X1 port map( A => n1177, B => DATAIN(3), S => n174, Z => n2893)
                           ;
   U1478 : MUX2_X1 port map( A => n1178, B => DATAIN(2), S => n174, Z => n2892)
                           ;
   U1479 : MUX2_X1 port map( A => n1179, B => DATAIN(1), S => n174, Z => n2891)
                           ;
   U1480 : MUX2_X1 port map( A => n1180, B => DATAIN(0), S => n174, Z => n2890)
                           ;
   U1481 : AND2_X1 port map( A1 => n1079, A2 => n836, ZN => n1149);
   U1482 : MUX2_X1 port map( A => n4126, B => DATAIN(31), S => n179, Z => n2889
                           );
   U1483 : MUX2_X1 port map( A => n4125, B => DATAIN(30), S => n179, Z => n2888
                           );
   U1484 : MUX2_X1 port map( A => n4124, B => DATAIN(29), S => n179, Z => n2887
                           );
   U1485 : MUX2_X1 port map( A => n4123, B => DATAIN(28), S => n179, Z => n2886
                           );
   U1486 : MUX2_X1 port map( A => n4122, B => DATAIN(27), S => n179, Z => n2885
                           );
   U1487 : MUX2_X1 port map( A => n4121, B => DATAIN(26), S => n179, Z => n2884
                           );
   U1488 : MUX2_X1 port map( A => n4120, B => DATAIN(25), S => n179, Z => n2883
                           );
   U1489 : MUX2_X1 port map( A => n4119, B => DATAIN(24), S => n179, Z => n2882
                           );
   U1490 : MUX2_X1 port map( A => n4118, B => DATAIN(23), S => n178, Z => n2881
                           );
   U1491 : MUX2_X1 port map( A => n4117, B => DATAIN(22), S => n178, Z => n2880
                           );
   U1492 : MUX2_X1 port map( A => n4116, B => DATAIN(21), S => n178, Z => n2879
                           );
   U1493 : MUX2_X1 port map( A => n4115, B => DATAIN(20), S => n178, Z => n2878
                           );
   U1494 : MUX2_X1 port map( A => n4114, B => DATAIN(19), S => n178, Z => n2877
                           );
   U1495 : MUX2_X1 port map( A => n4113, B => DATAIN(18), S => n178, Z => n2876
                           );
   U1496 : MUX2_X1 port map( A => n4112, B => DATAIN(17), S => n178, Z => n2875
                           );
   U1497 : MUX2_X1 port map( A => n4111, B => DATAIN(16), S => n178, Z => n2874
                           );
   U1498 : MUX2_X1 port map( A => n4110, B => DATAIN(15), S => n178, Z => n2873
                           );
   U1499 : MUX2_X1 port map( A => n4109, B => DATAIN(14), S => n178, Z => n2872
                           );
   U1500 : MUX2_X1 port map( A => n4108, B => DATAIN(13), S => n178, Z => n2871
                           );
   U1501 : MUX2_X1 port map( A => n4107, B => DATAIN(12), S => n178, Z => n2870
                           );
   U1502 : MUX2_X1 port map( A => n4106, B => DATAIN(11), S => n177, Z => n2869
                           );
   U1503 : MUX2_X1 port map( A => n4105, B => DATAIN(10), S => n177, Z => n2868
                           );
   U1504 : MUX2_X1 port map( A => n4104, B => DATAIN(9), S => n177, Z => n2867)
                           ;
   U1505 : MUX2_X1 port map( A => n4103, B => DATAIN(8), S => n177, Z => n2866)
                           ;
   U1506 : MUX2_X1 port map( A => n4102, B => DATAIN(7), S => n177, Z => n2865)
                           ;
   U1507 : MUX2_X1 port map( A => n4101, B => DATAIN(6), S => n177, Z => n2864)
                           ;
   U1508 : MUX2_X1 port map( A => n4100, B => DATAIN(5), S => n177, Z => n2863)
                           ;
   U1509 : MUX2_X1 port map( A => n4099, B => DATAIN(4), S => n177, Z => n2862)
                           ;
   U1510 : MUX2_X1 port map( A => n4098, B => DATAIN(3), S => n177, Z => n2861)
                           ;
   U1511 : MUX2_X1 port map( A => n4097, B => DATAIN(2), S => n177, Z => n2860)
                           ;
   U1512 : MUX2_X1 port map( A => n4096, B => DATAIN(1), S => n177, Z => n2859)
                           ;
   U1513 : MUX2_X1 port map( A => n4095, B => DATAIN(0), S => n177, Z => n2858)
                           ;
   U1514 : AND2_X1 port map( A1 => n1079, A2 => n870, ZN => n1181);
   U1515 : MUX2_X1 port map( A => n4094, B => DATAIN(31), S => n182, Z => n2857
                           );
   U1516 : MUX2_X1 port map( A => n4093, B => DATAIN(30), S => n182, Z => n2856
                           );
   U1517 : MUX2_X1 port map( A => n4092, B => DATAIN(29), S => n182, Z => n2855
                           );
   U1518 : MUX2_X1 port map( A => n4091, B => DATAIN(28), S => n182, Z => n2854
                           );
   U1519 : MUX2_X1 port map( A => n4090, B => DATAIN(27), S => n182, Z => n2853
                           );
   U1520 : MUX2_X1 port map( A => n4089, B => DATAIN(26), S => n182, Z => n2852
                           );
   U1521 : MUX2_X1 port map( A => n4088, B => DATAIN(25), S => n182, Z => n2851
                           );
   U1522 : MUX2_X1 port map( A => n4087, B => DATAIN(24), S => n182, Z => n2850
                           );
   U1523 : MUX2_X1 port map( A => n4086, B => DATAIN(23), S => n181, Z => n2849
                           );
   U1524 : MUX2_X1 port map( A => n4085, B => DATAIN(22), S => n181, Z => n2848
                           );
   U1525 : MUX2_X1 port map( A => n4084, B => DATAIN(21), S => n181, Z => n2847
                           );
   U1526 : MUX2_X1 port map( A => n4083, B => DATAIN(20), S => n181, Z => n2846
                           );
   U1527 : MUX2_X1 port map( A => n4082, B => DATAIN(19), S => n181, Z => n2845
                           );
   U1528 : MUX2_X1 port map( A => n4081, B => DATAIN(18), S => n181, Z => n2844
                           );
   U1529 : MUX2_X1 port map( A => n4080, B => DATAIN(17), S => n181, Z => n2843
                           );
   U1530 : MUX2_X1 port map( A => n4079, B => DATAIN(16), S => n181, Z => n2842
                           );
   U1531 : MUX2_X1 port map( A => n4078, B => DATAIN(15), S => n181, Z => n2841
                           );
   U1532 : MUX2_X1 port map( A => n4077, B => DATAIN(14), S => n181, Z => n2840
                           );
   U1533 : MUX2_X1 port map( A => n4076, B => DATAIN(13), S => n181, Z => n2839
                           );
   U1534 : MUX2_X1 port map( A => n4075, B => DATAIN(12), S => n181, Z => n2838
                           );
   U1535 : MUX2_X1 port map( A => n4074, B => DATAIN(11), S => n180, Z => n2837
                           );
   U1536 : MUX2_X1 port map( A => n4073, B => DATAIN(10), S => n180, Z => n2836
                           );
   U1537 : MUX2_X1 port map( A => n4072, B => DATAIN(9), S => n180, Z => n2835)
                           ;
   U1538 : MUX2_X1 port map( A => n4071, B => DATAIN(8), S => n180, Z => n2834)
                           ;
   U1539 : MUX2_X1 port map( A => n4070, B => DATAIN(7), S => n180, Z => n2833)
                           ;
   U1540 : MUX2_X1 port map( A => n4069, B => DATAIN(6), S => n180, Z => n2832)
                           ;
   U1541 : MUX2_X1 port map( A => n4068, B => DATAIN(5), S => n180, Z => n2831)
                           ;
   U1542 : MUX2_X1 port map( A => n4067, B => DATAIN(4), S => n180, Z => n2830)
                           ;
   U1543 : MUX2_X1 port map( A => n4066, B => DATAIN(3), S => n180, Z => n2829)
                           ;
   U1544 : MUX2_X1 port map( A => n4065, B => DATAIN(2), S => n180, Z => n2828)
                           ;
   U1545 : MUX2_X1 port map( A => n4064, B => DATAIN(1), S => n180, Z => n2827)
                           ;
   U1546 : MUX2_X1 port map( A => n4063, B => DATAIN(0), S => n180, Z => n2826)
                           ;
   U1547 : AND2_X1 port map( A1 => n1079, A2 => n872, ZN => n1182);
   U1548 : AND3_X1 port map( A1 => n875, A2 => n873, A3 => ADD_WR(4), ZN => 
                           n1079);
   U1549 : MUX2_X1 port map( A => n4062, B => DATAIN(31), S => n185, Z => n2825
                           );
   U1550 : MUX2_X1 port map( A => n4061, B => DATAIN(30), S => n185, Z => n2824
                           );
   U1551 : MUX2_X1 port map( A => n4060, B => DATAIN(29), S => n185, Z => n2823
                           );
   U1552 : MUX2_X1 port map( A => n4059, B => DATAIN(28), S => n185, Z => n2822
                           );
   U1553 : MUX2_X1 port map( A => n4058, B => DATAIN(27), S => n185, Z => n2821
                           );
   U1554 : MUX2_X1 port map( A => n4057, B => DATAIN(26), S => n185, Z => n2820
                           );
   U1555 : MUX2_X1 port map( A => n4056, B => DATAIN(25), S => n185, Z => n2819
                           );
   U1556 : MUX2_X1 port map( A => n4055, B => DATAIN(24), S => n185, Z => n2818
                           );
   U1557 : MUX2_X1 port map( A => n4054, B => DATAIN(23), S => n184, Z => n2817
                           );
   U1558 : MUX2_X1 port map( A => n4053, B => DATAIN(22), S => n184, Z => n2816
                           );
   U1559 : MUX2_X1 port map( A => n4052, B => DATAIN(21), S => n184, Z => n2815
                           );
   U1560 : MUX2_X1 port map( A => n4051, B => DATAIN(20), S => n184, Z => n2814
                           );
   U1561 : MUX2_X1 port map( A => n4050, B => DATAIN(19), S => n184, Z => n2813
                           );
   U1562 : MUX2_X1 port map( A => n4049, B => DATAIN(18), S => n184, Z => n2812
                           );
   U1563 : MUX2_X1 port map( A => n4048, B => DATAIN(17), S => n184, Z => n2811
                           );
   U1564 : MUX2_X1 port map( A => n4047, B => DATAIN(16), S => n184, Z => n2810
                           );
   U1565 : MUX2_X1 port map( A => n4046, B => DATAIN(15), S => n184, Z => n2809
                           );
   U1566 : MUX2_X1 port map( A => n4045, B => DATAIN(14), S => n184, Z => n2808
                           );
   U1567 : MUX2_X1 port map( A => n4044, B => DATAIN(13), S => n184, Z => n2807
                           );
   U1568 : MUX2_X1 port map( A => n4043, B => DATAIN(12), S => n184, Z => n2806
                           );
   U1569 : MUX2_X1 port map( A => n4042, B => DATAIN(11), S => n183, Z => n2805
                           );
   U1570 : MUX2_X1 port map( A => n4041, B => DATAIN(10), S => n183, Z => n2804
                           );
   U1571 : MUX2_X1 port map( A => n4040, B => DATAIN(9), S => n183, Z => n2803)
                           ;
   U1572 : MUX2_X1 port map( A => n4039, B => DATAIN(8), S => n183, Z => n2802)
                           ;
   U1573 : MUX2_X1 port map( A => n4038, B => DATAIN(7), S => n183, Z => n2801)
                           ;
   U1574 : MUX2_X1 port map( A => n4037, B => DATAIN(6), S => n183, Z => n2800)
                           ;
   U1575 : MUX2_X1 port map( A => n4036, B => DATAIN(5), S => n183, Z => n2799)
                           ;
   U1576 : MUX2_X1 port map( A => n4035, B => DATAIN(4), S => n183, Z => n2798)
                           ;
   U1577 : MUX2_X1 port map( A => n4034, B => DATAIN(3), S => n183, Z => n2797)
                           ;
   U1578 : MUX2_X1 port map( A => n4033, B => DATAIN(2), S => n183, Z => n2796)
                           ;
   U1579 : MUX2_X1 port map( A => n4032, B => DATAIN(1), S => n183, Z => n2795)
                           ;
   U1580 : MUX2_X1 port map( A => n4031, B => DATAIN(0), S => n183, Z => n2794)
                           ;
   U1581 : AND2_X1 port map( A1 => n1184, A2 => n910, ZN => n1183);
   U1582 : MUX2_X1 port map( A => n4030, B => DATAIN(31), S => n188, Z => n2793
                           );
   U1583 : MUX2_X1 port map( A => n4029, B => DATAIN(30), S => n188, Z => n2792
                           );
   U1584 : MUX2_X1 port map( A => n4028, B => DATAIN(29), S => n188, Z => n2791
                           );
   U1585 : MUX2_X1 port map( A => n4027, B => DATAIN(28), S => n188, Z => n2790
                           );
   U1586 : MUX2_X1 port map( A => n4026, B => DATAIN(27), S => n188, Z => n2789
                           );
   U1587 : MUX2_X1 port map( A => n4025, B => DATAIN(26), S => n188, Z => n2788
                           );
   U1588 : MUX2_X1 port map( A => n4024, B => DATAIN(25), S => n188, Z => n2787
                           );
   U1589 : MUX2_X1 port map( A => n4023, B => DATAIN(24), S => n188, Z => n2786
                           );
   U1590 : MUX2_X1 port map( A => n4022, B => DATAIN(23), S => n187, Z => n2785
                           );
   U1591 : MUX2_X1 port map( A => n4021, B => DATAIN(22), S => n187, Z => n2784
                           );
   U1592 : MUX2_X1 port map( A => n4020, B => DATAIN(21), S => n187, Z => n2783
                           );
   U1593 : MUX2_X1 port map( A => n4019, B => DATAIN(20), S => n187, Z => n2782
                           );
   U1594 : MUX2_X1 port map( A => n4018, B => DATAIN(19), S => n187, Z => n2781
                           );
   U1595 : MUX2_X1 port map( A => n4017, B => DATAIN(18), S => n187, Z => n2780
                           );
   U1596 : MUX2_X1 port map( A => n4016, B => DATAIN(17), S => n187, Z => n2779
                           );
   U1597 : MUX2_X1 port map( A => n4015, B => DATAIN(16), S => n187, Z => n2778
                           );
   U1598 : MUX2_X1 port map( A => n4014, B => DATAIN(15), S => n187, Z => n2777
                           );
   U1599 : MUX2_X1 port map( A => n4013, B => DATAIN(14), S => n187, Z => n2776
                           );
   U1600 : MUX2_X1 port map( A => n4012, B => DATAIN(13), S => n187, Z => n2775
                           );
   U1601 : MUX2_X1 port map( A => n4011, B => DATAIN(12), S => n187, Z => n2774
                           );
   U1602 : MUX2_X1 port map( A => n4010, B => DATAIN(11), S => n186, Z => n2773
                           );
   U1603 : MUX2_X1 port map( A => n4009, B => DATAIN(10), S => n186, Z => n2772
                           );
   U1604 : MUX2_X1 port map( A => n4008, B => DATAIN(9), S => n186, Z => n2771)
                           ;
   U1605 : MUX2_X1 port map( A => n4007, B => DATAIN(8), S => n186, Z => n2770)
                           ;
   U1606 : MUX2_X1 port map( A => n4006, B => DATAIN(7), S => n186, Z => n2769)
                           ;
   U1607 : MUX2_X1 port map( A => n4005, B => DATAIN(6), S => n186, Z => n2768)
                           ;
   U1608 : MUX2_X1 port map( A => n4004, B => DATAIN(5), S => n186, Z => n2767)
                           ;
   U1609 : MUX2_X1 port map( A => n4003, B => DATAIN(4), S => n186, Z => n2766)
                           ;
   U1610 : MUX2_X1 port map( A => n4002, B => DATAIN(3), S => n186, Z => n2765)
                           ;
   U1611 : MUX2_X1 port map( A => n4001, B => DATAIN(2), S => n186, Z => n2764)
                           ;
   U1612 : MUX2_X1 port map( A => n4000, B => DATAIN(1), S => n186, Z => n2763)
                           ;
   U1613 : MUX2_X1 port map( A => n3999, B => DATAIN(0), S => n186, Z => n2762)
                           ;
   U1614 : AND2_X1 port map( A1 => n1184, A2 => n763, ZN => n1185);
   U1615 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => n1186, ZN 
                           => n763);
   U1616 : MUX2_X1 port map( A => n1187, B => DATAIN(31), S => n191, Z => n2761
                           );
   U1617 : MUX2_X1 port map( A => n1189, B => DATAIN(30), S => n191, Z => n2760
                           );
   U1618 : MUX2_X1 port map( A => n1190, B => DATAIN(29), S => n191, Z => n2759
                           );
   U1619 : MUX2_X1 port map( A => n1191, B => DATAIN(28), S => n191, Z => n2758
                           );
   U1620 : MUX2_X1 port map( A => n1192, B => DATAIN(27), S => n191, Z => n2757
                           );
   U1621 : MUX2_X1 port map( A => n1193, B => DATAIN(26), S => n191, Z => n2756
                           );
   U1622 : MUX2_X1 port map( A => n1194, B => DATAIN(25), S => n191, Z => n2755
                           );
   U1623 : MUX2_X1 port map( A => n1195, B => DATAIN(24), S => n191, Z => n2754
                           );
   U1624 : MUX2_X1 port map( A => n1196, B => DATAIN(23), S => n190, Z => n2753
                           );
   U1625 : MUX2_X1 port map( A => n1197, B => DATAIN(22), S => n190, Z => n2752
                           );
   U1626 : MUX2_X1 port map( A => n1198, B => DATAIN(21), S => n190, Z => n2751
                           );
   U1627 : MUX2_X1 port map( A => n1199, B => DATAIN(20), S => n190, Z => n2750
                           );
   U1628 : MUX2_X1 port map( A => n1200, B => DATAIN(19), S => n190, Z => n2749
                           );
   U1629 : MUX2_X1 port map( A => n1201, B => DATAIN(18), S => n190, Z => n2748
                           );
   U1630 : MUX2_X1 port map( A => n1202, B => DATAIN(17), S => n190, Z => n2747
                           );
   U1631 : MUX2_X1 port map( A => n1203, B => DATAIN(16), S => n190, Z => n2746
                           );
   U1632 : MUX2_X1 port map( A => n1204, B => DATAIN(15), S => n190, Z => n2745
                           );
   U1633 : MUX2_X1 port map( A => n1205, B => DATAIN(14), S => n190, Z => n2744
                           );
   U1634 : MUX2_X1 port map( A => n1206, B => DATAIN(13), S => n190, Z => n2743
                           );
   U1635 : MUX2_X1 port map( A => n1207, B => DATAIN(12), S => n190, Z => n2742
                           );
   U1636 : MUX2_X1 port map( A => n1208, B => DATAIN(11), S => n189, Z => n2741
                           );
   U1637 : MUX2_X1 port map( A => n1209, B => DATAIN(10), S => n189, Z => n2740
                           );
   U1638 : MUX2_X1 port map( A => n1210, B => DATAIN(9), S => n189, Z => n2739)
                           ;
   U1639 : MUX2_X1 port map( A => n1211, B => DATAIN(8), S => n189, Z => n2738)
                           ;
   U1640 : MUX2_X1 port map( A => n1212, B => DATAIN(7), S => n189, Z => n2737)
                           ;
   U1641 : MUX2_X1 port map( A => n1213, B => DATAIN(6), S => n189, Z => n2736)
                           ;
   U1642 : MUX2_X1 port map( A => n1214, B => DATAIN(5), S => n189, Z => n2735)
                           ;
   U1643 : MUX2_X1 port map( A => n1215, B => DATAIN(4), S => n189, Z => n2734)
                           ;
   U1644 : MUX2_X1 port map( A => n1216, B => DATAIN(3), S => n189, Z => n2733)
                           ;
   U1645 : MUX2_X1 port map( A => n1217, B => DATAIN(2), S => n189, Z => n2732)
                           ;
   U1646 : MUX2_X1 port map( A => n1218, B => DATAIN(1), S => n189, Z => n2731)
                           ;
   U1647 : MUX2_X1 port map( A => n1219, B => DATAIN(0), S => n189, Z => n2730)
                           ;
   U1648 : AND2_X1 port map( A1 => n1184, A2 => n766, ZN => n1188);
   U1649 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(2), A3 => n1220, ZN 
                           => n766);
   U1650 : INV_X1 port map( A => n1221, ZN => n2729);
   U1651 : MUX2_X1 port map( A => n837, B => n593, S => n194, Z => n1221);
   U1652 : INV_X1 port map( A => n1223, ZN => n2728);
   U1653 : MUX2_X1 port map( A => n838, B => n592, S => n194, Z => n1223);
   U1654 : INV_X1 port map( A => n1224, ZN => n2727);
   U1655 : MUX2_X1 port map( A => n839, B => n591, S => n194, Z => n1224);
   U1656 : INV_X1 port map( A => n1225, ZN => n2726);
   U1657 : MUX2_X1 port map( A => n840, B => n590, S => n194, Z => n1225);
   U1658 : INV_X1 port map( A => n1226, ZN => n2725);
   U1659 : MUX2_X1 port map( A => n841, B => n589, S => n194, Z => n1226);
   U1660 : INV_X1 port map( A => n1227, ZN => n2724);
   U1661 : MUX2_X1 port map( A => n842, B => n588, S => n194, Z => n1227);
   U1662 : INV_X1 port map( A => n1228, ZN => n2723);
   U1663 : MUX2_X1 port map( A => n843, B => n587, S => n194, Z => n1228);
   U1664 : INV_X1 port map( A => n1229, ZN => n2722);
   U1665 : MUX2_X1 port map( A => n844, B => n586, S => n194, Z => n1229);
   U1666 : INV_X1 port map( A => n1230, ZN => n2721);
   U1667 : MUX2_X1 port map( A => n845, B => n585, S => n193, Z => n1230);
   U1668 : INV_X1 port map( A => n1231, ZN => n2720);
   U1669 : MUX2_X1 port map( A => n846, B => n584, S => n193, Z => n1231);
   U1670 : INV_X1 port map( A => n1232, ZN => n2719);
   U1671 : MUX2_X1 port map( A => n847, B => n583, S => n193, Z => n1232);
   U1672 : INV_X1 port map( A => n1233, ZN => n2718);
   U1673 : MUX2_X1 port map( A => n848, B => n582, S => n193, Z => n1233);
   U1674 : INV_X1 port map( A => n1234, ZN => n2717);
   U1675 : MUX2_X1 port map( A => n849, B => n581, S => n193, Z => n1234);
   U1676 : INV_X1 port map( A => n1235, ZN => n2716);
   U1677 : MUX2_X1 port map( A => n850, B => n580, S => n193, Z => n1235);
   U1678 : INV_X1 port map( A => n1236, ZN => n2715);
   U1679 : MUX2_X1 port map( A => n851, B => n579, S => n193, Z => n1236);
   U1680 : INV_X1 port map( A => n1237, ZN => n2714);
   U1681 : MUX2_X1 port map( A => n852, B => n578, S => n193, Z => n1237);
   U1682 : INV_X1 port map( A => n1238, ZN => n2713);
   U1683 : MUX2_X1 port map( A => n853, B => n577, S => n193, Z => n1238);
   U1684 : INV_X1 port map( A => n1239, ZN => n2712);
   U1685 : MUX2_X1 port map( A => n854, B => n576, S => n193, Z => n1239);
   U1686 : INV_X1 port map( A => n1240, ZN => n2711);
   U1687 : MUX2_X1 port map( A => n855, B => n575, S => n193, Z => n1240);
   U1688 : INV_X1 port map( A => n1241, ZN => n2710);
   U1689 : MUX2_X1 port map( A => n856, B => n574, S => n193, Z => n1241);
   U1690 : INV_X1 port map( A => n1242, ZN => n2709);
   U1691 : MUX2_X1 port map( A => n857, B => n573, S => n192, Z => n1242);
   U1692 : INV_X1 port map( A => n1243, ZN => n2708);
   U1693 : MUX2_X1 port map( A => n858, B => n572, S => n192, Z => n1243);
   U1694 : INV_X1 port map( A => n1244, ZN => n2707);
   U1695 : MUX2_X1 port map( A => n859, B => n571, S => n192, Z => n1244);
   U1696 : INV_X1 port map( A => n1245, ZN => n2706);
   U1697 : MUX2_X1 port map( A => n860, B => n570, S => n192, Z => n1245);
   U1698 : INV_X1 port map( A => n1246, ZN => n2705);
   U1699 : MUX2_X1 port map( A => n861, B => n569, S => n192, Z => n1246);
   U1700 : INV_X1 port map( A => n1247, ZN => n2704);
   U1701 : MUX2_X1 port map( A => n862, B => n568, S => n192, Z => n1247);
   U1702 : INV_X1 port map( A => n1248, ZN => n2703);
   U1703 : MUX2_X1 port map( A => n863, B => n567, S => n192, Z => n1248);
   U1704 : INV_X1 port map( A => n1249, ZN => n2702);
   U1705 : MUX2_X1 port map( A => n864, B => n566, S => n192, Z => n1249);
   U1706 : INV_X1 port map( A => n1250, ZN => n2701);
   U1707 : MUX2_X1 port map( A => n865, B => n565, S => n192, Z => n1250);
   U1708 : INV_X1 port map( A => n1251, ZN => n2700);
   U1709 : MUX2_X1 port map( A => n866, B => n564, S => n192, Z => n1251);
   U1710 : INV_X1 port map( A => n1252, ZN => n2699);
   U1711 : MUX2_X1 port map( A => n867, B => n563, S => n192, Z => n1252);
   U1712 : INV_X1 port map( A => n1253, ZN => n2698);
   U1713 : MUX2_X1 port map( A => n868, B => n562, S => n192, Z => n1253);
   U1714 : AND2_X1 port map( A1 => n1184, A2 => n768, ZN => n1222);
   U1715 : NOR3_X1 port map( A1 => n1186, A2 => ADD_WR(2), A3 => n1220, ZN => 
                           n768);
   U1716 : MUX2_X1 port map( A => n3998, B => DATAIN(31), S => n197, Z => n2697
                           );
   U1717 : MUX2_X1 port map( A => n3997, B => DATAIN(30), S => n197, Z => n2696
                           );
   U1718 : MUX2_X1 port map( A => n3996, B => DATAIN(29), S => n197, Z => n2695
                           );
   U1719 : MUX2_X1 port map( A => n3995, B => DATAIN(28), S => n197, Z => n2694
                           );
   U1720 : MUX2_X1 port map( A => n3994, B => DATAIN(27), S => n197, Z => n2693
                           );
   U1721 : MUX2_X1 port map( A => n3993, B => DATAIN(26), S => n197, Z => n2692
                           );
   U1722 : MUX2_X1 port map( A => n3992, B => DATAIN(25), S => n197, Z => n2691
                           );
   U1723 : MUX2_X1 port map( A => n3991, B => DATAIN(24), S => n197, Z => n2690
                           );
   U1724 : MUX2_X1 port map( A => n3990, B => DATAIN(23), S => n196, Z => n2689
                           );
   U1725 : MUX2_X1 port map( A => n3989, B => DATAIN(22), S => n196, Z => n2688
                           );
   U1726 : MUX2_X1 port map( A => n3988, B => DATAIN(21), S => n196, Z => n2687
                           );
   U1727 : MUX2_X1 port map( A => n3987, B => DATAIN(20), S => n196, Z => n2686
                           );
   U1728 : MUX2_X1 port map( A => n3986, B => DATAIN(19), S => n196, Z => n2685
                           );
   U1729 : MUX2_X1 port map( A => n3985, B => DATAIN(18), S => n196, Z => n2684
                           );
   U1730 : MUX2_X1 port map( A => n3984, B => DATAIN(17), S => n196, Z => n2683
                           );
   U1731 : MUX2_X1 port map( A => n3983, B => DATAIN(16), S => n196, Z => n2682
                           );
   U1732 : MUX2_X1 port map( A => n3982, B => DATAIN(15), S => n196, Z => n2681
                           );
   U1733 : MUX2_X1 port map( A => n3981, B => DATAIN(14), S => n196, Z => n2680
                           );
   U1734 : MUX2_X1 port map( A => n3980, B => DATAIN(13), S => n196, Z => n2679
                           );
   U1735 : MUX2_X1 port map( A => n3979, B => DATAIN(12), S => n196, Z => n2678
                           );
   U1736 : MUX2_X1 port map( A => n3978, B => DATAIN(11), S => n195, Z => n2677
                           );
   U1737 : MUX2_X1 port map( A => n3977, B => DATAIN(10), S => n195, Z => n2676
                           );
   U1738 : MUX2_X1 port map( A => n3976, B => DATAIN(9), S => n195, Z => n2675)
                           ;
   U1739 : MUX2_X1 port map( A => n3975, B => DATAIN(8), S => n195, Z => n2674)
                           ;
   U1740 : MUX2_X1 port map( A => n3974, B => DATAIN(7), S => n195, Z => n2673)
                           ;
   U1741 : MUX2_X1 port map( A => n3973, B => DATAIN(6), S => n195, Z => n2672)
                           ;
   U1742 : MUX2_X1 port map( A => n3972, B => DATAIN(5), S => n195, Z => n2671)
                           ;
   U1743 : MUX2_X1 port map( A => n3971, B => DATAIN(4), S => n195, Z => n2670)
                           ;
   U1744 : MUX2_X1 port map( A => n3970, B => DATAIN(3), S => n195, Z => n2669)
                           ;
   U1745 : MUX2_X1 port map( A => n3969, B => DATAIN(2), S => n195, Z => n2668)
                           ;
   U1746 : MUX2_X1 port map( A => n3968, B => DATAIN(1), S => n195, Z => n2667)
                           ;
   U1747 : MUX2_X1 port map( A => n3967, B => DATAIN(0), S => n195, Z => n2666)
                           ;
   U1748 : AND2_X1 port map( A1 => n1184, A2 => n802, ZN => n1254);
   U1749 : AND3_X1 port map( A1 => n1186, A2 => n1220, A3 => ADD_WR(2), ZN => 
                           n802);
   U1750 : MUX2_X1 port map( A => n3966, B => DATAIN(31), S => n200, Z => n2665
                           );
   U1751 : MUX2_X1 port map( A => n3965, B => DATAIN(30), S => n200, Z => n2664
                           );
   U1752 : MUX2_X1 port map( A => n3964, B => DATAIN(29), S => n200, Z => n2663
                           );
   U1753 : MUX2_X1 port map( A => n3963, B => DATAIN(28), S => n200, Z => n2662
                           );
   U1754 : MUX2_X1 port map( A => n3962, B => DATAIN(27), S => n200, Z => n2661
                           );
   U1755 : MUX2_X1 port map( A => n3961, B => DATAIN(26), S => n200, Z => n2660
                           );
   U1756 : MUX2_X1 port map( A => n3960, B => DATAIN(25), S => n200, Z => n2659
                           );
   U1757 : MUX2_X1 port map( A => n3959, B => DATAIN(24), S => n200, Z => n2658
                           );
   U1758 : MUX2_X1 port map( A => n3958, B => DATAIN(23), S => n199, Z => n2657
                           );
   U1759 : MUX2_X1 port map( A => n3957, B => DATAIN(22), S => n199, Z => n2656
                           );
   U1760 : MUX2_X1 port map( A => n3956, B => DATAIN(21), S => n199, Z => n2655
                           );
   U1761 : MUX2_X1 port map( A => n3955, B => DATAIN(20), S => n199, Z => n2654
                           );
   U1762 : MUX2_X1 port map( A => n3954, B => DATAIN(19), S => n199, Z => n2653
                           );
   U1763 : MUX2_X1 port map( A => n3953, B => DATAIN(18), S => n199, Z => n2652
                           );
   U1764 : MUX2_X1 port map( A => n3952, B => DATAIN(17), S => n199, Z => n2651
                           );
   U1765 : MUX2_X1 port map( A => n3951, B => DATAIN(16), S => n199, Z => n2650
                           );
   U1766 : MUX2_X1 port map( A => n3950, B => DATAIN(15), S => n199, Z => n2649
                           );
   U1767 : MUX2_X1 port map( A => n3949, B => DATAIN(14), S => n199, Z => n2648
                           );
   U1768 : MUX2_X1 port map( A => n3948, B => DATAIN(13), S => n199, Z => n2647
                           );
   U1769 : MUX2_X1 port map( A => n3947, B => DATAIN(12), S => n199, Z => n2646
                           );
   U1770 : MUX2_X1 port map( A => n3946, B => DATAIN(11), S => n198, Z => n2645
                           );
   U1771 : MUX2_X1 port map( A => n3945, B => DATAIN(10), S => n198, Z => n2644
                           );
   U1772 : MUX2_X1 port map( A => n3944, B => DATAIN(9), S => n198, Z => n2643)
                           ;
   U1773 : MUX2_X1 port map( A => n3943, B => DATAIN(8), S => n198, Z => n2642)
                           ;
   U1774 : MUX2_X1 port map( A => n3942, B => DATAIN(7), S => n198, Z => n2641)
                           ;
   U1775 : MUX2_X1 port map( A => n3941, B => DATAIN(6), S => n198, Z => n2640)
                           ;
   U1776 : MUX2_X1 port map( A => n3940, B => DATAIN(5), S => n198, Z => n2639)
                           ;
   U1777 : MUX2_X1 port map( A => n3939, B => DATAIN(4), S => n198, Z => n2638)
                           ;
   U1778 : MUX2_X1 port map( A => n3938, B => DATAIN(3), S => n198, Z => n2637)
                           ;
   U1779 : MUX2_X1 port map( A => n3937, B => DATAIN(2), S => n198, Z => n2636)
                           ;
   U1780 : MUX2_X1 port map( A => n3936, B => DATAIN(1), S => n198, Z => n2635)
                           ;
   U1781 : MUX2_X1 port map( A => n3935, B => DATAIN(0), S => n198, Z => n2634)
                           ;
   U1782 : AND2_X1 port map( A1 => n1184, A2 => n836, ZN => n1255);
   U1783 : AND3_X1 port map( A1 => ADD_WR(0), A2 => n1220, A3 => ADD_WR(2), ZN 
                           => n836);
   U1784 : INV_X1 port map( A => n1256, ZN => n2633);
   U1785 : MUX2_X1 port map( A => n933, B => n593, S => n203, Z => n1256);
   U1786 : INV_X1 port map( A => n1258, ZN => n2632);
   U1787 : MUX2_X1 port map( A => n934, B => n592, S => n203, Z => n1258);
   U1788 : INV_X1 port map( A => n1259, ZN => n2631);
   U1789 : MUX2_X1 port map( A => n935, B => n591, S => n203, Z => n1259);
   U1790 : INV_X1 port map( A => n1260, ZN => n2630);
   U1791 : MUX2_X1 port map( A => n936, B => n590, S => n203, Z => n1260);
   U1792 : INV_X1 port map( A => n1261, ZN => n2629);
   U1793 : MUX2_X1 port map( A => n937, B => n589, S => n203, Z => n1261);
   U1794 : INV_X1 port map( A => n1262, ZN => n2628);
   U1795 : MUX2_X1 port map( A => n938, B => n588, S => n203, Z => n1262);
   U1796 : INV_X1 port map( A => n1263, ZN => n2627);
   U1797 : MUX2_X1 port map( A => n939, B => n587, S => n203, Z => n1263);
   U1798 : INV_X1 port map( A => n1264, ZN => n2626);
   U1799 : MUX2_X1 port map( A => n940, B => n586, S => n203, Z => n1264);
   U1800 : INV_X1 port map( A => n1265, ZN => n2625);
   U1801 : MUX2_X1 port map( A => n941, B => n585, S => n202, Z => n1265);
   U1802 : INV_X1 port map( A => n1266, ZN => n2624);
   U1803 : MUX2_X1 port map( A => n942, B => n584, S => n202, Z => n1266);
   U1804 : INV_X1 port map( A => n1267, ZN => n2623);
   U1805 : MUX2_X1 port map( A => n943, B => n583, S => n202, Z => n1267);
   U1806 : INV_X1 port map( A => n1268, ZN => n2622);
   U1807 : MUX2_X1 port map( A => n944, B => n582, S => n202, Z => n1268);
   U1808 : INV_X1 port map( A => n1269, ZN => n2621);
   U1809 : MUX2_X1 port map( A => n945, B => n581, S => n202, Z => n1269);
   U1810 : INV_X1 port map( A => n1270, ZN => n2620);
   U1811 : MUX2_X1 port map( A => n946, B => n580, S => n202, Z => n1270);
   U1812 : INV_X1 port map( A => n1271, ZN => n2619);
   U1813 : MUX2_X1 port map( A => n947, B => n579, S => n202, Z => n1271);
   U1814 : INV_X1 port map( A => n1272, ZN => n2618);
   U1815 : MUX2_X1 port map( A => n948, B => n578, S => n202, Z => n1272);
   U1816 : INV_X1 port map( A => n1273, ZN => n2617);
   U1817 : MUX2_X1 port map( A => n949, B => n577, S => n202, Z => n1273);
   U1818 : INV_X1 port map( A => n1274, ZN => n2616);
   U1819 : MUX2_X1 port map( A => n950, B => n576, S => n202, Z => n1274);
   U1820 : INV_X1 port map( A => n1275, ZN => n2615);
   U1821 : MUX2_X1 port map( A => n951, B => n575, S => n202, Z => n1275);
   U1822 : INV_X1 port map( A => n1276, ZN => n2614);
   U1823 : MUX2_X1 port map( A => n952, B => n574, S => n202, Z => n1276);
   U1824 : INV_X1 port map( A => n1277, ZN => n2613);
   U1825 : MUX2_X1 port map( A => n953, B => n573, S => n201, Z => n1277);
   U1826 : INV_X1 port map( A => n1278, ZN => n2612);
   U1827 : MUX2_X1 port map( A => n954, B => n572, S => n201, Z => n1278);
   U1828 : INV_X1 port map( A => n1279, ZN => n2611);
   U1829 : MUX2_X1 port map( A => n955, B => n571, S => n201, Z => n1279);
   U1830 : INV_X1 port map( A => n1280, ZN => n2610);
   U1831 : MUX2_X1 port map( A => n956, B => n570, S => n201, Z => n1280);
   U1832 : INV_X1 port map( A => n1281, ZN => n2609);
   U1833 : MUX2_X1 port map( A => n957, B => n569, S => n201, Z => n1281);
   U1834 : INV_X1 port map( A => n1282, ZN => n2608);
   U1835 : MUX2_X1 port map( A => n958, B => n568, S => n201, Z => n1282);
   U1836 : INV_X1 port map( A => n1283, ZN => n2607);
   U1837 : MUX2_X1 port map( A => n959, B => n567, S => n201, Z => n1283);
   U1838 : INV_X1 port map( A => n1284, ZN => n2606);
   U1839 : MUX2_X1 port map( A => n960, B => n566, S => n201, Z => n1284);
   U1840 : INV_X1 port map( A => n1285, ZN => n2605);
   U1841 : MUX2_X1 port map( A => n961, B => n565, S => n201, Z => n1285);
   U1842 : INV_X1 port map( A => n1286, ZN => n2604);
   U1843 : MUX2_X1 port map( A => n962, B => n564, S => n201, Z => n1286);
   U1844 : INV_X1 port map( A => n1287, ZN => n2603);
   U1845 : MUX2_X1 port map( A => n963, B => n563, S => n201, Z => n1287);
   U1846 : INV_X1 port map( A => n1288, ZN => n2602);
   U1847 : MUX2_X1 port map( A => n964, B => n562, S => n201, Z => n1288);
   U1848 : AND2_X1 port map( A1 => n1184, A2 => n870, ZN => n1257);
   U1849 : AND3_X1 port map( A1 => ADD_WR(1), A2 => n1186, A3 => ADD_WR(2), ZN 
                           => n870);
   U1850 : MUX2_X1 port map( A => n1289, B => DATAIN(31), S => n206, Z => n2601
                           );
   U1851 : MUX2_X1 port map( A => n1291, B => DATAIN(30), S => n206, Z => n2600
                           );
   U1852 : MUX2_X1 port map( A => n1292, B => DATAIN(29), S => n206, Z => n2599
                           );
   U1853 : MUX2_X1 port map( A => n1293, B => DATAIN(28), S => n206, Z => n2598
                           );
   U1854 : MUX2_X1 port map( A => n1294, B => DATAIN(27), S => n206, Z => n2597
                           );
   U1855 : MUX2_X1 port map( A => n1295, B => DATAIN(26), S => n206, Z => n2596
                           );
   U1856 : MUX2_X1 port map( A => n1296, B => DATAIN(25), S => n206, Z => n2595
                           );
   U1857 : MUX2_X1 port map( A => n1297, B => DATAIN(24), S => n206, Z => n2594
                           );
   U1858 : MUX2_X1 port map( A => n1298, B => DATAIN(23), S => n205, Z => n2593
                           );
   U1859 : MUX2_X1 port map( A => n1299, B => DATAIN(22), S => n205, Z => n2592
                           );
   U1860 : MUX2_X1 port map( A => n1300, B => DATAIN(21), S => n205, Z => n2591
                           );
   U1861 : MUX2_X1 port map( A => n1301, B => DATAIN(20), S => n205, Z => n2590
                           );
   U1862 : MUX2_X1 port map( A => n1302, B => DATAIN(19), S => n205, Z => n2589
                           );
   U1863 : MUX2_X1 port map( A => n1303, B => DATAIN(18), S => n205, Z => n2588
                           );
   U1864 : MUX2_X1 port map( A => n1304, B => DATAIN(17), S => n205, Z => n2587
                           );
   U1865 : MUX2_X1 port map( A => n1305, B => DATAIN(16), S => n205, Z => n2586
                           );
   U1866 : MUX2_X1 port map( A => n1306, B => DATAIN(15), S => n205, Z => n2585
                           );
   U1867 : MUX2_X1 port map( A => n1307, B => DATAIN(14), S => n205, Z => n2584
                           );
   U1868 : MUX2_X1 port map( A => n1308, B => DATAIN(13), S => n205, Z => n2583
                           );
   U1869 : MUX2_X1 port map( A => n1309, B => DATAIN(12), S => n205, Z => n2582
                           );
   U1870 : MUX2_X1 port map( A => n1310, B => DATAIN(11), S => n204, Z => n2581
                           );
   U1871 : MUX2_X1 port map( A => n1311, B => DATAIN(10), S => n204, Z => n2580
                           );
   U1872 : MUX2_X1 port map( A => n1312, B => DATAIN(9), S => n204, Z => n2579)
                           ;
   U1873 : MUX2_X1 port map( A => n1313, B => DATAIN(8), S => n204, Z => n2578)
                           ;
   U1874 : MUX2_X1 port map( A => n1314, B => DATAIN(7), S => n204, Z => n2577)
                           ;
   U1875 : MUX2_X1 port map( A => n1315, B => DATAIN(6), S => n204, Z => n2576)
                           ;
   U1876 : MUX2_X1 port map( A => n1316, B => DATAIN(5), S => n204, Z => n2575)
                           ;
   U1877 : MUX2_X1 port map( A => n1317, B => DATAIN(4), S => n204, Z => n2574)
                           ;
   U1878 : MUX2_X1 port map( A => n1318, B => DATAIN(3), S => n204, Z => n2573)
                           ;
   U1879 : MUX2_X1 port map( A => n1319, B => DATAIN(2), S => n204, Z => n2572)
                           ;
   U1880 : MUX2_X1 port map( A => n1320, B => DATAIN(1), S => n204, Z => n2571)
                           ;
   U1881 : MUX2_X1 port map( A => n1321, B => DATAIN(0), S => n204, Z => n2570)
                           ;
   U1882 : AND2_X1 port map( A1 => n1184, A2 => n872, ZN => n1290);
   U1883 : AND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2),
                           ZN => n872);
   U1884 : AND3_X1 port map( A1 => ADD_WR(3), A2 => n875, A3 => ADD_WR(4), ZN 
                           => n1184);
   U1885 : NOR2_X1 port map( A1 => n1322, A2 => n1323, ZN => n875);
   U1886 : INV_X1 port map( A => ENABLE, ZN => n1322);
   U1887 : OAI222_X1 port map( A1 => n593, A2 => n209, B1 => n1325, B2 => n212,
                           C1 => n3934, C2 => n215, ZN => n2569);
   U1888 : NOR4_X1 port map( A1 => n1328, A2 => n1329, A3 => n1330, A4 => n1331
                           , ZN => n1325);
   U1889 : OAI221_X1 port map( B1 => n837, B2 => n218, C1 => n1333, C2 => n221,
                           A => n1335, ZN => n1331);
   U1890 : AOI22_X1 port map( A1 => n224, A2 => n4062, B1 => n225, B2 => n1187,
                           ZN => n1335);
   U1891 : OAI221_X1 port map( B1 => n1338, B2 => n294, C1 => n933, C2 => n297,
                           A => n1341, ZN => n1330);
   U1892 : AOI22_X1 port map( A1 => n300, A2 => n1289, B1 => n303, B2 => n4030,
                           ZN => n1341);
   U1893 : OAI211_X1 port map( C1 => n517, C2 => n306, A => n1345, B => n1346, 
                           ZN => n1329);
   U1894 : AOI221_X1 port map( B1 => n307, B2 => n1148, C1 => n312, C2 => n4158
                           , A => n1349, ZN => n1346);
   U1895 : OAI22_X1 port map( A1 => n613, A2 => n315, B1 => n1351, B2 => n318, 
                           ZN => n1349);
   U1896 : AOI22_X1 port map( A1 => n321, A2 => n4190, B1 => n324, B2 => n1046,
                           ZN => n1345);
   U1897 : NAND4_X1 port map( A1 => n1358, A2 => n1356, A3 => n1357, A4 => 
                           n1355, ZN => n1328);
   U1898 : AOI221_X1 port map( B1 => n327, B2 => n4222, C1 => n330, C2 => n4254
                           , A => n1361, ZN => n1358);
   U1899 : OAI22_X1 port map( A1 => n389, A2 => n333, B1 => n357, B2 => n20, ZN
                           => n1361);
   U1900 : AOI221_X1 port map( B1 => n336, B2 => n4286, C1 => n339, C2 => n4318
                           , A => n1366, ZN => n1357);
   U1901 : OAI22_X1 port map( A1 => n261, A2 => n342, B1 => n229, B2 => n343, 
                           ZN => n1366);
   U1902 : AOI221_X1 port map( B1 => n348, B2 => n769, C1 => n351, C2 => n803, 
                           A => n1371, ZN => n1356);
   U1903 : OAI22_X1 port map( A1 => n1372, A2 => n354, B1 => n1374, B2 => n421,
                           ZN => n1371);
   U1904 : AOI221_X1 port map( B1 => n423, B2 => n730, C1 => n427, C2 => n3966,
                           A => n1378, ZN => n1355);
   U1905 : OAI22_X1 port map( A1 => n1379, A2 => n430, B1 => n1381, B2 => n22, 
                           ZN => n1378);
   U1906 : OAI222_X1 port map( A1 => n592, A2 => n209, B1 => n1383, B2 => n212,
                           C1 => n3933, C2 => n215, ZN => n2568);
   U1907 : NOR4_X1 port map( A1 => n1384, A2 => n1385, A3 => n1386, A4 => n1387
                           , ZN => n1383);
   U1908 : OAI221_X1 port map( B1 => n838, B2 => n218, C1 => n1388, C2 => n221,
                           A => n1389, ZN => n1387);
   U1909 : AOI22_X1 port map( A1 => n224, A2 => n4061, B1 => n30, B2 => n1189, 
                           ZN => n1389);
   U1910 : OAI221_X1 port map( B1 => n1390, B2 => n294, C1 => n934, C2 => n297,
                           A => n1391, ZN => n1386);
   U1911 : AOI22_X1 port map( A1 => n300, A2 => n1291, B1 => n303, B2 => n4029,
                           ZN => n1391);
   U1912 : OAI211_X1 port map( C1 => n518, C2 => n306, A => n1392, B => n1393, 
                           ZN => n1385);
   U1913 : AOI221_X1 port map( B1 => n307, B2 => n1150, C1 => n312, C2 => n4157
                           , A => n1394, ZN => n1393);
   U1914 : OAI22_X1 port map( A1 => n614, A2 => n315, B1 => n1395, B2 => n318, 
                           ZN => n1394);
   U1915 : AOI22_X1 port map( A1 => n321, A2 => n4189, B1 => n324, B2 => n1048,
                           ZN => n1392);
   U1916 : NAND4_X1 port map( A1 => n1396, A2 => n1397, A3 => n1398, A4 => 
                           n1399, ZN => n1384);
   U1917 : AOI221_X1 port map( B1 => n327, B2 => n4221, C1 => n330, C2 => n4253
                           , A => n1400, ZN => n1399);
   U1918 : OAI22_X1 port map( A1 => n390, A2 => n32, B1 => n358, B2 => n21, ZN 
                           => n1400);
   U1919 : AOI221_X1 port map( B1 => n336, B2 => n4285, C1 => n339, C2 => n4317
                           , A => n1401, ZN => n1398);
   U1920 : OAI22_X1 port map( A1 => n262, A2 => n33, B1 => n230, B2 => n345, ZN
                           => n1401);
   U1921 : AOI221_X1 port map( B1 => n348, B2 => n771, C1 => n351, C2 => n805, 
                           A => n1402, ZN => n1397);
   U1922 : OAI22_X1 port map( A1 => n1403, A2 => n354, B1 => n1404, B2 => n421,
                           ZN => n1402);
   U1923 : AOI221_X1 port map( B1 => n423, B2 => n732, C1 => n427, C2 => n3965,
                           A => n1405, ZN => n1396);
   U1924 : OAI22_X1 port map( A1 => n1406, A2 => n430, B1 => n1407, B2 => n5, 
                           ZN => n1405);
   U1925 : OAI222_X1 port map( A1 => n591, A2 => n209, B1 => n1408, B2 => n212,
                           C1 => n3932, C2 => n215, ZN => n2567);
   U1926 : NOR4_X1 port map( A1 => n1409, A2 => n1410, A3 => n1411, A4 => n1412
                           , ZN => n1408);
   U1927 : OAI221_X1 port map( B1 => n839, B2 => n218, C1 => n1413, C2 => n221,
                           A => n1414, ZN => n1412);
   U1928 : AOI22_X1 port map( A1 => n224, A2 => n4060, B1 => n29, B2 => n1190, 
                           ZN => n1414);
   U1929 : OAI221_X1 port map( B1 => n1415, B2 => n294, C1 => n935, C2 => n297,
                           A => n1416, ZN => n1411);
   U1930 : AOI22_X1 port map( A1 => n300, A2 => n1292, B1 => n303, B2 => n4028,
                           ZN => n1416);
   U1931 : OAI211_X1 port map( C1 => n519, C2 => n306, A => n1417, B => n1418, 
                           ZN => n1410);
   U1932 : AOI221_X1 port map( B1 => n309, B2 => n1151, C1 => n312, C2 => n4156
                           , A => n1419, ZN => n1418);
   U1933 : OAI22_X1 port map( A1 => n615, A2 => n315, B1 => n1420, B2 => n318, 
                           ZN => n1419);
   U1934 : AOI22_X1 port map( A1 => n321, A2 => n4188, B1 => n324, B2 => n1049,
                           ZN => n1417);
   U1935 : NAND4_X1 port map( A1 => n1424, A2 => n1422, A3 => n1423, A4 => 
                           n1421, ZN => n1409);
   U1936 : AOI221_X1 port map( B1 => n327, B2 => n4220, C1 => n330, C2 => n4252
                           , A => n1425, ZN => n1424);
   U1937 : OAI22_X1 port map( A1 => n391, A2 => n332, B1 => n359, B2 => n21, ZN
                           => n1425);
   U1938 : AOI221_X1 port map( B1 => n336, B2 => n4284, C1 => n339, C2 => n4316
                           , A => n1426, ZN => n1423);
   U1939 : OAI22_X1 port map( A1 => n263, A2 => n34, B1 => n231, B2 => n343, ZN
                           => n1426);
   U1940 : AOI221_X1 port map( B1 => n348, B2 => n772, C1 => n351, C2 => n806, 
                           A => n1427, ZN => n1422);
   U1941 : OAI22_X1 port map( A1 => n1428, A2 => n354, B1 => n1429, B2 => n421,
                           ZN => n1427);
   U1942 : AOI221_X1 port map( B1 => n423, B2 => n733, C1 => n427, C2 => n3964,
                           A => n1430, ZN => n1421);
   U1943 : OAI22_X1 port map( A1 => n1431, A2 => n430, B1 => n1432, B2 => n5, 
                           ZN => n1430);
   U1944 : OAI222_X1 port map( A1 => n590, A2 => n209, B1 => n1433, B2 => n212,
                           C1 => n3931, C2 => n215, ZN => n2566);
   U1945 : NOR4_X1 port map( A1 => n1434, A2 => n1435, A3 => n1436, A4 => n1437
                           , ZN => n1433);
   U1946 : OAI221_X1 port map( B1 => n840, B2 => n218, C1 => n1438, C2 => n221,
                           A => n1439, ZN => n1437);
   U1947 : AOI22_X1 port map( A1 => n224, A2 => n4059, B1 => n227, B2 => n1191,
                           ZN => n1439);
   U1948 : OAI221_X1 port map( B1 => n1440, B2 => n294, C1 => n936, C2 => n297,
                           A => n1441, ZN => n1436);
   U1949 : AOI22_X1 port map( A1 => n300, A2 => n1293, B1 => n303, B2 => n4027,
                           ZN => n1441);
   U1950 : OAI211_X1 port map( C1 => n520, C2 => n306, A => n1442, B => n1443, 
                           ZN => n1435);
   U1951 : AOI221_X1 port map( B1 => n308, B2 => n1152, C1 => n312, C2 => n4155
                           , A => n1444, ZN => n1443);
   U1952 : OAI22_X1 port map( A1 => n616, A2 => n315, B1 => n1445, B2 => n318, 
                           ZN => n1444);
   U1953 : AOI22_X1 port map( A1 => n321, A2 => n4187, B1 => n324, B2 => n1050,
                           ZN => n1442);
   U1954 : NAND4_X1 port map( A1 => n1449, A2 => n1447, A3 => n1448, A4 => 
                           n1446, ZN => n1434);
   U1955 : AOI221_X1 port map( B1 => n327, B2 => n4219, C1 => n330, C2 => n4251
                           , A => n1450, ZN => n1449);
   U1956 : OAI22_X1 port map( A1 => n392, A2 => n31, B1 => n360, B2 => n20, ZN 
                           => n1450);
   U1957 : AOI221_X1 port map( B1 => n336, B2 => n4283, C1 => n339, C2 => n4315
                           , A => n1451, ZN => n1448);
   U1958 : OAI22_X1 port map( A1 => n264, A2 => n341, B1 => n232, B2 => n343, 
                           ZN => n1451);
   U1959 : AOI221_X1 port map( B1 => n348, B2 => n773, C1 => n351, C2 => n807, 
                           A => n1452, ZN => n1447);
   U1960 : OAI22_X1 port map( A1 => n1453, A2 => n354, B1 => n1454, B2 => n421,
                           ZN => n1452);
   U1961 : AOI221_X1 port map( B1 => n422, B2 => n734, C1 => n427, C2 => n3963,
                           A => n1455, ZN => n1446);
   U1962 : OAI22_X1 port map( A1 => n1456, A2 => n430, B1 => n1457, B2 => n23, 
                           ZN => n1455);
   U1963 : OAI222_X1 port map( A1 => n589, A2 => n209, B1 => n1458, B2 => n212,
                           C1 => n3930, C2 => n215, ZN => n2565);
   U1964 : NOR4_X1 port map( A1 => n1459, A2 => n1460, A3 => n1461, A4 => n1462
                           , ZN => n1458);
   U1965 : OAI221_X1 port map( B1 => n841, B2 => n218, C1 => n1463, C2 => n221,
                           A => n1464, ZN => n1462);
   U1966 : AOI22_X1 port map( A1 => n224, A2 => n4058, B1 => n225, B2 => n1192,
                           ZN => n1464);
   U1967 : OAI221_X1 port map( B1 => n1465, B2 => n294, C1 => n937, C2 => n297,
                           A => n1466, ZN => n1461);
   U1968 : AOI22_X1 port map( A1 => n300, A2 => n1294, B1 => n303, B2 => n4026,
                           ZN => n1466);
   U1969 : OAI211_X1 port map( C1 => n521, C2 => n306, A => n1467, B => n1468, 
                           ZN => n1460);
   U1970 : AOI221_X1 port map( B1 => n309, B2 => n1153, C1 => n312, C2 => n4154
                           , A => n1469, ZN => n1468);
   U1971 : OAI22_X1 port map( A1 => n617, A2 => n315, B1 => n1470, B2 => n318, 
                           ZN => n1469);
   U1972 : AOI22_X1 port map( A1 => n321, A2 => n4186, B1 => n324, B2 => n1051,
                           ZN => n1467);
   U1973 : NAND4_X1 port map( A1 => n1474, A2 => n1472, A3 => n1473, A4 => 
                           n1471, ZN => n1459);
   U1974 : AOI221_X1 port map( B1 => n327, B2 => n4218, C1 => n330, C2 => n4250
                           , A => n1475, ZN => n1474);
   U1975 : OAI22_X1 port map( A1 => n393, A2 => n331, B1 => n361, B2 => n20, ZN
                           => n1475);
   U1976 : AOI221_X1 port map( B1 => n336, B2 => n4282, C1 => n339, C2 => n4314
                           , A => n1476, ZN => n1473);
   U1977 : OAI22_X1 port map( A1 => n265, A2 => n340, B1 => n233, B2 => n345, 
                           ZN => n1476);
   U1978 : AOI221_X1 port map( B1 => n348, B2 => n774, C1 => n351, C2 => n808, 
                           A => n1477, ZN => n1472);
   U1979 : OAI22_X1 port map( A1 => n1478, A2 => n354, B1 => n1479, B2 => n421,
                           ZN => n1477);
   U1980 : AOI221_X1 port map( B1 => n423, B2 => n735, C1 => n427, C2 => n3962,
                           A => n1480, ZN => n1471);
   U1981 : OAI22_X1 port map( A1 => n1481, A2 => n430, B1 => n1482, B2 => n23, 
                           ZN => n1480);
   U1982 : OAI222_X1 port map( A1 => n588, A2 => n209, B1 => n1483, B2 => n212,
                           C1 => n3929, C2 => n215, ZN => n2564);
   U1983 : NOR4_X1 port map( A1 => n1484, A2 => n1485, A3 => n1486, A4 => n1487
                           , ZN => n1483);
   U1984 : OAI221_X1 port map( B1 => n842, B2 => n218, C1 => n1488, C2 => n221,
                           A => n1489, ZN => n1487);
   U1985 : AOI22_X1 port map( A1 => n224, A2 => n4057, B1 => n30, B2 => n1193, 
                           ZN => n1489);
   U1986 : OAI221_X1 port map( B1 => n1490, B2 => n294, C1 => n938, C2 => n297,
                           A => n1491, ZN => n1486);
   U1987 : AOI22_X1 port map( A1 => n300, A2 => n1295, B1 => n303, B2 => n4025,
                           ZN => n1491);
   U1988 : OAI211_X1 port map( C1 => n522, C2 => n306, A => n1492, B => n1493, 
                           ZN => n1485);
   U1989 : AOI221_X1 port map( B1 => n308, B2 => n1154, C1 => n312, C2 => n4153
                           , A => n1494, ZN => n1493);
   U1990 : OAI22_X1 port map( A1 => n618, A2 => n315, B1 => n1495, B2 => n318, 
                           ZN => n1494);
   U1991 : AOI22_X1 port map( A1 => n321, A2 => n4185, B1 => n324, B2 => n1052,
                           ZN => n1492);
   U1992 : NAND4_X1 port map( A1 => n1499, A2 => n1497, A3 => n1498, A4 => 
                           n1496, ZN => n1484);
   U1993 : AOI221_X1 port map( B1 => n327, B2 => n4217, C1 => n330, C2 => n4249
                           , A => n1500, ZN => n1499);
   U1994 : OAI22_X1 port map( A1 => n394, A2 => n333, B1 => n362, B2 => n20, ZN
                           => n1500);
   U1995 : AOI221_X1 port map( B1 => n336, B2 => n4281, C1 => n339, C2 => n4313
                           , A => n1501, ZN => n1498);
   U1996 : OAI22_X1 port map( A1 => n266, A2 => n342, B1 => n234, B2 => n345, 
                           ZN => n1501);
   U1997 : AOI221_X1 port map( B1 => n348, B2 => n775, C1 => n351, C2 => n809, 
                           A => n1502, ZN => n1497);
   U1998 : OAI22_X1 port map( A1 => n1503, A2 => n354, B1 => n1504, B2 => n421,
                           ZN => n1502);
   U1999 : AOI221_X1 port map( B1 => n422, B2 => n736, C1 => n427, C2 => n3961,
                           A => n1505, ZN => n1496);
   U2000 : OAI22_X1 port map( A1 => n1506, A2 => n430, B1 => n1507, B2 => n22, 
                           ZN => n1505);
   U2001 : OAI222_X1 port map( A1 => n587, A2 => n209, B1 => n1508, B2 => n212,
                           C1 => n3928, C2 => n215, ZN => n2563);
   U2002 : NOR4_X1 port map( A1 => n1509, A2 => n1510, A3 => n1511, A4 => n1512
                           , ZN => n1508);
   U2003 : OAI221_X1 port map( B1 => n843, B2 => n218, C1 => n1513, C2 => n221,
                           A => n1514, ZN => n1512);
   U2004 : AOI22_X1 port map( A1 => n224, A2 => n4056, B1 => n29, B2 => n1194, 
                           ZN => n1514);
   U2005 : OAI221_X1 port map( B1 => n1515, B2 => n294, C1 => n939, C2 => n297,
                           A => n1516, ZN => n1511);
   U2006 : AOI22_X1 port map( A1 => n300, A2 => n1296, B1 => n303, B2 => n4024,
                           ZN => n1516);
   U2007 : OAI211_X1 port map( C1 => n523, C2 => n306, A => n1517, B => n1518, 
                           ZN => n1510);
   U2008 : AOI221_X1 port map( B1 => n309, B2 => n1155, C1 => n312, C2 => n4152
                           , A => n1519, ZN => n1518);
   U2009 : OAI22_X1 port map( A1 => n619, A2 => n315, B1 => n1520, B2 => n318, 
                           ZN => n1519);
   U2010 : AOI22_X1 port map( A1 => n321, A2 => n4184, B1 => n324, B2 => n1053,
                           ZN => n1517);
   U2011 : NAND4_X1 port map( A1 => n1524, A2 => n1522, A3 => n1523, A4 => 
                           n1521, ZN => n1509);
   U2012 : AOI221_X1 port map( B1 => n327, B2 => n4216, C1 => n330, C2 => n4248
                           , A => n1525, ZN => n1524);
   U2013 : OAI22_X1 port map( A1 => n395, A2 => n332, B1 => n363, B2 => n21, ZN
                           => n1525);
   U2014 : AOI221_X1 port map( B1 => n336, B2 => n4280, C1 => n339, C2 => n4312
                           , A => n1526, ZN => n1523);
   U2015 : OAI22_X1 port map( A1 => n267, A2 => n33, B1 => n235, B2 => n343, ZN
                           => n1526);
   U2016 : AOI221_X1 port map( B1 => n348, B2 => n776, C1 => n351, C2 => n810, 
                           A => n1527, ZN => n1522);
   U2017 : OAI22_X1 port map( A1 => n1528, A2 => n354, B1 => n1529, B2 => n421,
                           ZN => n1527);
   U2018 : AOI221_X1 port map( B1 => n423, B2 => n737, C1 => n427, C2 => n3960,
                           A => n1530, ZN => n1521);
   U2019 : OAI22_X1 port map( A1 => n1531, A2 => n430, B1 => n1532, B2 => n23, 
                           ZN => n1530);
   U2020 : OAI222_X1 port map( A1 => n586, A2 => n209, B1 => n1533, B2 => n212,
                           C1 => n3927, C2 => n215, ZN => n2562);
   U2021 : NOR4_X1 port map( A1 => n1534, A2 => n1535, A3 => n1536, A4 => n1537
                           , ZN => n1533);
   U2022 : OAI221_X1 port map( B1 => n844, B2 => n218, C1 => n1538, C2 => n221,
                           A => n1539, ZN => n1537);
   U2023 : AOI22_X1 port map( A1 => n224, A2 => n4055, B1 => n227, B2 => n1195,
                           ZN => n1539);
   U2024 : OAI221_X1 port map( B1 => n1540, B2 => n294, C1 => n940, C2 => n297,
                           A => n1541, ZN => n1536);
   U2025 : AOI22_X1 port map( A1 => n300, A2 => n1297, B1 => n303, B2 => n4023,
                           ZN => n1541);
   U2026 : OAI211_X1 port map( C1 => n524, C2 => n306, A => n1542, B => n1543, 
                           ZN => n1535);
   U2027 : AOI221_X1 port map( B1 => n309, B2 => n1156, C1 => n312, C2 => n4151
                           , A => n1544, ZN => n1543);
   U2028 : OAI22_X1 port map( A1 => n620, A2 => n315, B1 => n1545, B2 => n318, 
                           ZN => n1544);
   U2029 : AOI22_X1 port map( A1 => n321, A2 => n4183, B1 => n324, B2 => n1054,
                           ZN => n1542);
   U2030 : NAND4_X1 port map( A1 => n1546, A2 => n1547, A3 => n1548, A4 => 
                           n1549, ZN => n1534);
   U2031 : AOI221_X1 port map( B1 => n327, B2 => n4215, C1 => n330, C2 => n4247
                           , A => n1550, ZN => n1549);
   U2032 : OAI22_X1 port map( A1 => n396, A2 => n331, B1 => n364, B2 => n21, ZN
                           => n1550);
   U2033 : AOI221_X1 port map( B1 => n336, B2 => n4279, C1 => n339, C2 => n4311
                           , A => n1551, ZN => n1548);
   U2034 : OAI22_X1 port map( A1 => n268, A2 => n34, B1 => n236, B2 => n345, ZN
                           => n1551);
   U2035 : AOI221_X1 port map( B1 => n348, B2 => n777, C1 => n351, C2 => n811, 
                           A => n1552, ZN => n1547);
   U2036 : OAI22_X1 port map( A1 => n1553, A2 => n354, B1 => n1554, B2 => n421,
                           ZN => n1552);
   U2037 : AOI221_X1 port map( B1 => n422, B2 => n738, C1 => n427, C2 => n3959,
                           A => n1555, ZN => n1546);
   U2038 : OAI22_X1 port map( A1 => n1556, A2 => n430, B1 => n1557, B2 => n22, 
                           ZN => n1555);
   U2039 : OAI222_X1 port map( A1 => n585, A2 => n208, B1 => n1558, B2 => n211,
                           C1 => n3926, C2 => n215, ZN => n2561);
   U2040 : NOR4_X1 port map( A1 => n1559, A2 => n1560, A3 => n1561, A4 => n1562
                           , ZN => n1558);
   U2041 : OAI221_X1 port map( B1 => n845, B2 => n217, C1 => n1563, C2 => n220,
                           A => n1564, ZN => n1562);
   U2042 : AOI22_X1 port map( A1 => n223, A2 => n4054, B1 => n225, B2 => n1196,
                           ZN => n1564);
   U2043 : OAI221_X1 port map( B1 => n1565, B2 => n293, C1 => n941, C2 => n296,
                           A => n1566, ZN => n1561);
   U2044 : AOI22_X1 port map( A1 => n299, A2 => n1298, B1 => n302, B2 => n4022,
                           ZN => n1566);
   U2045 : OAI211_X1 port map( C1 => n525, C2 => n305, A => n1567, B => n1568, 
                           ZN => n1560);
   U2046 : AOI221_X1 port map( B1 => n307, B2 => n1157, C1 => n311, C2 => n4150
                           , A => n1569, ZN => n1568);
   U2047 : OAI22_X1 port map( A1 => n621, A2 => n314, B1 => n1570, B2 => n317, 
                           ZN => n1569);
   U2048 : AOI22_X1 port map( A1 => n320, A2 => n4182, B1 => n323, B2 => n1055,
                           ZN => n1567);
   U2049 : NAND4_X1 port map( A1 => n1574, A2 => n1571, A3 => n1572, A4 => 
                           n1573, ZN => n1559);
   U2050 : AOI221_X1 port map( B1 => n326, B2 => n4214, C1 => n329, C2 => n4246
                           , A => n1575, ZN => n1574);
   U2051 : OAI22_X1 port map( A1 => n397, A2 => n31, B1 => n365, B2 => n21, ZN 
                           => n1575);
   U2052 : AOI221_X1 port map( B1 => n335, B2 => n4278, C1 => n338, C2 => n4310
                           , A => n1576, ZN => n1573);
   U2053 : OAI22_X1 port map( A1 => n269, A2 => n341, B1 => n237, B2 => n344, 
                           ZN => n1576);
   U2054 : AOI221_X1 port map( B1 => n347, B2 => n778, C1 => n350, C2 => n812, 
                           A => n1577, ZN => n1572);
   U2055 : OAI22_X1 port map( A1 => n1578, A2 => n353, B1 => n1579, B2 => n356,
                           ZN => n1577);
   U2056 : OAI22_X1 port map( A1 => n1581, A2 => n429, B1 => n1582, B2 => n5, 
                           ZN => n1580);
   U2057 : OAI222_X1 port map( A1 => n584, A2 => n208, B1 => n1583, B2 => n211,
                           C1 => n3925, C2 => n215, ZN => n2560);
   U2058 : OAI221_X1 port map( B1 => n846, B2 => n217, C1 => n1588, C2 => n220,
                           A => n1589, ZN => n1587);
   U2059 : AOI22_X1 port map( A1 => n223, A2 => n4053, B1 => n29, B2 => n1197, 
                           ZN => n1589);
   U2060 : OAI221_X1 port map( B1 => n1590, B2 => n293, C1 => n942, C2 => n296,
                           A => n1591, ZN => n1586);
   U2061 : AOI22_X1 port map( A1 => n299, A2 => n1299, B1 => n302, B2 => n4021,
                           ZN => n1591);
   U2062 : OAI211_X1 port map( C1 => n526, C2 => n305, A => n1592, B => n1593, 
                           ZN => n1585);
   U2063 : AOI221_X1 port map( B1 => n308, B2 => n1158, C1 => n311, C2 => n4149
                           , A => n1594, ZN => n1593);
   U2064 : OAI22_X1 port map( A1 => n622, A2 => n314, B1 => n1595, B2 => n317, 
                           ZN => n1594);
   U2065 : AOI22_X1 port map( A1 => n320, A2 => n4181, B1 => n323, B2 => n1056,
                           ZN => n1592);
   U2066 : NAND4_X1 port map( A1 => n1596, A2 => n1597, A3 => n1598, A4 => 
                           n1599, ZN => n1584);
   U2067 : AOI221_X1 port map( B1 => n326, B2 => n4213, C1 => n329, C2 => n4245
                           , A => n1600, ZN => n1599);
   U2068 : OAI22_X1 port map( A1 => n398, A2 => n332, B1 => n366, B2 => n21, ZN
                           => n1600);
   U2069 : AOI221_X1 port map( B1 => n335, B2 => n4277, C1 => n338, C2 => n4309
                           , A => n1601, ZN => n1598);
   U2070 : OAI22_X1 port map( A1 => n270, A2 => n341, B1 => n238, B2 => n345, 
                           ZN => n1601);
   U2071 : AOI221_X1 port map( B1 => n347, B2 => n779, C1 => n350, C2 => n813, 
                           A => n1602, ZN => n1597);
   U2072 : OAI22_X1 port map( A1 => n1603, A2 => n353, B1 => n1604, B2 => n356,
                           ZN => n1602);
   U2073 : AOI221_X1 port map( B1 => n422, B2 => n740, C1 => n426, C2 => n3957,
                           A => n1605, ZN => n1596);
   U2074 : OAI22_X1 port map( A1 => n1606, A2 => n429, B1 => n1607, B2 => n23, 
                           ZN => n1605);
   U2075 : OAI222_X1 port map( A1 => n583, A2 => n208, B1 => n1608, B2 => n211,
                           C1 => n3924, C2 => n214, ZN => n2559);
   U2076 : NOR4_X1 port map( A1 => n1609, A2 => n1610, A3 => n1611, A4 => n1612
                           , ZN => n1608);
   U2077 : OAI221_X1 port map( B1 => n847, B2 => n217, C1 => n1613, C2 => n220,
                           A => n1614, ZN => n1612);
   U2078 : AOI22_X1 port map( A1 => n223, A2 => n4052, B1 => n30, B2 => n1198, 
                           ZN => n1614);
   U2079 : OAI221_X1 port map( B1 => n1615, B2 => n293, C1 => n943, C2 => n296,
                           A => n1616, ZN => n1611);
   U2080 : AOI22_X1 port map( A1 => n299, A2 => n1300, B1 => n302, B2 => n4020,
                           ZN => n1616);
   U2081 : OAI211_X1 port map( C1 => n527, C2 => n305, A => n1617, B => n1618, 
                           ZN => n1610);
   U2082 : AOI221_X1 port map( B1 => n307, B2 => n1159, C1 => n311, C2 => n4148
                           , A => n1619, ZN => n1618);
   U2083 : OAI22_X1 port map( A1 => n623, A2 => n314, B1 => n1620, B2 => n317, 
                           ZN => n1619);
   U2084 : AOI22_X1 port map( A1 => n320, A2 => n4180, B1 => n323, B2 => n1057,
                           ZN => n1617);
   U2085 : NAND4_X1 port map( A1 => n1624, A2 => n1621, A3 => n1622, A4 => 
                           n1623, ZN => n1609);
   U2086 : AOI221_X1 port map( B1 => n326, B2 => n4212, C1 => n329, C2 => n4244
                           , A => n1625, ZN => n1624);
   U2087 : OAI22_X1 port map( A1 => n399, A2 => n332, B1 => n367, B2 => n20, ZN
                           => n1625);
   U2088 : AOI221_X1 port map( B1 => n335, B2 => n4276, C1 => n338, C2 => n4308
                           , A => n1626, ZN => n1623);
   U2089 : OAI22_X1 port map( A1 => n271, A2 => n340, B1 => n239, B2 => n344, 
                           ZN => n1626);
   U2090 : AOI221_X1 port map( B1 => n347, B2 => n780, C1 => n350, C2 => n814, 
                           A => n1627, ZN => n1622);
   U2091 : OAI22_X1 port map( A1 => n1628, A2 => n353, B1 => n1629, B2 => n356,
                           ZN => n1627);
   U2092 : OAI22_X1 port map( A1 => n1631, A2 => n429, B1 => n1632, B2 => n23, 
                           ZN => n1630);
   U2093 : OAI222_X1 port map( A1 => n582, A2 => n208, B1 => n1633, B2 => n211,
                           C1 => n3923, C2 => n214, ZN => n2558);
   U2094 : OAI221_X1 port map( B1 => n848, B2 => n217, C1 => n1638, C2 => n220,
                           A => n1639, ZN => n1637);
   U2095 : AOI22_X1 port map( A1 => n223, A2 => n4051, B1 => n227, B2 => n1199,
                           ZN => n1639);
   U2096 : OAI221_X1 port map( B1 => n1640, B2 => n293, C1 => n944, C2 => n296,
                           A => n1641, ZN => n1636);
   U2097 : AOI22_X1 port map( A1 => n299, A2 => n1301, B1 => n302, B2 => n4019,
                           ZN => n1641);
   U2098 : OAI211_X1 port map( C1 => n528, C2 => n305, A => n1642, B => n1643, 
                           ZN => n1635);
   U2099 : AOI221_X1 port map( B1 => n309, B2 => n1160, C1 => n311, C2 => n4147
                           , A => n1644, ZN => n1643);
   U2100 : OAI22_X1 port map( A1 => n624, A2 => n314, B1 => n1645, B2 => n317, 
                           ZN => n1644);
   U2101 : AOI22_X1 port map( A1 => n320, A2 => n4179, B1 => n323, B2 => n1058,
                           ZN => n1642);
   U2102 : NAND4_X1 port map( A1 => n1646, A2 => n1647, A3 => n1648, A4 => 
                           n1649, ZN => n1634);
   U2103 : AOI221_X1 port map( B1 => n326, B2 => n4211, C1 => n329, C2 => n4243
                           , A => n1650, ZN => n1649);
   U2104 : OAI22_X1 port map( A1 => n400, A2 => n333, B1 => n368, B2 => n20, ZN
                           => n1650);
   U2105 : AOI221_X1 port map( B1 => n335, B2 => n4275, C1 => n338, C2 => n4307
                           , A => n1651, ZN => n1648);
   U2106 : OAI22_X1 port map( A1 => n272, A2 => n340, B1 => n240, B2 => n343, 
                           ZN => n1651);
   U2107 : AOI221_X1 port map( B1 => n347, B2 => n781, C1 => n350, C2 => n815, 
                           A => n1652, ZN => n1647);
   U2108 : OAI22_X1 port map( A1 => n1653, A2 => n353, B1 => n1654, B2 => n356,
                           ZN => n1652);
   U2109 : AOI221_X1 port map( B1 => n423, B2 => n742, C1 => n426, C2 => n3955,
                           A => n1655, ZN => n1646);
   U2110 : OAI22_X1 port map( A1 => n1656, A2 => n429, B1 => n1657, B2 => n22, 
                           ZN => n1655);
   U2111 : OAI222_X1 port map( A1 => n581, A2 => n208, B1 => n1658, B2 => n211,
                           C1 => n3922, C2 => n214, ZN => n2557);
   U2112 : NOR4_X1 port map( A1 => n1659, A2 => n1660, A3 => n1661, A4 => n1662
                           , ZN => n1658);
   U2113 : OAI221_X1 port map( B1 => n849, B2 => n217, C1 => n1663, C2 => n220,
                           A => n1664, ZN => n1662);
   U2114 : AOI22_X1 port map( A1 => n223, A2 => n4050, B1 => n29, B2 => n1200, 
                           ZN => n1664);
   U2115 : OAI221_X1 port map( B1 => n1665, B2 => n293, C1 => n945, C2 => n296,
                           A => n1666, ZN => n1661);
   U2116 : AOI22_X1 port map( A1 => n299, A2 => n1302, B1 => n302, B2 => n4018,
                           ZN => n1666);
   U2117 : OAI211_X1 port map( C1 => n529, C2 => n305, A => n1667, B => n1668, 
                           ZN => n1660);
   U2118 : AOI221_X1 port map( B1 => n307, B2 => n1161, C1 => n311, C2 => n4146
                           , A => n1669, ZN => n1668);
   U2119 : OAI22_X1 port map( A1 => n625, A2 => n314, B1 => n1670, B2 => n317, 
                           ZN => n1669);
   U2120 : AOI22_X1 port map( A1 => n320, A2 => n4178, B1 => n323, B2 => n1059,
                           ZN => n1667);
   U2121 : NAND4_X1 port map( A1 => n1674, A2 => n1671, A3 => n1673, A4 => 
                           n1672, ZN => n1659);
   U2122 : AOI221_X1 port map( B1 => n326, B2 => n4210, C1 => n329, C2 => n4242
                           , A => n1675, ZN => n1674);
   U2123 : OAI22_X1 port map( A1 => n401, A2 => n333, B1 => n369, B2 => n20, ZN
                           => n1675);
   U2124 : AOI221_X1 port map( B1 => n335, B2 => n4274, C1 => n338, C2 => n4306
                           , A => n1676, ZN => n1673);
   U2125 : OAI22_X1 port map( A1 => n273, A2 => n342, B1 => n241, B2 => n344, 
                           ZN => n1676);
   U2126 : AOI221_X1 port map( B1 => n347, B2 => n782, C1 => n350, C2 => n816, 
                           A => n1677, ZN => n1672);
   U2127 : OAI22_X1 port map( A1 => n1678, A2 => n353, B1 => n1679, B2 => n356,
                           ZN => n1677);
   U2128 : OAI22_X1 port map( A1 => n1681, A2 => n429, B1 => n1682, B2 => n5, 
                           ZN => n1680);
   U2129 : OAI222_X1 port map( A1 => n580, A2 => n208, B1 => n1683, B2 => n211,
                           C1 => n3921, C2 => n214, ZN => n2556);
   U2130 : OAI221_X1 port map( B1 => n850, B2 => n217, C1 => n1688, C2 => n220,
                           A => n1689, ZN => n1687);
   U2131 : AOI22_X1 port map( A1 => n223, A2 => n4049, B1 => n225, B2 => n1201,
                           ZN => n1689);
   U2132 : OAI221_X1 port map( B1 => n1690, B2 => n293, C1 => n946, C2 => n296,
                           A => n1691, ZN => n1686);
   U2133 : AOI22_X1 port map( A1 => n299, A2 => n1303, B1 => n302, B2 => n4017,
                           ZN => n1691);
   U2134 : OAI211_X1 port map( C1 => n530, C2 => n305, A => n1692, B => n1693, 
                           ZN => n1685);
   U2135 : AOI221_X1 port map( B1 => n308, B2 => n1162, C1 => n311, C2 => n4145
                           , A => n1694, ZN => n1693);
   U2136 : OAI22_X1 port map( A1 => n626, A2 => n314, B1 => n1695, B2 => n317, 
                           ZN => n1694);
   U2137 : AOI22_X1 port map( A1 => n320, A2 => n4177, B1 => n323, B2 => n1060,
                           ZN => n1692);
   U2138 : NAND4_X1 port map( A1 => n1696, A2 => n1697, A3 => n1698, A4 => 
                           n1699, ZN => n1684);
   U2139 : AOI221_X1 port map( B1 => n326, B2 => n4209, C1 => n329, C2 => n4241
                           , A => n1700, ZN => n1699);
   U2140 : OAI22_X1 port map( A1 => n402, A2 => n32, B1 => n370, B2 => n20, ZN 
                           => n1700);
   U2141 : AOI221_X1 port map( B1 => n335, B2 => n4273, C1 => n338, C2 => n4305
                           , A => n1701, ZN => n1698);
   U2142 : OAI22_X1 port map( A1 => n274, A2 => n342, B1 => n242, B2 => n345, 
                           ZN => n1701);
   U2143 : AOI221_X1 port map( B1 => n347, B2 => n783, C1 => n350, C2 => n817, 
                           A => n1702, ZN => n1697);
   U2144 : OAI22_X1 port map( A1 => n1703, A2 => n353, B1 => n1704, B2 => n356,
                           ZN => n1702);
   U2145 : AOI221_X1 port map( B1 => n422, B2 => n744, C1 => n426, C2 => n3953,
                           A => n1705, ZN => n1696);
   U2146 : OAI22_X1 port map( A1 => n1706, A2 => n429, B1 => n1707, B2 => n23, 
                           ZN => n1705);
   U2147 : OAI222_X1 port map( A1 => n579, A2 => n208, B1 => n1708, B2 => n211,
                           C1 => n3920, C2 => n214, ZN => n2555);
   U2148 : NOR4_X1 port map( A1 => n1709, A2 => n1710, A3 => n1711, A4 => n1712
                           , ZN => n1708);
   U2149 : OAI221_X1 port map( B1 => n851, B2 => n217, C1 => n1713, C2 => n220,
                           A => n1714, ZN => n1712);
   U2150 : AOI22_X1 port map( A1 => n223, A2 => n4048, B1 => n227, B2 => n1202,
                           ZN => n1714);
   U2151 : OAI221_X1 port map( B1 => n1715, B2 => n293, C1 => n947, C2 => n296,
                           A => n1716, ZN => n1711);
   U2152 : AOI22_X1 port map( A1 => n299, A2 => n1304, B1 => n302, B2 => n4016,
                           ZN => n1716);
   U2153 : OAI211_X1 port map( C1 => n531, C2 => n305, A => n1717, B => n1718, 
                           ZN => n1710);
   U2154 : AOI221_X1 port map( B1 => n307, B2 => n1163, C1 => n311, C2 => n4144
                           , A => n1719, ZN => n1718);
   U2155 : OAI22_X1 port map( A1 => n627, A2 => n314, B1 => n1720, B2 => n317, 
                           ZN => n1719);
   U2156 : AOI22_X1 port map( A1 => n320, A2 => n4176, B1 => n323, B2 => n1061,
                           ZN => n1717);
   U2157 : NAND4_X1 port map( A1 => n1724, A2 => n1721, A3 => n1722, A4 => 
                           n1723, ZN => n1709);
   U2158 : AOI221_X1 port map( B1 => n326, B2 => n4208, C1 => n329, C2 => n4240
                           , A => n1725, ZN => n1724);
   U2159 : OAI22_X1 port map( A1 => n403, A2 => n32, B1 => n371, B2 => n21, ZN 
                           => n1725);
   U2160 : AOI221_X1 port map( B1 => n335, B2 => n4272, C1 => n338, C2 => n4304
                           , A => n1726, ZN => n1723);
   U2161 : OAI22_X1 port map( A1 => n275, A2 => n33, B1 => n243, B2 => n344, ZN
                           => n1726);
   U2162 : AOI221_X1 port map( B1 => n347, B2 => n784, C1 => n350, C2 => n818, 
                           A => n1727, ZN => n1722);
   U2163 : OAI22_X1 port map( A1 => n1728, A2 => n353, B1 => n1729, B2 => n356,
                           ZN => n1727);
   U2164 : OAI22_X1 port map( A1 => n1731, A2 => n429, B1 => n1732, B2 => n22, 
                           ZN => n1730);
   U2165 : OAI222_X1 port map( A1 => n578, A2 => n208, B1 => n1733, B2 => n211,
                           C1 => n3919, C2 => n214, ZN => n2554);
   U2166 : OAI221_X1 port map( B1 => n852, B2 => n217, C1 => n1738, C2 => n220,
                           A => n1739, ZN => n1737);
   U2167 : AOI22_X1 port map( A1 => n223, A2 => n4047, B1 => n225, B2 => n1203,
                           ZN => n1739);
   U2168 : OAI221_X1 port map( B1 => n1740, B2 => n293, C1 => n948, C2 => n296,
                           A => n1741, ZN => n1736);
   U2169 : AOI22_X1 port map( A1 => n299, A2 => n1305, B1 => n302, B2 => n4015,
                           ZN => n1741);
   U2170 : OAI211_X1 port map( C1 => n532, C2 => n305, A => n1742, B => n1743, 
                           ZN => n1735);
   U2171 : AOI221_X1 port map( B1 => n309, B2 => n1164, C1 => n311, C2 => n4143
                           , A => n1744, ZN => n1743);
   U2172 : OAI22_X1 port map( A1 => n628, A2 => n314, B1 => n1745, B2 => n317, 
                           ZN => n1744);
   U2173 : AOI22_X1 port map( A1 => n320, A2 => n4175, B1 => n323, B2 => n1062,
                           ZN => n1742);
   U2174 : NAND4_X1 port map( A1 => n1746, A2 => n1747, A3 => n1748, A4 => 
                           n1749, ZN => n1734);
   U2175 : AOI221_X1 port map( B1 => n326, B2 => n4207, C1 => n329, C2 => n4239
                           , A => n1750, ZN => n1749);
   U2176 : OAI22_X1 port map( A1 => n404, A2 => n32, B1 => n372, B2 => n21, ZN 
                           => n1750);
   U2177 : AOI221_X1 port map( B1 => n335, B2 => n4271, C1 => n338, C2 => n4303
                           , A => n1751, ZN => n1748);
   U2178 : OAI22_X1 port map( A1 => n276, A2 => n33, B1 => n244, B2 => n343, ZN
                           => n1751);
   U2179 : AOI221_X1 port map( B1 => n347, B2 => n785, C1 => n350, C2 => n819, 
                           A => n1752, ZN => n1747);
   U2180 : OAI22_X1 port map( A1 => n1753, A2 => n353, B1 => n1754, B2 => n356,
                           ZN => n1752);
   U2181 : AOI221_X1 port map( B1 => n423, B2 => n746, C1 => n426, C2 => n3951,
                           A => n1755, ZN => n1746);
   U2182 : OAI22_X1 port map( A1 => n1756, A2 => n429, B1 => n1757, B2 => n23, 
                           ZN => n1755);
   U2183 : OAI222_X1 port map( A1 => n577, A2 => n208, B1 => n1758, B2 => n211,
                           C1 => n3918, C2 => n214, ZN => n2553);
   U2184 : NOR4_X1 port map( A1 => n1759, A2 => n1760, A3 => n1761, A4 => n1762
                           , ZN => n1758);
   U2185 : OAI221_X1 port map( B1 => n853, B2 => n217, C1 => n1763, C2 => n220,
                           A => n1764, ZN => n1762);
   U2186 : AOI22_X1 port map( A1 => n223, A2 => n4046, B1 => n225, B2 => n1204,
                           ZN => n1764);
   U2187 : OAI221_X1 port map( B1 => n1765, B2 => n293, C1 => n949, C2 => n296,
                           A => n1766, ZN => n1761);
   U2188 : AOI22_X1 port map( A1 => n299, A2 => n1306, B1 => n302, B2 => n4014,
                           ZN => n1766);
   U2189 : OAI211_X1 port map( C1 => n533, C2 => n305, A => n1767, B => n1768, 
                           ZN => n1760);
   U2190 : AOI221_X1 port map( B1 => n307, B2 => n1165, C1 => n311, C2 => n4142
                           , A => n1769, ZN => n1768);
   U2191 : OAI22_X1 port map( A1 => n629, A2 => n314, B1 => n1770, B2 => n317, 
                           ZN => n1769);
   U2192 : AOI22_X1 port map( A1 => n320, A2 => n4174, B1 => n323, B2 => n1063,
                           ZN => n1767);
   U2193 : NAND4_X1 port map( A1 => n1774, A2 => n1771, A3 => n1772, A4 => 
                           n1773, ZN => n1759);
   U2194 : AOI221_X1 port map( B1 => n326, B2 => n4206, C1 => n329, C2 => n4238
                           , A => n1775, ZN => n1774);
   U2195 : OAI22_X1 port map( A1 => n405, A2 => n32, B1 => n373, B2 => n20, ZN 
                           => n1775);
   U2196 : AOI221_X1 port map( B1 => n335, B2 => n4270, C1 => n338, C2 => n4302
                           , A => n1776, ZN => n1773);
   U2197 : OAI22_X1 port map( A1 => n277, A2 => n34, B1 => n245, B2 => n344, ZN
                           => n1776);
   U2198 : AOI221_X1 port map( B1 => n347, B2 => n786, C1 => n350, C2 => n820, 
                           A => n1777, ZN => n1772);
   U2199 : OAI22_X1 port map( A1 => n1778, A2 => n353, B1 => n1779, B2 => n356,
                           ZN => n1777);
   U2200 : OAI22_X1 port map( A1 => n1781, A2 => n429, B1 => n1782, B2 => n22, 
                           ZN => n1780);
   U2201 : OAI222_X1 port map( A1 => n576, A2 => n208, B1 => n1783, B2 => n211,
                           C1 => n3917, C2 => n214, ZN => n2552);
   U2202 : OAI221_X1 port map( B1 => n854, B2 => n217, C1 => n1788, C2 => n220,
                           A => n1789, ZN => n1787);
   U2203 : AOI22_X1 port map( A1 => n223, A2 => n4045, B1 => n30, B2 => n1205, 
                           ZN => n1789);
   U2204 : OAI221_X1 port map( B1 => n1790, B2 => n293, C1 => n950, C2 => n296,
                           A => n1791, ZN => n1786);
   U2205 : AOI22_X1 port map( A1 => n299, A2 => n1307, B1 => n302, B2 => n4013,
                           ZN => n1791);
   U2206 : OAI211_X1 port map( C1 => n534, C2 => n305, A => n1792, B => n1793, 
                           ZN => n1785);
   U2207 : AOI221_X1 port map( B1 => n308, B2 => n1166, C1 => n311, C2 => n4141
                           , A => n1794, ZN => n1793);
   U2208 : OAI22_X1 port map( A1 => n630, A2 => n314, B1 => n1795, B2 => n317, 
                           ZN => n1794);
   U2209 : AOI22_X1 port map( A1 => n320, A2 => n4173, B1 => n323, B2 => n1064,
                           ZN => n1792);
   U2210 : NAND4_X1 port map( A1 => n1796, A2 => n1797, A3 => n1798, A4 => 
                           n1799, ZN => n1784);
   U2211 : AOI221_X1 port map( B1 => n326, B2 => n4205, C1 => n329, C2 => n4237
                           , A => n1800, ZN => n1799);
   U2212 : OAI22_X1 port map( A1 => n406, A2 => n31, B1 => n374, B2 => n21, ZN 
                           => n1800);
   U2213 : AOI221_X1 port map( B1 => n335, B2 => n4269, C1 => n338, C2 => n4301
                           , A => n1801, ZN => n1798);
   U2214 : OAI22_X1 port map( A1 => n278, A2 => n34, B1 => n246, B2 => n345, ZN
                           => n1801);
   U2215 : AOI221_X1 port map( B1 => n347, B2 => n787, C1 => n350, C2 => n821, 
                           A => n1802, ZN => n1797);
   U2216 : OAI22_X1 port map( A1 => n1803, A2 => n353, B1 => n1804, B2 => n356,
                           ZN => n1802);
   U2217 : AOI221_X1 port map( B1 => n422, B2 => n748, C1 => n426, C2 => n3949,
                           A => n1805, ZN => n1796);
   U2218 : OAI22_X1 port map( A1 => n1806, A2 => n429, B1 => n1807, B2 => n22, 
                           ZN => n1805);
   U2219 : OAI222_X1 port map( A1 => n575, A2 => n208, B1 => n1808, B2 => n211,
                           C1 => n3916, C2 => n214, ZN => n2551);
   U2220 : OAI221_X1 port map( B1 => n855, B2 => n217, C1 => n1813, C2 => n220,
                           A => n1814, ZN => n1812);
   U2221 : AOI22_X1 port map( A1 => n223, A2 => n4044, B1 => n226, B2 => n1206,
                           ZN => n1814);
   U2222 : OAI221_X1 port map( B1 => n1815, B2 => n293, C1 => n951, C2 => n296,
                           A => n1816, ZN => n1811);
   U2223 : AOI22_X1 port map( A1 => n299, A2 => n1308, B1 => n302, B2 => n4012,
                           ZN => n1816);
   U2224 : AOI221_X1 port map( B1 => n309, B2 => n1167, C1 => n311, C2 => n4140
                           , A => n1819, ZN => n1818);
   U2225 : OAI22_X1 port map( A1 => n631, A2 => n314, B1 => n1820, B2 => n317, 
                           ZN => n1819);
   U2226 : AOI22_X1 port map( A1 => n320, A2 => n4172, B1 => n323, B2 => n1065,
                           ZN => n1817);
   U2227 : NAND4_X1 port map( A1 => n1824, A2 => n1821, A3 => n1822, A4 => 
                           n1823, ZN => n1809);
   U2228 : AOI221_X1 port map( B1 => n326, B2 => n4204, C1 => n329, C2 => n4236
                           , A => n1825, ZN => n1824);
   U2229 : OAI22_X1 port map( A1 => n407, A2 => n332, B1 => n375, B2 => n20, ZN
                           => n1825);
   U2230 : AOI221_X1 port map( B1 => n335, B2 => n4268, C1 => n338, C2 => n4300
                           , A => n1826, ZN => n1823);
   U2231 : OAI22_X1 port map( A1 => n279, A2 => n341, B1 => n247, B2 => n344, 
                           ZN => n1826);
   U2232 : AOI221_X1 port map( B1 => n347, B2 => n788, C1 => n350, C2 => n822, 
                           A => n1827, ZN => n1822);
   U2233 : OAI22_X1 port map( A1 => n1828, A2 => n353, B1 => n1829, B2 => n356,
                           ZN => n1827);
   U2234 : OAI22_X1 port map( A1 => n1831, A2 => n429, B1 => n1832, B2 => n22, 
                           ZN => n1830);
   U2235 : OAI222_X1 port map( A1 => n574, A2 => n208, B1 => n1833, B2 => n211,
                           C1 => n3915, C2 => n214, ZN => n2550);
   U2236 : OAI221_X1 port map( B1 => n856, B2 => n217, C1 => n1838, C2 => n220,
                           A => n1839, ZN => n1837);
   U2237 : AOI22_X1 port map( A1 => n223, A2 => n4043, B1 => n29, B2 => n1207, 
                           ZN => n1839);
   U2238 : OAI221_X1 port map( B1 => n1840, B2 => n293, C1 => n952, C2 => n296,
                           A => n1841, ZN => n1836);
   U2239 : AOI22_X1 port map( A1 => n299, A2 => n1309, B1 => n302, B2 => n4011,
                           ZN => n1841);
   U2240 : OAI211_X1 port map( C1 => n536, C2 => n305, A => n1842, B => n1843, 
                           ZN => n1835);
   U2241 : AOI221_X1 port map( B1 => n309, B2 => n1168, C1 => n311, C2 => n4139
                           , A => n1844, ZN => n1843);
   U2242 : OAI22_X1 port map( A1 => n632, A2 => n314, B1 => n1845, B2 => n317, 
                           ZN => n1844);
   U2243 : AOI22_X1 port map( A1 => n320, A2 => n4171, B1 => n323, B2 => n1066,
                           ZN => n1842);
   U2244 : NAND4_X1 port map( A1 => n1846, A2 => n1847, A3 => n1848, A4 => 
                           n1849, ZN => n1834);
   U2245 : AOI221_X1 port map( B1 => n326, B2 => n4203, C1 => n329, C2 => n4235
                           , A => n1850, ZN => n1849);
   U2246 : OAI22_X1 port map( A1 => n408, A2 => n31, B1 => n376, B2 => n21, ZN 
                           => n1850);
   U2247 : AOI221_X1 port map( B1 => n335, B2 => n4267, C1 => n338, C2 => n4299
                           , A => n1851, ZN => n1848);
   U2248 : OAI22_X1 port map( A1 => n280, A2 => n341, B1 => n248, B2 => n343, 
                           ZN => n1851);
   U2249 : AOI221_X1 port map( B1 => n347, B2 => n789, C1 => n350, C2 => n823, 
                           A => n1852, ZN => n1847);
   U2250 : OAI22_X1 port map( A1 => n1853, A2 => n353, B1 => n1854, B2 => n356,
                           ZN => n1852);
   U2251 : AOI221_X1 port map( B1 => n423, B2 => n750, C1 => n426, C2 => n3947,
                           A => n1855, ZN => n1846);
   U2252 : OAI22_X1 port map( A1 => n1856, A2 => n429, B1 => n1857, B2 => n5, 
                           ZN => n1855);
   U2253 : OAI222_X1 port map( A1 => n573, A2 => n207, B1 => n1858, B2 => n210,
                           C1 => n3914, C2 => n214, ZN => n2549);
   U2254 : NOR4_X1 port map( A1 => n1859, A2 => n1860, A3 => n1861, A4 => n1862
                           , ZN => n1858);
   U2255 : OAI221_X1 port map( B1 => n857, B2 => n216, C1 => n1863, C2 => n219,
                           A => n1864, ZN => n1862);
   U2256 : AOI22_X1 port map( A1 => n222, A2 => n4042, B1 => n225, B2 => n1208,
                           ZN => n1864);
   U2257 : OAI221_X1 port map( B1 => n1865, B2 => n228, C1 => n953, C2 => n295,
                           A => n1866, ZN => n1861);
   U2258 : AOI22_X1 port map( A1 => n298, A2 => n1310, B1 => n301, B2 => n4010,
                           ZN => n1866);
   U2259 : OAI211_X1 port map( C1 => n537, C2 => n304, A => n1867, B => n1868, 
                           ZN => n1860);
   U2260 : AOI221_X1 port map( B1 => n307, B2 => n1169, C1 => n310, C2 => n4138
                           , A => n1869, ZN => n1868);
   U2261 : OAI22_X1 port map( A1 => n633, A2 => n313, B1 => n1870, B2 => n316, 
                           ZN => n1869);
   U2262 : AOI22_X1 port map( A1 => n319, A2 => n4170, B1 => n322, B2 => n1067,
                           ZN => n1867);
   U2263 : NAND4_X1 port map( A1 => n1872, A2 => n1873, A3 => n1871, A4 => 
                           n1874, ZN => n1859);
   U2264 : AOI221_X1 port map( B1 => n325, B2 => n4202, C1 => n328, C2 => n4234
                           , A => n1875, ZN => n1874);
   U2265 : OAI22_X1 port map( A1 => n409, A2 => n331, B1 => n377, B2 => n21, ZN
                           => n1875);
   U2266 : AOI221_X1 port map( B1 => n334, B2 => n4266, C1 => n337, C2 => n4298
                           , A => n1876, ZN => n1873);
   U2267 : OAI22_X1 port map( A1 => n281, A2 => n340, B1 => n249, B2 => n344, 
                           ZN => n1876);
   U2268 : AOI221_X1 port map( B1 => n346, B2 => n790, C1 => n349, C2 => n824, 
                           A => n1877, ZN => n1872);
   U2269 : OAI22_X1 port map( A1 => n1878, A2 => n352, B1 => n1879, B2 => n355,
                           ZN => n1877);
   U2270 : AOI221_X1 port map( B1 => n424, B2 => n751, C1 => n425, C2 => n3946,
                           A => n1880, ZN => n1871);
   U2271 : OAI22_X1 port map( A1 => n1881, A2 => n429, B1 => n1882, B2 => n5, 
                           ZN => n1880);
   U2272 : OAI222_X1 port map( A1 => n572, A2 => n207, B1 => n1883, B2 => n210,
                           C1 => n3913, C2 => n214, ZN => n2548);
   U2273 : OAI221_X1 port map( B1 => n858, B2 => n216, C1 => n1888, C2 => n219,
                           A => n1889, ZN => n1887);
   U2274 : AOI22_X1 port map( A1 => n222, A2 => n4041, B1 => n225, B2 => n1209,
                           ZN => n1889);
   U2275 : OAI221_X1 port map( B1 => n1890, B2 => n228, C1 => n954, C2 => n295,
                           A => n1891, ZN => n1886);
   U2276 : AOI22_X1 port map( A1 => n298, A2 => n1311, B1 => n301, B2 => n4009,
                           ZN => n1891);
   U2277 : OAI211_X1 port map( C1 => n538, C2 => n304, A => n1892, B => n1893, 
                           ZN => n1885);
   U2278 : AOI221_X1 port map( B1 => n308, B2 => n1170, C1 => n310, C2 => n4137
                           , A => n1894, ZN => n1893);
   U2279 : OAI22_X1 port map( A1 => n634, A2 => n313, B1 => n1895, B2 => n316, 
                           ZN => n1894);
   U2280 : AOI22_X1 port map( A1 => n319, A2 => n4169, B1 => n322, B2 => n1068,
                           ZN => n1892);
   U2281 : NAND4_X1 port map( A1 => n1896, A2 => n1897, A3 => n1898, A4 => 
                           n1899, ZN => n1884);
   U2282 : AOI221_X1 port map( B1 => n325, B2 => n4201, C1 => n328, C2 => n4233
                           , A => n1900, ZN => n1899);
   U2283 : OAI22_X1 port map( A1 => n410, A2 => n32, B1 => n378, B2 => n20, ZN 
                           => n1900);
   U2284 : AOI221_X1 port map( B1 => n334, B2 => n4265, C1 => n337, C2 => n4297
                           , A => n1901, ZN => n1898);
   U2285 : OAI22_X1 port map( A1 => n282, A2 => n340, B1 => n250, B2 => n345, 
                           ZN => n1901);
   U2286 : AOI221_X1 port map( B1 => n346, B2 => n791, C1 => n349, C2 => n825, 
                           A => n1902, ZN => n1897);
   U2287 : OAI22_X1 port map( A1 => n1903, A2 => n352, B1 => n1904, B2 => n355,
                           ZN => n1902);
   U2288 : AOI221_X1 port map( B1 => n422, B2 => n752, C1 => n425, C2 => n3945,
                           A => n1905, ZN => n1896);
   U2289 : OAI22_X1 port map( A1 => n1906, A2 => n428, B1 => n1907, B2 => n5, 
                           ZN => n1905);
   U2290 : OAI222_X1 port map( A1 => n571, A2 => n207, B1 => n1908, B2 => n210,
                           C1 => n3912, C2 => n213, ZN => n2547);
   U2291 : NOR4_X1 port map( A1 => n1909, A2 => n1910, A3 => n1911, A4 => n1912
                           , ZN => n1908);
   U2292 : OAI221_X1 port map( B1 => n859, B2 => n216, C1 => n1913, C2 => n219,
                           A => n1914, ZN => n1912);
   U2293 : AOI22_X1 port map( A1 => n222, A2 => n4040, B1 => n30, B2 => n1210, 
                           ZN => n1914);
   U2294 : OAI221_X1 port map( B1 => n1915, B2 => n228, C1 => n955, C2 => n295,
                           A => n1916, ZN => n1911);
   U2295 : AOI22_X1 port map( A1 => n298, A2 => n1312, B1 => n301, B2 => n4008,
                           ZN => n1916);
   U2296 : OAI211_X1 port map( C1 => n539, C2 => n304, A => n1917, B => n1918, 
                           ZN => n1910);
   U2297 : AOI221_X1 port map( B1 => n307, B2 => n1171, C1 => n310, C2 => n4136
                           , A => n1919, ZN => n1918);
   U2298 : OAI22_X1 port map( A1 => n635, A2 => n313, B1 => n1920, B2 => n316, 
                           ZN => n1919);
   U2299 : AOI22_X1 port map( A1 => n319, A2 => n4168, B1 => n322, B2 => n1069,
                           ZN => n1917);
   U2300 : NAND4_X1 port map( A1 => n1922, A2 => n1923, A3 => n1921, A4 => 
                           n1924, ZN => n1909);
   U2301 : AOI221_X1 port map( B1 => n325, B2 => n4200, C1 => n328, C2 => n4232
                           , A => n1925, ZN => n1924);
   U2302 : OAI22_X1 port map( A1 => n411, A2 => n331, B1 => n379, B2 => n20, ZN
                           => n1925);
   U2303 : AOI221_X1 port map( B1 => n334, B2 => n4264, C1 => n337, C2 => n4296
                           , A => n1926, ZN => n1923);
   U2304 : OAI22_X1 port map( A1 => n283, A2 => n342, B1 => n251, B2 => n344, 
                           ZN => n1926);
   U2305 : AOI221_X1 port map( B1 => n346, B2 => n792, C1 => n349, C2 => n826, 
                           A => n1927, ZN => n1922);
   U2306 : OAI22_X1 port map( A1 => n1928, A2 => n352, B1 => n1929, B2 => n355,
                           ZN => n1927);
   U2307 : AOI221_X1 port map( B1 => n424, B2 => n753, C1 => n425, C2 => n3944,
                           A => n1930, ZN => n1921);
   U2308 : OAI22_X1 port map( A1 => n1931, A2 => n428, B1 => n1932, B2 => n23, 
                           ZN => n1930);
   U2309 : OAI222_X1 port map( A1 => n570, A2 => n207, B1 => n1933, B2 => n210,
                           C1 => n3911, C2 => n213, ZN => n2546);
   U2310 : OAI221_X1 port map( B1 => n860, B2 => n216, C1 => n1938, C2 => n219,
                           A => n1939, ZN => n1937);
   U2311 : AOI22_X1 port map( A1 => n222, A2 => n4039, B1 => n30, B2 => n1211, 
                           ZN => n1939);
   U2312 : OAI221_X1 port map( B1 => n1940, B2 => n228, C1 => n956, C2 => n295,
                           A => n1941, ZN => n1936);
   U2313 : AOI22_X1 port map( A1 => n298, A2 => n1313, B1 => n301, B2 => n4007,
                           ZN => n1941);
   U2314 : OAI211_X1 port map( C1 => n540, C2 => n304, A => n1942, B => n1943, 
                           ZN => n1935);
   U2315 : AOI221_X1 port map( B1 => n309, B2 => n1172, C1 => n310, C2 => n4135
                           , A => n1944, ZN => n1943);
   U2316 : OAI22_X1 port map( A1 => n636, A2 => n313, B1 => n1945, B2 => n316, 
                           ZN => n1944);
   U2317 : AOI22_X1 port map( A1 => n319, A2 => n4167, B1 => n322, B2 => n1070,
                           ZN => n1942);
   U2318 : NAND4_X1 port map( A1 => n1946, A2 => n1947, A3 => n1948, A4 => 
                           n1949, ZN => n1934);
   U2319 : AOI221_X1 port map( B1 => n325, B2 => n4199, C1 => n328, C2 => n4231
                           , A => n1950, ZN => n1949);
   U2320 : OAI22_X1 port map( A1 => n412, A2 => n333, B1 => n380, B2 => n20, ZN
                           => n1950);
   U2321 : AOI221_X1 port map( B1 => n334, B2 => n4263, C1 => n337, C2 => n4295
                           , A => n1951, ZN => n1948);
   U2322 : OAI22_X1 port map( A1 => n284, A2 => n342, B1 => n252, B2 => n343, 
                           ZN => n1951);
   U2323 : AOI221_X1 port map( B1 => n346, B2 => n793, C1 => n349, C2 => n827, 
                           A => n1952, ZN => n1947);
   U2324 : OAI22_X1 port map( A1 => n1953, A2 => n352, B1 => n1954, B2 => n355,
                           ZN => n1952);
   U2325 : AOI221_X1 port map( B1 => n423, B2 => n754, C1 => n425, C2 => n3943,
                           A => n1955, ZN => n1946);
   U2326 : OAI22_X1 port map( A1 => n1956, A2 => n428, B1 => n1957, B2 => n23, 
                           ZN => n1955);
   U2327 : OAI222_X1 port map( A1 => n569, A2 => n207, B1 => n1958, B2 => n210,
                           C1 => n3910, C2 => n213, ZN => n2545);
   U2328 : NOR4_X1 port map( A1 => n1959, A2 => n1960, A3 => n1961, A4 => n1962
                           , ZN => n1958);
   U2329 : OAI221_X1 port map( B1 => n861, B2 => n216, C1 => n1963, C2 => n219,
                           A => n1964, ZN => n1962);
   U2330 : AOI22_X1 port map( A1 => n222, A2 => n4038, B1 => n29, B2 => n1212, 
                           ZN => n1964);
   U2331 : OAI221_X1 port map( B1 => n1965, B2 => n228, C1 => n957, C2 => n295,
                           A => n1966, ZN => n1961);
   U2332 : AOI22_X1 port map( A1 => n298, A2 => n1314, B1 => n301, B2 => n4006,
                           ZN => n1966);
   U2333 : OAI211_X1 port map( C1 => n541, C2 => n304, A => n1967, B => n1968, 
                           ZN => n1960);
   U2334 : AOI221_X1 port map( B1 => n307, B2 => n1173, C1 => n310, C2 => n4134
                           , A => n1969, ZN => n1968);
   U2335 : OAI22_X1 port map( A1 => n637, A2 => n313, B1 => n1970, B2 => n316, 
                           ZN => n1969);
   U2336 : AOI22_X1 port map( A1 => n319, A2 => n4166, B1 => n322, B2 => n1071,
                           ZN => n1967);
   U2337 : NAND4_X1 port map( A1 => n1972, A2 => n1973, A3 => n1971, A4 => 
                           n1974, ZN => n1959);
   U2338 : AOI221_X1 port map( B1 => n325, B2 => n4198, C1 => n328, C2 => n4230
                           , A => n1975, ZN => n1974);
   U2339 : OAI22_X1 port map( A1 => n413, A2 => n331, B1 => n381, B2 => n21, ZN
                           => n1975);
   U2340 : AOI221_X1 port map( B1 => n334, B2 => n4262, C1 => n337, C2 => n4294
                           , A => n1976, ZN => n1973);
   U2341 : OAI22_X1 port map( A1 => n285, A2 => n33, B1 => n253, B2 => n344, ZN
                           => n1976);
   U2342 : AOI221_X1 port map( B1 => n346, B2 => n794, C1 => n349, C2 => n828, 
                           A => n1977, ZN => n1972);
   U2343 : OAI22_X1 port map( A1 => n1978, A2 => n352, B1 => n1979, B2 => n355,
                           ZN => n1977);
   U2344 : AOI221_X1 port map( B1 => n424, B2 => n755, C1 => n425, C2 => n3942,
                           A => n1980, ZN => n1971);
   U2345 : OAI22_X1 port map( A1 => n1981, A2 => n428, B1 => n1982, B2 => n5, 
                           ZN => n1980);
   U2346 : OAI222_X1 port map( A1 => n568, A2 => n207, B1 => n1983, B2 => n210,
                           C1 => n3909, C2 => n213, ZN => n2544);
   U2347 : OAI221_X1 port map( B1 => n862, B2 => n216, C1 => n1988, C2 => n219,
                           A => n1989, ZN => n1987);
   U2348 : AOI22_X1 port map( A1 => n222, A2 => n4037, B1 => n29, B2 => n1213, 
                           ZN => n1989);
   U2349 : OAI221_X1 port map( B1 => n1990, B2 => n228, C1 => n958, C2 => n295,
                           A => n1991, ZN => n1986);
   U2350 : AOI22_X1 port map( A1 => n298, A2 => n1315, B1 => n301, B2 => n4005,
                           ZN => n1991);
   U2351 : OAI211_X1 port map( C1 => n542, C2 => n304, A => n1992, B => n1993, 
                           ZN => n1985);
   U2352 : AOI221_X1 port map( B1 => n308, B2 => n1174, C1 => n310, C2 => n4133
                           , A => n1994, ZN => n1993);
   U2353 : OAI22_X1 port map( A1 => n638, A2 => n313, B1 => n1995, B2 => n316, 
                           ZN => n1994);
   U2354 : AOI22_X1 port map( A1 => n319, A2 => n4165, B1 => n322, B2 => n1072,
                           ZN => n1992);
   U2355 : NAND4_X1 port map( A1 => n1996, A2 => n1997, A3 => n1998, A4 => 
                           n1999, ZN => n1984);
   U2356 : AOI221_X1 port map( B1 => n325, B2 => n4197, C1 => n328, C2 => n4229
                           , A => n2000, ZN => n1999);
   U2357 : OAI22_X1 port map( A1 => n414, A2 => n31, B1 => n382, B2 => n20, ZN 
                           => n2000);
   U2358 : AOI221_X1 port map( B1 => n334, B2 => n4261, C1 => n337, C2 => n4293
                           , A => n2001, ZN => n1998);
   U2359 : OAI22_X1 port map( A1 => n286, A2 => n33, B1 => n254, B2 => n345, ZN
                           => n2001);
   U2360 : AOI221_X1 port map( B1 => n346, B2 => n795, C1 => n349, C2 => n829, 
                           A => n2002, ZN => n1997);
   U2361 : OAI22_X1 port map( A1 => n2003, A2 => n352, B1 => n2004, B2 => n355,
                           ZN => n2002);
   U2362 : AOI221_X1 port map( B1 => n422, B2 => n756, C1 => n425, C2 => n3941,
                           A => n2005, ZN => n1996);
   U2363 : OAI22_X1 port map( A1 => n2006, A2 => n428, B1 => n2007, B2 => n23, 
                           ZN => n2005);
   U2364 : OAI222_X1 port map( A1 => n567, A2 => n207, B1 => n2008, B2 => n210,
                           C1 => n3908, C2 => n213, ZN => n2543);
   U2365 : NOR4_X1 port map( A1 => n2009, A2 => n2010, A3 => n2011, A4 => n2012
                           , ZN => n2008);
   U2366 : OAI221_X1 port map( B1 => n863, B2 => n216, C1 => n2013, C2 => n219,
                           A => n2014, ZN => n2012);
   U2367 : AOI22_X1 port map( A1 => n222, A2 => n4036, B1 => n227, B2 => n1214,
                           ZN => n2014);
   U2368 : OAI221_X1 port map( B1 => n2015, B2 => n228, C1 => n959, C2 => n295,
                           A => n2016, ZN => n2011);
   U2369 : AOI22_X1 port map( A1 => n298, A2 => n1316, B1 => n301, B2 => n4004,
                           ZN => n2016);
   U2370 : OAI211_X1 port map( C1 => n543, C2 => n304, A => n2017, B => n2018, 
                           ZN => n2010);
   U2371 : AOI221_X1 port map( B1 => n307, B2 => n1175, C1 => n310, C2 => n4132
                           , A => n2019, ZN => n2018);
   U2372 : OAI22_X1 port map( A1 => n639, A2 => n313, B1 => n2020, B2 => n316, 
                           ZN => n2019);
   U2373 : AOI22_X1 port map( A1 => n319, A2 => n4164, B1 => n322, B2 => n1073,
                           ZN => n2017);
   U2374 : NAND4_X1 port map( A1 => n2022, A2 => n2023, A3 => n2021, A4 => 
                           n2024, ZN => n2009);
   U2375 : AOI221_X1 port map( B1 => n325, B2 => n4196, C1 => n328, C2 => n4228
                           , A => n2025, ZN => n2024);
   U2376 : OAI22_X1 port map( A1 => n415, A2 => n331, B1 => n383, B2 => n20, ZN
                           => n2025);
   U2377 : AOI221_X1 port map( B1 => n334, B2 => n4260, C1 => n337, C2 => n4292
                           , A => n2026, ZN => n2023);
   U2378 : OAI22_X1 port map( A1 => n287, A2 => n34, B1 => n255, B2 => n344, ZN
                           => n2026);
   U2379 : AOI221_X1 port map( B1 => n346, B2 => n796, C1 => n349, C2 => n830, 
                           A => n2027, ZN => n2022);
   U2380 : OAI22_X1 port map( A1 => n2028, A2 => n352, B1 => n2029, B2 => n355,
                           ZN => n2027);
   U2381 : AOI221_X1 port map( B1 => n424, B2 => n757, C1 => n425, C2 => n3940,
                           A => n2030, ZN => n2021);
   U2382 : OAI22_X1 port map( A1 => n2031, A2 => n428, B1 => n2032, B2 => n22, 
                           ZN => n2030);
   U2383 : OAI222_X1 port map( A1 => n566, A2 => n207, B1 => n2033, B2 => n210,
                           C1 => n3907, C2 => n213, ZN => n2542);
   U2384 : OAI221_X1 port map( B1 => n864, B2 => n216, C1 => n2038, C2 => n219,
                           A => n2039, ZN => n2037);
   U2385 : AOI22_X1 port map( A1 => n222, A2 => n4035, B1 => n227, B2 => n1215,
                           ZN => n2039);
   U2386 : OAI221_X1 port map( B1 => n2040, B2 => n228, C1 => n960, C2 => n295,
                           A => n2041, ZN => n2036);
   U2387 : AOI22_X1 port map( A1 => n298, A2 => n1317, B1 => n301, B2 => n4003,
                           ZN => n2041);
   U2388 : OAI211_X1 port map( C1 => n544, C2 => n304, A => n2042, B => n2043, 
                           ZN => n2035);
   U2389 : AOI221_X1 port map( B1 => n309, B2 => n1176, C1 => n310, C2 => n4131
                           , A => n2044, ZN => n2043);
   U2390 : OAI22_X1 port map( A1 => n640, A2 => n313, B1 => n2045, B2 => n316, 
                           ZN => n2044);
   U2391 : AOI22_X1 port map( A1 => n319, A2 => n4163, B1 => n322, B2 => n1074,
                           ZN => n2042);
   U2392 : NAND4_X1 port map( A1 => n2046, A2 => n2047, A3 => n2048, A4 => 
                           n2049, ZN => n2034);
   U2393 : AOI221_X1 port map( B1 => n325, B2 => n4195, C1 => n328, C2 => n4227
                           , A => n2050, ZN => n2049);
   U2394 : OAI22_X1 port map( A1 => n416, A2 => n332, B1 => n384, B2 => n21, ZN
                           => n2050);
   U2395 : AOI221_X1 port map( B1 => n334, B2 => n4259, C1 => n337, C2 => n4291
                           , A => n2051, ZN => n2048);
   U2396 : OAI22_X1 port map( A1 => n288, A2 => n34, B1 => n256, B2 => n343, ZN
                           => n2051);
   U2397 : AOI221_X1 port map( B1 => n346, B2 => n797, C1 => n349, C2 => n831, 
                           A => n2052, ZN => n2047);
   U2398 : OAI22_X1 port map( A1 => n2053, A2 => n352, B1 => n2054, B2 => n355,
                           ZN => n2052);
   U2399 : AOI221_X1 port map( B1 => n423, B2 => n758, C1 => n425, C2 => n3939,
                           A => n2055, ZN => n2046);
   U2400 : OAI22_X1 port map( A1 => n2056, A2 => n428, B1 => n2057, B2 => n5, 
                           ZN => n2055);
   U2401 : OAI222_X1 port map( A1 => n565, A2 => n207, B1 => n2058, B2 => n210,
                           C1 => n3906, C2 => n213, ZN => n2541);
   U2402 : OAI221_X1 port map( B1 => n865, B2 => n216, C1 => n2063, C2 => n219,
                           A => n2064, ZN => n2062);
   U2403 : AOI22_X1 port map( A1 => n222, A2 => n4034, B1 => n226, B2 => n1216,
                           ZN => n2064);
   U2404 : OAI221_X1 port map( B1 => n2065, B2 => n228, C1 => n961, C2 => n295,
                           A => n2066, ZN => n2061);
   U2405 : AOI22_X1 port map( A1 => n298, A2 => n1318, B1 => n301, B2 => n4002,
                           ZN => n2066);
   U2406 : OAI211_X1 port map( C1 => n545, C2 => n304, A => n2067, B => n2068, 
                           ZN => n2060);
   U2407 : AOI221_X1 port map( B1 => n308, B2 => n1177, C1 => n310, C2 => n4130
                           , A => n2069, ZN => n2068);
   U2408 : OAI22_X1 port map( A1 => n641, A2 => n313, B1 => n2070, B2 => n316, 
                           ZN => n2069);
   U2409 : AOI22_X1 port map( A1 => n319, A2 => n4162, B1 => n322, B2 => n1075,
                           ZN => n2067);
   U2410 : NAND4_X1 port map( A1 => n2071, A2 => n2074, A3 => n2072, A4 => 
                           n2073, ZN => n2059);
   U2411 : OAI22_X1 port map( A1 => n417, A2 => n333, B1 => n385, B2 => n21, ZN
                           => n2075);
   U2412 : AOI221_X1 port map( B1 => n334, B2 => n4258, C1 => n337, C2 => n4290
                           , A => n2076, ZN => n2073);
   U2413 : OAI22_X1 port map( A1 => n289, A2 => n341, B1 => n257, B2 => n344, 
                           ZN => n2076);
   U2414 : AOI221_X1 port map( B1 => n346, B2 => n798, C1 => n349, C2 => n832, 
                           A => n2077, ZN => n2072);
   U2415 : OAI22_X1 port map( A1 => n2078, A2 => n352, B1 => n2079, B2 => n355,
                           ZN => n2077);
   U2416 : AOI221_X1 port map( B1 => n422, B2 => n759, C1 => n425, C2 => n3938,
                           A => n2080, ZN => n2071);
   U2417 : OAI22_X1 port map( A1 => n2081, A2 => n428, B1 => n2082, B2 => n5, 
                           ZN => n2080);
   U2418 : OAI222_X1 port map( A1 => n564, A2 => n207, B1 => n2083, B2 => n210,
                           C1 => n3905, C2 => n213, ZN => n2540);
   U2419 : OAI221_X1 port map( B1 => n866, B2 => n216, C1 => n2088, C2 => n219,
                           A => n2089, ZN => n2087);
   U2420 : AOI22_X1 port map( A1 => n222, A2 => n4033, B1 => n227, B2 => n1217,
                           ZN => n2089);
   U2421 : OAI221_X1 port map( B1 => n2090, B2 => n228, C1 => n962, C2 => n295,
                           A => n2091, ZN => n2086);
   U2422 : AOI22_X1 port map( A1 => n298, A2 => n1319, B1 => n301, B2 => n4001,
                           ZN => n2091);
   U2423 : OAI211_X1 port map( C1 => n546, C2 => n304, A => n2092, B => n2093, 
                           ZN => n2085);
   U2424 : AOI221_X1 port map( B1 => n308, B2 => n1178, C1 => n310, C2 => n4129
                           , A => n2094, ZN => n2093);
   U2425 : OAI22_X1 port map( A1 => n642, A2 => n313, B1 => n2095, B2 => n316, 
                           ZN => n2094);
   U2426 : AOI22_X1 port map( A1 => n319, A2 => n4161, B1 => n322, B2 => n1076,
                           ZN => n2092);
   U2427 : NAND4_X1 port map( A1 => n2096, A2 => n2097, A3 => n2098, A4 => 
                           n2099, ZN => n2084);
   U2428 : AOI221_X1 port map( B1 => n325, B2 => n4193, C1 => n328, C2 => n4225
                           , A => n2100, ZN => n2099);
   U2429 : OAI22_X1 port map( A1 => n418, A2 => n31, B1 => n386, B2 => n21, ZN 
                           => n2100);
   U2430 : AOI221_X1 port map( B1 => n334, B2 => n4257, C1 => n337, C2 => n4289
                           , A => n2101, ZN => n2098);
   U2431 : OAI22_X1 port map( A1 => n290, A2 => n341, B1 => n258, B2 => n343, 
                           ZN => n2101);
   U2432 : OAI22_X1 port map( A1 => n2103, A2 => n352, B1 => n2104, B2 => n355,
                           ZN => n2102);
   U2433 : AOI221_X1 port map( B1 => n423, B2 => n760, C1 => n425, C2 => n3937,
                           A => n2105, ZN => n2096);
   U2434 : OAI22_X1 port map( A1 => n2106, A2 => n428, B1 => n2107, B2 => n23, 
                           ZN => n2105);
   U2435 : OAI222_X1 port map( A1 => n563, A2 => n207, B1 => n2108, B2 => n210,
                           C1 => n3904, C2 => n213, ZN => n2539);
   U2436 : OAI221_X1 port map( B1 => n867, B2 => n216, C1 => n2113, C2 => n219,
                           A => n2114, ZN => n2112);
   U2437 : AOI22_X1 port map( A1 => n222, A2 => n4032, B1 => n226, B2 => n1218,
                           ZN => n2114);
   U2438 : OAI221_X1 port map( B1 => n2115, B2 => n228, C1 => n963, C2 => n295,
                           A => n2116, ZN => n2111);
   U2439 : AOI22_X1 port map( A1 => n298, A2 => n1320, B1 => n301, B2 => n4000,
                           ZN => n2116);
   U2440 : AOI221_X1 port map( B1 => n308, B2 => n1179, C1 => n310, C2 => n4128
                           , A => n2119, ZN => n2118);
   U2441 : OAI22_X1 port map( A1 => n643, A2 => n313, B1 => n2120, B2 => n316, 
                           ZN => n2119);
   U2442 : AOI22_X1 port map( A1 => n319, A2 => n4160, B1 => n322, B2 => n1077,
                           ZN => n2117);
   U2443 : NAND4_X1 port map( A1 => n2121, A2 => n2122, A3 => n2124, A4 => 
                           n2123, ZN => n2109);
   U2444 : AOI221_X1 port map( B1 => n325, B2 => n4192, C1 => n328, C2 => n4224
                           , A => n2125, ZN => n2124);
   U2445 : OAI22_X1 port map( A1 => n419, A2 => n332, B1 => n387, B2 => n21, ZN
                           => n2125);
   U2446 : AOI221_X1 port map( B1 => n334, B2 => n4256, C1 => n337, C2 => n4288
                           , A => n2126, ZN => n2123);
   U2447 : OAI22_X1 port map( A1 => n291, A2 => n340, B1 => n259, B2 => n343, 
                           ZN => n2126);
   U2448 : OAI22_X1 port map( A1 => n2128, A2 => n352, B1 => n2129, B2 => n355,
                           ZN => n2127);
   U2449 : AOI221_X1 port map( B1 => n422, B2 => n761, C1 => n425, C2 => n3936,
                           A => n2130, ZN => n2121);
   U2450 : OAI22_X1 port map( A1 => n2131, A2 => n428, B1 => n2132, B2 => n22, 
                           ZN => n2130);
   U2451 : OAI222_X1 port map( A1 => n562, A2 => n207, B1 => n2133, B2 => n210,
                           C1 => n3903, C2 => n213, ZN => n2538);
   U2452 : NAND2_X1 port map( A1 => n213, A2 => n2134, ZN => n1326);
   U2453 : OAI221_X1 port map( B1 => n868, B2 => n216, C1 => n2139, C2 => n219,
                           A => n2140, ZN => n2138);
   U2454 : AOI22_X1 port map( A1 => n222, A2 => n4031, B1 => n226, B2 => n1219,
                           ZN => n2140);
   U2455 : AND2_X1 port map( A1 => n2141, A2 => n2142, ZN => n1337);
   U2456 : AND2_X1 port map( A1 => n2141, A2 => n2143, ZN => n1336);
   U2457 : NAND2_X1 port map( A1 => n2144, A2 => n2145, ZN => n1334);
   U2458 : NAND2_X1 port map( A1 => n2146, A2 => n2142, ZN => n1332);
   U2459 : OAI221_X1 port map( B1 => n2147, B2 => n228, C1 => n964, C2 => n295,
                           A => n2148, ZN => n2137);
   U2460 : AOI22_X1 port map( A1 => n298, A2 => n1321, B1 => n301, B2 => n3999,
                           ZN => n2148);
   U2461 : AND2_X1 port map( A1 => n2146, A2 => n2143, ZN => n1343);
   U2462 : AND2_X1 port map( A1 => n2146, A2 => n2145, ZN => n1342);
   U2463 : NAND2_X1 port map( A1 => n54, A2 => n2145, ZN => n1340);
   U2464 : NAND2_X1 port map( A1 => n54, A2 => n85, ZN => n1339);
   U2465 : NOR3_X1 port map( A1 => n2151, A2 => ADD_RS2(0), A3 => n2150, ZN => 
                           n2141);
   U2466 : OAI211_X1 port map( C1 => n548, C2 => n304, A => n2152, B => n2153, 
                           ZN => n2136);
   U2467 : AOI221_X1 port map( B1 => n309, B2 => n1180, C1 => n310, C2 => n4127
                           , A => n2154, ZN => n2153);
   U2468 : OAI22_X1 port map( A1 => n644, A2 => n313, B1 => n2155, B2 => n316, 
                           ZN => n2154);
   U2469 : NAND2_X1 port map( A1 => n2156, A2 => n2145, ZN => n1352);
   U2470 : NAND2_X1 port map( A1 => n2149, A2 => n2156, ZN => n1350);
   U2471 : AND2_X1 port map( A1 => n2144, A2 => n2142, ZN => n1348);
   U2472 : AND2_X1 port map( A1 => n2149, A2 => n2144, ZN => n1347);
   U2473 : AOI22_X1 port map( A1 => n319, A2 => n4159, B1 => n322, B2 => n1078,
                           ZN => n2152);
   U2474 : AND2_X1 port map( A1 => n26, A2 => n18, ZN => n1354);
   U2475 : AND2_X1 port map( A1 => n26, A2 => n2142, ZN => n1353);
   U2476 : NOR3_X1 port map( A1 => ADD_RS2(0), A2 => n86, A3 => ADD_RS2(3), ZN 
                           => n2156);
   U2477 : NAND2_X1 port map( A1 => n2144, A2 => n18, ZN => n1344);
   U2478 : NOR3_X1 port map( A1 => n80, A2 => n2150, A3 => n77, ZN => n2144);
   U2479 : NAND4_X1 port map( A1 => n2157, A2 => n2158, A3 => n2160, A4 => 
                           n2159, ZN => n2135);
   U2480 : AOI221_X1 port map( B1 => n325, B2 => n4191, C1 => n328, C2 => n4223
                           , A => n2161, ZN => n2160);
   U2481 : OAI22_X1 port map( A1 => n420, A2 => n333, B1 => n388, B2 => n20, ZN
                           => n2161);
   U2482 : NAND2_X1 port map( A1 => n2162, A2 => n2149, ZN => n1363);
   U2483 : NAND2_X1 port map( A1 => n2163, A2 => n2149, ZN => n1362);
   U2484 : AND2_X1 port map( A1 => n19, A2 => n2145, ZN => n1360);
   U2485 : AND2_X1 port map( A1 => n2145, A2 => n35, ZN => n1359);
   U2486 : AOI221_X1 port map( B1 => n334, B2 => n4255, C1 => n337, C2 => n4287
                           , A => n2164, ZN => n2159);
   U2487 : OAI22_X1 port map( A1 => n292, A2 => n340, B1 => n260, B2 => n345, 
                           ZN => n2164);
   U2488 : NAND2_X1 port map( A1 => n2162, A2 => n2143, ZN => n1368);
   U2489 : NAND2_X1 port map( A1 => n2163, A2 => n2143, ZN => n1367);
   U2490 : AND2_X1 port map( A1 => n2142, A2 => n19, ZN => n1365);
   U2491 : NOR3_X1 port map( A1 => n2151, A2 => ADD_RS2(4), A3 => ADD_RS2(0), 
                           ZN => n2162);
   U2492 : AND2_X1 port map( A1 => n2142, A2 => n35, ZN => n1364);
   U2493 : NOR3_X1 port map( A1 => n77, A2 => ADD_RS2(4), A3 => n2151, ZN => 
                           n2163);
   U2494 : OAI22_X1 port map( A1 => n2166, A2 => n352, B1 => n2167, B2 => n355,
                           ZN => n2165);
   U2495 : NAND2_X1 port map( A1 => n2168, A2 => n2145, ZN => n1375);
   U2496 : NAND2_X1 port map( A1 => n2169, A2 => n2145, ZN => n1373);
   U2497 : AND2_X1 port map( A1 => n79, A2 => n78, ZN => n1370);
   U2498 : AND2_X1 port map( A1 => n2169, A2 => n78, ZN => n1369);
   U2499 : AOI221_X1 port map( B1 => n422, B2 => n762, C1 => n425, C2 => n3935,
                           A => n2170, ZN => n2157);
   U2500 : OAI22_X1 port map( A1 => n2171, A2 => n428, B1 => n2172, B2 => n22, 
                           ZN => n2170);
   U2501 : NAND2_X1 port map( A1 => n2168, A2 => n2142, ZN => n1382);
   U2502 : NAND2_X1 port map( A1 => n2169, A2 => n2142, ZN => n1380);
   U2503 : NOR3_X1 port map( A1 => ADD_RS2(0), A2 => ADD_RS2(4), A3 => 
                           ADD_RS2(3), ZN => n2169);
   U2504 : AND2_X1 port map( A1 => n2146, A2 => n85, ZN => n1377);
   U2505 : NOR2_X1 port map( A1 => n2173, A2 => ADD_RS2(1), ZN => n2149);
   U2506 : INV_X1 port map( A => ADD_RS2(2), ZN => n2173);
   U2507 : NOR3_X1 port map( A1 => n2150, A2 => n2151, A3 => n77, ZN => n2146);
   U2508 : INV_X1 port map( A => ADD_RS2(3), ZN => n2151);
   U2509 : INV_X1 port map( A => ADD_RS2(4), ZN => n2150);
   U2510 : AND2_X1 port map( A1 => n79, A2 => n2143, ZN => n1376);
   U2511 : NOR2_X1 port map( A1 => ADD_RS2(1), A2 => ADD_RS2(2), ZN => n2143);
   U2512 : NAND2_X1 port map( A1 => n2174, A2 => n213, ZN => n1324);
   U2513 : AND3_X1 port map( A1 => RD2, A2 => ENABLE, A3 => n715, ZN => n1327);
   U2514 : INV_X1 port map( A => n2134, ZN => n2174);
   U2515 : NAND4_X1 port map( A1 => n2175, A2 => n2176, A3 => n2177, A4 => 
                           n2178, ZN => n2134);
   U2516 : NOR3_X1 port map( A1 => n2179, A2 => n1323, A3 => n2180, ZN => n2178
                           );
   U2517 : XNOR2_X1 port map( A => n1220, B => n4, ZN => n2180);
   U2518 : XNOR2_X1 port map( A => n1186, B => n1, ZN => n2179);
   U2519 : XNOR2_X1 port map( A => ADD_WR(3), B => n80, ZN => n2177);
   U2520 : XNOR2_X1 port map( A => ADD_WR(4), B => ADD_RS2(4), ZN => n2176);
   U2521 : XNOR2_X1 port map( A => ADD_RS2(2), B => ADD_WR(2), ZN => n2175);
   U2522 : OAI222_X1 port map( A1 => n593, A2 => n433, B1 => n2182, B2 => n436,
                           C1 => n3902, C2 => n439, ZN => n2537);
   U2523 : NOR4_X1 port map( A1 => n2185, A2 => n2186, A3 => n2187, A4 => n2188
                           , ZN => n2182);
   U2524 : OAI221_X1 port map( B1 => n837, B2 => n442, C1 => n1333, C2 => n445,
                           A => n2191, ZN => n2188);
   U2525 : AOI22_X1 port map( A1 => n448, A2 => n4062, B1 => n451, B2 => n1187,
                           ZN => n2191);
   U2526 : OAI221_X1 port map( B1 => n1338, B2 => n454, C1 => n933, C2 => n457,
                           A => n2196, ZN => n2187);
   U2527 : AOI22_X1 port map( A1 => n460, A2 => n1289, B1 => n463, B2 => n4030,
                           ZN => n2196);
   U2528 : OAI211_X1 port map( C1 => n517, C2 => n466, A => n2200, B => n2201, 
                           ZN => n2186);
   U2529 : AOI221_X1 port map( B1 => n469, B2 => n1148, C1 => n472, C2 => n4158
                           , A => n2204, ZN => n2201);
   U2530 : OAI22_X1 port map( A1 => n613, A2 => n475, B1 => n1351, B2 => n476, 
                           ZN => n2204);
   U2531 : AOI22_X1 port map( A1 => n481, A2 => n4190, B1 => n484, B2 => n1046,
                           ZN => n2200);
   U2532 : NAND4_X1 port map( A1 => n2209, A2 => n2210, A3 => n2211, A4 => 
                           n2212, ZN => n2185);
   U2533 : AOI221_X1 port map( B1 => n487, B2 => n4222, C1 => n490, C2 => n4254
                           , A => n2215, ZN => n2212);
   U2534 : OAI22_X1 port map( A1 => n389, A2 => n493, B1 => n357, B2 => n496, 
                           ZN => n2215);
   U2535 : AOI221_X1 port map( B1 => n499, B2 => n4286, C1 => n502, C2 => n4318
                           , A => n2220, ZN => n2211);
   U2536 : OAI22_X1 port map( A1 => n261, A2 => n505, B1 => n229, B2 => n24, ZN
                           => n2220);
   U2537 : AOI221_X1 port map( B1 => n508, B2 => n769, C1 => n511, C2 => n803, 
                           A => n2225, ZN => n2210);
   U2538 : OAI22_X1 port map( A1 => n1372, A2 => n514, B1 => n1374, B2 => n549,
                           ZN => n2225);
   U2539 : AOI221_X1 port map( B1 => n552, B2 => n730, C1 => n555, C2 => n3966,
                           A => n2230, ZN => n2209);
   U2540 : OAI22_X1 port map( A1 => n1379, A2 => n558, B1 => n1381, B2 => n561,
                           ZN => n2230);
   U2541 : OAI222_X1 port map( A1 => n592, A2 => n433, B1 => n2233, B2 => n436,
                           C1 => n3901, C2 => n439, ZN => n2536);
   U2542 : NOR4_X1 port map( A1 => n2234, A2 => n2235, A3 => n2236, A4 => n2237
                           , ZN => n2233);
   U2543 : OAI221_X1 port map( B1 => n838, B2 => n442, C1 => n1388, C2 => n445,
                           A => n2238, ZN => n2237);
   U2544 : AOI22_X1 port map( A1 => n448, A2 => n4061, B1 => n451, B2 => n1189,
                           ZN => n2238);
   U2545 : OAI221_X1 port map( B1 => n1390, B2 => n454, C1 => n934, C2 => n457,
                           A => n2239, ZN => n2236);
   U2546 : AOI22_X1 port map( A1 => n460, A2 => n1291, B1 => n463, B2 => n4029,
                           ZN => n2239);
   U2547 : OAI211_X1 port map( C1 => n518, C2 => n466, A => n2240, B => n2241, 
                           ZN => n2235);
   U2548 : AOI221_X1 port map( B1 => n469, B2 => n1150, C1 => n472, C2 => n4157
                           , A => n2242, ZN => n2241);
   U2549 : OAI22_X1 port map( A1 => n614, A2 => n473, B1 => n1395, B2 => n477, 
                           ZN => n2242);
   U2550 : AOI22_X1 port map( A1 => n481, A2 => n4189, B1 => n484, B2 => n1048,
                           ZN => n2240);
   U2551 : NAND4_X1 port map( A1 => n2243, A2 => n2244, A3 => n2245, A4 => 
                           n2246, ZN => n2234);
   U2552 : AOI221_X1 port map( B1 => n487, B2 => n4221, C1 => n490, C2 => n4253
                           , A => n2247, ZN => n2246);
   U2553 : OAI22_X1 port map( A1 => n390, A2 => n493, B1 => n358, B2 => n496, 
                           ZN => n2247);
   U2554 : AOI221_X1 port map( B1 => n499, B2 => n4285, C1 => n502, C2 => n4317
                           , A => n2248, ZN => n2245);
   U2555 : OAI22_X1 port map( A1 => n262, A2 => n505, B1 => n230, B2 => n25, ZN
                           => n2248);
   U2556 : AOI221_X1 port map( B1 => n508, B2 => n771, C1 => n511, C2 => n805, 
                           A => n2249, ZN => n2244);
   U2557 : OAI22_X1 port map( A1 => n1403, A2 => n514, B1 => n1404, B2 => n549,
                           ZN => n2249);
   U2558 : AOI221_X1 port map( B1 => n552, B2 => n732, C1 => n555, C2 => n3965,
                           A => n2250, ZN => n2243);
   U2559 : OAI22_X1 port map( A1 => n1406, A2 => n558, B1 => n1407, B2 => n561,
                           ZN => n2250);
   U2560 : OAI222_X1 port map( A1 => n591, A2 => n433, B1 => n2251, B2 => n436,
                           C1 => n3900, C2 => n439, ZN => n2535);
   U2561 : NOR4_X1 port map( A1 => n2252, A2 => n2253, A3 => n2254, A4 => n2255
                           , ZN => n2251);
   U2562 : OAI221_X1 port map( B1 => n839, B2 => n442, C1 => n1413, C2 => n445,
                           A => n2256, ZN => n2255);
   U2563 : AOI22_X1 port map( A1 => n448, A2 => n4060, B1 => n451, B2 => n1190,
                           ZN => n2256);
   U2564 : OAI221_X1 port map( B1 => n1415, B2 => n454, C1 => n935, C2 => n457,
                           A => n2257, ZN => n2254);
   U2565 : AOI22_X1 port map( A1 => n460, A2 => n1292, B1 => n463, B2 => n4028,
                           ZN => n2257);
   U2566 : OAI211_X1 port map( C1 => n519, C2 => n466, A => n2258, B => n2259, 
                           ZN => n2253);
   U2567 : AOI221_X1 port map( B1 => n469, B2 => n1151, C1 => n472, C2 => n4156
                           , A => n2260, ZN => n2259);
   U2568 : OAI22_X1 port map( A1 => n615, A2 => n28, B1 => n1420, B2 => n478, 
                           ZN => n2260);
   U2569 : AOI22_X1 port map( A1 => n481, A2 => n4188, B1 => n484, B2 => n1049,
                           ZN => n2258);
   U2570 : NAND4_X1 port map( A1 => n2261, A2 => n2262, A3 => n2263, A4 => 
                           n2264, ZN => n2252);
   U2571 : AOI221_X1 port map( B1 => n487, B2 => n4220, C1 => n490, C2 => n4252
                           , A => n2265, ZN => n2264);
   U2572 : OAI22_X1 port map( A1 => n391, A2 => n493, B1 => n359, B2 => n496, 
                           ZN => n2265);
   U2573 : AOI221_X1 port map( B1 => n499, B2 => n4284, C1 => n502, C2 => n4316
                           , A => n2266, ZN => n2263);
   U2574 : OAI22_X1 port map( A1 => n263, A2 => n505, B1 => n231, B2 => n24, ZN
                           => n2266);
   U2575 : AOI221_X1 port map( B1 => n508, B2 => n772, C1 => n511, C2 => n806, 
                           A => n2267, ZN => n2262);
   U2576 : OAI22_X1 port map( A1 => n1428, A2 => n514, B1 => n1429, B2 => n549,
                           ZN => n2267);
   U2577 : AOI221_X1 port map( B1 => n552, B2 => n733, C1 => n555, C2 => n3964,
                           A => n2268, ZN => n2261);
   U2578 : OAI22_X1 port map( A1 => n1431, A2 => n558, B1 => n1432, B2 => n561,
                           ZN => n2268);
   U2579 : OAI222_X1 port map( A1 => n590, A2 => n433, B1 => n2269, B2 => n436,
                           C1 => n3899, C2 => n439, ZN => n2534);
   U2580 : NOR4_X1 port map( A1 => n2270, A2 => n2271, A3 => n2272, A4 => n2273
                           , ZN => n2269);
   U2581 : OAI221_X1 port map( B1 => n840, B2 => n442, C1 => n1438, C2 => n445,
                           A => n2274, ZN => n2273);
   U2582 : AOI22_X1 port map( A1 => n448, A2 => n4059, B1 => n451, B2 => n1191,
                           ZN => n2274);
   U2583 : OAI221_X1 port map( B1 => n1440, B2 => n454, C1 => n936, C2 => n457,
                           A => n2275, ZN => n2272);
   U2584 : AOI22_X1 port map( A1 => n460, A2 => n1293, B1 => n463, B2 => n4027,
                           ZN => n2275);
   U2585 : OAI211_X1 port map( C1 => n520, C2 => n466, A => n2276, B => n2277, 
                           ZN => n2271);
   U2586 : AOI221_X1 port map( B1 => n469, B2 => n1152, C1 => n472, C2 => n4155
                           , A => n2278, ZN => n2277);
   U2587 : OAI22_X1 port map( A1 => n616, A2 => n27, B1 => n1445, B2 => n476, 
                           ZN => n2278);
   U2588 : AOI22_X1 port map( A1 => n481, A2 => n4187, B1 => n484, B2 => n1050,
                           ZN => n2276);
   U2589 : NAND4_X1 port map( A1 => n2279, A2 => n2280, A3 => n2281, A4 => 
                           n2282, ZN => n2270);
   U2590 : AOI221_X1 port map( B1 => n487, B2 => n4219, C1 => n490, C2 => n4251
                           , A => n2283, ZN => n2282);
   U2591 : OAI22_X1 port map( A1 => n392, A2 => n493, B1 => n360, B2 => n496, 
                           ZN => n2283);
   U2592 : AOI221_X1 port map( B1 => n499, B2 => n4283, C1 => n502, C2 => n4315
                           , A => n2284, ZN => n2281);
   U2593 : OAI22_X1 port map( A1 => n264, A2 => n505, B1 => n232, B2 => n25, ZN
                           => n2284);
   U2594 : AOI221_X1 port map( B1 => n508, B2 => n773, C1 => n511, C2 => n807, 
                           A => n2285, ZN => n2280);
   U2595 : OAI22_X1 port map( A1 => n1453, A2 => n514, B1 => n1454, B2 => n549,
                           ZN => n2285);
   U2596 : AOI221_X1 port map( B1 => n552, B2 => n734, C1 => n555, C2 => n3963,
                           A => n2286, ZN => n2279);
   U2597 : OAI22_X1 port map( A1 => n1456, A2 => n558, B1 => n1457, B2 => n561,
                           ZN => n2286);
   U2598 : OAI222_X1 port map( A1 => n589, A2 => n433, B1 => n2287, B2 => n436,
                           C1 => n3898, C2 => n439, ZN => n2533);
   U2599 : NOR4_X1 port map( A1 => n2288, A2 => n2289, A3 => n2290, A4 => n2291
                           , ZN => n2287);
   U2600 : OAI221_X1 port map( B1 => n841, B2 => n442, C1 => n1463, C2 => n445,
                           A => n2292, ZN => n2291);
   U2601 : AOI22_X1 port map( A1 => n448, A2 => n4058, B1 => n451, B2 => n1192,
                           ZN => n2292);
   U2602 : OAI221_X1 port map( B1 => n1465, B2 => n454, C1 => n937, C2 => n457,
                           A => n2293, ZN => n2290);
   U2603 : AOI22_X1 port map( A1 => n460, A2 => n1294, B1 => n463, B2 => n4026,
                           ZN => n2293);
   U2604 : OAI211_X1 port map( C1 => n521, C2 => n466, A => n2294, B => n2295, 
                           ZN => n2289);
   U2605 : AOI221_X1 port map( B1 => n469, B2 => n1153, C1 => n472, C2 => n4154
                           , A => n2296, ZN => n2295);
   U2606 : OAI22_X1 port map( A1 => n617, A2 => n475, B1 => n1470, B2 => n478, 
                           ZN => n2296);
   U2607 : AOI22_X1 port map( A1 => n481, A2 => n4186, B1 => n484, B2 => n1051,
                           ZN => n2294);
   U2608 : NAND4_X1 port map( A1 => n2297, A2 => n2298, A3 => n2299, A4 => 
                           n2300, ZN => n2288);
   U2609 : AOI221_X1 port map( B1 => n487, B2 => n4218, C1 => n490, C2 => n4250
                           , A => n2301, ZN => n2300);
   U2610 : OAI22_X1 port map( A1 => n393, A2 => n493, B1 => n361, B2 => n496, 
                           ZN => n2301);
   U2611 : AOI221_X1 port map( B1 => n499, B2 => n4282, C1 => n502, C2 => n4314
                           , A => n2302, ZN => n2299);
   U2612 : OAI22_X1 port map( A1 => n265, A2 => n505, B1 => n233, B2 => n24, ZN
                           => n2302);
   U2613 : AOI221_X1 port map( B1 => n508, B2 => n774, C1 => n511, C2 => n808, 
                           A => n2303, ZN => n2298);
   U2614 : OAI22_X1 port map( A1 => n1478, A2 => n514, B1 => n1479, B2 => n549,
                           ZN => n2303);
   U2615 : AOI221_X1 port map( B1 => n552, B2 => n735, C1 => n555, C2 => n3962,
                           A => n2304, ZN => n2297);
   U2616 : OAI22_X1 port map( A1 => n1481, A2 => n558, B1 => n1482, B2 => n561,
                           ZN => n2304);
   U2617 : OAI222_X1 port map( A1 => n588, A2 => n433, B1 => n2305, B2 => n436,
                           C1 => n3897, C2 => n439, ZN => n2532);
   U2618 : NOR4_X1 port map( A1 => n2306, A2 => n2307, A3 => n2308, A4 => n2309
                           , ZN => n2305);
   U2619 : OAI221_X1 port map( B1 => n842, B2 => n442, C1 => n1488, C2 => n445,
                           A => n2310, ZN => n2309);
   U2620 : AOI22_X1 port map( A1 => n448, A2 => n4057, B1 => n451, B2 => n1193,
                           ZN => n2310);
   U2621 : OAI221_X1 port map( B1 => n1490, B2 => n454, C1 => n938, C2 => n457,
                           A => n2311, ZN => n2308);
   U2622 : AOI22_X1 port map( A1 => n460, A2 => n1295, B1 => n463, B2 => n4025,
                           ZN => n2311);
   U2623 : OAI211_X1 port map( C1 => n522, C2 => n466, A => n2312, B => n2313, 
                           ZN => n2307);
   U2624 : AOI221_X1 port map( B1 => n469, B2 => n1154, C1 => n472, C2 => n4153
                           , A => n2314, ZN => n2313);
   U2625 : OAI22_X1 port map( A1 => n618, A2 => n473, B1 => n1495, B2 => n478, 
                           ZN => n2314);
   U2626 : AOI22_X1 port map( A1 => n481, A2 => n4185, B1 => n484, B2 => n1052,
                           ZN => n2312);
   U2627 : NAND4_X1 port map( A1 => n2315, A2 => n2316, A3 => n2317, A4 => 
                           n2318, ZN => n2306);
   U2628 : AOI221_X1 port map( B1 => n487, B2 => n4217, C1 => n490, C2 => n4249
                           , A => n2319, ZN => n2318);
   U2629 : OAI22_X1 port map( A1 => n394, A2 => n493, B1 => n362, B2 => n496, 
                           ZN => n2319);
   U2630 : AOI221_X1 port map( B1 => n499, B2 => n4281, C1 => n502, C2 => n4313
                           , A => n2320, ZN => n2317);
   U2631 : OAI22_X1 port map( A1 => n266, A2 => n505, B1 => n234, B2 => n25, ZN
                           => n2320);
   U2632 : AOI221_X1 port map( B1 => n508, B2 => n775, C1 => n511, C2 => n809, 
                           A => n2321, ZN => n2316);
   U2633 : OAI22_X1 port map( A1 => n1503, A2 => n514, B1 => n1504, B2 => n549,
                           ZN => n2321);
   U2634 : AOI221_X1 port map( B1 => n552, B2 => n736, C1 => n555, C2 => n3961,
                           A => n2322, ZN => n2315);
   U2635 : OAI22_X1 port map( A1 => n1506, A2 => n558, B1 => n1507, B2 => n561,
                           ZN => n2322);
   U2636 : OAI222_X1 port map( A1 => n587, A2 => n433, B1 => n2323, B2 => n436,
                           C1 => n3896, C2 => n439, ZN => n2531);
   U2637 : NOR4_X1 port map( A1 => n2324, A2 => n2325, A3 => n2326, A4 => n2327
                           , ZN => n2323);
   U2638 : OAI221_X1 port map( B1 => n843, B2 => n442, C1 => n1513, C2 => n445,
                           A => n2328, ZN => n2327);
   U2639 : AOI22_X1 port map( A1 => n448, A2 => n4056, B1 => n451, B2 => n1194,
                           ZN => n2328);
   U2640 : OAI221_X1 port map( B1 => n1515, B2 => n454, C1 => n939, C2 => n457,
                           A => n2329, ZN => n2326);
   U2641 : AOI22_X1 port map( A1 => n460, A2 => n1296, B1 => n463, B2 => n4024,
                           ZN => n2329);
   U2642 : OAI211_X1 port map( C1 => n523, C2 => n466, A => n2330, B => n2331, 
                           ZN => n2325);
   U2643 : AOI221_X1 port map( B1 => n469, B2 => n1155, C1 => n472, C2 => n4152
                           , A => n2332, ZN => n2331);
   U2644 : OAI22_X1 port map( A1 => n619, A2 => n28, B1 => n1520, B2 => n476, 
                           ZN => n2332);
   U2645 : AOI22_X1 port map( A1 => n481, A2 => n4184, B1 => n484, B2 => n1053,
                           ZN => n2330);
   U2646 : NAND4_X1 port map( A1 => n2333, A2 => n2334, A3 => n2335, A4 => 
                           n2336, ZN => n2324);
   U2647 : AOI221_X1 port map( B1 => n487, B2 => n4216, C1 => n490, C2 => n4248
                           , A => n2337, ZN => n2336);
   U2648 : OAI22_X1 port map( A1 => n395, A2 => n493, B1 => n363, B2 => n496, 
                           ZN => n2337);
   U2649 : AOI221_X1 port map( B1 => n499, B2 => n4280, C1 => n502, C2 => n4312
                           , A => n2338, ZN => n2335);
   U2650 : OAI22_X1 port map( A1 => n267, A2 => n505, B1 => n235, B2 => n24, ZN
                           => n2338);
   U2651 : AOI221_X1 port map( B1 => n508, B2 => n776, C1 => n511, C2 => n810, 
                           A => n2339, ZN => n2334);
   U2652 : OAI22_X1 port map( A1 => n1528, A2 => n514, B1 => n1529, B2 => n549,
                           ZN => n2339);
   U2653 : AOI221_X1 port map( B1 => n552, B2 => n737, C1 => n555, C2 => n3960,
                           A => n2340, ZN => n2333);
   U2654 : OAI22_X1 port map( A1 => n1531, A2 => n558, B1 => n1532, B2 => n561,
                           ZN => n2340);
   U2655 : OAI222_X1 port map( A1 => n586, A2 => n433, B1 => n2341, B2 => n436,
                           C1 => n3895, C2 => n439, ZN => n2530);
   U2656 : NOR4_X1 port map( A1 => n2342, A2 => n2343, A3 => n2344, A4 => n2345
                           , ZN => n2341);
   U2657 : OAI221_X1 port map( B1 => n844, B2 => n442, C1 => n1538, C2 => n445,
                           A => n2346, ZN => n2345);
   U2658 : AOI22_X1 port map( A1 => n448, A2 => n4055, B1 => n451, B2 => n1195,
                           ZN => n2346);
   U2659 : OAI221_X1 port map( B1 => n1540, B2 => n454, C1 => n940, C2 => n457,
                           A => n2347, ZN => n2344);
   U2660 : AOI22_X1 port map( A1 => n460, A2 => n1297, B1 => n463, B2 => n4023,
                           ZN => n2347);
   U2661 : OAI211_X1 port map( C1 => n524, C2 => n466, A => n2348, B => n2349, 
                           ZN => n2343);
   U2662 : AOI221_X1 port map( B1 => n469, B2 => n1156, C1 => n472, C2 => n4151
                           , A => n2350, ZN => n2349);
   U2663 : OAI22_X1 port map( A1 => n620, A2 => n27, B1 => n1545, B2 => n478, 
                           ZN => n2350);
   U2664 : AOI22_X1 port map( A1 => n481, A2 => n4183, B1 => n484, B2 => n1054,
                           ZN => n2348);
   U2665 : NAND4_X1 port map( A1 => n2351, A2 => n2352, A3 => n2353, A4 => 
                           n2354, ZN => n2342);
   U2666 : AOI221_X1 port map( B1 => n487, B2 => n4215, C1 => n490, C2 => n4247
                           , A => n2355, ZN => n2354);
   U2667 : OAI22_X1 port map( A1 => n396, A2 => n493, B1 => n364, B2 => n496, 
                           ZN => n2355);
   U2668 : AOI221_X1 port map( B1 => n499, B2 => n4279, C1 => n502, C2 => n4311
                           , A => n2356, ZN => n2353);
   U2669 : OAI22_X1 port map( A1 => n268, A2 => n505, B1 => n236, B2 => n25, ZN
                           => n2356);
   U2670 : AOI221_X1 port map( B1 => n508, B2 => n777, C1 => n511, C2 => n811, 
                           A => n2357, ZN => n2352);
   U2671 : OAI22_X1 port map( A1 => n1553, A2 => n514, B1 => n1554, B2 => n549,
                           ZN => n2357);
   U2672 : AOI221_X1 port map( B1 => n552, B2 => n738, C1 => n555, C2 => n3959,
                           A => n2358, ZN => n2351);
   U2673 : OAI22_X1 port map( A1 => n1556, A2 => n558, B1 => n1557, B2 => n561,
                           ZN => n2358);
   U2674 : OAI222_X1 port map( A1 => n585, A2 => n432, B1 => n2359, B2 => n435,
                           C1 => n3894, C2 => n439, ZN => n2529);
   U2675 : NOR4_X1 port map( A1 => n2360, A2 => n2361, A3 => n2362, A4 => n2363
                           , ZN => n2359);
   U2676 : OAI221_X1 port map( B1 => n845, B2 => n441, C1 => n1563, C2 => n444,
                           A => n2364, ZN => n2363);
   U2677 : AOI22_X1 port map( A1 => n447, A2 => n4054, B1 => n450, B2 => n1196,
                           ZN => n2364);
   U2678 : OAI221_X1 port map( B1 => n1565, B2 => n453, C1 => n941, C2 => n456,
                           A => n2365, ZN => n2362);
   U2679 : AOI22_X1 port map( A1 => n459, A2 => n1298, B1 => n462, B2 => n4022,
                           ZN => n2365);
   U2680 : OAI211_X1 port map( C1 => n525, C2 => n465, A => n2366, B => n2367, 
                           ZN => n2361);
   U2681 : AOI221_X1 port map( B1 => n468, B2 => n1157, C1 => n471, C2 => n4150
                           , A => n2368, ZN => n2367);
   U2682 : OAI22_X1 port map( A1 => n621, A2 => n474, B1 => n1570, B2 => n477, 
                           ZN => n2368);
   U2683 : AOI22_X1 port map( A1 => n480, A2 => n4182, B1 => n483, B2 => n1055,
                           ZN => n2366);
   U2684 : NAND4_X1 port map( A1 => n2369, A2 => n2372, A3 => n2371, A4 => 
                           n2370, ZN => n2360);
   U2685 : AOI221_X1 port map( B1 => n486, B2 => n4214, C1 => n489, C2 => n4246
                           , A => n2373, ZN => n2372);
   U2686 : OAI22_X1 port map( A1 => n397, A2 => n492, B1 => n365, B2 => n496, 
                           ZN => n2373);
   U2687 : AOI221_X1 port map( B1 => n498, B2 => n4278, C1 => n501, C2 => n4310
                           , A => n2374, ZN => n2371);
   U2688 : OAI22_X1 port map( A1 => n269, A2 => n504, B1 => n237, B2 => n25, ZN
                           => n2374);
   U2689 : AOI221_X1 port map( B1 => n507, B2 => n778, C1 => n510, C2 => n812, 
                           A => n2375, ZN => n2370);
   U2690 : OAI22_X1 port map( A1 => n1578, A2 => n513, B1 => n1579, B2 => n549,
                           ZN => n2375);
   U2691 : AOI221_X1 port map( B1 => n551, B2 => n739, C1 => n554, C2 => n3958,
                           A => n2376, ZN => n2369);
   U2692 : OAI22_X1 port map( A1 => n1581, A2 => n557, B1 => n1582, B2 => n560,
                           ZN => n2376);
   U2693 : OAI222_X1 port map( A1 => n584, A2 => n432, B1 => n2377, B2 => n435,
                           C1 => n3893, C2 => n439, ZN => n2528);
   U2694 : NOR4_X1 port map( A1 => n2378, A2 => n2379, A3 => n2380, A4 => n2381
                           , ZN => n2377);
   U2695 : OAI221_X1 port map( B1 => n846, B2 => n441, C1 => n1588, C2 => n444,
                           A => n2382, ZN => n2381);
   U2696 : AOI22_X1 port map( A1 => n447, A2 => n4053, B1 => n450, B2 => n1197,
                           ZN => n2382);
   U2697 : OAI221_X1 port map( B1 => n1590, B2 => n453, C1 => n942, C2 => n456,
                           A => n2383, ZN => n2380);
   U2698 : AOI22_X1 port map( A1 => n459, A2 => n1299, B1 => n462, B2 => n4021,
                           ZN => n2383);
   U2699 : OAI211_X1 port map( C1 => n526, C2 => n465, A => n2384, B => n2385, 
                           ZN => n2379);
   U2700 : AOI221_X1 port map( B1 => n468, B2 => n1158, C1 => n471, C2 => n4149
                           , A => n2386, ZN => n2385);
   U2701 : OAI22_X1 port map( A1 => n622, A2 => n474, B1 => n1595, B2 => n477, 
                           ZN => n2386);
   U2702 : AOI22_X1 port map( A1 => n480, A2 => n4181, B1 => n483, B2 => n1056,
                           ZN => n2384);
   U2703 : NAND4_X1 port map( A1 => n2387, A2 => n2390, A3 => n2389, A4 => 
                           n2388, ZN => n2378);
   U2704 : AOI221_X1 port map( B1 => n486, B2 => n4213, C1 => n489, C2 => n4245
                           , A => n2391, ZN => n2390);
   U2705 : OAI22_X1 port map( A1 => n398, A2 => n492, B1 => n366, B2 => n495, 
                           ZN => n2391);
   U2706 : AOI221_X1 port map( B1 => n498, B2 => n4277, C1 => n501, C2 => n4309
                           , A => n2392, ZN => n2389);
   U2707 : OAI22_X1 port map( A1 => n270, A2 => n504, B1 => n238, B2 => n24, ZN
                           => n2392);
   U2708 : AOI221_X1 port map( B1 => n507, B2 => n779, C1 => n510, C2 => n813, 
                           A => n2393, ZN => n2388);
   U2709 : OAI22_X1 port map( A1 => n1603, A2 => n513, B1 => n1604, B2 => n516,
                           ZN => n2393);
   U2710 : AOI221_X1 port map( B1 => n551, B2 => n740, C1 => n554, C2 => n3957,
                           A => n2394, ZN => n2387);
   U2711 : OAI22_X1 port map( A1 => n1606, A2 => n557, B1 => n1607, B2 => n560,
                           ZN => n2394);
   U2712 : OAI222_X1 port map( A1 => n583, A2 => n432, B1 => n2395, B2 => n435,
                           C1 => n3892, C2 => n438, ZN => n2527);
   U2713 : NOR4_X1 port map( A1 => n2396, A2 => n2397, A3 => n2398, A4 => n2399
                           , ZN => n2395);
   U2714 : OAI221_X1 port map( B1 => n847, B2 => n441, C1 => n1613, C2 => n444,
                           A => n2400, ZN => n2399);
   U2715 : AOI22_X1 port map( A1 => n447, A2 => n4052, B1 => n450, B2 => n1198,
                           ZN => n2400);
   U2716 : OAI221_X1 port map( B1 => n1615, B2 => n453, C1 => n943, C2 => n456,
                           A => n2401, ZN => n2398);
   U2717 : AOI22_X1 port map( A1 => n459, A2 => n1300, B1 => n462, B2 => n4020,
                           ZN => n2401);
   U2718 : OAI211_X1 port map( C1 => n527, C2 => n465, A => n2402, B => n2403, 
                           ZN => n2397);
   U2719 : AOI221_X1 port map( B1 => n468, B2 => n1159, C1 => n471, C2 => n4148
                           , A => n2404, ZN => n2403);
   U2720 : OAI22_X1 port map( A1 => n623, A2 => n474, B1 => n1620, B2 => n477, 
                           ZN => n2404);
   U2721 : AOI22_X1 port map( A1 => n480, A2 => n4180, B1 => n483, B2 => n1057,
                           ZN => n2402);
   U2722 : NAND4_X1 port map( A1 => n2405, A2 => n2408, A3 => n2407, A4 => 
                           n2406, ZN => n2396);
   U2723 : AOI221_X1 port map( B1 => n486, B2 => n4212, C1 => n489, C2 => n4244
                           , A => n2409, ZN => n2408);
   U2724 : OAI22_X1 port map( A1 => n399, A2 => n492, B1 => n367, B2 => n495, 
                           ZN => n2409);
   U2725 : AOI221_X1 port map( B1 => n498, B2 => n4276, C1 => n501, C2 => n4308
                           , A => n2410, ZN => n2407);
   U2726 : OAI22_X1 port map( A1 => n271, A2 => n504, B1 => n239, B2 => n25, ZN
                           => n2410);
   U2727 : AOI221_X1 port map( B1 => n507, B2 => n780, C1 => n510, C2 => n814, 
                           A => n2411, ZN => n2406);
   U2728 : OAI22_X1 port map( A1 => n1628, A2 => n513, B1 => n1629, B2 => n516,
                           ZN => n2411);
   U2729 : AOI221_X1 port map( B1 => n551, B2 => n741, C1 => n554, C2 => n3956,
                           A => n2412, ZN => n2405);
   U2730 : OAI22_X1 port map( A1 => n1631, A2 => n557, B1 => n1632, B2 => n560,
                           ZN => n2412);
   U2731 : OAI222_X1 port map( A1 => n582, A2 => n432, B1 => n2413, B2 => n435,
                           C1 => n3891, C2 => n438, ZN => n2526);
   U2732 : NOR4_X1 port map( A1 => n2414, A2 => n2415, A3 => n2416, A4 => n2417
                           , ZN => n2413);
   U2733 : OAI221_X1 port map( B1 => n848, B2 => n441, C1 => n1638, C2 => n444,
                           A => n2418, ZN => n2417);
   U2734 : AOI22_X1 port map( A1 => n447, A2 => n4051, B1 => n450, B2 => n1199,
                           ZN => n2418);
   U2735 : OAI221_X1 port map( B1 => n1640, B2 => n453, C1 => n944, C2 => n456,
                           A => n2419, ZN => n2416);
   U2736 : AOI22_X1 port map( A1 => n459, A2 => n1301, B1 => n462, B2 => n4019,
                           ZN => n2419);
   U2737 : OAI211_X1 port map( C1 => n528, C2 => n465, A => n2420, B => n2421, 
                           ZN => n2415);
   U2738 : AOI221_X1 port map( B1 => n468, B2 => n1160, C1 => n471, C2 => n4147
                           , A => n2422, ZN => n2421);
   U2739 : OAI22_X1 port map( A1 => n624, A2 => n475, B1 => n1645, B2 => n477, 
                           ZN => n2422);
   U2740 : AOI22_X1 port map( A1 => n480, A2 => n4179, B1 => n483, B2 => n1058,
                           ZN => n2420);
   U2741 : NAND4_X1 port map( A1 => n2423, A2 => n2426, A3 => n2425, A4 => 
                           n2424, ZN => n2414);
   U2742 : AOI221_X1 port map( B1 => n486, B2 => n4211, C1 => n489, C2 => n4243
                           , A => n2427, ZN => n2426);
   U2743 : OAI22_X1 port map( A1 => n400, A2 => n492, B1 => n368, B2 => n495, 
                           ZN => n2427);
   U2744 : AOI221_X1 port map( B1 => n498, B2 => n4275, C1 => n501, C2 => n4307
                           , A => n2428, ZN => n2425);
   U2745 : OAI22_X1 port map( A1 => n272, A2 => n504, B1 => n240, B2 => n24, ZN
                           => n2428);
   U2746 : AOI221_X1 port map( B1 => n507, B2 => n781, C1 => n510, C2 => n815, 
                           A => n2429, ZN => n2424);
   U2747 : OAI22_X1 port map( A1 => n1653, A2 => n513, B1 => n1654, B2 => n516,
                           ZN => n2429);
   U2748 : AOI221_X1 port map( B1 => n551, B2 => n742, C1 => n554, C2 => n3955,
                           A => n2430, ZN => n2423);
   U2749 : OAI22_X1 port map( A1 => n1656, A2 => n557, B1 => n1657, B2 => n560,
                           ZN => n2430);
   U2750 : OAI222_X1 port map( A1 => n581, A2 => n432, B1 => n2431, B2 => n435,
                           C1 => n3890, C2 => n438, ZN => n2525);
   U2751 : NOR4_X1 port map( A1 => n2432, A2 => n2433, A3 => n2434, A4 => n2435
                           , ZN => n2431);
   U2752 : OAI221_X1 port map( B1 => n849, B2 => n441, C1 => n1663, C2 => n444,
                           A => n2436, ZN => n2435);
   U2753 : AOI22_X1 port map( A1 => n447, A2 => n4050, B1 => n450, B2 => n1200,
                           ZN => n2436);
   U2754 : OAI221_X1 port map( B1 => n1665, B2 => n453, C1 => n945, C2 => n456,
                           A => n2437, ZN => n2434);
   U2755 : AOI22_X1 port map( A1 => n459, A2 => n1302, B1 => n462, B2 => n4018,
                           ZN => n2437);
   U2756 : OAI211_X1 port map( C1 => n529, C2 => n465, A => n2438, B => n2439, 
                           ZN => n2433);
   U2757 : AOI221_X1 port map( B1 => n468, B2 => n1161, C1 => n471, C2 => n4146
                           , A => n2440, ZN => n2439);
   U2758 : OAI22_X1 port map( A1 => n625, A2 => n473, B1 => n1670, B2 => n477, 
                           ZN => n2440);
   U2759 : AOI22_X1 port map( A1 => n480, A2 => n4178, B1 => n483, B2 => n1059,
                           ZN => n2438);
   U2760 : NAND4_X1 port map( A1 => n2441, A2 => n2444, A3 => n2443, A4 => 
                           n2442, ZN => n2432);
   U2761 : AOI221_X1 port map( B1 => n486, B2 => n4210, C1 => n489, C2 => n4242
                           , A => n2445, ZN => n2444);
   U2762 : OAI22_X1 port map( A1 => n401, A2 => n492, B1 => n369, B2 => n495, 
                           ZN => n2445);
   U2763 : AOI221_X1 port map( B1 => n498, B2 => n4274, C1 => n501, C2 => n4306
                           , A => n2446, ZN => n2443);
   U2764 : OAI22_X1 port map( A1 => n273, A2 => n504, B1 => n241, B2 => n25, ZN
                           => n2446);
   U2765 : AOI221_X1 port map( B1 => n507, B2 => n782, C1 => n510, C2 => n816, 
                           A => n2447, ZN => n2442);
   U2766 : OAI22_X1 port map( A1 => n1678, A2 => n513, B1 => n1679, B2 => n516,
                           ZN => n2447);
   U2767 : AOI221_X1 port map( B1 => n551, B2 => n743, C1 => n554, C2 => n3954,
                           A => n2448, ZN => n2441);
   U2768 : OAI22_X1 port map( A1 => n1681, A2 => n557, B1 => n1682, B2 => n560,
                           ZN => n2448);
   U2769 : OAI222_X1 port map( A1 => n580, A2 => n432, B1 => n2449, B2 => n435,
                           C1 => n3889, C2 => n438, ZN => n2524);
   U2770 : NOR4_X1 port map( A1 => n2450, A2 => n2451, A3 => n2452, A4 => n2453
                           , ZN => n2449);
   U2771 : OAI221_X1 port map( B1 => n850, B2 => n441, C1 => n1688, C2 => n444,
                           A => n2454, ZN => n2453);
   U2772 : AOI22_X1 port map( A1 => n447, A2 => n4049, B1 => n450, B2 => n1201,
                           ZN => n2454);
   U2773 : OAI221_X1 port map( B1 => n1690, B2 => n453, C1 => n946, C2 => n456,
                           A => n2455, ZN => n2452);
   U2774 : AOI22_X1 port map( A1 => n459, A2 => n1303, B1 => n462, B2 => n4017,
                           ZN => n2455);
   U2775 : OAI211_X1 port map( C1 => n530, C2 => n465, A => n2456, B => n2457, 
                           ZN => n2451);
   U2776 : AOI221_X1 port map( B1 => n468, B2 => n1162, C1 => n471, C2 => n4145
                           , A => n2458, ZN => n2457);
   U2777 : OAI22_X1 port map( A1 => n626, A2 => n28, B1 => n1695, B2 => n477, 
                           ZN => n2458);
   U2778 : AOI22_X1 port map( A1 => n480, A2 => n4177, B1 => n483, B2 => n1060,
                           ZN => n2456);
   U2779 : NAND4_X1 port map( A1 => n2459, A2 => n2462, A3 => n2461, A4 => 
                           n2460, ZN => n2450);
   U2780 : AOI221_X1 port map( B1 => n486, B2 => n4209, C1 => n489, C2 => n4241
                           , A => n2463, ZN => n2462);
   U2781 : OAI22_X1 port map( A1 => n402, A2 => n492, B1 => n370, B2 => n495, 
                           ZN => n2463);
   U2782 : AOI221_X1 port map( B1 => n498, B2 => n4273, C1 => n501, C2 => n4305
                           , A => n2464, ZN => n2461);
   U2783 : OAI22_X1 port map( A1 => n274, A2 => n504, B1 => n242, B2 => n24, ZN
                           => n2464);
   U2784 : AOI221_X1 port map( B1 => n507, B2 => n783, C1 => n510, C2 => n817, 
                           A => n2465, ZN => n2460);
   U2785 : OAI22_X1 port map( A1 => n1703, A2 => n513, B1 => n1704, B2 => n516,
                           ZN => n2465);
   U2786 : AOI221_X1 port map( B1 => n551, B2 => n744, C1 => n554, C2 => n3953,
                           A => n2466, ZN => n2459);
   U2787 : OAI22_X1 port map( A1 => n1706, A2 => n557, B1 => n1707, B2 => n560,
                           ZN => n2466);
   U2788 : OAI222_X1 port map( A1 => n579, A2 => n432, B1 => n2467, B2 => n435,
                           C1 => n3888, C2 => n438, ZN => n2523);
   U2789 : OAI221_X1 port map( B1 => n851, B2 => n441, C1 => n1713, C2 => n444,
                           A => n2472, ZN => n2471);
   U2790 : AOI22_X1 port map( A1 => n447, A2 => n4048, B1 => n450, B2 => n1202,
                           ZN => n2472);
   U2791 : OAI221_X1 port map( B1 => n1715, B2 => n453, C1 => n947, C2 => n456,
                           A => n2473, ZN => n2470);
   U2792 : AOI22_X1 port map( A1 => n459, A2 => n1304, B1 => n462, B2 => n4016,
                           ZN => n2473);
   U2793 : OAI211_X1 port map( C1 => n531, C2 => n465, A => n2474, B => n2475, 
                           ZN => n2469);
   U2794 : AOI221_X1 port map( B1 => n468, B2 => n1163, C1 => n471, C2 => n4144
                           , A => n2476, ZN => n2475);
   U2795 : OAI22_X1 port map( A1 => n627, A2 => n27, B1 => n1720, B2 => n476, 
                           ZN => n2476);
   U2796 : AOI22_X1 port map( A1 => n480, A2 => n4176, B1 => n483, B2 => n1061,
                           ZN => n2474);
   U2797 : NAND4_X1 port map( A1 => n2477, A2 => n2480, A3 => n2479, A4 => 
                           n2478, ZN => n2468);
   U2798 : AOI221_X1 port map( B1 => n486, B2 => n4208, C1 => n489, C2 => n4240
                           , A => n2481, ZN => n2480);
   U2799 : OAI22_X1 port map( A1 => n403, A2 => n492, B1 => n371, B2 => n495, 
                           ZN => n2481);
   U2800 : AOI221_X1 port map( B1 => n498, B2 => n4272, C1 => n501, C2 => n4304
                           , A => n2482, ZN => n2479);
   U2801 : OAI22_X1 port map( A1 => n275, A2 => n504, B1 => n243, B2 => n24, ZN
                           => n2482);
   U2802 : AOI221_X1 port map( B1 => n507, B2 => n784, C1 => n510, C2 => n818, 
                           A => n2483, ZN => n2478);
   U2803 : OAI22_X1 port map( A1 => n1728, A2 => n513, B1 => n1729, B2 => n516,
                           ZN => n2483);
   U2804 : AOI221_X1 port map( B1 => n551, B2 => n745, C1 => n554, C2 => n3952,
                           A => n2484, ZN => n2477);
   U2805 : OAI22_X1 port map( A1 => n1731, A2 => n557, B1 => n1732, B2 => n560,
                           ZN => n2484);
   U2806 : OAI222_X1 port map( A1 => n578, A2 => n432, B1 => n2485, B2 => n435,
                           C1 => n3887, C2 => n438, ZN => n2522);
   U2807 : OAI221_X1 port map( B1 => n852, B2 => n441, C1 => n1738, C2 => n444,
                           A => n2490, ZN => n2489);
   U2808 : AOI22_X1 port map( A1 => n447, A2 => n4047, B1 => n450, B2 => n1203,
                           ZN => n2490);
   U2809 : OAI221_X1 port map( B1 => n1740, B2 => n453, C1 => n948, C2 => n456,
                           A => n2491, ZN => n2488);
   U2810 : AOI22_X1 port map( A1 => n459, A2 => n1305, B1 => n462, B2 => n4015,
                           ZN => n2491);
   U2811 : OAI211_X1 port map( C1 => n532, C2 => n465, A => n2492, B => n2493, 
                           ZN => n2487);
   U2812 : AOI221_X1 port map( B1 => n468, B2 => n1164, C1 => n471, C2 => n4143
                           , A => n2494, ZN => n2493);
   U2813 : OAI22_X1 port map( A1 => n628, A2 => n27, B1 => n1745, B2 => n478, 
                           ZN => n2494);
   U2814 : AOI22_X1 port map( A1 => n480, A2 => n4175, B1 => n483, B2 => n1062,
                           ZN => n2492);
   U2815 : NAND4_X1 port map( A1 => n2495, A2 => n2498, A3 => n2497, A4 => 
                           n2496, ZN => n2486);
   U2816 : AOI221_X1 port map( B1 => n486, B2 => n4207, C1 => n489, C2 => n4239
                           , A => n2499, ZN => n2498);
   U2817 : OAI22_X1 port map( A1 => n404, A2 => n492, B1 => n372, B2 => n495, 
                           ZN => n2499);
   U2818 : AOI221_X1 port map( B1 => n498, B2 => n4271, C1 => n501, C2 => n4303
                           , A => n2500, ZN => n2497);
   U2819 : OAI22_X1 port map( A1 => n276, A2 => n504, B1 => n244, B2 => n25, ZN
                           => n2500);
   U2820 : AOI221_X1 port map( B1 => n507, B2 => n785, C1 => n510, C2 => n819, 
                           A => n2501, ZN => n2496);
   U2821 : OAI22_X1 port map( A1 => n1753, A2 => n513, B1 => n1754, B2 => n516,
                           ZN => n2501);
   U2822 : AOI221_X1 port map( B1 => n551, B2 => n746, C1 => n554, C2 => n3951,
                           A => n2502, ZN => n2495);
   U2823 : OAI22_X1 port map( A1 => n1756, A2 => n557, B1 => n1757, B2 => n560,
                           ZN => n2502);
   U2824 : OAI222_X1 port map( A1 => n577, A2 => n432, B1 => n2503, B2 => n435,
                           C1 => n3886, C2 => n438, ZN => n2521);
   U2825 : OAI221_X1 port map( B1 => n853, B2 => n441, C1 => n1763, C2 => n444,
                           A => n3564, ZN => n3563);
   U2826 : AOI22_X1 port map( A1 => n447, A2 => n4046, B1 => n450, B2 => n1204,
                           ZN => n3564);
   U2827 : OAI221_X1 port map( B1 => n1765, B2 => n453, C1 => n949, C2 => n456,
                           A => n3565, ZN => n3562);
   U2828 : AOI22_X1 port map( A1 => n459, A2 => n1306, B1 => n462, B2 => n4014,
                           ZN => n3565);
   U2829 : OAI211_X1 port map( C1 => n533, C2 => n465, A => n3566, B => n3567, 
                           ZN => n2505);
   U2830 : AOI221_X1 port map( B1 => n468, B2 => n1165, C1 => n471, C2 => n4142
                           , A => n3568, ZN => n3567);
   U2831 : OAI22_X1 port map( A1 => n629, A2 => n475, B1 => n1770, B2 => n476, 
                           ZN => n3568);
   U2832 : AOI22_X1 port map( A1 => n480, A2 => n4174, B1 => n483, B2 => n1063,
                           ZN => n3566);
   U2833 : NAND4_X1 port map( A1 => n3569, A2 => n3572, A3 => n3571, A4 => 
                           n3570, ZN => n2504);
   U2834 : AOI221_X1 port map( B1 => n486, B2 => n4206, C1 => n489, C2 => n4238
                           , A => n3573, ZN => n3572);
   U2835 : OAI22_X1 port map( A1 => n405, A2 => n492, B1 => n373, B2 => n495, 
                           ZN => n3573);
   U2836 : AOI221_X1 port map( B1 => n498, B2 => n4270, C1 => n501, C2 => n4302
                           , A => n3574, ZN => n3571);
   U2837 : OAI22_X1 port map( A1 => n277, A2 => n504, B1 => n245, B2 => n24, ZN
                           => n3574);
   U2838 : AOI221_X1 port map( B1 => n507, B2 => n786, C1 => n510, C2 => n820, 
                           A => n3575, ZN => n3570);
   U2839 : OAI22_X1 port map( A1 => n1778, A2 => n513, B1 => n1779, B2 => n516,
                           ZN => n3575);
   U2840 : AOI221_X1 port map( B1 => n551, B2 => n747, C1 => n554, C2 => n3950,
                           A => n3576, ZN => n3569);
   U2841 : OAI22_X1 port map( A1 => n1781, A2 => n557, B1 => n1782, B2 => n560,
                           ZN => n3576);
   U2842 : OAI222_X1 port map( A1 => n576, A2 => n432, B1 => n3577, B2 => n435,
                           C1 => n3885, C2 => n438, ZN => n2520);
   U2843 : OAI221_X1 port map( B1 => n854, B2 => n441, C1 => n1788, C2 => n444,
                           A => n3582, ZN => n3581);
   U2844 : AOI22_X1 port map( A1 => n447, A2 => n4045, B1 => n450, B2 => n1205,
                           ZN => n3582);
   U2845 : OAI221_X1 port map( B1 => n1790, B2 => n453, C1 => n950, C2 => n456,
                           A => n3583, ZN => n3580);
   U2846 : AOI22_X1 port map( A1 => n459, A2 => n1307, B1 => n462, B2 => n4013,
                           ZN => n3583);
   U2847 : OAI211_X1 port map( C1 => n534, C2 => n465, A => n3584, B => n3585, 
                           ZN => n3579);
   U2848 : AOI221_X1 port map( B1 => n468, B2 => n1166, C1 => n471, C2 => n4141
                           , A => n3586, ZN => n3585);
   U2849 : OAI22_X1 port map( A1 => n630, A2 => n473, B1 => n1795, B2 => n478, 
                           ZN => n3586);
   U2850 : AOI22_X1 port map( A1 => n480, A2 => n4173, B1 => n483, B2 => n1064,
                           ZN => n3584);
   U2851 : NAND4_X1 port map( A1 => n3587, A2 => n3590, A3 => n3589, A4 => 
                           n3588, ZN => n3578);
   U2852 : AOI221_X1 port map( B1 => n486, B2 => n4205, C1 => n489, C2 => n4237
                           , A => n3591, ZN => n3590);
   U2853 : OAI22_X1 port map( A1 => n406, A2 => n492, B1 => n374, B2 => n495, 
                           ZN => n3591);
   U2854 : AOI221_X1 port map( B1 => n498, B2 => n4269, C1 => n501, C2 => n4301
                           , A => n3592, ZN => n3589);
   U2855 : OAI22_X1 port map( A1 => n278, A2 => n504, B1 => n246, B2 => n25, ZN
                           => n3592);
   U2856 : AOI221_X1 port map( B1 => n507, B2 => n787, C1 => n510, C2 => n821, 
                           A => n3593, ZN => n3588);
   U2857 : OAI22_X1 port map( A1 => n1803, A2 => n513, B1 => n1804, B2 => n516,
                           ZN => n3593);
   U2858 : AOI221_X1 port map( B1 => n551, B2 => n748, C1 => n554, C2 => n3949,
                           A => n3594, ZN => n3587);
   U2859 : OAI22_X1 port map( A1 => n1806, A2 => n557, B1 => n1807, B2 => n560,
                           ZN => n3594);
   U2860 : OAI222_X1 port map( A1 => n575, A2 => n432, B1 => n3595, B2 => n435,
                           C1 => n3884, C2 => n438, ZN => n2519);
   U2861 : OAI221_X1 port map( B1 => n855, B2 => n441, C1 => n1813, C2 => n444,
                           A => n3600, ZN => n3599);
   U2862 : AOI22_X1 port map( A1 => n447, A2 => n4044, B1 => n450, B2 => n1206,
                           ZN => n3600);
   U2863 : OAI221_X1 port map( B1 => n1815, B2 => n453, C1 => n951, C2 => n456,
                           A => n3601, ZN => n3598);
   U2864 : AOI22_X1 port map( A1 => n459, A2 => n1308, B1 => n462, B2 => n4012,
                           ZN => n3601);
   U2865 : OAI211_X1 port map( C1 => n535, C2 => n465, A => n3602, B => n3603, 
                           ZN => n3597);
   U2866 : AOI221_X1 port map( B1 => n468, B2 => n1167, C1 => n471, C2 => n4140
                           , A => n3604, ZN => n3603);
   U2867 : OAI22_X1 port map( A1 => n631, A2 => n475, B1 => n1820, B2 => n476, 
                           ZN => n3604);
   U2868 : AOI22_X1 port map( A1 => n480, A2 => n4172, B1 => n483, B2 => n1065,
                           ZN => n3602);
   U2869 : NAND4_X1 port map( A1 => n3605, A2 => n3608, A3 => n3607, A4 => 
                           n3606, ZN => n3596);
   U2870 : AOI221_X1 port map( B1 => n486, B2 => n4204, C1 => n489, C2 => n4236
                           , A => n3609, ZN => n3608);
   U2871 : OAI22_X1 port map( A1 => n407, A2 => n492, B1 => n375, B2 => n495, 
                           ZN => n3609);
   U2872 : AOI221_X1 port map( B1 => n498, B2 => n4268, C1 => n501, C2 => n4300
                           , A => n3610, ZN => n3607);
   U2873 : OAI22_X1 port map( A1 => n279, A2 => n504, B1 => n247, B2 => n24, ZN
                           => n3610);
   U2874 : AOI221_X1 port map( B1 => n507, B2 => n788, C1 => n510, C2 => n822, 
                           A => n3611, ZN => n3606);
   U2875 : OAI22_X1 port map( A1 => n1828, A2 => n513, B1 => n1829, B2 => n516,
                           ZN => n3611);
   U2876 : AOI221_X1 port map( B1 => n551, B2 => n749, C1 => n554, C2 => n3948,
                           A => n3612, ZN => n3605);
   U2877 : OAI22_X1 port map( A1 => n1831, A2 => n557, B1 => n1832, B2 => n560,
                           ZN => n3612);
   U2878 : OAI222_X1 port map( A1 => n574, A2 => n432, B1 => n3613, B2 => n435,
                           C1 => n3883, C2 => n438, ZN => n2518);
   U2879 : OAI221_X1 port map( B1 => n856, B2 => n441, C1 => n1838, C2 => n444,
                           A => n3618, ZN => n3617);
   U2880 : AOI22_X1 port map( A1 => n447, A2 => n4043, B1 => n450, B2 => n1207,
                           ZN => n3618);
   U2881 : OAI221_X1 port map( B1 => n1840, B2 => n453, C1 => n952, C2 => n456,
                           A => n3619, ZN => n3616);
   U2882 : AOI22_X1 port map( A1 => n459, A2 => n1309, B1 => n462, B2 => n4011,
                           ZN => n3619);
   U2883 : OAI211_X1 port map( C1 => n536, C2 => n465, A => n3620, B => n3621, 
                           ZN => n3615);
   U2884 : AOI221_X1 port map( B1 => n468, B2 => n1168, C1 => n471, C2 => n4139
                           , A => n3622, ZN => n3621);
   U2885 : OAI22_X1 port map( A1 => n632, A2 => n473, B1 => n1845, B2 => n478, 
                           ZN => n3622);
   U2886 : AOI22_X1 port map( A1 => n480, A2 => n4171, B1 => n483, B2 => n1066,
                           ZN => n3620);
   U2887 : NAND4_X1 port map( A1 => n3623, A2 => n3626, A3 => n3625, A4 => 
                           n3624, ZN => n3614);
   U2888 : AOI221_X1 port map( B1 => n486, B2 => n4203, C1 => n489, C2 => n4235
                           , A => n3627, ZN => n3626);
   U2889 : OAI22_X1 port map( A1 => n408, A2 => n492, B1 => n376, B2 => n495, 
                           ZN => n3627);
   U2890 : AOI221_X1 port map( B1 => n498, B2 => n4267, C1 => n501, C2 => n4299
                           , A => n3628, ZN => n3625);
   U2891 : OAI22_X1 port map( A1 => n280, A2 => n504, B1 => n248, B2 => n25, ZN
                           => n3628);
   U2892 : AOI221_X1 port map( B1 => n507, B2 => n789, C1 => n510, C2 => n823, 
                           A => n3629, ZN => n3624);
   U2893 : OAI22_X1 port map( A1 => n1853, A2 => n513, B1 => n1854, B2 => n516,
                           ZN => n3629);
   U2894 : AOI221_X1 port map( B1 => n551, B2 => n750, C1 => n554, C2 => n3947,
                           A => n3630, ZN => n3623);
   U2895 : OAI22_X1 port map( A1 => n1856, A2 => n557, B1 => n1857, B2 => n560,
                           ZN => n3630);
   U2896 : OAI222_X1 port map( A1 => n573, A2 => n431, B1 => n3631, B2 => n434,
                           C1 => n3882, C2 => n438, ZN => n2517);
   U2897 : NOR4_X1 port map( A1 => n3632, A2 => n3633, A3 => n3634, A4 => n3635
                           , ZN => n3631);
   U2898 : OAI221_X1 port map( B1 => n857, B2 => n440, C1 => n1863, C2 => n443,
                           A => n3636, ZN => n3635);
   U2899 : AOI22_X1 port map( A1 => n446, A2 => n4042, B1 => n449, B2 => n1208,
                           ZN => n3636);
   U2900 : OAI221_X1 port map( B1 => n1865, B2 => n452, C1 => n953, C2 => n455,
                           A => n3637, ZN => n3634);
   U2901 : AOI22_X1 port map( A1 => n458, A2 => n1310, B1 => n461, B2 => n4010,
                           ZN => n3637);
   U2902 : OAI211_X1 port map( C1 => n537, C2 => n464, A => n3638, B => n3639, 
                           ZN => n3633);
   U2903 : AOI221_X1 port map( B1 => n467, B2 => n1169, C1 => n470, C2 => n4138
                           , A => n3640, ZN => n3639);
   U2904 : OAI22_X1 port map( A1 => n633, A2 => n474, B1 => n1870, B2 => n477, 
                           ZN => n3640);
   U2905 : AOI22_X1 port map( A1 => n479, A2 => n4170, B1 => n482, B2 => n1067,
                           ZN => n3638);
   U2906 : NAND4_X1 port map( A1 => n3641, A2 => n3642, A3 => n3643, A4 => 
                           n3644, ZN => n3632);
   U2907 : AOI221_X1 port map( B1 => n485, B2 => n4202, C1 => n488, C2 => n4234
                           , A => n3645, ZN => n3644);
   U2908 : OAI22_X1 port map( A1 => n409, A2 => n491, B1 => n377, B2 => n494, 
                           ZN => n3645);
   U2909 : AOI221_X1 port map( B1 => n497, B2 => n4266, C1 => n500, C2 => n4298
                           , A => n3646, ZN => n3643);
   U2910 : OAI22_X1 port map( A1 => n281, A2 => n503, B1 => n249, B2 => n24, ZN
                           => n3646);
   U2911 : OAI22_X1 port map( A1 => n1878, A2 => n512, B1 => n1879, B2 => n515,
                           ZN => n3647);
   U2912 : AOI221_X1 port map( B1 => n550, B2 => n751, C1 => n553, C2 => n3946,
                           A => n3648, ZN => n3641);
   U2913 : OAI22_X1 port map( A1 => n1881, A2 => n556, B1 => n1882, B2 => n559,
                           ZN => n3648);
   U2914 : OAI222_X1 port map( A1 => n572, A2 => n431, B1 => n3649, B2 => n434,
                           C1 => n3881, C2 => n438, ZN => n2516);
   U2915 : NOR4_X1 port map( A1 => n3650, A2 => n3651, A3 => n3652, A4 => n3653
                           , ZN => n3649);
   U2916 : OAI221_X1 port map( B1 => n858, B2 => n440, C1 => n1888, C2 => n443,
                           A => n3654, ZN => n3653);
   U2917 : AOI22_X1 port map( A1 => n446, A2 => n4041, B1 => n449, B2 => n1209,
                           ZN => n3654);
   U2918 : OAI221_X1 port map( B1 => n1890, B2 => n452, C1 => n954, C2 => n455,
                           A => n3655, ZN => n3652);
   U2919 : AOI22_X1 port map( A1 => n458, A2 => n1311, B1 => n461, B2 => n4009,
                           ZN => n3655);
   U2920 : OAI211_X1 port map( C1 => n538, C2 => n464, A => n3656, B => n3657, 
                           ZN => n3651);
   U2921 : AOI221_X1 port map( B1 => n467, B2 => n1170, C1 => n470, C2 => n4137
                           , A => n3658, ZN => n3657);
   U2922 : OAI22_X1 port map( A1 => n634, A2 => n474, B1 => n1895, B2 => n477, 
                           ZN => n3658);
   U2923 : AOI22_X1 port map( A1 => n479, A2 => n4169, B1 => n482, B2 => n1068,
                           ZN => n3656);
   U2924 : NAND4_X1 port map( A1 => n3659, A2 => n3660, A3 => n3661, A4 => 
                           n3662, ZN => n3650);
   U2925 : AOI221_X1 port map( B1 => n485, B2 => n4201, C1 => n488, C2 => n4233
                           , A => n3663, ZN => n3662);
   U2926 : OAI22_X1 port map( A1 => n410, A2 => n491, B1 => n378, B2 => n494, 
                           ZN => n3663);
   U2927 : AOI221_X1 port map( B1 => n497, B2 => n4265, C1 => n500, C2 => n4297
                           , A => n3664, ZN => n3661);
   U2928 : OAI22_X1 port map( A1 => n282, A2 => n503, B1 => n250, B2 => n25, ZN
                           => n3664);
   U2929 : OAI22_X1 port map( A1 => n1903, A2 => n512, B1 => n1904, B2 => n515,
                           ZN => n3665);
   U2930 : AOI221_X1 port map( B1 => n550, B2 => n752, C1 => n553, C2 => n3945,
                           A => n3666, ZN => n3659);
   U2931 : OAI22_X1 port map( A1 => n1906, A2 => n556, B1 => n1907, B2 => n559,
                           ZN => n3666);
   U2932 : OAI222_X1 port map( A1 => n571, A2 => n431, B1 => n3667, B2 => n434,
                           C1 => n3880, C2 => n437, ZN => n2515);
   U2933 : OAI221_X1 port map( B1 => n859, B2 => n440, C1 => n1913, C2 => n443,
                           A => n3672, ZN => n3671);
   U2934 : AOI22_X1 port map( A1 => n446, A2 => n4040, B1 => n449, B2 => n1210,
                           ZN => n3672);
   U2935 : OAI221_X1 port map( B1 => n1915, B2 => n452, C1 => n955, C2 => n455,
                           A => n3673, ZN => n3670);
   U2936 : AOI22_X1 port map( A1 => n458, A2 => n1312, B1 => n461, B2 => n4008,
                           ZN => n3673);
   U2937 : OAI211_X1 port map( C1 => n539, C2 => n464, A => n3674, B => n3675, 
                           ZN => n3669);
   U2938 : AOI221_X1 port map( B1 => n467, B2 => n1171, C1 => n470, C2 => n4136
                           , A => n3676, ZN => n3675);
   U2939 : OAI22_X1 port map( A1 => n635, A2 => n475, B1 => n1920, B2 => n476, 
                           ZN => n3676);
   U2940 : AOI22_X1 port map( A1 => n479, A2 => n4168, B1 => n482, B2 => n1069,
                           ZN => n3674);
   U2941 : NAND4_X1 port map( A1 => n3677, A2 => n3678, A3 => n3679, A4 => 
                           n3680, ZN => n3668);
   U2942 : AOI221_X1 port map( B1 => n485, B2 => n4200, C1 => n488, C2 => n4232
                           , A => n3681, ZN => n3680);
   U2943 : OAI22_X1 port map( A1 => n411, A2 => n491, B1 => n379, B2 => n494, 
                           ZN => n3681);
   U2944 : AOI221_X1 port map( B1 => n497, B2 => n4264, C1 => n500, C2 => n4296
                           , A => n3682, ZN => n3679);
   U2945 : OAI22_X1 port map( A1 => n283, A2 => n503, B1 => n251, B2 => n24, ZN
                           => n3682);
   U2946 : AOI221_X1 port map( B1 => n506, B2 => n792, C1 => n509, C2 => n826, 
                           A => n3683, ZN => n3678);
   U2947 : OAI22_X1 port map( A1 => n1928, A2 => n512, B1 => n1929, B2 => n515,
                           ZN => n3683);
   U2948 : AOI221_X1 port map( B1 => n550, B2 => n753, C1 => n553, C2 => n3944,
                           A => n3684, ZN => n3677);
   U2949 : OAI22_X1 port map( A1 => n1931, A2 => n556, B1 => n1932, B2 => n559,
                           ZN => n3684);
   U2950 : OAI222_X1 port map( A1 => n570, A2 => n431, B1 => n3685, B2 => n434,
                           C1 => n3879, C2 => n437, ZN => n2514);
   U2951 : OAI221_X1 port map( B1 => n860, B2 => n440, C1 => n1938, C2 => n443,
                           A => n3690, ZN => n3689);
   U2952 : AOI22_X1 port map( A1 => n446, A2 => n4039, B1 => n449, B2 => n1211,
                           ZN => n3690);
   U2953 : OAI221_X1 port map( B1 => n1940, B2 => n452, C1 => n956, C2 => n455,
                           A => n3691, ZN => n3688);
   U2954 : AOI22_X1 port map( A1 => n458, A2 => n1313, B1 => n461, B2 => n4007,
                           ZN => n3691);
   U2955 : OAI211_X1 port map( C1 => n540, C2 => n464, A => n3692, B => n3693, 
                           ZN => n3687);
   U2956 : AOI221_X1 port map( B1 => n467, B2 => n1172, C1 => n470, C2 => n4135
                           , A => n3694, ZN => n3693);
   U2957 : OAI22_X1 port map( A1 => n636, A2 => n475, B1 => n1945, B2 => n478, 
                           ZN => n3694);
   U2958 : AOI22_X1 port map( A1 => n479, A2 => n4167, B1 => n482, B2 => n1070,
                           ZN => n3692);
   U2959 : NAND4_X1 port map( A1 => n3695, A2 => n3696, A3 => n3697, A4 => 
                           n3698, ZN => n3686);
   U2960 : AOI221_X1 port map( B1 => n485, B2 => n4199, C1 => n488, C2 => n4231
                           , A => n3699, ZN => n3698);
   U2961 : OAI22_X1 port map( A1 => n412, A2 => n491, B1 => n380, B2 => n494, 
                           ZN => n3699);
   U2962 : AOI221_X1 port map( B1 => n497, B2 => n4263, C1 => n500, C2 => n4295
                           , A => n3700, ZN => n3697);
   U2963 : OAI22_X1 port map( A1 => n284, A2 => n503, B1 => n252, B2 => n25, ZN
                           => n3700);
   U2964 : OAI22_X1 port map( A1 => n1953, A2 => n512, B1 => n1954, B2 => n515,
                           ZN => n3701);
   U2965 : AOI221_X1 port map( B1 => n550, B2 => n754, C1 => n553, C2 => n3943,
                           A => n3702, ZN => n3695);
   U2966 : OAI22_X1 port map( A1 => n1956, A2 => n556, B1 => n1957, B2 => n559,
                           ZN => n3702);
   U2967 : OAI222_X1 port map( A1 => n569, A2 => n431, B1 => n3703, B2 => n434,
                           C1 => n3878, C2 => n437, ZN => n2513);
   U2968 : NOR4_X1 port map( A1 => n3704, A2 => n3705, A3 => n3706, A4 => n3707
                           , ZN => n3703);
   U2969 : OAI221_X1 port map( B1 => n861, B2 => n440, C1 => n1963, C2 => n443,
                           A => n3708, ZN => n3707);
   U2970 : AOI22_X1 port map( A1 => n446, A2 => n4038, B1 => n449, B2 => n1212,
                           ZN => n3708);
   U2971 : OAI221_X1 port map( B1 => n1965, B2 => n452, C1 => n957, C2 => n455,
                           A => n3709, ZN => n3706);
   U2972 : AOI22_X1 port map( A1 => n458, A2 => n1314, B1 => n461, B2 => n4006,
                           ZN => n3709);
   U2973 : OAI211_X1 port map( C1 => n541, C2 => n464, A => n3710, B => n3711, 
                           ZN => n3705);
   U2974 : AOI221_X1 port map( B1 => n467, B2 => n1173, C1 => n470, C2 => n4134
                           , A => n3712, ZN => n3711);
   U2975 : OAI22_X1 port map( A1 => n637, A2 => n474, B1 => n1970, B2 => n477, 
                           ZN => n3712);
   U2976 : AOI22_X1 port map( A1 => n479, A2 => n4166, B1 => n482, B2 => n1071,
                           ZN => n3710);
   U2977 : NAND4_X1 port map( A1 => n3713, A2 => n3714, A3 => n3715, A4 => 
                           n3716, ZN => n3704);
   U2978 : AOI221_X1 port map( B1 => n485, B2 => n4198, C1 => n488, C2 => n4230
                           , A => n3717, ZN => n3716);
   U2979 : OAI22_X1 port map( A1 => n413, A2 => n491, B1 => n381, B2 => n494, 
                           ZN => n3717);
   U2980 : AOI221_X1 port map( B1 => n497, B2 => n4262, C1 => n500, C2 => n4294
                           , A => n3718, ZN => n3715);
   U2981 : OAI22_X1 port map( A1 => n285, A2 => n503, B1 => n253, B2 => n24, ZN
                           => n3718);
   U2982 : OAI22_X1 port map( A1 => n1978, A2 => n512, B1 => n1979, B2 => n515,
                           ZN => n3719);
   U2983 : AOI221_X1 port map( B1 => n550, B2 => n755, C1 => n553, C2 => n3942,
                           A => n3720, ZN => n3713);
   U2984 : OAI22_X1 port map( A1 => n1981, A2 => n556, B1 => n1982, B2 => n559,
                           ZN => n3720);
   U2985 : OAI222_X1 port map( A1 => n568, A2 => n431, B1 => n3721, B2 => n434,
                           C1 => n3877, C2 => n437, ZN => n2512);
   U2986 : OAI221_X1 port map( B1 => n862, B2 => n440, C1 => n1988, C2 => n443,
                           A => n3726, ZN => n3725);
   U2987 : AOI22_X1 port map( A1 => n446, A2 => n4037, B1 => n449, B2 => n1213,
                           ZN => n3726);
   U2988 : OAI221_X1 port map( B1 => n1990, B2 => n452, C1 => n958, C2 => n455,
                           A => n3727, ZN => n3724);
   U2989 : AOI22_X1 port map( A1 => n458, A2 => n1315, B1 => n461, B2 => n4005,
                           ZN => n3727);
   U2990 : OAI211_X1 port map( C1 => n542, C2 => n464, A => n3728, B => n3729, 
                           ZN => n3723);
   U2991 : AOI221_X1 port map( B1 => n467, B2 => n1174, C1 => n470, C2 => n4133
                           , A => n3730, ZN => n3729);
   U2992 : OAI22_X1 port map( A1 => n638, A2 => n28, B1 => n1995, B2 => n476, 
                           ZN => n3730);
   U2993 : AOI22_X1 port map( A1 => n479, A2 => n4165, B1 => n482, B2 => n1072,
                           ZN => n3728);
   U2994 : NAND4_X1 port map( A1 => n3731, A2 => n3732, A3 => n3733, A4 => 
                           n3734, ZN => n3722);
   U2995 : AOI221_X1 port map( B1 => n485, B2 => n4197, C1 => n488, C2 => n4229
                           , A => n3735, ZN => n3734);
   U2996 : OAI22_X1 port map( A1 => n414, A2 => n491, B1 => n382, B2 => n494, 
                           ZN => n3735);
   U2997 : AOI221_X1 port map( B1 => n497, B2 => n4261, C1 => n500, C2 => n4293
                           , A => n3736, ZN => n3733);
   U2998 : OAI22_X1 port map( A1 => n286, A2 => n503, B1 => n254, B2 => n24, ZN
                           => n3736);
   U2999 : OAI22_X1 port map( A1 => n2003, A2 => n512, B1 => n2004, B2 => n515,
                           ZN => n3737);
   U3000 : AOI221_X1 port map( B1 => n550, B2 => n756, C1 => n553, C2 => n3941,
                           A => n3738, ZN => n3731);
   U3001 : OAI22_X1 port map( A1 => n2006, A2 => n556, B1 => n2007, B2 => n559,
                           ZN => n3738);
   U3002 : OAI222_X1 port map( A1 => n567, A2 => n431, B1 => n3739, B2 => n434,
                           C1 => n3876, C2 => n437, ZN => n2511);
   U3003 : OAI221_X1 port map( B1 => n863, B2 => n440, C1 => n2013, C2 => n443,
                           A => n3744, ZN => n3743);
   U3004 : AOI22_X1 port map( A1 => n446, A2 => n4036, B1 => n449, B2 => n1214,
                           ZN => n3744);
   U3005 : OAI221_X1 port map( B1 => n2015, B2 => n452, C1 => n959, C2 => n455,
                           A => n3745, ZN => n3742);
   U3006 : AOI22_X1 port map( A1 => n458, A2 => n1316, B1 => n461, B2 => n4004,
                           ZN => n3745);
   U3007 : OAI211_X1 port map( C1 => n543, C2 => n464, A => n3746, B => n3747, 
                           ZN => n3741);
   U3008 : AOI221_X1 port map( B1 => n467, B2 => n1175, C1 => n470, C2 => n4132
                           , A => n3748, ZN => n3747);
   U3009 : OAI22_X1 port map( A1 => n639, A2 => n27, B1 => n2020, B2 => n478, 
                           ZN => n3748);
   U3010 : AOI22_X1 port map( A1 => n479, A2 => n4164, B1 => n482, B2 => n1073,
                           ZN => n3746);
   U3011 : NAND4_X1 port map( A1 => n3749, A2 => n3750, A3 => n3751, A4 => 
                           n3752, ZN => n3740);
   U3012 : AOI221_X1 port map( B1 => n485, B2 => n4196, C1 => n488, C2 => n4228
                           , A => n3753, ZN => n3752);
   U3013 : OAI22_X1 port map( A1 => n415, A2 => n491, B1 => n383, B2 => n494, 
                           ZN => n3753);
   U3014 : AOI221_X1 port map( B1 => n497, B2 => n4260, C1 => n500, C2 => n4292
                           , A => n3754, ZN => n3751);
   U3015 : OAI22_X1 port map( A1 => n287, A2 => n503, B1 => n255, B2 => n25, ZN
                           => n3754);
   U3016 : OAI22_X1 port map( A1 => n2028, A2 => n512, B1 => n2029, B2 => n515,
                           ZN => n3755);
   U3017 : AOI221_X1 port map( B1 => n550, B2 => n757, C1 => n553, C2 => n3940,
                           A => n3756, ZN => n3749);
   U3018 : OAI22_X1 port map( A1 => n2031, A2 => n556, B1 => n2032, B2 => n559,
                           ZN => n3756);
   U3019 : OAI222_X1 port map( A1 => n566, A2 => n431, B1 => n3757, B2 => n434,
                           C1 => n3875, C2 => n437, ZN => n2510);
   U3020 : OAI221_X1 port map( B1 => n864, B2 => n440, C1 => n2038, C2 => n443,
                           A => n3762, ZN => n3761);
   U3021 : AOI22_X1 port map( A1 => n446, A2 => n4035, B1 => n449, B2 => n1215,
                           ZN => n3762);
   U3022 : OAI221_X1 port map( B1 => n2040, B2 => n452, C1 => n960, C2 => n455,
                           A => n3763, ZN => n3760);
   U3023 : AOI22_X1 port map( A1 => n458, A2 => n1317, B1 => n461, B2 => n4003,
                           ZN => n3763);
   U3024 : OAI211_X1 port map( C1 => n544, C2 => n464, A => n3764, B => n3765, 
                           ZN => n3759);
   U3025 : AOI221_X1 port map( B1 => n467, B2 => n1176, C1 => n470, C2 => n4131
                           , A => n3766, ZN => n3765);
   U3026 : OAI22_X1 port map( A1 => n640, A2 => n473, B1 => n2045, B2 => n476, 
                           ZN => n3766);
   U3027 : AOI22_X1 port map( A1 => n479, A2 => n4163, B1 => n482, B2 => n1074,
                           ZN => n3764);
   U3028 : NAND4_X1 port map( A1 => n3767, A2 => n3768, A3 => n3769, A4 => 
                           n3770, ZN => n3758);
   U3029 : AOI221_X1 port map( B1 => n485, B2 => n4195, C1 => n488, C2 => n4227
                           , A => n3771, ZN => n3770);
   U3030 : OAI22_X1 port map( A1 => n416, A2 => n491, B1 => n384, B2 => n494, 
                           ZN => n3771);
   U3031 : AOI221_X1 port map( B1 => n497, B2 => n4259, C1 => n500, C2 => n4291
                           , A => n3772, ZN => n3769);
   U3032 : OAI22_X1 port map( A1 => n288, A2 => n503, B1 => n256, B2 => n24, ZN
                           => n3772);
   U3033 : AOI221_X1 port map( B1 => n506, B2 => n797, C1 => n509, C2 => n831, 
                           A => n3773, ZN => n3768);
   U3034 : OAI22_X1 port map( A1 => n2053, A2 => n512, B1 => n2054, B2 => n515,
                           ZN => n3773);
   U3035 : AOI221_X1 port map( B1 => n550, B2 => n758, C1 => n553, C2 => n3939,
                           A => n3774, ZN => n3767);
   U3036 : OAI22_X1 port map( A1 => n2056, A2 => n556, B1 => n2057, B2 => n559,
                           ZN => n3774);
   U3037 : OAI222_X1 port map( A1 => n565, A2 => n431, B1 => n3775, B2 => n434,
                           C1 => n3874, C2 => n437, ZN => n2509);
   U3038 : OAI221_X1 port map( B1 => n865, B2 => n440, C1 => n2063, C2 => n443,
                           A => n3780, ZN => n3779);
   U3039 : AOI22_X1 port map( A1 => n446, A2 => n4034, B1 => n449, B2 => n1216,
                           ZN => n3780);
   U3040 : OAI221_X1 port map( B1 => n2065, B2 => n452, C1 => n961, C2 => n455,
                           A => n3781, ZN => n3778);
   U3041 : AOI22_X1 port map( A1 => n458, A2 => n1318, B1 => n461, B2 => n4002,
                           ZN => n3781);
   U3042 : OAI211_X1 port map( C1 => n545, C2 => n464, A => n3782, B => n3783, 
                           ZN => n3777);
   U3043 : AOI221_X1 port map( B1 => n467, B2 => n1177, C1 => n470, C2 => n4130
                           , A => n3784, ZN => n3783);
   U3044 : OAI22_X1 port map( A1 => n641, A2 => n28, B1 => n2070, B2 => n478, 
                           ZN => n3784);
   U3045 : AOI22_X1 port map( A1 => n479, A2 => n4162, B1 => n482, B2 => n1075,
                           ZN => n3782);
   U3046 : NAND4_X1 port map( A1 => n3785, A2 => n3786, A3 => n3787, A4 => 
                           n3788, ZN => n3776);
   U3047 : AOI221_X1 port map( B1 => n485, B2 => n4194, C1 => n488, C2 => n4226
                           , A => n3789, ZN => n3788);
   U3048 : OAI22_X1 port map( A1 => n417, A2 => n491, B1 => n385, B2 => n494, 
                           ZN => n3789);
   U3049 : AOI221_X1 port map( B1 => n497, B2 => n4258, C1 => n500, C2 => n4290
                           , A => n3790, ZN => n3787);
   U3050 : OAI22_X1 port map( A1 => n289, A2 => n503, B1 => n257, B2 => n25, ZN
                           => n3790);
   U3051 : AOI221_X1 port map( B1 => n506, B2 => n798, C1 => n509, C2 => n832, 
                           A => n3791, ZN => n3786);
   U3052 : OAI22_X1 port map( A1 => n2078, A2 => n512, B1 => n2079, B2 => n515,
                           ZN => n3791);
   U3053 : AOI221_X1 port map( B1 => n550, B2 => n759, C1 => n553, C2 => n3938,
                           A => n3792, ZN => n3785);
   U3054 : OAI22_X1 port map( A1 => n2081, A2 => n556, B1 => n2082, B2 => n559,
                           ZN => n3792);
   U3055 : OAI222_X1 port map( A1 => n564, A2 => n431, B1 => n3793, B2 => n434,
                           C1 => n3873, C2 => n437, ZN => n2508);
   U3056 : OAI221_X1 port map( B1 => n866, B2 => n440, C1 => n2088, C2 => n443,
                           A => n3798, ZN => n3797);
   U3057 : AOI22_X1 port map( A1 => n446, A2 => n4033, B1 => n449, B2 => n1217,
                           ZN => n3798);
   U3058 : OAI221_X1 port map( B1 => n2090, B2 => n452, C1 => n962, C2 => n455,
                           A => n3799, ZN => n3796);
   U3059 : AOI22_X1 port map( A1 => n458, A2 => n1319, B1 => n461, B2 => n4001,
                           ZN => n3799);
   U3060 : OAI211_X1 port map( C1 => n546, C2 => n464, A => n3800, B => n3801, 
                           ZN => n3795);
   U3061 : AOI221_X1 port map( B1 => n467, B2 => n1178, C1 => n470, C2 => n4129
                           , A => n3802, ZN => n3801);
   U3062 : OAI22_X1 port map( A1 => n642, A2 => n27, B1 => n2095, B2 => n476, 
                           ZN => n3802);
   U3063 : AOI22_X1 port map( A1 => n479, A2 => n4161, B1 => n482, B2 => n1076,
                           ZN => n3800);
   U3064 : NAND4_X1 port map( A1 => n3803, A2 => n3804, A3 => n3805, A4 => 
                           n3806, ZN => n3794);
   U3065 : AOI221_X1 port map( B1 => n485, B2 => n4193, C1 => n488, C2 => n4225
                           , A => n3807, ZN => n3806);
   U3066 : OAI22_X1 port map( A1 => n418, A2 => n491, B1 => n386, B2 => n494, 
                           ZN => n3807);
   U3067 : AOI221_X1 port map( B1 => n497, B2 => n4257, C1 => n500, C2 => n4289
                           , A => n3808, ZN => n3805);
   U3068 : OAI22_X1 port map( A1 => n290, A2 => n503, B1 => n258, B2 => n24, ZN
                           => n3808);
   U3069 : OAI22_X1 port map( A1 => n2103, A2 => n512, B1 => n2104, B2 => n515,
                           ZN => n3809);
   U3070 : AOI221_X1 port map( B1 => n550, B2 => n760, C1 => n553, C2 => n3937,
                           A => n3810, ZN => n3803);
   U3071 : OAI22_X1 port map( A1 => n2106, A2 => n556, B1 => n2107, B2 => n559,
                           ZN => n3810);
   U3072 : OAI222_X1 port map( A1 => n563, A2 => n431, B1 => n3811, B2 => n434,
                           C1 => n3872, C2 => n437, ZN => n2507);
   U3073 : OAI221_X1 port map( B1 => n867, B2 => n440, C1 => n2113, C2 => n443,
                           A => n3816, ZN => n3815);
   U3074 : AOI22_X1 port map( A1 => n446, A2 => n4032, B1 => n449, B2 => n1218,
                           ZN => n3816);
   U3075 : OAI221_X1 port map( B1 => n2115, B2 => n452, C1 => n963, C2 => n455,
                           A => n3817, ZN => n3814);
   U3076 : AOI22_X1 port map( A1 => n458, A2 => n1320, B1 => n461, B2 => n4000,
                           ZN => n3817);
   U3077 : OAI211_X1 port map( C1 => n547, C2 => n464, A => n3818, B => n3819, 
                           ZN => n3813);
   U3078 : AOI221_X1 port map( B1 => n467, B2 => n1179, C1 => n470, C2 => n4128
                           , A => n3820, ZN => n3819);
   U3079 : OAI22_X1 port map( A1 => n643, A2 => n475, B1 => n2120, B2 => n478, 
                           ZN => n3820);
   U3080 : AOI22_X1 port map( A1 => n479, A2 => n4160, B1 => n482, B2 => n1077,
                           ZN => n3818);
   U3081 : NAND4_X1 port map( A1 => n3821, A2 => n3822, A3 => n3823, A4 => 
                           n3824, ZN => n3812);
   U3082 : AOI221_X1 port map( B1 => n485, B2 => n4192, C1 => n488, C2 => n4224
                           , A => n3825, ZN => n3824);
   U3083 : OAI22_X1 port map( A1 => n419, A2 => n491, B1 => n387, B2 => n494, 
                           ZN => n3825);
   U3084 : AOI221_X1 port map( B1 => n497, B2 => n4256, C1 => n500, C2 => n4288
                           , A => n3826, ZN => n3823);
   U3085 : OAI22_X1 port map( A1 => n291, A2 => n503, B1 => n259, B2 => n25, ZN
                           => n3826);
   U3086 : AOI221_X1 port map( B1 => n506, B2 => n800, C1 => n509, C2 => n834, 
                           A => n3827, ZN => n3822);
   U3087 : OAI22_X1 port map( A1 => n2128, A2 => n512, B1 => n2129, B2 => n515,
                           ZN => n3827);
   U3088 : AOI221_X1 port map( B1 => n550, B2 => n761, C1 => n553, C2 => n3936,
                           A => n3828, ZN => n3821);
   U3089 : OAI22_X1 port map( A1 => n2131, A2 => n556, B1 => n2132, B2 => n559,
                           ZN => n3828);
   U3090 : OAI222_X1 port map( A1 => n562, A2 => n431, B1 => n3829, B2 => n434,
                           C1 => n3871, C2 => n437, ZN => n2506);
   U3091 : NAND2_X1 port map( A1 => n437, A2 => n3830, ZN => n2183);
   U3092 : NOR4_X1 port map( A1 => n3831, A2 => n3832, A3 => n3833, A4 => n3834
                           , ZN => n3829);
   U3093 : OAI221_X1 port map( B1 => n868, B2 => n440, C1 => n2139, C2 => n443,
                           A => n3835, ZN => n3834);
   U3094 : AOI22_X1 port map( A1 => n446, A2 => n4031, B1 => n449, B2 => n1219,
                           ZN => n3835);
   U3095 : AND2_X1 port map( A1 => n3836, A2 => n3837, ZN => n2193);
   U3096 : AND2_X1 port map( A1 => n3836, A2 => n3838, ZN => n2192);
   U3097 : NAND2_X1 port map( A1 => n3839, A2 => n3840, ZN => n2190);
   U3098 : NAND2_X1 port map( A1 => n3841, A2 => n3837, ZN => n2189);
   U3099 : OAI221_X1 port map( B1 => n2147, B2 => n452, C1 => n964, C2 => n455,
                           A => n3842, ZN => n3833);
   U3100 : AOI22_X1 port map( A1 => n458, A2 => n1321, B1 => n461, B2 => n3999,
                           ZN => n3842);
   U3101 : AND2_X1 port map( A1 => n3841, A2 => n3838, ZN => n2198);
   U3102 : AND2_X1 port map( A1 => n3841, A2 => n3840, ZN => n2197);
   U3103 : NAND2_X1 port map( A1 => n3836, A2 => n3840, ZN => n2195);
   U3104 : NAND2_X1 port map( A1 => n3836, A2 => n113, ZN => n2194);
   U3105 : NOR3_X1 port map( A1 => n55, A2 => ADD_RS1(0), A3 => n3844, ZN => 
                           n3836);
   U3106 : OAI211_X1 port map( C1 => n548, C2 => n464, A => n3845, B => n3846, 
                           ZN => n3832);
   U3107 : OAI22_X1 port map( A1 => n644, A2 => n28, B1 => n2155, B2 => n476, 
                           ZN => n3847);
   U3108 : NAND2_X1 port map( A1 => n2, A2 => n3840, ZN => n2206);
   U3109 : NAND2_X1 port map( A1 => n3848, A2 => n3843, ZN => n2205);
   U3110 : AND2_X1 port map( A1 => n3839, A2 => n3837, ZN => n2203);
   U3111 : AND2_X1 port map( A1 => n3839, A2 => n113, ZN => n2202);
   U3112 : AOI22_X1 port map( A1 => n479, A2 => n4159, B1 => n482, B2 => n1078,
                           ZN => n3845);
   U3113 : AND2_X1 port map( A1 => n58, A2 => n3838, ZN => n2208);
   U3114 : AND2_X1 port map( A1 => n58, A2 => n3837, ZN => n2207);
   U3115 : NOR3_X1 port map( A1 => ADD_RS1(0), A2 => ADD_RS1(3), A3 => n56, ZN 
                           => n3848);
   U3116 : NAND2_X1 port map( A1 => n3839, A2 => n3838, ZN => n2199);
   U3117 : NOR3_X1 port map( A1 => n83, A2 => ADD_RS1(3), A3 => n55, ZN => 
                           n3839);
   U3118 : NAND4_X1 port map( A1 => n3849, A2 => n3850, A3 => n3851, A4 => 
                           n3852, ZN => n3831);
   U3119 : AOI221_X1 port map( B1 => n485, B2 => n4191, C1 => n488, C2 => n4223
                           , A => n3853, ZN => n3852);
   U3120 : OAI22_X1 port map( A1 => n420, A2 => n491, B1 => n388, B2 => n494, 
                           ZN => n3853);
   U3121 : NAND2_X1 port map( A1 => n3843, A2 => n3854, ZN => n2217);
   U3122 : NAND2_X1 port map( A1 => n113, A2 => n3855, ZN => n2216);
   U3123 : AND2_X1 port map( A1 => n36, A2 => n3840, ZN => n2214);
   U3124 : AND2_X1 port map( A1 => n3840, A2 => n3855, ZN => n2213);
   U3125 : AOI221_X1 port map( B1 => n497, B2 => n4255, C1 => n500, C2 => n4287
                           , A => n3856, ZN => n3851);
   U3126 : OAI22_X1 port map( A1 => n292, A2 => n503, B1 => n260, B2 => n25, ZN
                           => n3856);
   U3127 : NAND2_X1 port map( A1 => n3838, A2 => n3854, ZN => n2222);
   U3128 : NAND2_X1 port map( A1 => n3838, A2 => n3855, ZN => n2221);
   U3129 : AND2_X1 port map( A1 => n3837, A2 => n36, ZN => n2219);
   U3130 : NOR3_X1 port map( A1 => ADD_RS1(0), A2 => ADD_RS1(4), A3 => n3844, 
                           ZN => n3854);
   U3131 : AND2_X1 port map( A1 => n3837, A2 => n3855, ZN => n2218);
   U3132 : OAI22_X1 port map( A1 => n2166, A2 => n512, B1 => n2167, B2 => n515,
                           ZN => n3857);
   U3133 : NAND2_X1 port map( A1 => n3858, A2 => n3840, ZN => n2227);
   U3134 : NAND2_X1 port map( A1 => n3859, A2 => n3840, ZN => n2226);
   U3135 : AND2_X1 port map( A1 => n3, A2 => n113, ZN => n2224);
   U3136 : AND2_X1 port map( A1 => n3859, A2 => n113, ZN => n2223);
   U3137 : OAI22_X1 port map( A1 => n2171, A2 => n556, B1 => n2172, B2 => n559,
                           ZN => n3860);
   U3138 : NAND2_X1 port map( A1 => n3858, A2 => n3837, ZN => n2232);
   U3139 : NAND2_X1 port map( A1 => n3859, A2 => n3837, ZN => n2231);
   U3140 : AND2_X1 port map( A1 => ADD_RS1(1), A2 => n3861, ZN => n3837);
   U3141 : NOR3_X1 port map( A1 => ADD_RS1(3), A2 => ADD_RS1(4), A3 => 
                           ADD_RS1(0), ZN => n3859);
   U3142 : AND2_X1 port map( A1 => n3841, A2 => n113, ZN => n2229);
   U3143 : NOR2_X1 port map( A1 => n3861, A2 => ADD_RS1(1), ZN => n3843);
   U3144 : INV_X1 port map( A => ADD_RS1(2), ZN => n3861);
   U3145 : NOR3_X1 port map( A1 => n56, A2 => n84, A3 => n3844, ZN => n3841);
   U3146 : INV_X1 port map( A => ADD_RS1(3), ZN => n3844);
   U3147 : AND2_X1 port map( A1 => n3, A2 => n3838, ZN => n2228);
   U3148 : NOR2_X1 port map( A1 => ADD_RS1(1), A2 => n57, ZN => n3838);
   U3149 : NOR3_X1 port map( A1 => ADD_RS1(3), A2 => ADD_RS1(4), A3 => n84, ZN 
                           => n3858);
   U3150 : NAND2_X1 port map( A1 => n3862, A2 => n437, ZN => n2181);
   U3151 : AND3_X1 port map( A1 => n715, A2 => ENABLE, A3 => RD1, ZN => n2184);
   U3152 : INV_X1 port map( A => n3830, ZN => n3862);
   U3153 : NAND4_X1 port map( A1 => n3863, A2 => n3864, A3 => n3865, A4 => 
                           n3866, ZN => n3830);
   U3154 : NOR3_X1 port map( A1 => n3867, A2 => n1323, A3 => n3868, ZN => n3866
                           );
   U3155 : XNOR2_X1 port map( A => n1220, B => ADD_RS1(1), ZN => n3868);
   U3156 : INV_X1 port map( A => ADD_WR(1), ZN => n1220);
   U3157 : OAI21_X1 port map( B1 => n3869, B2 => n3870, A => WR, ZN => n1323);
   U3158 : NAND2_X1 port map( A1 => n873, A2 => n874, ZN => n3870);
   U3159 : INV_X1 port map( A => ADD_WR(4), ZN => n874);
   U3160 : INV_X1 port map( A => ADD_WR(3), ZN => n873);
   U3161 : INV_X1 port map( A => n910, ZN => n3869);
   U3162 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => ADD_WR(0),
                           ZN => n910);
   U3163 : XNOR2_X1 port map( A => ADD_RS1(0), B => n1186, ZN => n3867);
   U3164 : INV_X1 port map( A => ADD_WR(0), ZN => n1186);
   U3165 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS1(3), ZN => n3865);
   U3166 : XNOR2_X1 port map( A => ADD_WR(4), B => ADD_RS1(4), ZN => n3864);
   U3167 : XNOR2_X1 port map( A => n57, B => ADD_WR(2), ZN => n3863);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT5_0 is

   port( A, B : in std_logic_vector (4 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (4 downto 0));

end mux21_NBIT5_0;

architecture SYN_bhv of mux21_NBIT5_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8, n9, n10, n11, n1, n2, n3 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => S, Z => n1);
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : INV_X1 port map( A => n7, ZN => Z(4));
   U4 : AOI22_X1 port map( A1 => A(4), A2 => n3, B1 => n2, B2 => B(4), ZN => n7
                           );
   U5 : INV_X1 port map( A => n10, ZN => Z(1));
   U6 : INV_X1 port map( A => n9, ZN => Z(2));
   U7 : INV_X1 port map( A => n8, ZN => Z(3));
   U8 : AOI22_X1 port map( A1 => A(3), A2 => n3, B1 => B(3), B2 => n1, ZN => n8
                           );
   U9 : INV_X1 port map( A => n11, ZN => Z(0));
   U10 : AOI22_X1 port map( A1 => A(1), A2 => n3, B1 => B(1), B2 => n1, ZN => 
                           n10);
   U11 : AOI22_X1 port map( A1 => A(2), A2 => n3, B1 => B(2), B2 => n1, ZN => 
                           n9);
   U12 : AOI22_X1 port map( A1 => A(0), A2 => n3, B1 => B(0), B2 => n1, ZN => 
                           n11);
   U13 : INV_X1 port map( A => n2, ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N5_0 is

   port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in std_logic; 
         DOUT : out std_logic_vector (4 downto 0));

end regn_N5_0;

architecture SYN_bhv of regn_N5_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15 : 
      std_logic;

begin
   
   DOUT_reg_4_inst : DFFR_X1 port map( D => n15, CK => CLK, RN => RST, Q => 
                           DOUT(4), QN => n10);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n14, CK => CLK, RN => RST, Q => 
                           DOUT(3), QN => n9);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n13, CK => CLK, RN => RST, Q => 
                           DOUT(2), QN => n8);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n12, CK => CLK, RN => RST, Q => 
                           DOUT(1), QN => n7);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n11, CK => CLK, RN => RST, Q => 
                           DOUT(0), QN => n6);
   U2 : OAI21_X1 port map( B1 => n7, B2 => EN, A => n2, ZN => n12);
   U3 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n2);
   U4 : OAI21_X1 port map( B1 => n8, B2 => EN, A => n3, ZN => n13);
   U5 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n3);
   U6 : OAI21_X1 port map( B1 => n9, B2 => EN, A => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n4);
   U8 : OAI21_X1 port map( B1 => n10, B2 => EN, A => n5, ZN => n15);
   U9 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n5);
   U10 : OAI21_X1 port map( B1 => n6, B2 => EN, A => n1, ZN => n11);
   U11 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n1);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity instruction_decomposition is

   port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype : in
         std_logic;  ADD_RS1, ADD_RS2, ADD_WR : out std_logic_vector (4 downto 
         0);  IMM : out std_logic_vector (31 downto 0);  RD1, RD2 : out 
         std_logic);

end instruction_decomposition;

architecture SYN_bhv of instruction_decomposition is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal IMM_24_port, IMM_23_port, IMM_22_port, IMM_21_port, IMM_20_port, 
      IMM_19_port, IMM_18_port, IMM_17_port, IMM_16_port, IMM_15_port, 
      IMM_14_port, IMM_13_port, IMM_12_port, IMM_11_port, IMM_10_port, 
      IMM_9_port, IMM_8_port, IMM_7_port, IMM_6_port, IMM_5_port, IMM_4_port, 
      IMM_3_port, IMM_2_port, IMM_1_port, IMM_0_port, RD1_port, n25, n26, n27, 
      n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n1, n2, n3, n4, n5, n6,
      n7, IMM_31_port, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, 
      n20, n21, n22, n23, n24, n38, n39, n40, n41, n42 : std_logic;

begin
   IMM <= ( IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, 
      IMM_31_port, IMM_31_port, IMM_24_port, IMM_23_port, IMM_22_port, 
      IMM_21_port, IMM_20_port, IMM_19_port, IMM_18_port, IMM_17_port, 
      IMM_16_port, IMM_15_port, IMM_14_port, IMM_13_port, IMM_12_port, 
      IMM_11_port, IMM_10_port, IMM_9_port, IMM_8_port, IMM_7_port, IMM_6_port,
      IMM_5_port, IMM_4_port, IMM_3_port, IMM_2_port, IMM_1_port, IMM_0_port );
   RD1 <= RD1_port;
   
   U42 : NOR2_X2 port map( A1 => n5, A2 => n20, ZN => ADD_RS2(4));
   U44 : NOR2_X2 port map( A1 => n6, A2 => n22, ZN => ADD_RS2(2));
   U46 : NOR2_X2 port map( A1 => n3, A2 => n24, ZN => ADD_RS2(0));
   U54 : NOR2_X2 port map( A1 => n4, A2 => n19, ZN => ADD_RS1(0));
   U80 : NAND3_X1 port map( A1 => n11, A2 => INST_IN(26), A3 => INST_IN(30), ZN
                           => n34);
   U81 : XOR2_X1 port map( A => INST_IN(26), B => n15, Z => n36);
   U3 : AND2_X1 port map( A1 => n2, A2 => INST_IN(22), ZN => ADD_RS1(1));
   U4 : AND2_X1 port map( A1 => n2, A2 => INST_IN(24), ZN => ADD_RS1(3));
   U5 : AND2_X1 port map( A1 => n2, A2 => INST_IN(25), ZN => ADD_RS1(4));
   U6 : AND2_X2 port map( A1 => n13, A2 => n35, ZN => n3);
   U7 : CLKBUF_X1 port map( A => Itype, Z => n1);
   U8 : AND2_X1 port map( A1 => RD1_port, A2 => INST_IN(23), ZN => ADD_RS1(2));
   U9 : OR2_X1 port map( A1 => Rtype, A2 => Itype, ZN => n2);
   U10 : OR2_X1 port map( A1 => Rtype, A2 => Itype, ZN => RD1_port);
   U11 : AND2_X1 port map( A1 => n13, A2 => n35, ZN => n5);
   U12 : INV_X1 port map( A => n30, ZN => n12);
   U13 : INV_X1 port map( A => n31, ZN => n11);
   U14 : INV_X1 port map( A => Rtype, ZN => n13);
   U15 : OAI221_X1 port map( B1 => n31, B2 => n24, C1 => n42, C2 => n13, A => 
                           n7, ZN => ADD_WR(0));
   U16 : OAI221_X1 port map( B1 => n31, B2 => n23, C1 => n41, C2 => n13, A => 
                           n7, ZN => ADD_WR(1));
   U17 : OAI221_X1 port map( B1 => n31, B2 => n22, C1 => n40, C2 => n13, A => 
                           n7, ZN => ADD_WR(2));
   U18 : OAI221_X1 port map( B1 => n31, B2 => n21, C1 => n39, C2 => n13, A => 
                           n7, ZN => ADD_WR(3));
   U19 : OAI221_X1 port map( B1 => n31, B2 => n20, C1 => n38, C2 => n13, A => 
                           n7, ZN => ADD_WR(4));
   U20 : NAND2_X1 port map( A1 => n11, A2 => INST_IN(15), ZN => n29);
   U21 : INV_X1 port map( A => n25, ZN => IMM_31_port);
   U22 : OAI21_X1 port map( B1 => n26, B2 => n27, A => n13, ZN => n25);
   U23 : INV_X1 port map( A => n32, ZN => n7);
   U24 : OAI21_X1 port map( B1 => n33, B2 => n34, A => n28, ZN => n32);
   U25 : INV_X1 port map( A => INST_IN(16), ZN => n24);
   U26 : INV_X1 port map( A => INST_IN(20), ZN => n20);
   U27 : INV_X1 port map( A => INST_IN(18), ZN => n22);
   U28 : INV_X1 port map( A => INST_IN(15), ZN => n38);
   U29 : INV_X1 port map( A => INST_IN(19), ZN => n21);
   U30 : INV_X1 port map( A => INST_IN(17), ZN => n23);
   U31 : INV_X1 port map( A => INST_IN(21), ZN => n19);
   U32 : INV_X1 port map( A => INST_IN(11), ZN => n42);
   U33 : INV_X1 port map( A => INST_IN(12), ZN => n41);
   U34 : INV_X1 port map( A => INST_IN(13), ZN => n40);
   U35 : INV_X1 port map( A => INST_IN(14), ZN => n39);
   U36 : OAI21_X1 port map( B1 => n28, B2 => n24, A => n29, ZN => IMM_16_port);
   U37 : OAI21_X1 port map( B1 => n28, B2 => n23, A => n29, ZN => IMM_17_port);
   U38 : OAI21_X1 port map( B1 => n28, B2 => n22, A => n29, ZN => IMM_18_port);
   U39 : OAI21_X1 port map( B1 => n28, B2 => n21, A => n29, ZN => IMM_19_port);
   U40 : OAI21_X1 port map( B1 => n28, B2 => n20, A => n29, ZN => IMM_20_port);
   U41 : OAI21_X1 port map( B1 => n28, B2 => n19, A => n29, ZN => IMM_21_port);
   U43 : OAI21_X1 port map( B1 => n28, B2 => n18, A => n29, ZN => IMM_22_port);
   U45 : OAI21_X1 port map( B1 => n28, B2 => n17, A => n29, ZN => IMM_23_port);
   U47 : OAI21_X1 port map( B1 => n28, B2 => n16, A => n29, ZN => IMM_24_port);
   U48 : NOR2_X1 port map( A1 => n30, A2 => n42, ZN => IMM_11_port);
   U49 : NOR2_X1 port map( A1 => n30, A2 => n41, ZN => IMM_12_port);
   U50 : NOR2_X1 port map( A1 => n30, A2 => n40, ZN => IMM_13_port);
   U51 : NOR2_X1 port map( A1 => n30, A2 => n39, ZN => IMM_14_port);
   U52 : NOR2_X1 port map( A1 => n30, A2 => n38, ZN => IMM_15_port);
   U53 : AND2_X1 port map( A1 => INST_IN(1), A2 => n12, ZN => IMM_1_port);
   U55 : AND2_X1 port map( A1 => INST_IN(3), A2 => n12, ZN => IMM_3_port);
   U56 : AND2_X1 port map( A1 => INST_IN(2), A2 => n12, ZN => IMM_2_port);
   U57 : AND2_X1 port map( A1 => INST_IN(5), A2 => n12, ZN => IMM_5_port);
   U58 : AND2_X1 port map( A1 => INST_IN(4), A2 => n12, ZN => IMM_4_port);
   U59 : AND2_X1 port map( A1 => INST_IN(6), A2 => n12, ZN => IMM_6_port);
   U60 : AND2_X1 port map( A1 => INST_IN(7), A2 => n12, ZN => IMM_7_port);
   U61 : AND2_X1 port map( A1 => INST_IN(8), A2 => n12, ZN => IMM_8_port);
   U62 : AND2_X1 port map( A1 => INST_IN(9), A2 => n12, ZN => IMM_9_port);
   U63 : AND2_X1 port map( A1 => INST_IN(10), A2 => n12, ZN => IMM_10_port);
   U64 : AND2_X1 port map( A1 => INST_IN(0), A2 => n12, ZN => IMM_0_port);
   U65 : INV_X1 port map( A => INST_IN(23), ZN => n17);
   U66 : INV_X1 port map( A => n3, ZN => RD2);
   U67 : INV_X1 port map( A => RD1_port, ZN => n4);
   U68 : AND2_X1 port map( A1 => n13, A2 => n35, ZN => n6);
   U69 : INV_X1 port map( A => INST_IN(22), ZN => n18);
   U70 : NOR2_X1 port map( A1 => n5, A2 => n23, ZN => ADD_RS2(1));
   U71 : NOR2_X1 port map( A1 => n6, A2 => n21, ZN => ADD_RS2(3));
   U72 : INV_X1 port map( A => RD1_port, ZN => n9);
   U73 : INV_X1 port map( A => INST_IN(24), ZN => n16);
   U74 : NAND2_X1 port map( A1 => Jtype, A2 => n9, ZN => n28);
   U75 : NAND2_X1 port map( A1 => n1, A2 => n13, ZN => n31);
   U76 : OAI21_X1 port map( B1 => n1, B2 => Jtype, A => n13, ZN => n30);
   U77 : INV_X1 port map( A => INST_IN(29), ZN => n14);
   U78 : NOR2_X1 port map( A1 => n10, A2 => n38, ZN => n27);
   U79 : AND3_X1 port map( A1 => Jtype, A2 => n10, A3 => INST_IN(25), ZN => n26
                           );
   U82 : INV_X1 port map( A => n1, ZN => n10);
   U83 : INV_X1 port map( A => INST_IN(27), ZN => n15);
   U84 : NOR3_X1 port map( A1 => n14, A2 => INST_IN(30), A3 => INST_IN(28), ZN 
                           => n37);
   U85 : OR4_X1 port map( A1 => n15, A2 => INST_IN(28), A3 => INST_IN(29), A4 
                           => INST_IN(31), ZN => n33);
   U86 : NAND4_X1 port map( A1 => Itype, A2 => INST_IN(31), A3 => n36, A4 => 
                           n37, ZN => n35);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity instruction_type is

   port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype : 
         out std_logic);

end instruction_type;

architecture SYN_bhv of instruction_type is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, 
      n21, n1, n2, n3, n4, n5, n6, n22, n23, n24, n25, n26, n27, n28 : 
      std_logic;

begin
   
   U24 : OAI33_X1 port map( A1 => n15, A2 => n25, A3 => n11, B1 => n16, B2 => 
                           n1, B3 => INST_IN(28), ZN => n14);
   U1 : INV_X1 port map( A => n17, ZN => n23);
   U2 : NOR2_X1 port map( A1 => n7, A2 => n28, ZN => Rtype);
   U3 : NOR2_X1 port map( A1 => n27, A2 => n7, ZN => Jtype);
   U4 : INV_X1 port map( A => n25, ZN => n1);
   U5 : NOR2_X1 port map( A1 => INST_IN(27), A2 => INST_IN(26), ZN => n2);
   U6 : NOR2_X1 port map( A1 => INST_IN(27), A2 => INST_IN(26), ZN => n8);
   U7 : OR2_X1 port map( A1 => n9, A2 => n27, ZN => n3);
   U8 : OR2_X1 port map( A1 => n10, A2 => n11, ZN => n4);
   U9 : NAND3_X1 port map( A1 => n12, A2 => n4, A3 => n3, ZN => Itype);
   U10 : OR2_X1 port map( A1 => INST_IN(29), A2 => INST_IN(30), ZN => n5);
   U11 : NAND2_X1 port map( A1 => n5, A2 => n20, ZN => n18);
   U12 : CLKBUF_X1 port map( A => INST_IN(31), Z => n6);
   U13 : INV_X1 port map( A => n2, ZN => n28);
   U14 : INV_X1 port map( A => INST_IN(29), ZN => n26);
   U15 : NAND2_X1 port map( A1 => INST_IN(26), A2 => n27, ZN => n11);
   U16 : INV_X1 port map( A => INST_IN(30), ZN => n25);
   U17 : AOI21_X1 port map( B1 => INST_IN(26), B2 => INST_IN(27), A => n8, ZN 
                           => n16);
   U18 : INV_X1 port map( A => INST_IN(27), ZN => n27);
   U19 : AND2_X1 port map( A1 => INST_IN(28), A2 => INST_IN(30), ZN => n22);
   U20 : NOR2_X1 port map( A1 => n22, A2 => n20, ZN => n19);
   U21 : NAND2_X1 port map( A1 => INST_IN(29), A2 => INST_IN(28), ZN => n15);
   U22 : NAND4_X1 port map( A1 => INST_IN(30), A2 => INST_IN(28), A3 => n26, A4
                           => n24, ZN => n17);
   U23 : NAND2_X1 port map( A1 => n24, A2 => INST_IN(29), ZN => n20);
   U25 : NAND2_X1 port map( A1 => n10, A2 => n17, ZN => n13);
   U26 : NOR3_X1 port map( A1 => n21, A2 => n23, A3 => n19, ZN => n9);
   U27 : AOI211_X1 port map( C1 => n6, C2 => n26, A => n25, B => INST_IN(28), 
                           ZN => n21);
   U28 : OR4_X1 port map( A1 => INST_IN(28), A2 => INST_IN(29), A3 => n1, A4 =>
                           INST_IN(31), ZN => n7);
   U29 : AOI21_X1 port map( B1 => INST_IN(28), B2 => n18, A => n19, ZN => n10);
   U30 : INV_X1 port map( A => INST_IN(31), ZN => n24);
   U31 : AOI22_X1 port map( A1 => n13, A2 => n2, B1 => n6, B2 => n14, ZN => n12
                           );

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity regn_N32_0 is

   port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in std_logic;
         DOUT : out std_logic_vector (31 downto 0));

end regn_N32_0;

architecture SYN_bhv of regn_N32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DOUT_15_port, DOUT_14_port, DOUT_13_port, DOUT_12_port, DOUT_11_port,
      DOUT_10_port, DOUT_9_port, DOUT_8_port, DOUT_7_port, DOUT_6_port, 
      DOUT_5_port, DOUT_4_port, DOUT_3_port, DOUT_2_port, DOUT_1_port, 
      DOUT_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
      n15, n16, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, n93, n94, n95, n96, n17, n18, n19, DOUT_16_port, DOUT_17_port
      , DOUT_18_port, DOUT_19_port, DOUT_20_port, DOUT_21_port, DOUT_22_port, 
      DOUT_23_port, DOUT_24_port, DOUT_25_port, DOUT_26_port, DOUT_27_port, 
      DOUT_28_port, DOUT_29_port, DOUT_30_port, DOUT_31_port, n_1966, n_1967, 
      n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, 
      n_1977, n_1978, n_1979, n_1980, n_1981 : std_logic;

begin
   DOUT <= ( DOUT_31_port, DOUT_30_port, DOUT_29_port, DOUT_28_port, 
      DOUT_27_port, DOUT_26_port, DOUT_25_port, DOUT_24_port, DOUT_23_port, 
      DOUT_22_port, DOUT_21_port, DOUT_20_port, DOUT_19_port, DOUT_18_port, 
      DOUT_17_port, DOUT_16_port, DOUT_15_port, DOUT_14_port, DOUT_13_port, 
      DOUT_12_port, DOUT_11_port, DOUT_10_port, DOUT_9_port, DOUT_8_port, 
      DOUT_7_port, DOUT_6_port, DOUT_5_port, DOUT_4_port, DOUT_3_port, 
      DOUT_2_port, DOUT_1_port, DOUT_0_port );
   
   DOUT_reg_31_inst : DFFR_X1 port map( D => n96, CK => CLK, RN => n19, Q => 
                           DOUT_31_port, QN => n_1966);
   DOUT_reg_30_inst : DFFR_X1 port map( D => n95, CK => CLK, RN => n19, Q => 
                           DOUT_30_port, QN => n_1967);
   DOUT_reg_29_inst : DFFR_X1 port map( D => n94, CK => CLK, RN => n19, Q => 
                           DOUT_29_port, QN => n_1968);
   DOUT_reg_28_inst : DFFR_X1 port map( D => n93, CK => CLK, RN => n19, Q => 
                           DOUT_28_port, QN => n_1969);
   DOUT_reg_27_inst : DFFR_X1 port map( D => n92, CK => CLK, RN => n19, Q => 
                           DOUT_27_port, QN => n_1970);
   DOUT_reg_26_inst : DFFR_X1 port map( D => n91, CK => CLK, RN => n19, Q => 
                           DOUT_26_port, QN => n_1971);
   DOUT_reg_25_inst : DFFR_X1 port map( D => n90, CK => CLK, RN => n19, Q => 
                           DOUT_25_port, QN => n_1972);
   DOUT_reg_24_inst : DFFR_X1 port map( D => n89, CK => CLK, RN => n19, Q => 
                           DOUT_24_port, QN => n_1973);
   DOUT_reg_23_inst : DFFR_X1 port map( D => n88, CK => CLK, RN => n18, Q => 
                           DOUT_23_port, QN => n_1974);
   DOUT_reg_22_inst : DFFR_X1 port map( D => n87, CK => CLK, RN => n18, Q => 
                           DOUT_22_port, QN => n_1975);
   DOUT_reg_21_inst : DFFR_X1 port map( D => n86, CK => CLK, RN => n18, Q => 
                           DOUT_21_port, QN => n_1976);
   DOUT_reg_20_inst : DFFR_X1 port map( D => n85, CK => CLK, RN => n18, Q => 
                           DOUT_20_port, QN => n_1977);
   DOUT_reg_19_inst : DFFR_X1 port map( D => n84, CK => CLK, RN => n18, Q => 
                           DOUT_19_port, QN => n_1978);
   DOUT_reg_18_inst : DFFR_X1 port map( D => n83, CK => CLK, RN => n18, Q => 
                           DOUT_18_port, QN => n_1979);
   DOUT_reg_17_inst : DFFR_X1 port map( D => n82, CK => CLK, RN => n18, Q => 
                           DOUT_17_port, QN => n_1980);
   DOUT_reg_16_inst : DFFR_X1 port map( D => n81, CK => CLK, RN => n18, Q => 
                           DOUT_16_port, QN => n_1981);
   DOUT_reg_15_inst : DFFR_X1 port map( D => n80, CK => CLK, RN => n18, Q => 
                           DOUT_15_port, QN => n48);
   DOUT_reg_14_inst : DFFR_X1 port map( D => n79, CK => CLK, RN => n18, Q => 
                           DOUT_14_port, QN => n47);
   DOUT_reg_13_inst : DFFR_X1 port map( D => n78, CK => CLK, RN => n18, Q => 
                           DOUT_13_port, QN => n46);
   DOUT_reg_12_inst : DFFR_X1 port map( D => n77, CK => CLK, RN => n18, Q => 
                           DOUT_12_port, QN => n45);
   DOUT_reg_11_inst : DFFR_X1 port map( D => n76, CK => CLK, RN => n17, Q => 
                           DOUT_11_port, QN => n44);
   DOUT_reg_10_inst : DFFR_X1 port map( D => n75, CK => CLK, RN => n17, Q => 
                           DOUT_10_port, QN => n43);
   DOUT_reg_9_inst : DFFR_X1 port map( D => n74, CK => CLK, RN => n17, Q => 
                           DOUT_9_port, QN => n42);
   DOUT_reg_8_inst : DFFR_X1 port map( D => n73, CK => CLK, RN => n17, Q => 
                           DOUT_8_port, QN => n41);
   DOUT_reg_7_inst : DFFR_X1 port map( D => n72, CK => CLK, RN => n17, Q => 
                           DOUT_7_port, QN => n40);
   DOUT_reg_6_inst : DFFR_X1 port map( D => n71, CK => CLK, RN => n17, Q => 
                           DOUT_6_port, QN => n39);
   DOUT_reg_5_inst : DFFR_X1 port map( D => n70, CK => CLK, RN => n17, Q => 
                           DOUT_5_port, QN => n38);
   DOUT_reg_4_inst : DFFR_X1 port map( D => n69, CK => CLK, RN => n17, Q => 
                           DOUT_4_port, QN => n37);
   DOUT_reg_3_inst : DFFR_X1 port map( D => n68, CK => CLK, RN => n17, Q => 
                           DOUT_3_port, QN => n36);
   DOUT_reg_2_inst : DFFR_X1 port map( D => n67, CK => CLK, RN => n17, Q => 
                           DOUT_2_port, QN => n35);
   DOUT_reg_1_inst : DFFR_X1 port map( D => n66, CK => CLK, RN => n17, Q => 
                           DOUT_1_port, QN => n34);
   DOUT_reg_0_inst : DFFR_X1 port map( D => n65, CK => CLK, RN => n17, Q => 
                           DOUT_0_port, QN => n33);
   U2 : BUF_X1 port map( A => RST, Z => n17);
   U3 : BUF_X1 port map( A => RST, Z => n18);
   U4 : BUF_X1 port map( A => RST, Z => n19);
   U5 : OAI21_X1 port map( B1 => n44, B2 => EN, A => n12, ZN => n76);
   U6 : NAND2_X1 port map( A1 => DIN(11), A2 => EN, ZN => n12);
   U7 : OAI21_X1 port map( B1 => n46, B2 => EN, A => n14, ZN => n78);
   U8 : NAND2_X1 port map( A1 => DIN(13), A2 => EN, ZN => n14);
   U9 : OAI21_X1 port map( B1 => n47, B2 => EN, A => n15, ZN => n79);
   U10 : NAND2_X1 port map( A1 => DIN(14), A2 => EN, ZN => n15);
   U11 : OAI21_X1 port map( B1 => n34, B2 => EN, A => n2, ZN => n66);
   U12 : NAND2_X1 port map( A1 => DIN(1), A2 => EN, ZN => n2);
   U13 : OAI21_X1 port map( B1 => n35, B2 => EN, A => n3, ZN => n67);
   U14 : NAND2_X1 port map( A1 => DIN(2), A2 => EN, ZN => n3);
   U15 : OAI21_X1 port map( B1 => n36, B2 => EN, A => n4, ZN => n68);
   U16 : NAND2_X1 port map( A1 => DIN(3), A2 => EN, ZN => n4);
   U17 : OAI21_X1 port map( B1 => n37, B2 => EN, A => n5, ZN => n69);
   U18 : NAND2_X1 port map( A1 => DIN(4), A2 => EN, ZN => n5);
   U19 : OAI21_X1 port map( B1 => n38, B2 => EN, A => n6, ZN => n70);
   U20 : NAND2_X1 port map( A1 => DIN(5), A2 => EN, ZN => n6);
   U21 : OAI21_X1 port map( B1 => n39, B2 => EN, A => n7, ZN => n71);
   U22 : NAND2_X1 port map( A1 => DIN(6), A2 => EN, ZN => n7);
   U23 : OAI21_X1 port map( B1 => n41, B2 => EN, A => n9, ZN => n73);
   U24 : NAND2_X1 port map( A1 => DIN(8), A2 => EN, ZN => n9);
   U25 : OAI21_X1 port map( B1 => n43, B2 => EN, A => n11, ZN => n75);
   U26 : NAND2_X1 port map( A1 => DIN(10), A2 => EN, ZN => n11);
   U27 : OAI21_X1 port map( B1 => n45, B2 => EN, A => n13, ZN => n77);
   U28 : NAND2_X1 port map( A1 => DIN(12), A2 => EN, ZN => n13);
   U29 : OAI21_X1 port map( B1 => n42, B2 => EN, A => n10, ZN => n74);
   U30 : NAND2_X1 port map( A1 => DIN(9), A2 => EN, ZN => n10);
   U31 : OAI21_X1 port map( B1 => n33, B2 => EN, A => n1, ZN => n65);
   U32 : NAND2_X1 port map( A1 => EN, A2 => DIN(0), ZN => n1);
   U33 : OAI21_X1 port map( B1 => n48, B2 => EN, A => n16, ZN => n80);
   U34 : NAND2_X1 port map( A1 => DIN(15), A2 => EN, ZN => n16);
   U35 : NAND2_X1 port map( A1 => DIN(7), A2 => EN, ZN => n8);
   U36 : OAI21_X1 port map( B1 => n40, B2 => EN, A => n8, ZN => n72);
   U37 : MUX2_X1 port map( A => DOUT_16_port, B => DIN(16), S => EN, Z => n81);
   U38 : MUX2_X1 port map( A => DOUT_17_port, B => DIN(17), S => EN, Z => n82);
   U39 : MUX2_X1 port map( A => DOUT_18_port, B => DIN(18), S => EN, Z => n83);
   U40 : MUX2_X1 port map( A => DOUT_19_port, B => DIN(19), S => EN, Z => n84);
   U41 : MUX2_X1 port map( A => DOUT_20_port, B => DIN(20), S => EN, Z => n85);
   U42 : MUX2_X1 port map( A => DOUT_21_port, B => DIN(21), S => EN, Z => n86);
   U43 : MUX2_X1 port map( A => DOUT_22_port, B => DIN(22), S => EN, Z => n87);
   U44 : MUX2_X1 port map( A => DOUT_23_port, B => DIN(23), S => EN, Z => n88);
   U45 : MUX2_X1 port map( A => DOUT_24_port, B => DIN(24), S => EN, Z => n89);
   U46 : MUX2_X1 port map( A => DOUT_25_port, B => DIN(25), S => EN, Z => n90);
   U47 : MUX2_X1 port map( A => DOUT_26_port, B => DIN(26), S => EN, Z => n91);
   U48 : MUX2_X1 port map( A => DOUT_27_port, B => DIN(27), S => EN, Z => n92);
   U49 : MUX2_X1 port map( A => DOUT_28_port, B => DIN(28), S => EN, Z => n93);
   U50 : MUX2_X1 port map( A => DOUT_29_port, B => DIN(29), S => EN, Z => n94);
   U51 : MUX2_X1 port map( A => DOUT_30_port, B => DIN(30), S => EN, Z => n95);
   U52 : MUX2_X1 port map( A => DOUT_31_port, B => DIN(31), S => EN, Z => n96);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity mux21_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : out 
         std_logic_vector (31 downto 0));

end mux21_NBIT32_0;

architecture SYN_bhv of mux21_NBIT32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n43, n54, n59, n60, n61, n62, n63,
      n64, n65, n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => n2);
   U2 : INV_X1 port map( A => n7, ZN => n1);
   U3 : BUF_X1 port map( A => n8, Z => n5);
   U4 : BUF_X1 port map( A => n8, Z => n6);
   U5 : BUF_X1 port map( A => n8, Z => n3);
   U6 : BUF_X1 port map( A => n8, Z => n4);
   U7 : BUF_X1 port map( A => n8, Z => n7);
   U8 : INV_X1 port map( A => S, ZN => n8);
   U9 : INV_X1 port map( A => n63, ZN => Z(11));
   U10 : AOI22_X1 port map( A1 => A(11), A2 => n3, B1 => B(11), B2 => n2, ZN =>
                           n63);
   U11 : INV_X1 port map( A => n61, ZN => Z(13));
   U12 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => B(13), B2 => n1, ZN =>
                           n61);
   U13 : INV_X1 port map( A => n60, ZN => Z(14));
   U14 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => B(14), B2 => n1, ZN =>
                           n60);
   U15 : INV_X1 port map( A => n54, ZN => Z(1));
   U16 : AOI22_X1 port map( A1 => A(1), A2 => n4, B1 => B(1), B2 => n1, ZN => 
                           n54);
   U17 : INV_X1 port map( A => n43, ZN => Z(2));
   U18 : AOI22_X1 port map( A1 => A(2), A2 => n5, B1 => B(2), B2 => n1, ZN => 
                           n43);
   U19 : INV_X1 port map( A => n40, ZN => Z(3));
   U20 : AOI22_X1 port map( A1 => A(3), A2 => n5, B1 => B(3), B2 => n1, ZN => 
                           n40);
   U21 : INV_X1 port map( A => n39, ZN => Z(4));
   U22 : AOI22_X1 port map( A1 => A(4), A2 => n5, B1 => B(4), B2 => n1, ZN => 
                           n39);
   U23 : INV_X1 port map( A => n38, ZN => Z(5));
   U24 : AOI22_X1 port map( A1 => A(5), A2 => n5, B1 => B(5), B2 => n1, ZN => 
                           n38);
   U25 : INV_X1 port map( A => n37, ZN => Z(6));
   U26 : AOI22_X1 port map( A1 => A(6), A2 => n6, B1 => B(6), B2 => n1, ZN => 
                           n37);
   U27 : INV_X1 port map( A => n35, ZN => Z(8));
   U28 : AOI22_X1 port map( A1 => A(8), A2 => n6, B1 => B(8), B2 => n1, ZN => 
                           n35);
   U29 : INV_X1 port map( A => n64, ZN => Z(10));
   U30 : AOI22_X1 port map( A1 => A(10), A2 => n3, B1 => B(10), B2 => n2, ZN =>
                           n64);
   U31 : INV_X1 port map( A => n62, ZN => Z(12));
   U32 : AOI22_X1 port map( A1 => A(12), A2 => n3, B1 => B(12), B2 => n1, ZN =>
                           n62);
   U33 : INV_X1 port map( A => n34, ZN => Z(9));
   U34 : AOI22_X1 port map( A1 => A(9), A2 => n6, B1 => n2, B2 => B(9), ZN => 
                           n34);
   U35 : INV_X1 port map( A => n65, ZN => Z(0));
   U36 : AOI22_X1 port map( A1 => A(0), A2 => n3, B1 => B(0), B2 => n2, ZN => 
                           n65);
   U37 : INV_X1 port map( A => n59, ZN => Z(15));
   U38 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => B(15), B2 => n1, ZN =>
                           n59);
   U39 : INV_X1 port map( A => n36, ZN => Z(7));
   U40 : AOI22_X1 port map( A1 => A(7), A2 => n6, B1 => B(7), B2 => n1, ZN => 
                           n36);
   U41 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Z(16));
   U42 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Z(17));
   U43 : MUX2_X1 port map( A => A(18), B => B(18), S => n1, Z => Z(18));
   U44 : MUX2_X1 port map( A => A(19), B => B(19), S => S, Z => Z(19));
   U45 : MUX2_X1 port map( A => A(20), B => B(20), S => S, Z => Z(20));
   U46 : MUX2_X1 port map( A => A(21), B => B(21), S => S, Z => Z(21));
   U47 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Z(22));
   U48 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Z(23));
   U49 : MUX2_X1 port map( A => A(24), B => B(24), S => n2, Z => Z(24));
   U50 : MUX2_X1 port map( A => A(25), B => B(25), S => n2, Z => Z(25));
   U51 : MUX2_X1 port map( A => A(26), B => B(26), S => n2, Z => Z(26));
   U52 : MUX2_X1 port map( A => A(27), B => B(27), S => n2, Z => Z(27));
   U53 : MUX2_X1 port map( A => A(28), B => B(28), S => n2, Z => Z(28));
   U54 : MUX2_X1 port map( A => A(29), B => B(29), S => n2, Z => Z(29));
   U55 : MUX2_X1 port map( A => A(30), B => B(30), S => n2, Z => Z(30));
   U56 : MUX2_X1 port map( A => A(31), B => B(31), S => n2, Z => Z(31));

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity HazardDetection is

   port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : in std_logic_vector (4
         downto 0);  DRAM_R : in std_logic;  INS_IN, PC_IN : in 
         std_logic_vector (31 downto 0);  Bubble : out std_logic;  HDU_INS_OUT,
         HDU_PC_OUT, HDU_NPC_OUT : out std_logic_vector (31 downto 0));

end HazardDetection;

architecture SYN_arch of HazardDetection is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component HazardDetection_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n7, n8, n11, n1, n2, n3, n4, n5, n6, n9, n10, n12, n13, n14, n15, n16
      , n_1982 : std_logic;

begin
   HDU_INS_OUT <= ( INS_IN(31), INS_IN(30), INS_IN(29), INS_IN(28), INS_IN(27),
      INS_IN(26), INS_IN(25), INS_IN(24), INS_IN(23), INS_IN(22), INS_IN(21), 
      INS_IN(20), INS_IN(19), INS_IN(18), INS_IN(17), INS_IN(16), INS_IN(15), 
      INS_IN(14), INS_IN(13), INS_IN(12), INS_IN(11), INS_IN(10), INS_IN(9), 
      INS_IN(8), INS_IN(7), INS_IN(6), INS_IN(5), INS_IN(4), INS_IN(3), 
      INS_IN(2), INS_IN(1), INS_IN(0) );
   HDU_PC_OUT <= ( PC_IN(31), PC_IN(30), PC_IN(29), PC_IN(28), PC_IN(27), 
      PC_IN(26), PC_IN(25), PC_IN(24), PC_IN(23), PC_IN(22), PC_IN(21), 
      PC_IN(20), PC_IN(19), PC_IN(18), PC_IN(17), PC_IN(16), PC_IN(15), 
      PC_IN(14), PC_IN(13), PC_IN(12), PC_IN(11), PC_IN(10), PC_IN(9), PC_IN(8)
      , PC_IN(7), PC_IN(6), PC_IN(5), PC_IN(4), PC_IN(3), PC_IN(2), PC_IN(1), 
      PC_IN(0) );
   
   n7 <= '0';
   n8 <= '1';
   n11 <= '0';
   add_32 : HazardDetection_DW01_add_0 port map( A(31) => PC_IN(31), A(30) => 
                           PC_IN(30), A(29) => PC_IN(29), A(28) => PC_IN(28), 
                           A(27) => PC_IN(27), A(26) => PC_IN(26), A(25) => 
                           PC_IN(25), A(24) => PC_IN(24), A(23) => PC_IN(23), 
                           A(22) => PC_IN(22), A(21) => PC_IN(21), A(20) => 
                           PC_IN(20), A(19) => PC_IN(19), A(18) => PC_IN(18), 
                           A(17) => PC_IN(17), A(16) => PC_IN(16), A(15) => 
                           PC_IN(15), A(14) => PC_IN(14), A(13) => PC_IN(13), 
                           A(12) => PC_IN(12), A(11) => PC_IN(11), A(10) => 
                           PC_IN(10), A(9) => PC_IN(9), A(8) => PC_IN(8), A(7) 
                           => PC_IN(7), A(6) => PC_IN(6), A(5) => PC_IN(5), 
                           A(4) => PC_IN(4), A(3) => PC_IN(3), A(2) => PC_IN(2)
                           , A(1) => PC_IN(1), A(0) => PC_IN(0), B(31) => n7, 
                           B(30) => n7, B(29) => n7, B(28) => n7, B(27) => n7, 
                           B(26) => n7, B(25) => n7, B(24) => n7, B(23) => n7, 
                           B(22) => n7, B(21) => n7, B(20) => n7, B(19) => n7, 
                           B(18) => n7, B(17) => n7, B(16) => n7, B(15) => n7, 
                           B(14) => n7, B(13) => n7, B(12) => n7, B(11) => n7, 
                           B(10) => n7, B(9) => n7, B(8) => n7, B(7) => n7, 
                           B(6) => n7, B(5) => n7, B(4) => n7, B(3) => n7, B(2)
                           => n8, B(1) => n7, B(0) => n7, CI => n11, SUM(31) =>
                           HDU_NPC_OUT(31), SUM(30) => HDU_NPC_OUT(30), SUM(29)
                           => HDU_NPC_OUT(29), SUM(28) => HDU_NPC_OUT(28), 
                           SUM(27) => HDU_NPC_OUT(27), SUM(26) => 
                           HDU_NPC_OUT(26), SUM(25) => HDU_NPC_OUT(25), SUM(24)
                           => HDU_NPC_OUT(24), SUM(23) => HDU_NPC_OUT(23), 
                           SUM(22) => HDU_NPC_OUT(22), SUM(21) => 
                           HDU_NPC_OUT(21), SUM(20) => HDU_NPC_OUT(20), SUM(19)
                           => HDU_NPC_OUT(19), SUM(18) => HDU_NPC_OUT(18), 
                           SUM(17) => HDU_NPC_OUT(17), SUM(16) => 
                           HDU_NPC_OUT(16), SUM(15) => HDU_NPC_OUT(15), SUM(14)
                           => HDU_NPC_OUT(14), SUM(13) => HDU_NPC_OUT(13), 
                           SUM(12) => HDU_NPC_OUT(12), SUM(11) => 
                           HDU_NPC_OUT(11), SUM(10) => HDU_NPC_OUT(10), SUM(9) 
                           => HDU_NPC_OUT(9), SUM(8) => HDU_NPC_OUT(8), SUM(7) 
                           => HDU_NPC_OUT(7), SUM(6) => HDU_NPC_OUT(6), SUM(5) 
                           => HDU_NPC_OUT(5), SUM(4) => HDU_NPC_OUT(4), SUM(3) 
                           => HDU_NPC_OUT(3), SUM(2) => HDU_NPC_OUT(2), SUM(1) 
                           => HDU_NPC_OUT(1), SUM(0) => HDU_NPC_OUT(0), CO => 
                           n_1982);
   U4 : AND3_X1 port map( A1 => DRAM_R, A2 => n1, A3 => RST, ZN => Bubble);
   U5 : OAI33_X1 port map( A1 => n2, A2 => n3, A3 => n4, B1 => n5, B2 => n6, B3
                           => n9, ZN => n1);
   U6 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RS2(4), Z => n9);
   U8 : XOR2_X1 port map( A => ADD_WR(2), B => ADD_RS2(2), Z => n6);
   U9 : NAND3_X1 port map( A1 => n10, A2 => n12, A3 => n13, ZN => n5);
   U11 : XNOR2_X1 port map( A => ADD_WR(0), B => ADD_RS2(0), ZN => n13);
   U12 : XNOR2_X1 port map( A => ADD_WR(1), B => ADD_RS2(1), ZN => n12);
   U13 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS2(3), ZN => n10);
   U14 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RS1(4), Z => n4);
   U15 : XOR2_X1 port map( A => ADD_WR(2), B => ADD_RS1(2), Z => n3);
   U16 : NAND3_X1 port map( A1 => n14, A2 => n15, A3 => n16, ZN => n2);
   U17 : XNOR2_X1 port map( A => ADD_WR(0), B => ADD_RS1(0), ZN => n16);
   U18 : XNOR2_X1 port map( A => ADD_WR(1), B => ADD_RS1(1), ZN => n15);
   U19 : XNOR2_X1 port map( A => ADD_WR(3), B => ADD_RS1(3), ZN => n14);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Writeback is

   port( WB_MUX_SEL : in std_logic;  DATA_IN, ALU_RES_IN : in std_logic_vector 
         (31 downto 0);  ADD_WR_IN : in std_logic_vector (4 downto 0);  
         DATA_OUT : out std_logic_vector (31 downto 0);  ADD_WR_OUT : out 
         std_logic_vector (4 downto 0));

end Writeback;

architecture SYN_struct of Writeback is

   component mux21_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;

begin
   ADD_WR_OUT <= ( ADD_WR_IN(4), ADD_WR_IN(3), ADD_WR_IN(2), ADD_WR_IN(1), 
      ADD_WR_IN(0) );
   
   WBmux : mux21_NBIT32_3 port map( A(31) => ALU_RES_IN(31), A(30) => 
                           ALU_RES_IN(30), A(29) => ALU_RES_IN(29), A(28) => 
                           ALU_RES_IN(28), A(27) => ALU_RES_IN(27), A(26) => 
                           ALU_RES_IN(26), A(25) => ALU_RES_IN(25), A(24) => 
                           ALU_RES_IN(24), A(23) => ALU_RES_IN(23), A(22) => 
                           ALU_RES_IN(22), A(21) => ALU_RES_IN(21), A(20) => 
                           ALU_RES_IN(20), A(19) => ALU_RES_IN(19), A(18) => 
                           ALU_RES_IN(18), A(17) => ALU_RES_IN(17), A(16) => 
                           ALU_RES_IN(16), A(15) => ALU_RES_IN(15), A(14) => 
                           ALU_RES_IN(14), A(13) => ALU_RES_IN(13), A(12) => 
                           ALU_RES_IN(12), A(11) => ALU_RES_IN(11), A(10) => 
                           ALU_RES_IN(10), A(9) => ALU_RES_IN(9), A(8) => 
                           ALU_RES_IN(8), A(7) => ALU_RES_IN(7), A(6) => 
                           ALU_RES_IN(6), A(5) => ALU_RES_IN(5), A(4) => 
                           ALU_RES_IN(4), A(3) => ALU_RES_IN(3), A(2) => 
                           ALU_RES_IN(2), A(1) => ALU_RES_IN(1), A(0) => 
                           ALU_RES_IN(0), B(31) => DATA_IN(31), B(30) => 
                           DATA_IN(30), B(29) => DATA_IN(29), B(28) => 
                           DATA_IN(28), B(27) => DATA_IN(27), B(26) => 
                           DATA_IN(26), B(25) => DATA_IN(25), B(24) => 
                           DATA_IN(24), B(23) => DATA_IN(23), B(22) => 
                           DATA_IN(22), B(21) => DATA_IN(21), B(20) => 
                           DATA_IN(20), B(19) => DATA_IN(19), B(18) => 
                           DATA_IN(18), B(17) => DATA_IN(17), B(16) => 
                           DATA_IN(16), B(15) => DATA_IN(15), B(14) => 
                           DATA_IN(14), B(13) => DATA_IN(13), B(12) => 
                           DATA_IN(12), B(11) => DATA_IN(11), B(10) => 
                           DATA_IN(10), B(9) => DATA_IN(9), B(8) => DATA_IN(8),
                           B(7) => DATA_IN(7), B(6) => DATA_IN(6), B(5) => 
                           DATA_IN(5), B(4) => DATA_IN(4), B(3) => DATA_IN(3), 
                           B(2) => DATA_IN(2), B(1) => DATA_IN(1), B(0) => 
                           DATA_IN(0), S => WB_MUX_SEL, Z(31) => DATA_OUT(31), 
                           Z(30) => DATA_OUT(30), Z(29) => DATA_OUT(29), Z(28) 
                           => DATA_OUT(28), Z(27) => DATA_OUT(27), Z(26) => 
                           DATA_OUT(26), Z(25) => DATA_OUT(25), Z(24) => 
                           DATA_OUT(24), Z(23) => DATA_OUT(23), Z(22) => 
                           DATA_OUT(22), Z(21) => DATA_OUT(21), Z(20) => 
                           DATA_OUT(20), Z(19) => DATA_OUT(19), Z(18) => 
                           DATA_OUT(18), Z(17) => DATA_OUT(17), Z(16) => 
                           DATA_OUT(16), Z(15) => DATA_OUT(15), Z(14) => 
                           DATA_OUT(14), Z(13) => DATA_OUT(13), Z(12) => 
                           DATA_OUT(12), Z(11) => DATA_OUT(11), Z(10) => 
                           DATA_OUT(10), Z(9) => DATA_OUT(9), Z(8) => 
                           DATA_OUT(8), Z(7) => DATA_OUT(7), Z(6) => 
                           DATA_OUT(6), Z(5) => DATA_OUT(5), Z(4) => 
                           DATA_OUT(4), Z(3) => DATA_OUT(3), Z(2) => 
                           DATA_OUT(2), Z(1) => DATA_OUT(1), Z(0) => 
                           DATA_OUT(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Memory is

   port( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN : in std_logic;  PC_SEL : in
         std_logic_vector (1 downto 0);  NPC_IN, NPC_ABS, NPC_REL, ALU_RES_IN, 
         B_IN : in std_logic_vector (31 downto 0);  ADD_WR_IN : in 
         std_logic_vector (4 downto 0);  DRAM_DATA_IN : in std_logic_vector (31
         downto 0);  LOAD_TYPE_IN : in std_logic_vector (1 downto 0);  
         STORE_TYPE_IN : in std_logic;  PC_OUT : out std_logic_vector (31 
         downto 0);  DRAM_R_OUT, DRAM_W_OUT : out std_logic;  DRAM_ADDR_OUT, 
         DRAM_DATA_OUT, DATA_OUT, ALU_RES_OUT, OP_MEM : out std_logic_vector 
         (31 downto 0);  ADD_WR_MEM, ADD_WR_OUT : out std_logic_vector (4 
         downto 0);  LOAD_TYPE_OUT : out std_logic_vector (1 downto 0);  
         STORE_TYPE_OUT : out std_logic);

end Memory;

architecture SYN_struct of Memory is

   component mux41_NBIT32_2
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component regn_N32_1
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N5_1
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   signal X_Logic0_port : std_logic;

begin
   DRAM_R_OUT <= DRAM_R_IN;
   DRAM_W_OUT <= DRAM_W_IN;
   DRAM_ADDR_OUT <= ( ALU_RES_IN(31), ALU_RES_IN(30), ALU_RES_IN(29), 
      ALU_RES_IN(28), ALU_RES_IN(27), ALU_RES_IN(26), ALU_RES_IN(25), 
      ALU_RES_IN(24), ALU_RES_IN(23), ALU_RES_IN(22), ALU_RES_IN(21), 
      ALU_RES_IN(20), ALU_RES_IN(19), ALU_RES_IN(18), ALU_RES_IN(17), 
      ALU_RES_IN(16), ALU_RES_IN(15), ALU_RES_IN(14), ALU_RES_IN(13), 
      ALU_RES_IN(12), ALU_RES_IN(11), ALU_RES_IN(10), ALU_RES_IN(9), 
      ALU_RES_IN(8), ALU_RES_IN(7), ALU_RES_IN(6), ALU_RES_IN(5), ALU_RES_IN(4)
      , ALU_RES_IN(3), ALU_RES_IN(2), ALU_RES_IN(1), ALU_RES_IN(0) );
   DRAM_DATA_OUT <= ( B_IN(31), B_IN(30), B_IN(29), B_IN(28), B_IN(27), 
      B_IN(26), B_IN(25), B_IN(24), B_IN(23), B_IN(22), B_IN(21), B_IN(20), 
      B_IN(19), B_IN(18), B_IN(17), B_IN(16), B_IN(15), B_IN(14), B_IN(13), 
      B_IN(12), B_IN(11), B_IN(10), B_IN(9), B_IN(8), B_IN(7), B_IN(6), B_IN(5)
      , B_IN(4), B_IN(3), B_IN(2), B_IN(1), B_IN(0) );
   DATA_OUT <= ( DRAM_DATA_IN(31), DRAM_DATA_IN(30), DRAM_DATA_IN(29), 
      DRAM_DATA_IN(28), DRAM_DATA_IN(27), DRAM_DATA_IN(26), DRAM_DATA_IN(25), 
      DRAM_DATA_IN(24), DRAM_DATA_IN(23), DRAM_DATA_IN(22), DRAM_DATA_IN(21), 
      DRAM_DATA_IN(20), DRAM_DATA_IN(19), DRAM_DATA_IN(18), DRAM_DATA_IN(17), 
      DRAM_DATA_IN(16), DRAM_DATA_IN(15), DRAM_DATA_IN(14), DRAM_DATA_IN(13), 
      DRAM_DATA_IN(12), DRAM_DATA_IN(11), DRAM_DATA_IN(10), DRAM_DATA_IN(9), 
      DRAM_DATA_IN(8), DRAM_DATA_IN(7), DRAM_DATA_IN(6), DRAM_DATA_IN(5), 
      DRAM_DATA_IN(4), DRAM_DATA_IN(3), DRAM_DATA_IN(2), DRAM_DATA_IN(1), 
      DRAM_DATA_IN(0) );
   OP_MEM <= ( ALU_RES_IN(31), ALU_RES_IN(30), ALU_RES_IN(29), ALU_RES_IN(28), 
      ALU_RES_IN(27), ALU_RES_IN(26), ALU_RES_IN(25), ALU_RES_IN(24), 
      ALU_RES_IN(23), ALU_RES_IN(22), ALU_RES_IN(21), ALU_RES_IN(20), 
      ALU_RES_IN(19), ALU_RES_IN(18), ALU_RES_IN(17), ALU_RES_IN(16), 
      ALU_RES_IN(15), ALU_RES_IN(14), ALU_RES_IN(13), ALU_RES_IN(12), 
      ALU_RES_IN(11), ALU_RES_IN(10), ALU_RES_IN(9), ALU_RES_IN(8), 
      ALU_RES_IN(7), ALU_RES_IN(6), ALU_RES_IN(5), ALU_RES_IN(4), ALU_RES_IN(3)
      , ALU_RES_IN(2), ALU_RES_IN(1), ALU_RES_IN(0) );
   ADD_WR_MEM <= ( ADD_WR_IN(4), ADD_WR_IN(3), ADD_WR_IN(2), ADD_WR_IN(1), 
      ADD_WR_IN(0) );
   LOAD_TYPE_OUT <= ( LOAD_TYPE_IN(1), LOAD_TYPE_IN(0) );
   STORE_TYPE_OUT <= STORE_TYPE_IN;
   
   X_Logic0_port <= '0';
   reg0 : regn_N5_1 port map( DIN(4) => ADD_WR_IN(4), DIN(3) => ADD_WR_IN(3), 
                           DIN(2) => ADD_WR_IN(2), DIN(1) => ADD_WR_IN(1), 
                           DIN(0) => ADD_WR_IN(0), CLK => CLK, EN => MEM_EN_IN,
                           RST => RST, DOUT(4) => ADD_WR_OUT(4), DOUT(3) => 
                           ADD_WR_OUT(3), DOUT(2) => ADD_WR_OUT(2), DOUT(1) => 
                           ADD_WR_OUT(1), DOUT(0) => ADD_WR_OUT(0));
   reg1 : regn_N32_1 port map( DIN(31) => ALU_RES_IN(31), DIN(30) => 
                           ALU_RES_IN(30), DIN(29) => ALU_RES_IN(29), DIN(28) 
                           => ALU_RES_IN(28), DIN(27) => ALU_RES_IN(27), 
                           DIN(26) => ALU_RES_IN(26), DIN(25) => ALU_RES_IN(25)
                           , DIN(24) => ALU_RES_IN(24), DIN(23) => 
                           ALU_RES_IN(23), DIN(22) => ALU_RES_IN(22), DIN(21) 
                           => ALU_RES_IN(21), DIN(20) => ALU_RES_IN(20), 
                           DIN(19) => ALU_RES_IN(19), DIN(18) => ALU_RES_IN(18)
                           , DIN(17) => ALU_RES_IN(17), DIN(16) => 
                           ALU_RES_IN(16), DIN(15) => ALU_RES_IN(15), DIN(14) 
                           => ALU_RES_IN(14), DIN(13) => ALU_RES_IN(13), 
                           DIN(12) => ALU_RES_IN(12), DIN(11) => ALU_RES_IN(11)
                           , DIN(10) => ALU_RES_IN(10), DIN(9) => ALU_RES_IN(9)
                           , DIN(8) => ALU_RES_IN(8), DIN(7) => ALU_RES_IN(7), 
                           DIN(6) => ALU_RES_IN(6), DIN(5) => ALU_RES_IN(5), 
                           DIN(4) => ALU_RES_IN(4), DIN(3) => ALU_RES_IN(3), 
                           DIN(2) => ALU_RES_IN(2), DIN(1) => ALU_RES_IN(1), 
                           DIN(0) => ALU_RES_IN(0), CLK => CLK, EN => MEM_EN_IN
                           , RST => RST, DOUT(31) => ALU_RES_OUT(31), DOUT(30) 
                           => ALU_RES_OUT(30), DOUT(29) => ALU_RES_OUT(29), 
                           DOUT(28) => ALU_RES_OUT(28), DOUT(27) => 
                           ALU_RES_OUT(27), DOUT(26) => ALU_RES_OUT(26), 
                           DOUT(25) => ALU_RES_OUT(25), DOUT(24) => 
                           ALU_RES_OUT(24), DOUT(23) => ALU_RES_OUT(23), 
                           DOUT(22) => ALU_RES_OUT(22), DOUT(21) => 
                           ALU_RES_OUT(21), DOUT(20) => ALU_RES_OUT(20), 
                           DOUT(19) => ALU_RES_OUT(19), DOUT(18) => 
                           ALU_RES_OUT(18), DOUT(17) => ALU_RES_OUT(17), 
                           DOUT(16) => ALU_RES_OUT(16), DOUT(15) => 
                           ALU_RES_OUT(15), DOUT(14) => ALU_RES_OUT(14), 
                           DOUT(13) => ALU_RES_OUT(13), DOUT(12) => 
                           ALU_RES_OUT(12), DOUT(11) => ALU_RES_OUT(11), 
                           DOUT(10) => ALU_RES_OUT(10), DOUT(9) => 
                           ALU_RES_OUT(9), DOUT(8) => ALU_RES_OUT(8), DOUT(7) 
                           => ALU_RES_OUT(7), DOUT(6) => ALU_RES_OUT(6), 
                           DOUT(5) => ALU_RES_OUT(5), DOUT(4) => ALU_RES_OUT(4)
                           , DOUT(3) => ALU_RES_OUT(3), DOUT(2) => 
                           ALU_RES_OUT(2), DOUT(1) => ALU_RES_OUT(1), DOUT(0) 
                           => ALU_RES_OUT(0));
   PCsel : mux41_NBIT32_2 port map( A(31) => NPC_IN(31), A(30) => NPC_IN(30), 
                           A(29) => NPC_IN(29), A(28) => NPC_IN(28), A(27) => 
                           NPC_IN(27), A(26) => NPC_IN(26), A(25) => NPC_IN(25)
                           , A(24) => NPC_IN(24), A(23) => NPC_IN(23), A(22) =>
                           NPC_IN(22), A(21) => NPC_IN(21), A(20) => NPC_IN(20)
                           , A(19) => NPC_IN(19), A(18) => NPC_IN(18), A(17) =>
                           NPC_IN(17), A(16) => NPC_IN(16), A(15) => NPC_IN(15)
                           , A(14) => NPC_IN(14), A(13) => NPC_IN(13), A(12) =>
                           NPC_IN(12), A(11) => NPC_IN(11), A(10) => NPC_IN(10)
                           , A(9) => NPC_IN(9), A(8) => NPC_IN(8), A(7) => 
                           NPC_IN(7), A(6) => NPC_IN(6), A(5) => NPC_IN(5), 
                           A(4) => NPC_IN(4), A(3) => NPC_IN(3), A(2) => 
                           NPC_IN(2), A(1) => NPC_IN(1), A(0) => NPC_IN(0), 
                           B(31) => NPC_REL(31), B(30) => NPC_REL(30), B(29) =>
                           NPC_REL(29), B(28) => NPC_REL(28), B(27) => 
                           NPC_REL(27), B(26) => NPC_REL(26), B(25) => 
                           NPC_REL(25), B(24) => NPC_REL(24), B(23) => 
                           NPC_REL(23), B(22) => NPC_REL(22), B(21) => 
                           NPC_REL(21), B(20) => NPC_REL(20), B(19) => 
                           NPC_REL(19), B(18) => NPC_REL(18), B(17) => 
                           NPC_REL(17), B(16) => NPC_REL(16), B(15) => 
                           NPC_REL(15), B(14) => NPC_REL(14), B(13) => 
                           NPC_REL(13), B(12) => NPC_REL(12), B(11) => 
                           NPC_REL(11), B(10) => NPC_REL(10), B(9) => 
                           NPC_REL(9), B(8) => NPC_REL(8), B(7) => NPC_REL(7), 
                           B(6) => NPC_REL(6), B(5) => NPC_REL(5), B(4) => 
                           NPC_REL(4), B(3) => NPC_REL(3), B(2) => NPC_REL(2), 
                           B(1) => NPC_REL(1), B(0) => NPC_REL(0), C(31) => 
                           NPC_ABS(31), C(30) => NPC_ABS(30), C(29) => 
                           NPC_ABS(29), C(28) => NPC_ABS(28), C(27) => 
                           NPC_ABS(27), C(26) => NPC_ABS(26), C(25) => 
                           NPC_ABS(25), C(24) => NPC_ABS(24), C(23) => 
                           NPC_ABS(23), C(22) => NPC_ABS(22), C(21) => 
                           NPC_ABS(21), C(20) => NPC_ABS(20), C(19) => 
                           NPC_ABS(19), C(18) => NPC_ABS(18), C(17) => 
                           NPC_ABS(17), C(16) => NPC_ABS(16), C(15) => 
                           NPC_ABS(15), C(14) => NPC_ABS(14), C(13) => 
                           NPC_ABS(13), C(12) => NPC_ABS(12), C(11) => 
                           NPC_ABS(11), C(10) => NPC_ABS(10), C(9) => 
                           NPC_ABS(9), C(8) => NPC_ABS(8), C(7) => NPC_ABS(7), 
                           C(6) => NPC_ABS(6), C(5) => NPC_ABS(5), C(4) => 
                           NPC_ABS(4), C(3) => NPC_ABS(3), C(2) => NPC_ABS(2), 
                           C(1) => NPC_ABS(1), C(0) => NPC_ABS(0), D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => X_Logic0_port, D(25) => 
                           X_Logic0_port, D(24) => X_Logic0_port, D(23) => 
                           X_Logic0_port, D(22) => X_Logic0_port, D(21) => 
                           X_Logic0_port, D(20) => X_Logic0_port, D(19) => 
                           X_Logic0_port, D(18) => X_Logic0_port, D(17) => 
                           X_Logic0_port, D(16) => X_Logic0_port, D(15) => 
                           X_Logic0_port, D(14) => X_Logic0_port, D(13) => 
                           X_Logic0_port, D(12) => X_Logic0_port, D(11) => 
                           X_Logic0_port, D(10) => X_Logic0_port, D(9) => 
                           X_Logic0_port, D(8) => X_Logic0_port, D(7) => 
                           X_Logic0_port, D(6) => X_Logic0_port, D(5) => 
                           X_Logic0_port, D(4) => X_Logic0_port, D(3) => 
                           X_Logic0_port, D(2) => X_Logic0_port, D(1) => 
                           X_Logic0_port, D(0) => X_Logic0_port, S(1) => 
                           PC_SEL(1), S(0) => PC_SEL(0), Z(31) => PC_OUT(31), 
                           Z(30) => PC_OUT(30), Z(29) => PC_OUT(29), Z(28) => 
                           PC_OUT(28), Z(27) => PC_OUT(27), Z(26) => PC_OUT(26)
                           , Z(25) => PC_OUT(25), Z(24) => PC_OUT(24), Z(23) =>
                           PC_OUT(23), Z(22) => PC_OUT(22), Z(21) => PC_OUT(21)
                           , Z(20) => PC_OUT(20), Z(19) => PC_OUT(19), Z(18) =>
                           PC_OUT(18), Z(17) => PC_OUT(17), Z(16) => PC_OUT(16)
                           , Z(15) => PC_OUT(15), Z(14) => PC_OUT(14), Z(13) =>
                           PC_OUT(13), Z(12) => PC_OUT(12), Z(11) => PC_OUT(11)
                           , Z(10) => PC_OUT(10), Z(9) => PC_OUT(9), Z(8) => 
                           PC_OUT(8), Z(7) => PC_OUT(7), Z(6) => PC_OUT(6), 
                           Z(5) => PC_OUT(5), Z(4) => PC_OUT(4), Z(3) => 
                           PC_OUT(3), Z(2) => PC_OUT(2), Z(1) => PC_OUT(1), 
                           Z(0) => PC_OUT(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity ff_0 is

   port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);

end ff_0;

architecture SYN_bhv of ff_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   Q_reg : DFFR_X1 port map( D => n3, CK => CLK, RN => RST, Q => Q, QN => n2);
   U2 : OAI21_X1 port map( B1 => n2, B2 => EN, A => n1, ZN => n3);
   U3 : NAND2_X1 port map( A1 => EN, A2 => D, ZN => n1);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Execute is

   port( CLK, RST, MUX_A_SEL : in std_logic;  MUX_B_SEL : in std_logic_vector 
         (1 downto 0);  ALU_OPC : in std_logic_vector (0 to 4);  ALU_OUTREG_EN 
         : in std_logic;  JUMP_TYPE : in std_logic_vector (1 downto 0);  PC_IN,
         A_IN, B_IN, IMM_IN : in std_logic_vector (31 downto 0);  ADD_WR_IN, 
         ADD_RS1_IN, ADD_RS2_IN, ADD_WR_MEM, ADD_WR_WB : in std_logic_vector (4
         downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;  OP_MEM, OP_WB : in 
         std_logic_vector (31 downto 0);  PC_SEL : out std_logic_vector (1 
         downto 0);  ZERO_FLAG : out std_logic;  NPC_ABS, NPC_REL, ALU_RES, 
         B_OUT : out std_logic_vector (31 downto 0);  ADD_WR_OUT : out 
         std_logic_vector (4 downto 0));

end Execute;

architecture SYN_struct of Execute is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component Execute_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component Execute_DW01_add_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component regn_N32_2
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_3
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N5_2
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N32_4
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_5
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component ALU_NBIT32
      port( OP1, OP2 : in std_logic_vector (31 downto 0);  ALU_OPC : in 
            std_logic_vector (0 to 4);  ALU_RES : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux41_NBIT32_3
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux21_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux41_NBIT32_4
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux41_NBIT32_0
      port( A, B, C, D : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (1 downto 0);  Z : out std_logic_vector (31 downto
            0));
   end component;
   
   component FWD_Unit
      port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB : in 
            std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB : in std_logic;
            FWDA, FWDB : out std_logic_vector (1 downto 0));
   end component;
   
   component regn_N2
      port( DIN : in std_logic_vector (1 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (1 downto 0));
   end component;
   
   component ff_1
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Branch_Cond_Unit_NBIT32
      port( RST : in std_logic;  A : in std_logic_vector (31 downto 0);  
            ALU_OPC : in std_logic_vector (0 to 4);  JUMP_TYPE : in 
            std_logic_vector (1 downto 0);  PC_SEL : out std_logic_vector (1 
            downto 0);  ZERO : out std_logic);
   end component;
   
   signal ZERO_FLAG_port, sig_RST, sig_NPC_ABS_31_port, sig_NPC_ABS_30_port, 
      sig_NPC_ABS_29_port, sig_NPC_ABS_28_port, sig_NPC_ABS_27_port, 
      sig_NPC_ABS_26_port, sig_NPC_ABS_25_port, sig_NPC_ABS_24_port, 
      sig_NPC_ABS_23_port, sig_NPC_ABS_22_port, sig_NPC_ABS_21_port, 
      sig_NPC_ABS_20_port, sig_NPC_ABS_19_port, sig_NPC_ABS_18_port, 
      sig_NPC_ABS_17_port, sig_NPC_ABS_16_port, sig_NPC_ABS_15_port, 
      sig_NPC_ABS_14_port, sig_NPC_ABS_13_port, sig_NPC_ABS_12_port, 
      sig_NPC_ABS_11_port, sig_NPC_ABS_10_port, sig_NPC_ABS_9_port, 
      sig_NPC_ABS_8_port, sig_NPC_ABS_7_port, sig_NPC_ABS_6_port, 
      sig_NPC_ABS_5_port, sig_NPC_ABS_4_port, sig_NPC_ABS_3_port, 
      sig_NPC_ABS_2_port, sig_NPC_ABS_1_port, sig_NPC_ABS_0_port, 
      sig_NPC_REL_31_port, sig_NPC_REL_30_port, sig_NPC_REL_29_port, 
      sig_NPC_REL_28_port, sig_NPC_REL_27_port, sig_NPC_REL_26_port, 
      sig_NPC_REL_25_port, sig_NPC_REL_24_port, sig_NPC_REL_23_port, 
      sig_NPC_REL_22_port, sig_NPC_REL_21_port, sig_NPC_REL_20_port, 
      sig_NPC_REL_19_port, sig_NPC_REL_18_port, sig_NPC_REL_17_port, 
      sig_NPC_REL_16_port, sig_NPC_REL_15_port, sig_NPC_REL_14_port, 
      sig_NPC_REL_13_port, sig_NPC_REL_12_port, sig_NPC_REL_11_port, 
      sig_NPC_REL_10_port, sig_NPC_REL_9_port, sig_NPC_REL_8_port, 
      sig_NPC_REL_7_port, sig_NPC_REL_6_port, sig_NPC_REL_5_port, 
      sig_NPC_REL_4_port, sig_NPC_REL_3_port, sig_NPC_REL_2_port, 
      sig_NPC_REL_1_port, sig_NPC_REL_0_port, sig_PC_SEL_1_port, 
      sig_PC_SEL_0_port, sig_ZERO_FLAG, FWDA_1_port, FWDA_0_port, FWDB_1_port, 
      FWDB_0_port, OP2_FW_31_port, OP2_FW_30_port, OP2_FW_29_port, 
      OP2_FW_28_port, OP2_FW_27_port, OP2_FW_26_port, OP2_FW_25_port, 
      OP2_FW_24_port, OP2_FW_23_port, OP2_FW_22_port, OP2_FW_21_port, 
      OP2_FW_20_port, OP2_FW_19_port, OP2_FW_18_port, OP2_FW_17_port, 
      OP2_FW_16_port, OP2_FW_15_port, OP2_FW_14_port, OP2_FW_13_port, 
      OP2_FW_12_port, OP2_FW_11_port, OP2_FW_10_port, OP2_FW_9_port, 
      OP2_FW_8_port, OP2_FW_7_port, OP2_FW_6_port, OP2_FW_5_port, OP2_FW_4_port
      , OP2_FW_3_port, OP2_FW_2_port, OP2_FW_1_port, OP2_FW_0_port, 
      sig_OP1_31_port, sig_OP1_30_port, sig_OP1_29_port, sig_OP1_28_port, 
      sig_OP1_27_port, sig_OP1_26_port, sig_OP1_25_port, sig_OP1_24_port, 
      sig_OP1_23_port, sig_OP1_22_port, sig_OP1_21_port, sig_OP1_20_port, 
      sig_OP1_19_port, sig_OP1_18_port, sig_OP1_17_port, sig_OP1_16_port, 
      sig_OP1_15_port, sig_OP1_14_port, sig_OP1_13_port, sig_OP1_12_port, 
      sig_OP1_11_port, sig_OP1_10_port, sig_OP1_9_port, sig_OP1_8_port, 
      sig_OP1_7_port, sig_OP1_6_port, sig_OP1_5_port, sig_OP1_4_port, 
      sig_OP1_3_port, sig_OP1_2_port, sig_OP1_1_port, sig_OP1_0_port, 
      sig_OP2_31_port, sig_OP2_30_port, sig_OP2_29_port, sig_OP2_28_port, 
      sig_OP2_27_port, sig_OP2_26_port, sig_OP2_25_port, sig_OP2_24_port, 
      sig_OP2_23_port, sig_OP2_22_port, sig_OP2_21_port, sig_OP2_20_port, 
      sig_OP2_19_port, sig_OP2_18_port, sig_OP2_17_port, sig_OP2_16_port, 
      sig_OP2_15_port, sig_OP2_14_port, sig_OP2_13_port, sig_OP2_12_port, 
      sig_OP2_11_port, sig_OP2_10_port, sig_OP2_9_port, sig_OP2_8_port, 
      sig_OP2_7_port, sig_OP2_6_port, sig_OP2_5_port, sig_OP2_4_port, 
      sig_OP2_3_port, sig_OP2_2_port, sig_OP2_1_port, sig_OP2_0_port, 
      sig_ALU_RES_31_port, sig_ALU_RES_30_port, sig_ALU_RES_29_port, 
      sig_ALU_RES_28_port, sig_ALU_RES_27_port, sig_ALU_RES_26_port, 
      sig_ALU_RES_25_port, sig_ALU_RES_24_port, sig_ALU_RES_23_port, 
      sig_ALU_RES_22_port, sig_ALU_RES_21_port, sig_ALU_RES_20_port, 
      sig_ALU_RES_19_port, sig_ALU_RES_18_port, sig_ALU_RES_17_port, 
      sig_ALU_RES_16_port, sig_ALU_RES_15_port, sig_ALU_RES_14_port, 
      sig_ALU_RES_13_port, sig_ALU_RES_12_port, sig_ALU_RES_11_port, 
      sig_ALU_RES_10_port, sig_ALU_RES_9_port, sig_ALU_RES_8_port, 
      sig_ALU_RES_7_port, sig_ALU_RES_6_port, sig_ALU_RES_5_port, 
      sig_ALU_RES_4_port, sig_ALU_RES_3_port, sig_ALU_RES_2_port, 
      sig_ALU_RES_1_port, sig_ALU_RES_0_port, N9, N8, N7, N6, N5, N4, N31, N30,
      N3, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N2, N19, N18, N17, 
      N16, N15, N14, N13, N12, N11, N10, N1, N0, n1_port, n2_port, n3_port, 
      n4_port, n5_port, n6_port, n7_port, n_1983, n_1984 : std_logic;

begin
   ZERO_FLAG <= ZERO_FLAG_port;
   
   n7_port <= '1';
   n6_port <= '0';
   Branch_Cond : Branch_Cond_Unit_NBIT32 port map( RST => sig_RST, A(31) => 
                           sig_NPC_ABS_31_port, A(30) => sig_NPC_ABS_30_port, 
                           A(29) => sig_NPC_ABS_29_port, A(28) => 
                           sig_NPC_ABS_28_port, A(27) => sig_NPC_ABS_27_port, 
                           A(26) => sig_NPC_ABS_26_port, A(25) => 
                           sig_NPC_ABS_25_port, A(24) => sig_NPC_ABS_24_port, 
                           A(23) => sig_NPC_ABS_23_port, A(22) => 
                           sig_NPC_ABS_22_port, A(21) => sig_NPC_ABS_21_port, 
                           A(20) => sig_NPC_ABS_20_port, A(19) => 
                           sig_NPC_ABS_19_port, A(18) => sig_NPC_ABS_18_port, 
                           A(17) => sig_NPC_ABS_17_port, A(16) => 
                           sig_NPC_ABS_16_port, A(15) => sig_NPC_ABS_15_port, 
                           A(14) => sig_NPC_ABS_14_port, A(13) => 
                           sig_NPC_ABS_13_port, A(12) => sig_NPC_ABS_12_port, 
                           A(11) => sig_NPC_ABS_11_port, A(10) => 
                           sig_NPC_ABS_10_port, A(9) => sig_NPC_ABS_9_port, 
                           A(8) => sig_NPC_ABS_8_port, A(7) => 
                           sig_NPC_ABS_7_port, A(6) => sig_NPC_ABS_6_port, A(5)
                           => sig_NPC_ABS_5_port, A(4) => sig_NPC_ABS_4_port, 
                           A(3) => sig_NPC_ABS_3_port, A(2) => 
                           sig_NPC_ABS_2_port, A(1) => sig_NPC_ABS_1_port, A(0)
                           => sig_NPC_ABS_0_port, ALU_OPC(0) => ALU_OPC(0), 
                           ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => ALU_OPC(2), 
                           ALU_OPC(3) => ALU_OPC(3), ALU_OPC(4) => ALU_OPC(4), 
                           JUMP_TYPE(1) => JUMP_TYPE(1), JUMP_TYPE(0) => 
                           JUMP_TYPE(0), PC_SEL(1) => sig_PC_SEL_1_port, 
                           PC_SEL(0) => sig_PC_SEL_0_port, ZERO => 
                           sig_ZERO_FLAG);
   ff0 : ff_1 port map( D => sig_ZERO_FLAG, CLK => CLK, EN => n7_port, RST => 
                           RST, Q => ZERO_FLAG_port);
   reg0 : regn_N2 port map( DIN(1) => sig_PC_SEL_1_port, DIN(0) => 
                           sig_PC_SEL_0_port, CLK => CLK, EN => n7_port, RST =>
                           RST, DOUT(1) => PC_SEL(1), DOUT(0) => PC_SEL(0));
   FWD : FWD_Unit port map( RST => sig_RST, ADD_RS1(4) => ADD_RS1_IN(4), 
                           ADD_RS1(3) => ADD_RS1_IN(3), ADD_RS1(2) => 
                           ADD_RS1_IN(2), ADD_RS1(1) => ADD_RS1_IN(1), 
                           ADD_RS1(0) => ADD_RS1_IN(0), ADD_RS2(4) => 
                           ADD_RS2_IN(4), ADD_RS2(3) => ADD_RS2_IN(3), 
                           ADD_RS2(2) => ADD_RS2_IN(2), ADD_RS2(1) => 
                           ADD_RS2_IN(1), ADD_RS2(0) => ADD_RS2_IN(0), 
                           ADD_WR_MEM(4) => ADD_WR_MEM(4), ADD_WR_MEM(3) => 
                           ADD_WR_MEM(3), ADD_WR_MEM(2) => ADD_WR_MEM(2), 
                           ADD_WR_MEM(1) => ADD_WR_MEM(1), ADD_WR_MEM(0) => 
                           ADD_WR_MEM(0), ADD_WR_WB(4) => ADD_WR_WB(4), 
                           ADD_WR_WB(3) => ADD_WR_WB(3), ADD_WR_WB(2) => 
                           ADD_WR_WB(2), ADD_WR_WB(1) => ADD_WR_WB(1), 
                           ADD_WR_WB(0) => ADD_WR_WB(0), RF_WE_MEM => RF_WE_MEM
                           , RF_WE_WB => RF_WE_WB, FWDA(1) => FWDA_1_port, 
                           FWDA(0) => FWDA_0_port, FWDB(1) => FWDB_1_port, 
                           FWDB(0) => FWDB_0_port);
   FW1 : mux41_NBIT32_0 port map( A(31) => A_IN(31), A(30) => A_IN(30), A(29) 
                           => A_IN(29), A(28) => A_IN(28), A(27) => A_IN(27), 
                           A(26) => A_IN(26), A(25) => A_IN(25), A(24) => 
                           A_IN(24), A(23) => A_IN(23), A(22) => A_IN(22), 
                           A(21) => A_IN(21), A(20) => A_IN(20), A(19) => 
                           A_IN(19), A(18) => A_IN(18), A(17) => A_IN(17), 
                           A(16) => A_IN(16), A(15) => A_IN(15), A(14) => 
                           A_IN(14), A(13) => A_IN(13), A(12) => A_IN(12), 
                           A(11) => A_IN(11), A(10) => A_IN(10), A(9) => 
                           A_IN(9), A(8) => A_IN(8), A(7) => A_IN(7), A(6) => 
                           A_IN(6), A(5) => A_IN(5), A(4) => A_IN(4), A(3) => 
                           A_IN(3), A(2) => A_IN(2), A(1) => A_IN(1), A(0) => 
                           A_IN(0), B(31) => OP_WB(31), B(30) => OP_WB(30), 
                           B(29) => OP_WB(29), B(28) => OP_WB(28), B(27) => 
                           OP_WB(27), B(26) => OP_WB(26), B(25) => OP_WB(25), 
                           B(24) => OP_WB(24), B(23) => OP_WB(23), B(22) => 
                           OP_WB(22), B(21) => OP_WB(21), B(20) => OP_WB(20), 
                           B(19) => OP_WB(19), B(18) => OP_WB(18), B(17) => 
                           OP_WB(17), B(16) => OP_WB(16), B(15) => OP_WB(15), 
                           B(14) => OP_WB(14), B(13) => OP_WB(13), B(12) => 
                           OP_WB(12), B(11) => OP_WB(11), B(10) => OP_WB(10), 
                           B(9) => OP_WB(9), B(8) => OP_WB(8), B(7) => OP_WB(7)
                           , B(6) => OP_WB(6), B(5) => OP_WB(5), B(4) => 
                           OP_WB(4), B(3) => OP_WB(3), B(2) => OP_WB(2), B(1) 
                           => OP_WB(1), B(0) => OP_WB(0), C(31) => OP_MEM(31), 
                           C(30) => OP_MEM(30), C(29) => OP_MEM(29), C(28) => 
                           OP_MEM(28), C(27) => OP_MEM(27), C(26) => OP_MEM(26)
                           , C(25) => OP_MEM(25), C(24) => OP_MEM(24), C(23) =>
                           OP_MEM(23), C(22) => OP_MEM(22), C(21) => OP_MEM(21)
                           , C(20) => OP_MEM(20), C(19) => OP_MEM(19), C(18) =>
                           OP_MEM(18), C(17) => OP_MEM(17), C(16) => OP_MEM(16)
                           , C(15) => OP_MEM(15), C(14) => OP_MEM(14), C(13) =>
                           OP_MEM(13), C(12) => OP_MEM(12), C(11) => OP_MEM(11)
                           , C(10) => OP_MEM(10), C(9) => OP_MEM(9), C(8) => 
                           OP_MEM(8), C(7) => OP_MEM(7), C(6) => OP_MEM(6), 
                           C(5) => OP_MEM(5), C(4) => OP_MEM(4), C(3) => 
                           OP_MEM(3), C(2) => OP_MEM(2), C(1) => OP_MEM(1), 
                           C(0) => OP_MEM(0), D(31) => A_IN(31), D(30) => 
                           A_IN(30), D(29) => A_IN(29), D(28) => A_IN(28), 
                           D(27) => A_IN(27), D(26) => A_IN(26), D(25) => 
                           A_IN(25), D(24) => A_IN(24), D(23) => A_IN(23), 
                           D(22) => A_IN(22), D(21) => A_IN(21), D(20) => 
                           A_IN(20), D(19) => A_IN(19), D(18) => A_IN(18), 
                           D(17) => A_IN(17), D(16) => A_IN(16), D(15) => 
                           A_IN(15), D(14) => A_IN(14), D(13) => A_IN(13), 
                           D(12) => A_IN(12), D(11) => A_IN(11), D(10) => 
                           A_IN(10), D(9) => A_IN(9), D(8) => A_IN(8), D(7) => 
                           A_IN(7), D(6) => A_IN(6), D(5) => A_IN(5), D(4) => 
                           A_IN(4), D(3) => A_IN(3), D(2) => A_IN(2), D(1) => 
                           A_IN(1), D(0) => A_IN(0), S(1) => FWDA_1_port, S(0) 
                           => FWDA_0_port, Z(31) => sig_NPC_ABS_31_port, Z(30) 
                           => sig_NPC_ABS_30_port, Z(29) => sig_NPC_ABS_29_port
                           , Z(28) => sig_NPC_ABS_28_port, Z(27) => 
                           sig_NPC_ABS_27_port, Z(26) => sig_NPC_ABS_26_port, 
                           Z(25) => sig_NPC_ABS_25_port, Z(24) => 
                           sig_NPC_ABS_24_port, Z(23) => sig_NPC_ABS_23_port, 
                           Z(22) => sig_NPC_ABS_22_port, Z(21) => 
                           sig_NPC_ABS_21_port, Z(20) => sig_NPC_ABS_20_port, 
                           Z(19) => sig_NPC_ABS_19_port, Z(18) => 
                           sig_NPC_ABS_18_port, Z(17) => sig_NPC_ABS_17_port, 
                           Z(16) => sig_NPC_ABS_16_port, Z(15) => 
                           sig_NPC_ABS_15_port, Z(14) => sig_NPC_ABS_14_port, 
                           Z(13) => sig_NPC_ABS_13_port, Z(12) => 
                           sig_NPC_ABS_12_port, Z(11) => sig_NPC_ABS_11_port, 
                           Z(10) => sig_NPC_ABS_10_port, Z(9) => 
                           sig_NPC_ABS_9_port, Z(8) => sig_NPC_ABS_8_port, Z(7)
                           => sig_NPC_ABS_7_port, Z(6) => sig_NPC_ABS_6_port, 
                           Z(5) => sig_NPC_ABS_5_port, Z(4) => 
                           sig_NPC_ABS_4_port, Z(3) => sig_NPC_ABS_3_port, Z(2)
                           => sig_NPC_ABS_2_port, Z(1) => sig_NPC_ABS_1_port, 
                           Z(0) => sig_NPC_ABS_0_port);
   FW2 : mux41_NBIT32_4 port map( A(31) => B_IN(31), A(30) => B_IN(30), A(29) 
                           => B_IN(29), A(28) => B_IN(28), A(27) => B_IN(27), 
                           A(26) => B_IN(26), A(25) => B_IN(25), A(24) => 
                           B_IN(24), A(23) => B_IN(23), A(22) => B_IN(22), 
                           A(21) => B_IN(21), A(20) => B_IN(20), A(19) => 
                           B_IN(19), A(18) => B_IN(18), A(17) => B_IN(17), 
                           A(16) => B_IN(16), A(15) => B_IN(15), A(14) => 
                           B_IN(14), A(13) => B_IN(13), A(12) => B_IN(12), 
                           A(11) => B_IN(11), A(10) => B_IN(10), A(9) => 
                           B_IN(9), A(8) => B_IN(8), A(7) => B_IN(7), A(6) => 
                           B_IN(6), A(5) => B_IN(5), A(4) => B_IN(4), A(3) => 
                           B_IN(3), A(2) => B_IN(2), A(1) => B_IN(1), A(0) => 
                           B_IN(0), B(31) => OP_WB(31), B(30) => OP_WB(30), 
                           B(29) => OP_WB(29), B(28) => OP_WB(28), B(27) => 
                           OP_WB(27), B(26) => OP_WB(26), B(25) => OP_WB(25), 
                           B(24) => OP_WB(24), B(23) => OP_WB(23), B(22) => 
                           OP_WB(22), B(21) => OP_WB(21), B(20) => OP_WB(20), 
                           B(19) => OP_WB(19), B(18) => OP_WB(18), B(17) => 
                           OP_WB(17), B(16) => OP_WB(16), B(15) => OP_WB(15), 
                           B(14) => OP_WB(14), B(13) => OP_WB(13), B(12) => 
                           OP_WB(12), B(11) => OP_WB(11), B(10) => OP_WB(10), 
                           B(9) => OP_WB(9), B(8) => OP_WB(8), B(7) => OP_WB(7)
                           , B(6) => OP_WB(6), B(5) => OP_WB(5), B(4) => 
                           OP_WB(4), B(3) => OP_WB(3), B(2) => OP_WB(2), B(1) 
                           => OP_WB(1), B(0) => OP_WB(0), C(31) => OP_MEM(31), 
                           C(30) => OP_MEM(30), C(29) => OP_MEM(29), C(28) => 
                           OP_MEM(28), C(27) => OP_MEM(27), C(26) => OP_MEM(26)
                           , C(25) => OP_MEM(25), C(24) => OP_MEM(24), C(23) =>
                           OP_MEM(23), C(22) => OP_MEM(22), C(21) => OP_MEM(21)
                           , C(20) => OP_MEM(20), C(19) => OP_MEM(19), C(18) =>
                           OP_MEM(18), C(17) => OP_MEM(17), C(16) => OP_MEM(16)
                           , C(15) => OP_MEM(15), C(14) => OP_MEM(14), C(13) =>
                           OP_MEM(13), C(12) => OP_MEM(12), C(11) => OP_MEM(11)
                           , C(10) => OP_MEM(10), C(9) => OP_MEM(9), C(8) => 
                           OP_MEM(8), C(7) => OP_MEM(7), C(6) => OP_MEM(6), 
                           C(5) => OP_MEM(5), C(4) => OP_MEM(4), C(3) => 
                           OP_MEM(3), C(2) => OP_MEM(2), C(1) => OP_MEM(1), 
                           C(0) => OP_MEM(0), D(31) => B_IN(31), D(30) => 
                           B_IN(30), D(29) => B_IN(29), D(28) => B_IN(28), 
                           D(27) => B_IN(27), D(26) => B_IN(26), D(25) => 
                           B_IN(25), D(24) => B_IN(24), D(23) => B_IN(23), 
                           D(22) => B_IN(22), D(21) => B_IN(21), D(20) => 
                           B_IN(20), D(19) => B_IN(19), D(18) => B_IN(18), 
                           D(17) => B_IN(17), D(16) => B_IN(16), D(15) => 
                           B_IN(15), D(14) => B_IN(14), D(13) => B_IN(13), 
                           D(12) => B_IN(12), D(11) => B_IN(11), D(10) => 
                           B_IN(10), D(9) => B_IN(9), D(8) => B_IN(8), D(7) => 
                           B_IN(7), D(6) => B_IN(6), D(5) => B_IN(5), D(4) => 
                           B_IN(4), D(3) => B_IN(3), D(2) => B_IN(2), D(1) => 
                           B_IN(1), D(0) => B_IN(0), S(1) => FWDB_1_port, S(0) 
                           => FWDB_0_port, Z(31) => OP2_FW_31_port, Z(30) => 
                           OP2_FW_30_port, Z(29) => OP2_FW_29_port, Z(28) => 
                           OP2_FW_28_port, Z(27) => OP2_FW_27_port, Z(26) => 
                           OP2_FW_26_port, Z(25) => OP2_FW_25_port, Z(24) => 
                           OP2_FW_24_port, Z(23) => OP2_FW_23_port, Z(22) => 
                           OP2_FW_22_port, Z(21) => OP2_FW_21_port, Z(20) => 
                           OP2_FW_20_port, Z(19) => OP2_FW_19_port, Z(18) => 
                           OP2_FW_18_port, Z(17) => OP2_FW_17_port, Z(16) => 
                           OP2_FW_16_port, Z(15) => OP2_FW_15_port, Z(14) => 
                           OP2_FW_14_port, Z(13) => OP2_FW_13_port, Z(12) => 
                           OP2_FW_12_port, Z(11) => OP2_FW_11_port, Z(10) => 
                           OP2_FW_10_port, Z(9) => OP2_FW_9_port, Z(8) => 
                           OP2_FW_8_port, Z(7) => OP2_FW_7_port, Z(6) => 
                           OP2_FW_6_port, Z(5) => OP2_FW_5_port, Z(4) => 
                           OP2_FW_4_port, Z(3) => OP2_FW_3_port, Z(2) => 
                           OP2_FW_2_port, Z(1) => OP2_FW_1_port, Z(0) => 
                           OP2_FW_0_port);
   muxA : mux21_NBIT32_4 port map( A(31) => sig_NPC_ABS_31_port, A(30) => 
                           sig_NPC_ABS_30_port, A(29) => sig_NPC_ABS_29_port, 
                           A(28) => sig_NPC_ABS_28_port, A(27) => 
                           sig_NPC_ABS_27_port, A(26) => sig_NPC_ABS_26_port, 
                           A(25) => sig_NPC_ABS_25_port, A(24) => 
                           sig_NPC_ABS_24_port, A(23) => sig_NPC_ABS_23_port, 
                           A(22) => sig_NPC_ABS_22_port, A(21) => 
                           sig_NPC_ABS_21_port, A(20) => sig_NPC_ABS_20_port, 
                           A(19) => sig_NPC_ABS_19_port, A(18) => 
                           sig_NPC_ABS_18_port, A(17) => sig_NPC_ABS_17_port, 
                           A(16) => sig_NPC_ABS_16_port, A(15) => 
                           sig_NPC_ABS_15_port, A(14) => sig_NPC_ABS_14_port, 
                           A(13) => sig_NPC_ABS_13_port, A(12) => 
                           sig_NPC_ABS_12_port, A(11) => sig_NPC_ABS_11_port, 
                           A(10) => sig_NPC_ABS_10_port, A(9) => 
                           sig_NPC_ABS_9_port, A(8) => sig_NPC_ABS_8_port, A(7)
                           => sig_NPC_ABS_7_port, A(6) => sig_NPC_ABS_6_port, 
                           A(5) => sig_NPC_ABS_5_port, A(4) => 
                           sig_NPC_ABS_4_port, A(3) => sig_NPC_ABS_3_port, A(2)
                           => sig_NPC_ABS_2_port, A(1) => sig_NPC_ABS_1_port, 
                           A(0) => sig_NPC_ABS_0_port, B(31) => PC_IN(31), 
                           B(30) => PC_IN(30), B(29) => PC_IN(29), B(28) => 
                           PC_IN(28), B(27) => PC_IN(27), B(26) => PC_IN(26), 
                           B(25) => PC_IN(25), B(24) => PC_IN(24), B(23) => 
                           PC_IN(23), B(22) => PC_IN(22), B(21) => PC_IN(21), 
                           B(20) => PC_IN(20), B(19) => PC_IN(19), B(18) => 
                           PC_IN(18), B(17) => PC_IN(17), B(16) => PC_IN(16), 
                           B(15) => PC_IN(15), B(14) => PC_IN(14), B(13) => 
                           PC_IN(13), B(12) => PC_IN(12), B(11) => PC_IN(11), 
                           B(10) => PC_IN(10), B(9) => PC_IN(9), B(8) => 
                           PC_IN(8), B(7) => PC_IN(7), B(6) => PC_IN(6), B(5) 
                           => PC_IN(5), B(4) => PC_IN(4), B(3) => PC_IN(3), 
                           B(2) => PC_IN(2), B(1) => PC_IN(1), B(0) => PC_IN(0)
                           , S => MUX_A_SEL, Z(31) => sig_OP1_31_port, Z(30) =>
                           sig_OP1_30_port, Z(29) => sig_OP1_29_port, Z(28) => 
                           sig_OP1_28_port, Z(27) => sig_OP1_27_port, Z(26) => 
                           sig_OP1_26_port, Z(25) => sig_OP1_25_port, Z(24) => 
                           sig_OP1_24_port, Z(23) => sig_OP1_23_port, Z(22) => 
                           sig_OP1_22_port, Z(21) => sig_OP1_21_port, Z(20) => 
                           sig_OP1_20_port, Z(19) => sig_OP1_19_port, Z(18) => 
                           sig_OP1_18_port, Z(17) => sig_OP1_17_port, Z(16) => 
                           sig_OP1_16_port, Z(15) => sig_OP1_15_port, Z(14) => 
                           sig_OP1_14_port, Z(13) => sig_OP1_13_port, Z(12) => 
                           sig_OP1_12_port, Z(11) => sig_OP1_11_port, Z(10) => 
                           sig_OP1_10_port, Z(9) => sig_OP1_9_port, Z(8) => 
                           sig_OP1_8_port, Z(7) => sig_OP1_7_port, Z(6) => 
                           sig_OP1_6_port, Z(5) => sig_OP1_5_port, Z(4) => 
                           sig_OP1_4_port, Z(3) => sig_OP1_3_port, Z(2) => 
                           sig_OP1_2_port, Z(1) => sig_OP1_1_port, Z(0) => 
                           sig_OP1_0_port);
   muxB : mux41_NBIT32_3 port map( A(31) => OP2_FW_31_port, A(30) => 
                           OP2_FW_30_port, A(29) => OP2_FW_29_port, A(28) => 
                           OP2_FW_28_port, A(27) => OP2_FW_27_port, A(26) => 
                           OP2_FW_26_port, A(25) => OP2_FW_25_port, A(24) => 
                           OP2_FW_24_port, A(23) => OP2_FW_23_port, A(22) => 
                           OP2_FW_22_port, A(21) => OP2_FW_21_port, A(20) => 
                           OP2_FW_20_port, A(19) => OP2_FW_19_port, A(18) => 
                           OP2_FW_18_port, A(17) => OP2_FW_17_port, A(16) => 
                           OP2_FW_16_port, A(15) => OP2_FW_15_port, A(14) => 
                           OP2_FW_14_port, A(13) => OP2_FW_13_port, A(12) => 
                           OP2_FW_12_port, A(11) => OP2_FW_11_port, A(10) => 
                           OP2_FW_10_port, A(9) => OP2_FW_9_port, A(8) => 
                           OP2_FW_8_port, A(7) => OP2_FW_7_port, A(6) => 
                           OP2_FW_6_port, A(5) => OP2_FW_5_port, A(4) => 
                           OP2_FW_4_port, A(3) => OP2_FW_3_port, A(2) => 
                           OP2_FW_2_port, A(1) => OP2_FW_1_port, A(0) => 
                           OP2_FW_0_port, B(31) => IMM_IN(31), B(30) => 
                           IMM_IN(30), B(29) => IMM_IN(29), B(28) => IMM_IN(28)
                           , B(27) => IMM_IN(27), B(26) => IMM_IN(26), B(25) =>
                           IMM_IN(25), B(24) => IMM_IN(24), B(23) => IMM_IN(23)
                           , B(22) => IMM_IN(22), B(21) => IMM_IN(21), B(20) =>
                           IMM_IN(20), B(19) => IMM_IN(19), B(18) => IMM_IN(18)
                           , B(17) => IMM_IN(17), B(16) => IMM_IN(16), B(15) =>
                           IMM_IN(15), B(14) => IMM_IN(14), B(13) => IMM_IN(13)
                           , B(12) => IMM_IN(12), B(11) => IMM_IN(11), B(10) =>
                           IMM_IN(10), B(9) => IMM_IN(9), B(8) => IMM_IN(8), 
                           B(7) => IMM_IN(7), B(6) => IMM_IN(6), B(5) => 
                           IMM_IN(5), B(4) => IMM_IN(4), B(3) => IMM_IN(3), 
                           B(2) => IMM_IN(2), B(1) => IMM_IN(1), B(0) => 
                           IMM_IN(0), C(31) => n6_port, C(30) => n6_port, C(29)
                           => n6_port, C(28) => n6_port, C(27) => n6_port, 
                           C(26) => n6_port, C(25) => n6_port, C(24) => n6_port
                           , C(23) => n6_port, C(22) => n6_port, C(21) => 
                           n6_port, C(20) => n6_port, C(19) => n6_port, C(18) 
                           => n6_port, C(17) => n6_port, C(16) => n6_port, 
                           C(15) => n6_port, C(14) => n6_port, C(13) => n6_port
                           , C(12) => n6_port, C(11) => n6_port, C(10) => 
                           n6_port, C(9) => n6_port, C(8) => n6_port, C(7) => 
                           n6_port, C(6) => n6_port, C(5) => n6_port, C(4) => 
                           n6_port, C(3) => n6_port, C(2) => n7_port, C(1) => 
                           n6_port, C(0) => n6_port, D(31) => n6_port, D(30) =>
                           n6_port, D(29) => n6_port, D(28) => n6_port, D(27) 
                           => n6_port, D(26) => n6_port, D(25) => n6_port, 
                           D(24) => n6_port, D(23) => n6_port, D(22) => n6_port
                           , D(21) => n6_port, D(20) => n6_port, D(19) => 
                           n6_port, D(18) => n6_port, D(17) => n6_port, D(16) 
                           => n6_port, D(15) => n6_port, D(14) => n6_port, 
                           D(13) => n6_port, D(12) => n6_port, D(11) => n6_port
                           , D(10) => n6_port, D(9) => n6_port, D(8) => n6_port
                           , D(7) => n6_port, D(6) => n6_port, D(5) => n6_port,
                           D(4) => n6_port, D(3) => n6_port, D(2) => n6_port, 
                           D(1) => n6_port, D(0) => n6_port, S(1) => 
                           MUX_B_SEL(1), S(0) => MUX_B_SEL(0), Z(31) => 
                           sig_OP2_31_port, Z(30) => sig_OP2_30_port, Z(29) => 
                           sig_OP2_29_port, Z(28) => sig_OP2_28_port, Z(27) => 
                           sig_OP2_27_port, Z(26) => sig_OP2_26_port, Z(25) => 
                           sig_OP2_25_port, Z(24) => sig_OP2_24_port, Z(23) => 
                           sig_OP2_23_port, Z(22) => sig_OP2_22_port, Z(21) => 
                           sig_OP2_21_port, Z(20) => sig_OP2_20_port, Z(19) => 
                           sig_OP2_19_port, Z(18) => sig_OP2_18_port, Z(17) => 
                           sig_OP2_17_port, Z(16) => sig_OP2_16_port, Z(15) => 
                           sig_OP2_15_port, Z(14) => sig_OP2_14_port, Z(13) => 
                           sig_OP2_13_port, Z(12) => sig_OP2_12_port, Z(11) => 
                           sig_OP2_11_port, Z(10) => sig_OP2_10_port, Z(9) => 
                           sig_OP2_9_port, Z(8) => sig_OP2_8_port, Z(7) => 
                           sig_OP2_7_port, Z(6) => sig_OP2_6_port, Z(5) => 
                           sig_OP2_5_port, Z(4) => sig_OP2_4_port, Z(3) => 
                           sig_OP2_3_port, Z(2) => sig_OP2_2_port, Z(1) => 
                           sig_OP2_1_port, Z(0) => sig_OP2_0_port);
   alu0 : ALU_NBIT32 port map( OP1(31) => sig_OP1_31_port, OP1(30) => 
                           sig_OP1_30_port, OP1(29) => sig_OP1_29_port, OP1(28)
                           => sig_OP1_28_port, OP1(27) => sig_OP1_27_port, 
                           OP1(26) => sig_OP1_26_port, OP1(25) => 
                           sig_OP1_25_port, OP1(24) => sig_OP1_24_port, OP1(23)
                           => sig_OP1_23_port, OP1(22) => sig_OP1_22_port, 
                           OP1(21) => sig_OP1_21_port, OP1(20) => 
                           sig_OP1_20_port, OP1(19) => sig_OP1_19_port, OP1(18)
                           => sig_OP1_18_port, OP1(17) => sig_OP1_17_port, 
                           OP1(16) => sig_OP1_16_port, OP1(15) => 
                           sig_OP1_15_port, OP1(14) => sig_OP1_14_port, OP1(13)
                           => sig_OP1_13_port, OP1(12) => sig_OP1_12_port, 
                           OP1(11) => sig_OP1_11_port, OP1(10) => 
                           sig_OP1_10_port, OP1(9) => sig_OP1_9_port, OP1(8) =>
                           sig_OP1_8_port, OP1(7) => sig_OP1_7_port, OP1(6) => 
                           sig_OP1_6_port, OP1(5) => sig_OP1_5_port, OP1(4) => 
                           sig_OP1_4_port, OP1(3) => sig_OP1_3_port, OP1(2) => 
                           sig_OP1_2_port, OP1(1) => sig_OP1_1_port, OP1(0) => 
                           sig_OP1_0_port, OP2(31) => sig_OP2_31_port, OP2(30) 
                           => sig_OP2_30_port, OP2(29) => sig_OP2_29_port, 
                           OP2(28) => sig_OP2_28_port, OP2(27) => 
                           sig_OP2_27_port, OP2(26) => sig_OP2_26_port, OP2(25)
                           => sig_OP2_25_port, OP2(24) => sig_OP2_24_port, 
                           OP2(23) => sig_OP2_23_port, OP2(22) => 
                           sig_OP2_22_port, OP2(21) => sig_OP2_21_port, OP2(20)
                           => sig_OP2_20_port, OP2(19) => sig_OP2_19_port, 
                           OP2(18) => sig_OP2_18_port, OP2(17) => 
                           sig_OP2_17_port, OP2(16) => sig_OP2_16_port, OP2(15)
                           => sig_OP2_15_port, OP2(14) => sig_OP2_14_port, 
                           OP2(13) => sig_OP2_13_port, OP2(12) => 
                           sig_OP2_12_port, OP2(11) => sig_OP2_11_port, OP2(10)
                           => sig_OP2_10_port, OP2(9) => sig_OP2_9_port, OP2(8)
                           => sig_OP2_8_port, OP2(7) => sig_OP2_7_port, OP2(6) 
                           => sig_OP2_6_port, OP2(5) => sig_OP2_5_port, OP2(4) 
                           => sig_OP2_4_port, OP2(3) => sig_OP2_3_port, OP2(2) 
                           => sig_OP2_2_port, OP2(1) => sig_OP2_1_port, OP2(0) 
                           => sig_OP2_0_port, ALU_OPC(0) => ALU_OPC(0), 
                           ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => ALU_OPC(2), 
                           ALU_OPC(3) => ALU_OPC(3), ALU_OPC(4) => ALU_OPC(4), 
                           ALU_RES(31) => sig_ALU_RES_31_port, ALU_RES(30) => 
                           sig_ALU_RES_30_port, ALU_RES(29) => 
                           sig_ALU_RES_29_port, ALU_RES(28) => 
                           sig_ALU_RES_28_port, ALU_RES(27) => 
                           sig_ALU_RES_27_port, ALU_RES(26) => 
                           sig_ALU_RES_26_port, ALU_RES(25) => 
                           sig_ALU_RES_25_port, ALU_RES(24) => 
                           sig_ALU_RES_24_port, ALU_RES(23) => 
                           sig_ALU_RES_23_port, ALU_RES(22) => 
                           sig_ALU_RES_22_port, ALU_RES(21) => 
                           sig_ALU_RES_21_port, ALU_RES(20) => 
                           sig_ALU_RES_20_port, ALU_RES(19) => 
                           sig_ALU_RES_19_port, ALU_RES(18) => 
                           sig_ALU_RES_18_port, ALU_RES(17) => 
                           sig_ALU_RES_17_port, ALU_RES(16) => 
                           sig_ALU_RES_16_port, ALU_RES(15) => 
                           sig_ALU_RES_15_port, ALU_RES(14) => 
                           sig_ALU_RES_14_port, ALU_RES(13) => 
                           sig_ALU_RES_13_port, ALU_RES(12) => 
                           sig_ALU_RES_12_port, ALU_RES(11) => 
                           sig_ALU_RES_11_port, ALU_RES(10) => 
                           sig_ALU_RES_10_port, ALU_RES(9) => 
                           sig_ALU_RES_9_port, ALU_RES(8) => sig_ALU_RES_8_port
                           , ALU_RES(7) => sig_ALU_RES_7_port, ALU_RES(6) => 
                           sig_ALU_RES_6_port, ALU_RES(5) => sig_ALU_RES_5_port
                           , ALU_RES(4) => sig_ALU_RES_4_port, ALU_RES(3) => 
                           sig_ALU_RES_3_port, ALU_RES(2) => sig_ALU_RES_2_port
                           , ALU_RES(1) => sig_ALU_RES_1_port, ALU_RES(0) => 
                           sig_ALU_RES_0_port);
   alureg : regn_N32_5 port map( DIN(31) => sig_ALU_RES_31_port, DIN(30) => 
                           sig_ALU_RES_30_port, DIN(29) => sig_ALU_RES_29_port,
                           DIN(28) => sig_ALU_RES_28_port, DIN(27) => 
                           sig_ALU_RES_27_port, DIN(26) => sig_ALU_RES_26_port,
                           DIN(25) => sig_ALU_RES_25_port, DIN(24) => 
                           sig_ALU_RES_24_port, DIN(23) => sig_ALU_RES_23_port,
                           DIN(22) => sig_ALU_RES_22_port, DIN(21) => 
                           sig_ALU_RES_21_port, DIN(20) => sig_ALU_RES_20_port,
                           DIN(19) => sig_ALU_RES_19_port, DIN(18) => 
                           sig_ALU_RES_18_port, DIN(17) => sig_ALU_RES_17_port,
                           DIN(16) => sig_ALU_RES_16_port, DIN(15) => 
                           sig_ALU_RES_15_port, DIN(14) => sig_ALU_RES_14_port,
                           DIN(13) => sig_ALU_RES_13_port, DIN(12) => 
                           sig_ALU_RES_12_port, DIN(11) => sig_ALU_RES_11_port,
                           DIN(10) => sig_ALU_RES_10_port, DIN(9) => 
                           sig_ALU_RES_9_port, DIN(8) => sig_ALU_RES_8_port, 
                           DIN(7) => sig_ALU_RES_7_port, DIN(6) => 
                           sig_ALU_RES_6_port, DIN(5) => sig_ALU_RES_5_port, 
                           DIN(4) => sig_ALU_RES_4_port, DIN(3) => 
                           sig_ALU_RES_3_port, DIN(2) => sig_ALU_RES_2_port, 
                           DIN(1) => sig_ALU_RES_1_port, DIN(0) => 
                           sig_ALU_RES_0_port, CLK => CLK, EN => ALU_OUTREG_EN,
                           RST => RST, DOUT(31) => ALU_RES(31), DOUT(30) => 
                           ALU_RES(30), DOUT(29) => ALU_RES(29), DOUT(28) => 
                           ALU_RES(28), DOUT(27) => ALU_RES(27), DOUT(26) => 
                           ALU_RES(26), DOUT(25) => ALU_RES(25), DOUT(24) => 
                           ALU_RES(24), DOUT(23) => ALU_RES(23), DOUT(22) => 
                           ALU_RES(22), DOUT(21) => ALU_RES(21), DOUT(20) => 
                           ALU_RES(20), DOUT(19) => ALU_RES(19), DOUT(18) => 
                           ALU_RES(18), DOUT(17) => ALU_RES(17), DOUT(16) => 
                           ALU_RES(16), DOUT(15) => ALU_RES(15), DOUT(14) => 
                           ALU_RES(14), DOUT(13) => ALU_RES(13), DOUT(12) => 
                           ALU_RES(12), DOUT(11) => ALU_RES(11), DOUT(10) => 
                           ALU_RES(10), DOUT(9) => ALU_RES(9), DOUT(8) => 
                           ALU_RES(8), DOUT(7) => ALU_RES(7), DOUT(6) => 
                           ALU_RES(6), DOUT(5) => ALU_RES(5), DOUT(4) => 
                           ALU_RES(4), DOUT(3) => ALU_RES(3), DOUT(2) => 
                           ALU_RES(2), DOUT(1) => ALU_RES(1), DOUT(0) => 
                           ALU_RES(0));
   B_reg : regn_N32_4 port map( DIN(31) => OP2_FW_31_port, DIN(30) => 
                           OP2_FW_30_port, DIN(29) => OP2_FW_29_port, DIN(28) 
                           => OP2_FW_28_port, DIN(27) => OP2_FW_27_port, 
                           DIN(26) => OP2_FW_26_port, DIN(25) => OP2_FW_25_port
                           , DIN(24) => OP2_FW_24_port, DIN(23) => 
                           OP2_FW_23_port, DIN(22) => OP2_FW_22_port, DIN(21) 
                           => OP2_FW_21_port, DIN(20) => OP2_FW_20_port, 
                           DIN(19) => OP2_FW_19_port, DIN(18) => OP2_FW_18_port
                           , DIN(17) => OP2_FW_17_port, DIN(16) => 
                           OP2_FW_16_port, DIN(15) => OP2_FW_15_port, DIN(14) 
                           => OP2_FW_14_port, DIN(13) => OP2_FW_13_port, 
                           DIN(12) => OP2_FW_12_port, DIN(11) => OP2_FW_11_port
                           , DIN(10) => OP2_FW_10_port, DIN(9) => OP2_FW_9_port
                           , DIN(8) => OP2_FW_8_port, DIN(7) => OP2_FW_7_port, 
                           DIN(6) => OP2_FW_6_port, DIN(5) => OP2_FW_5_port, 
                           DIN(4) => OP2_FW_4_port, DIN(3) => OP2_FW_3_port, 
                           DIN(2) => OP2_FW_2_port, DIN(1) => OP2_FW_1_port, 
                           DIN(0) => OP2_FW_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => B_OUT(31), 
                           DOUT(30) => B_OUT(30), DOUT(29) => B_OUT(29), 
                           DOUT(28) => B_OUT(28), DOUT(27) => B_OUT(27), 
                           DOUT(26) => B_OUT(26), DOUT(25) => B_OUT(25), 
                           DOUT(24) => B_OUT(24), DOUT(23) => B_OUT(23), 
                           DOUT(22) => B_OUT(22), DOUT(21) => B_OUT(21), 
                           DOUT(20) => B_OUT(20), DOUT(19) => B_OUT(19), 
                           DOUT(18) => B_OUT(18), DOUT(17) => B_OUT(17), 
                           DOUT(16) => B_OUT(16), DOUT(15) => B_OUT(15), 
                           DOUT(14) => B_OUT(14), DOUT(13) => B_OUT(13), 
                           DOUT(12) => B_OUT(12), DOUT(11) => B_OUT(11), 
                           DOUT(10) => B_OUT(10), DOUT(9) => B_OUT(9), DOUT(8) 
                           => B_OUT(8), DOUT(7) => B_OUT(7), DOUT(6) => 
                           B_OUT(6), DOUT(5) => B_OUT(5), DOUT(4) => B_OUT(4), 
                           DOUT(3) => B_OUT(3), DOUT(2) => B_OUT(2), DOUT(1) =>
                           B_OUT(1), DOUT(0) => B_OUT(0));
   ADD_WR_reg : regn_N5_2 port map( DIN(4) => ADD_WR_IN(4), DIN(3) => 
                           ADD_WR_IN(3), DIN(2) => ADD_WR_IN(2), DIN(1) => 
                           ADD_WR_IN(1), DIN(0) => ADD_WR_IN(0), CLK => CLK, EN
                           => n7_port, RST => RST, DOUT(4) => ADD_WR_OUT(4), 
                           DOUT(3) => ADD_WR_OUT(3), DOUT(2) => ADD_WR_OUT(2), 
                           DOUT(1) => ADD_WR_OUT(1), DOUT(0) => ADD_WR_OUT(0));
   NPC_ABS_reg : regn_N32_3 port map( DIN(31) => sig_NPC_ABS_31_port, DIN(30) 
                           => sig_NPC_ABS_30_port, DIN(29) => 
                           sig_NPC_ABS_29_port, DIN(28) => sig_NPC_ABS_28_port,
                           DIN(27) => sig_NPC_ABS_27_port, DIN(26) => 
                           sig_NPC_ABS_26_port, DIN(25) => sig_NPC_ABS_25_port,
                           DIN(24) => sig_NPC_ABS_24_port, DIN(23) => 
                           sig_NPC_ABS_23_port, DIN(22) => sig_NPC_ABS_22_port,
                           DIN(21) => sig_NPC_ABS_21_port, DIN(20) => 
                           sig_NPC_ABS_20_port, DIN(19) => sig_NPC_ABS_19_port,
                           DIN(18) => sig_NPC_ABS_18_port, DIN(17) => 
                           sig_NPC_ABS_17_port, DIN(16) => sig_NPC_ABS_16_port,
                           DIN(15) => sig_NPC_ABS_15_port, DIN(14) => 
                           sig_NPC_ABS_14_port, DIN(13) => sig_NPC_ABS_13_port,
                           DIN(12) => sig_NPC_ABS_12_port, DIN(11) => 
                           sig_NPC_ABS_11_port, DIN(10) => sig_NPC_ABS_10_port,
                           DIN(9) => sig_NPC_ABS_9_port, DIN(8) => 
                           sig_NPC_ABS_8_port, DIN(7) => sig_NPC_ABS_7_port, 
                           DIN(6) => sig_NPC_ABS_6_port, DIN(5) => 
                           sig_NPC_ABS_5_port, DIN(4) => sig_NPC_ABS_4_port, 
                           DIN(3) => sig_NPC_ABS_3_port, DIN(2) => 
                           sig_NPC_ABS_2_port, DIN(1) => sig_NPC_ABS_1_port, 
                           DIN(0) => sig_NPC_ABS_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => NPC_ABS(31), 
                           DOUT(30) => NPC_ABS(30), DOUT(29) => NPC_ABS(29), 
                           DOUT(28) => NPC_ABS(28), DOUT(27) => NPC_ABS(27), 
                           DOUT(26) => NPC_ABS(26), DOUT(25) => NPC_ABS(25), 
                           DOUT(24) => NPC_ABS(24), DOUT(23) => NPC_ABS(23), 
                           DOUT(22) => NPC_ABS(22), DOUT(21) => NPC_ABS(21), 
                           DOUT(20) => NPC_ABS(20), DOUT(19) => NPC_ABS(19), 
                           DOUT(18) => NPC_ABS(18), DOUT(17) => NPC_ABS(17), 
                           DOUT(16) => NPC_ABS(16), DOUT(15) => NPC_ABS(15), 
                           DOUT(14) => NPC_ABS(14), DOUT(13) => NPC_ABS(13), 
                           DOUT(12) => NPC_ABS(12), DOUT(11) => NPC_ABS(11), 
                           DOUT(10) => NPC_ABS(10), DOUT(9) => NPC_ABS(9), 
                           DOUT(8) => NPC_ABS(8), DOUT(7) => NPC_ABS(7), 
                           DOUT(6) => NPC_ABS(6), DOUT(5) => NPC_ABS(5), 
                           DOUT(4) => NPC_ABS(4), DOUT(3) => NPC_ABS(3), 
                           DOUT(2) => NPC_ABS(2), DOUT(1) => NPC_ABS(1), 
                           DOUT(0) => NPC_ABS(0));
   NPC_REL_reg : regn_N32_2 port map( DIN(31) => sig_NPC_REL_31_port, DIN(30) 
                           => sig_NPC_REL_30_port, DIN(29) => 
                           sig_NPC_REL_29_port, DIN(28) => sig_NPC_REL_28_port,
                           DIN(27) => sig_NPC_REL_27_port, DIN(26) => 
                           sig_NPC_REL_26_port, DIN(25) => sig_NPC_REL_25_port,
                           DIN(24) => sig_NPC_REL_24_port, DIN(23) => 
                           sig_NPC_REL_23_port, DIN(22) => sig_NPC_REL_22_port,
                           DIN(21) => sig_NPC_REL_21_port, DIN(20) => 
                           sig_NPC_REL_20_port, DIN(19) => sig_NPC_REL_19_port,
                           DIN(18) => sig_NPC_REL_18_port, DIN(17) => 
                           sig_NPC_REL_17_port, DIN(16) => sig_NPC_REL_16_port,
                           DIN(15) => sig_NPC_REL_15_port, DIN(14) => 
                           sig_NPC_REL_14_port, DIN(13) => sig_NPC_REL_13_port,
                           DIN(12) => sig_NPC_REL_12_port, DIN(11) => 
                           sig_NPC_REL_11_port, DIN(10) => sig_NPC_REL_10_port,
                           DIN(9) => sig_NPC_REL_9_port, DIN(8) => 
                           sig_NPC_REL_8_port, DIN(7) => sig_NPC_REL_7_port, 
                           DIN(6) => sig_NPC_REL_6_port, DIN(5) => 
                           sig_NPC_REL_5_port, DIN(4) => sig_NPC_REL_4_port, 
                           DIN(3) => sig_NPC_REL_3_port, DIN(2) => 
                           sig_NPC_REL_2_port, DIN(1) => sig_NPC_REL_1_port, 
                           DIN(0) => sig_NPC_REL_0_port, CLK => CLK, EN => 
                           ALU_OUTREG_EN, RST => RST, DOUT(31) => NPC_REL(31), 
                           DOUT(30) => NPC_REL(30), DOUT(29) => NPC_REL(29), 
                           DOUT(28) => NPC_REL(28), DOUT(27) => NPC_REL(27), 
                           DOUT(26) => NPC_REL(26), DOUT(25) => NPC_REL(25), 
                           DOUT(24) => NPC_REL(24), DOUT(23) => NPC_REL(23), 
                           DOUT(22) => NPC_REL(22), DOUT(21) => NPC_REL(21), 
                           DOUT(20) => NPC_REL(20), DOUT(19) => NPC_REL(19), 
                           DOUT(18) => NPC_REL(18), DOUT(17) => NPC_REL(17), 
                           DOUT(16) => NPC_REL(16), DOUT(15) => NPC_REL(15), 
                           DOUT(14) => NPC_REL(14), DOUT(13) => NPC_REL(13), 
                           DOUT(12) => NPC_REL(12), DOUT(11) => NPC_REL(11), 
                           DOUT(10) => NPC_REL(10), DOUT(9) => NPC_REL(9), 
                           DOUT(8) => NPC_REL(8), DOUT(7) => NPC_REL(7), 
                           DOUT(6) => NPC_REL(6), DOUT(5) => NPC_REL(5), 
                           DOUT(4) => NPC_REL(4), DOUT(3) => NPC_REL(3), 
                           DOUT(2) => NPC_REL(2), DOUT(1) => NPC_REL(1), 
                           DOUT(0) => NPC_REL(0));
   add_1_root_add_0_root_add_122_2 : Execute_DW01_add_1 port map( A(31) => 
                           n2_port, A(30) => n2_port, A(29) => n2_port, A(28) 
                           => n2_port, A(27) => n2_port, A(26) => n2_port, 
                           A(25) => n2_port, A(24) => n2_port, A(23) => n2_port
                           , A(22) => n2_port, A(21) => n2_port, A(20) => 
                           n2_port, A(19) => n2_port, A(18) => n2_port, A(17) 
                           => n2_port, A(16) => n2_port, A(15) => n2_port, 
                           A(14) => n2_port, A(13) => n2_port, A(12) => n2_port
                           , A(11) => n2_port, A(10) => n2_port, A(9) => 
                           n2_port, A(8) => n2_port, A(7) => n2_port, A(6) => 
                           n2_port, A(5) => n2_port, A(4) => n2_port, A(3) => 
                           n2_port, A(2) => n3_port, A(1) => n2_port, A(0) => 
                           n2_port, B(31) => IMM_IN(31), B(30) => IMM_IN(30), 
                           B(29) => IMM_IN(29), B(28) => IMM_IN(28), B(27) => 
                           IMM_IN(27), B(26) => IMM_IN(26), B(25) => IMM_IN(25)
                           , B(24) => IMM_IN(24), B(23) => IMM_IN(23), B(22) =>
                           IMM_IN(22), B(21) => IMM_IN(21), B(20) => IMM_IN(20)
                           , B(19) => IMM_IN(19), B(18) => IMM_IN(18), B(17) =>
                           IMM_IN(17), B(16) => IMM_IN(16), B(15) => IMM_IN(15)
                           , B(14) => IMM_IN(14), B(13) => IMM_IN(13), B(12) =>
                           IMM_IN(12), B(11) => IMM_IN(11), B(10) => IMM_IN(10)
                           , B(9) => IMM_IN(9), B(8) => IMM_IN(8), B(7) => 
                           IMM_IN(7), B(6) => IMM_IN(6), B(5) => IMM_IN(5), 
                           B(4) => IMM_IN(4), B(3) => IMM_IN(3), B(2) => 
                           IMM_IN(2), B(1) => IMM_IN(1), B(0) => IMM_IN(0), CI 
                           => n4_port, SUM(31) => N31, SUM(30) => N30, SUM(29) 
                           => N29, SUM(28) => N28, SUM(27) => N27, SUM(26) => 
                           N26, SUM(25) => N25, SUM(24) => N24, SUM(23) => N23,
                           SUM(22) => N22, SUM(21) => N21, SUM(20) => N20, 
                           SUM(19) => N19, SUM(18) => N18, SUM(17) => N17, 
                           SUM(16) => N16, SUM(15) => N15, SUM(14) => N14, 
                           SUM(13) => N13, SUM(12) => N12, SUM(11) => N11, 
                           SUM(10) => N10, SUM(9) => N9, SUM(8) => N8, SUM(7) 
                           => N7, SUM(6) => N6, SUM(5) => N5, SUM(4) => N4, 
                           SUM(3) => N3, SUM(2) => N2, SUM(1) => N1, SUM(0) => 
                           N0, CO => n_1983);
   add_0_root_add_0_root_add_122_2 : Execute_DW01_add_0 port map( A(31) => 
                           PC_IN(31), A(30) => PC_IN(30), A(29) => PC_IN(29), 
                           A(28) => PC_IN(28), A(27) => PC_IN(27), A(26) => 
                           PC_IN(26), A(25) => PC_IN(25), A(24) => PC_IN(24), 
                           A(23) => PC_IN(23), A(22) => PC_IN(22), A(21) => 
                           PC_IN(21), A(20) => PC_IN(20), A(19) => PC_IN(19), 
                           A(18) => PC_IN(18), A(17) => PC_IN(17), A(16) => 
                           PC_IN(16), A(15) => PC_IN(15), A(14) => PC_IN(14), 
                           A(13) => PC_IN(13), A(12) => PC_IN(12), A(11) => 
                           PC_IN(11), A(10) => PC_IN(10), A(9) => PC_IN(9), 
                           A(8) => PC_IN(8), A(7) => PC_IN(7), A(6) => PC_IN(6)
                           , A(5) => PC_IN(5), A(4) => PC_IN(4), A(3) => 
                           PC_IN(3), A(2) => PC_IN(2), A(1) => PC_IN(1), A(0) 
                           => PC_IN(0), B(31) => N31, B(30) => N30, B(29) => 
                           N29, B(28) => N28, B(27) => N27, B(26) => N26, B(25)
                           => N25, B(24) => N24, B(23) => N23, B(22) => N22, 
                           B(21) => N21, B(20) => N20, B(19) => N19, B(18) => 
                           N18, B(17) => N17, B(16) => N16, B(15) => N15, B(14)
                           => N14, B(13) => N13, B(12) => N12, B(11) => N11, 
                           B(10) => N10, B(9) => N9, B(8) => N8, B(7) => N7, 
                           B(6) => N6, B(5) => N5, B(4) => N4, B(3) => N3, B(2)
                           => N2, B(1) => N1, B(0) => N0, CI => n5_port, 
                           SUM(31) => sig_NPC_REL_31_port, SUM(30) => 
                           sig_NPC_REL_30_port, SUM(29) => sig_NPC_REL_29_port,
                           SUM(28) => sig_NPC_REL_28_port, SUM(27) => 
                           sig_NPC_REL_27_port, SUM(26) => sig_NPC_REL_26_port,
                           SUM(25) => sig_NPC_REL_25_port, SUM(24) => 
                           sig_NPC_REL_24_port, SUM(23) => sig_NPC_REL_23_port,
                           SUM(22) => sig_NPC_REL_22_port, SUM(21) => 
                           sig_NPC_REL_21_port, SUM(20) => sig_NPC_REL_20_port,
                           SUM(19) => sig_NPC_REL_19_port, SUM(18) => 
                           sig_NPC_REL_18_port, SUM(17) => sig_NPC_REL_17_port,
                           SUM(16) => sig_NPC_REL_16_port, SUM(15) => 
                           sig_NPC_REL_15_port, SUM(14) => sig_NPC_REL_14_port,
                           SUM(13) => sig_NPC_REL_13_port, SUM(12) => 
                           sig_NPC_REL_12_port, SUM(11) => sig_NPC_REL_11_port,
                           SUM(10) => sig_NPC_REL_10_port, SUM(9) => 
                           sig_NPC_REL_9_port, SUM(8) => sig_NPC_REL_8_port, 
                           SUM(7) => sig_NPC_REL_7_port, SUM(6) => 
                           sig_NPC_REL_6_port, SUM(5) => sig_NPC_REL_5_port, 
                           SUM(4) => sig_NPC_REL_4_port, SUM(3) => 
                           sig_NPC_REL_3_port, SUM(2) => sig_NPC_REL_2_port, 
                           SUM(1) => sig_NPC_REL_1_port, SUM(0) => 
                           sig_NPC_REL_0_port, CO => n_1984);
   U3 : NOR2_X1 port map( A1 => ZERO_FLAG_port, A2 => n1_port, ZN => sig_RST);
   U4 : INV_X1 port map( A => RST, ZN => n1_port);
   n2_port <= '0';
   n3_port <= '1';
   n4_port <= '0';
   n5_port <= '0';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Decode is

   port( CLK, RST, Bubble, RF_WE, ZERO_FLAG : in std_logic;  PC_IN, INS_IN : in
         std_logic_vector (31 downto 0);  ADD_WR : in std_logic_vector (4 
         downto 0);  DATA_WR_IN : in std_logic_vector (31 downto 0);  PC_OUT, 
         A_OUT, B_OUT, IMM_OUT : out std_logic_vector (31 downto 0);  
         ADD_RS1_HDU, ADD_RS2_HDU, ADD_WR_OUT, ADD_RS1_OUT, ADD_RS2_OUT : out 
         std_logic_vector (4 downto 0));

end Decode;

architecture SYN_struct of Decode is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component register_file_NBIT_ADD5_NBIT_DATA32
      port( CLK, RST, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RS1, 
            ADD_RS2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component mux21_NBIT5_1
      port( A, B : in std_logic_vector (4 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component mux21_NBIT5_2
      port( A, B : in std_logic_vector (4 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component mux21_NBIT5_0
      port( A, B : in std_logic_vector (4 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N5_3
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N5_4
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N5_0
      port( DIN : in std_logic_vector (4 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (4 downto 0));
   end component;
   
   component regn_N32_6
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_7
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component instruction_decomposition
      port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype :
            in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : out std_logic_vector (4 
            downto 0);  IMM : out std_logic_vector (31 downto 0);  RD1, RD2 : 
            out std_logic);
   end component;
   
   component instruction_type
      port( INST_IN : in std_logic_vector (31 downto 0);  Rtype, Itype, Jtype :
            out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, ADD_RS1_HDU_4_port, n13, n14, n15, 
      ADD_RS1_HDU_0_port, n16, n17, n18, n19, n20, sig_RST, sig_Rtype, 
      sig_Itype, sig_Jtype, sig_ADD_WR_4_port, sig_ADD_WR_3_port, 
      sig_ADD_WR_2_port, sig_ADD_WR_1_port, sig_ADD_WR_0_port, sig_IMM_31_port,
      sig_IMM_30_port, sig_IMM_29_port, sig_IMM_28_port, sig_IMM_27_port, 
      sig_IMM_26_port, sig_IMM_25_port, sig_IMM_24_port, sig_IMM_23_port, 
      sig_IMM_22_port, sig_IMM_21_port, sig_IMM_20_port, sig_IMM_19_port, 
      sig_IMM_18_port, sig_IMM_17_port, sig_IMM_16_port, sig_IMM_15_port, 
      sig_IMM_14_port, sig_IMM_13_port, sig_IMM_12_port, sig_IMM_11_port, 
      sig_IMM_10_port, sig_IMM_9_port, sig_IMM_8_port, sig_IMM_7_port, 
      sig_IMM_6_port, sig_IMM_5_port, sig_IMM_4_port, sig_IMM_3_port, 
      sig_IMM_2_port, sig_IMM_1_port, sig_IMM_0_port, RD1, RD2, 
      sig_ADD_WRHAZ_4_port, sig_ADD_WRHAZ_3_port, sig_ADD_WRHAZ_2_port, 
      sig_ADD_WRHAZ_1_port, sig_ADD_WRHAZ_0_port, sig_ADD_RS1HAZ_4_port, 
      sig_ADD_RS1HAZ_3_port, sig_ADD_RS1HAZ_2_port, sig_ADD_RS1HAZ_1_port, 
      sig_ADD_RS1HAZ_0_port, sig_ADD_RS2HAZ_4_port, sig_ADD_RS2HAZ_3_port, 
      sig_ADD_RS2HAZ_2_port, sig_ADD_RS2HAZ_1_port, sig_ADD_RS2HAZ_0_port, 
      ADD_RS2_HDU_2_port, ADD_RS1_HDU_2_port, ADD_RS2_HDU_1_port, 
      ADD_RS1_HDU_1_port, ADD_RS2_HDU_0_port, n6, n7, ADD_RS2_HDU_4_port, 
      ADD_RS2_HDU_3_port, ADD_RS1_HDU_3_port, n11, n12 : std_logic;

begin
   ADD_RS1_HDU <= ( ADD_RS1_HDU_4_port, ADD_RS1_HDU_3_port, ADD_RS1_HDU_2_port,
      ADD_RS1_HDU_1_port, ADD_RS1_HDU_0_port );
   ADD_RS2_HDU <= ( ADD_RS2_HDU_4_port, ADD_RS2_HDU_3_port, ADD_RS2_HDU_2_port,
      ADD_RS2_HDU_1_port, ADD_RS2_HDU_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   U3 : NOR2_X2 port map( A1 => ZERO_FLAG, A2 => n12, ZN => sig_RST);
   ins_type : instruction_type port map( INST_IN(31) => INS_IN(31), INST_IN(30)
                           => INS_IN(30), INST_IN(29) => INS_IN(29), 
                           INST_IN(28) => INS_IN(28), INST_IN(27) => INS_IN(27)
                           , INST_IN(26) => INS_IN(26), INST_IN(25) => 
                           INS_IN(25), INST_IN(24) => INS_IN(24), INST_IN(23) 
                           => INS_IN(23), INST_IN(22) => INS_IN(22), 
                           INST_IN(21) => INS_IN(21), INST_IN(20) => INS_IN(20)
                           , INST_IN(19) => INS_IN(19), INST_IN(18) => 
                           INS_IN(18), INST_IN(17) => INS_IN(17), INST_IN(16) 
                           => INS_IN(16), INST_IN(15) => INS_IN(15), 
                           INST_IN(14) => INS_IN(14), INST_IN(13) => INS_IN(13)
                           , INST_IN(12) => INS_IN(12), INST_IN(11) => 
                           INS_IN(11), INST_IN(10) => INS_IN(10), INST_IN(9) =>
                           INS_IN(9), INST_IN(8) => INS_IN(8), INST_IN(7) => 
                           INS_IN(7), INST_IN(6) => INS_IN(6), INST_IN(5) => 
                           INS_IN(5), INST_IN(4) => INS_IN(4), INST_IN(3) => 
                           INS_IN(3), INST_IN(2) => INS_IN(2), INST_IN(1) => 
                           INS_IN(1), INST_IN(0) => INS_IN(0), Rtype => 
                           sig_Rtype, Itype => sig_Itype, Jtype => sig_Jtype);
   ins_dec : instruction_decomposition port map( INST_IN(31) => INS_IN(31), 
                           INST_IN(30) => n7, INST_IN(29) => n6, INST_IN(28) =>
                           INS_IN(28), INST_IN(27) => INS_IN(27), INST_IN(26) 
                           => INS_IN(26), INST_IN(25) => INS_IN(25), 
                           INST_IN(24) => INS_IN(24), INST_IN(23) => INS_IN(23)
                           , INST_IN(22) => INS_IN(22), INST_IN(21) => 
                           INS_IN(21), INST_IN(20) => INS_IN(20), INST_IN(19) 
                           => INS_IN(19), INST_IN(18) => INS_IN(18), 
                           INST_IN(17) => INS_IN(17), INST_IN(16) => INS_IN(16)
                           , INST_IN(15) => INS_IN(15), INST_IN(14) => 
                           INS_IN(14), INST_IN(13) => INS_IN(13), INST_IN(12) 
                           => INS_IN(12), INST_IN(11) => INS_IN(11), 
                           INST_IN(10) => INS_IN(10), INST_IN(9) => INS_IN(9), 
                           INST_IN(8) => INS_IN(8), INST_IN(7) => INS_IN(7), 
                           INST_IN(6) => INS_IN(6), INST_IN(5) => INS_IN(5), 
                           INST_IN(4) => INS_IN(4), INST_IN(3) => INS_IN(3), 
                           INST_IN(2) => INS_IN(2), INST_IN(1) => INS_IN(1), 
                           INST_IN(0) => INS_IN(0), Rtype => sig_Rtype, Itype 
                           => sig_Itype, Jtype => sig_Jtype, ADD_RS1(4) => 
                           ADD_RS1_HDU_4_port, ADD_RS1(3) => n13, ADD_RS1(2) =>
                           n14, ADD_RS1(1) => n15, ADD_RS1(0) => 
                           ADD_RS1_HDU_0_port, ADD_RS2(4) => n16, ADD_RS2(3) =>
                           n17, ADD_RS2(2) => n18, ADD_RS2(1) => n19, 
                           ADD_RS2(0) => n20, ADD_WR(4) => sig_ADD_WR_4_port, 
                           ADD_WR(3) => sig_ADD_WR_3_port, ADD_WR(2) => 
                           sig_ADD_WR_2_port, ADD_WR(1) => sig_ADD_WR_1_port, 
                           ADD_WR(0) => sig_ADD_WR_0_port, IMM(31) => 
                           sig_IMM_31_port, IMM(30) => sig_IMM_30_port, IMM(29)
                           => sig_IMM_29_port, IMM(28) => sig_IMM_28_port, 
                           IMM(27) => sig_IMM_27_port, IMM(26) => 
                           sig_IMM_26_port, IMM(25) => sig_IMM_25_port, IMM(24)
                           => sig_IMM_24_port, IMM(23) => sig_IMM_23_port, 
                           IMM(22) => sig_IMM_22_port, IMM(21) => 
                           sig_IMM_21_port, IMM(20) => sig_IMM_20_port, IMM(19)
                           => sig_IMM_19_port, IMM(18) => sig_IMM_18_port, 
                           IMM(17) => sig_IMM_17_port, IMM(16) => 
                           sig_IMM_16_port, IMM(15) => sig_IMM_15_port, IMM(14)
                           => sig_IMM_14_port, IMM(13) => sig_IMM_13_port, 
                           IMM(12) => sig_IMM_12_port, IMM(11) => 
                           sig_IMM_11_port, IMM(10) => sig_IMM_10_port, IMM(9) 
                           => sig_IMM_9_port, IMM(8) => sig_IMM_8_port, IMM(7) 
                           => sig_IMM_7_port, IMM(6) => sig_IMM_6_port, IMM(5) 
                           => sig_IMM_5_port, IMM(4) => sig_IMM_4_port, IMM(3) 
                           => sig_IMM_3_port, IMM(2) => sig_IMM_2_port, IMM(1) 
                           => sig_IMM_1_port, IMM(0) => sig_IMM_0_port, RD1 => 
                           RD1, RD2 => RD2);
   regPC : regn_N32_7 port map( DIN(31) => PC_IN(31), DIN(30) => PC_IN(30), 
                           DIN(29) => PC_IN(29), DIN(28) => PC_IN(28), DIN(27) 
                           => PC_IN(27), DIN(26) => PC_IN(26), DIN(25) => 
                           PC_IN(25), DIN(24) => PC_IN(24), DIN(23) => 
                           PC_IN(23), DIN(22) => PC_IN(22), DIN(21) => 
                           PC_IN(21), DIN(20) => PC_IN(20), DIN(19) => 
                           PC_IN(19), DIN(18) => PC_IN(18), DIN(17) => 
                           PC_IN(17), DIN(16) => PC_IN(16), DIN(15) => 
                           PC_IN(15), DIN(14) => PC_IN(14), DIN(13) => 
                           PC_IN(13), DIN(12) => PC_IN(12), DIN(11) => 
                           PC_IN(11), DIN(10) => PC_IN(10), DIN(9) => PC_IN(9),
                           DIN(8) => PC_IN(8), DIN(7) => PC_IN(7), DIN(6) => 
                           PC_IN(6), DIN(5) => PC_IN(5), DIN(4) => PC_IN(4), 
                           DIN(3) => PC_IN(3), DIN(2) => PC_IN(2), DIN(1) => 
                           PC_IN(1), DIN(0) => PC_IN(0), CLK => CLK, EN => 
                           X_Logic1_port, RST => sig_RST, DOUT(31) => 
                           PC_OUT(31), DOUT(30) => PC_OUT(30), DOUT(29) => 
                           PC_OUT(29), DOUT(28) => PC_OUT(28), DOUT(27) => 
                           PC_OUT(27), DOUT(26) => PC_OUT(26), DOUT(25) => 
                           PC_OUT(25), DOUT(24) => PC_OUT(24), DOUT(23) => 
                           PC_OUT(23), DOUT(22) => PC_OUT(22), DOUT(21) => 
                           PC_OUT(21), DOUT(20) => PC_OUT(20), DOUT(19) => 
                           PC_OUT(19), DOUT(18) => PC_OUT(18), DOUT(17) => 
                           PC_OUT(17), DOUT(16) => PC_OUT(16), DOUT(15) => 
                           PC_OUT(15), DOUT(14) => PC_OUT(14), DOUT(13) => 
                           PC_OUT(13), DOUT(12) => PC_OUT(12), DOUT(11) => 
                           PC_OUT(11), DOUT(10) => PC_OUT(10), DOUT(9) => 
                           PC_OUT(9), DOUT(8) => PC_OUT(8), DOUT(7) => 
                           PC_OUT(7), DOUT(6) => PC_OUT(6), DOUT(5) => 
                           PC_OUT(5), DOUT(4) => PC_OUT(4), DOUT(3) => 
                           PC_OUT(3), DOUT(2) => PC_OUT(2), DOUT(1) => 
                           PC_OUT(1), DOUT(0) => PC_OUT(0));
   regIMM : regn_N32_6 port map( DIN(31) => sig_IMM_31_port, DIN(30) => 
                           sig_IMM_30_port, DIN(29) => sig_IMM_29_port, DIN(28)
                           => sig_IMM_28_port, DIN(27) => sig_IMM_27_port, 
                           DIN(26) => sig_IMM_26_port, DIN(25) => 
                           sig_IMM_25_port, DIN(24) => sig_IMM_24_port, DIN(23)
                           => sig_IMM_23_port, DIN(22) => sig_IMM_22_port, 
                           DIN(21) => sig_IMM_21_port, DIN(20) => 
                           sig_IMM_20_port, DIN(19) => sig_IMM_19_port, DIN(18)
                           => sig_IMM_18_port, DIN(17) => sig_IMM_17_port, 
                           DIN(16) => sig_IMM_16_port, DIN(15) => 
                           sig_IMM_15_port, DIN(14) => sig_IMM_14_port, DIN(13)
                           => sig_IMM_13_port, DIN(12) => sig_IMM_12_port, 
                           DIN(11) => sig_IMM_11_port, DIN(10) => 
                           sig_IMM_10_port, DIN(9) => sig_IMM_9_port, DIN(8) =>
                           sig_IMM_8_port, DIN(7) => sig_IMM_7_port, DIN(6) => 
                           sig_IMM_6_port, DIN(5) => sig_IMM_5_port, DIN(4) => 
                           sig_IMM_4_port, DIN(3) => sig_IMM_3_port, DIN(2) => 
                           sig_IMM_2_port, DIN(1) => sig_IMM_1_port, DIN(0) => 
                           sig_IMM_0_port, CLK => CLK, EN => X_Logic1_port, RST
                           => sig_RST, DOUT(31) => IMM_OUT(31), DOUT(30) => 
                           IMM_OUT(30), DOUT(29) => IMM_OUT(29), DOUT(28) => 
                           IMM_OUT(28), DOUT(27) => IMM_OUT(27), DOUT(26) => 
                           IMM_OUT(26), DOUT(25) => IMM_OUT(25), DOUT(24) => 
                           IMM_OUT(24), DOUT(23) => IMM_OUT(23), DOUT(22) => 
                           IMM_OUT(22), DOUT(21) => IMM_OUT(21), DOUT(20) => 
                           IMM_OUT(20), DOUT(19) => IMM_OUT(19), DOUT(18) => 
                           IMM_OUT(18), DOUT(17) => IMM_OUT(17), DOUT(16) => 
                           IMM_OUT(16), DOUT(15) => IMM_OUT(15), DOUT(14) => 
                           IMM_OUT(14), DOUT(13) => IMM_OUT(13), DOUT(12) => 
                           IMM_OUT(12), DOUT(11) => IMM_OUT(11), DOUT(10) => 
                           IMM_OUT(10), DOUT(9) => IMM_OUT(9), DOUT(8) => 
                           IMM_OUT(8), DOUT(7) => IMM_OUT(7), DOUT(6) => 
                           IMM_OUT(6), DOUT(5) => IMM_OUT(5), DOUT(4) => 
                           IMM_OUT(4), DOUT(3) => IMM_OUT(3), DOUT(2) => 
                           IMM_OUT(2), DOUT(1) => IMM_OUT(1), DOUT(0) => 
                           IMM_OUT(0));
   regWR : regn_N5_0 port map( DIN(4) => sig_ADD_WRHAZ_4_port, DIN(3) => 
                           sig_ADD_WRHAZ_3_port, DIN(2) => sig_ADD_WRHAZ_2_port
                           , DIN(1) => sig_ADD_WRHAZ_1_port, DIN(0) => 
                           sig_ADD_WRHAZ_0_port, CLK => CLK, EN => 
                           X_Logic1_port, RST => sig_RST, DOUT(4) => 
                           ADD_WR_OUT(4), DOUT(3) => ADD_WR_OUT(3), DOUT(2) => 
                           ADD_WR_OUT(2), DOUT(1) => ADD_WR_OUT(1), DOUT(0) => 
                           ADD_WR_OUT(0));
   regRS1 : regn_N5_4 port map( DIN(4) => sig_ADD_RS1HAZ_4_port, DIN(3) => 
                           sig_ADD_RS1HAZ_3_port, DIN(2) => 
                           sig_ADD_RS1HAZ_2_port, DIN(1) => 
                           sig_ADD_RS1HAZ_1_port, DIN(0) => 
                           sig_ADD_RS1HAZ_0_port, CLK => CLK, EN => 
                           X_Logic1_port, RST => sig_RST, DOUT(4) => 
                           ADD_RS1_OUT(4), DOUT(3) => ADD_RS1_OUT(3), DOUT(2) 
                           => ADD_RS1_OUT(2), DOUT(1) => ADD_RS1_OUT(1), 
                           DOUT(0) => ADD_RS1_OUT(0));
   regRS2 : regn_N5_3 port map( DIN(4) => sig_ADD_RS2HAZ_4_port, DIN(3) => 
                           sig_ADD_RS2HAZ_3_port, DIN(2) => 
                           sig_ADD_RS2HAZ_2_port, DIN(1) => 
                           sig_ADD_RS2HAZ_1_port, DIN(0) => 
                           sig_ADD_RS2HAZ_0_port, CLK => CLK, EN => 
                           X_Logic1_port, RST => sig_RST, DOUT(4) => 
                           ADD_RS2_OUT(4), DOUT(3) => ADD_RS2_OUT(3), DOUT(2) 
                           => ADD_RS2_OUT(2), DOUT(1) => ADD_RS2_OUT(1), 
                           DOUT(0) => ADD_RS2_OUT(0));
   muxRS1 : mux21_NBIT5_0 port map( A(4) => ADD_RS1_HDU_4_port, A(3) => 
                           ADD_RS1_HDU_3_port, A(2) => ADD_RS1_HDU_2_port, A(1)
                           => ADD_RS1_HDU_1_port, A(0) => ADD_RS1_HDU_0_port, 
                           B(4) => X_Logic0_port, B(3) => X_Logic0_port, B(2) 
                           => X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, S => n11, Z(4) => 
                           sig_ADD_RS1HAZ_4_port, Z(3) => sig_ADD_RS1HAZ_3_port
                           , Z(2) => sig_ADD_RS1HAZ_2_port, Z(1) => 
                           sig_ADD_RS1HAZ_1_port, Z(0) => sig_ADD_RS1HAZ_0_port
                           );
   muxRS2 : mux21_NBIT5_2 port map( A(4) => ADD_RS2_HDU_4_port, A(3) => 
                           ADD_RS2_HDU_3_port, A(2) => ADD_RS2_HDU_2_port, A(1)
                           => ADD_RS2_HDU_1_port, A(0) => ADD_RS2_HDU_0_port, 
                           B(4) => X_Logic0_port, B(3) => X_Logic0_port, B(2) 
                           => X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, S => n11, Z(4) => 
                           sig_ADD_RS2HAZ_4_port, Z(3) => sig_ADD_RS2HAZ_3_port
                           , Z(2) => sig_ADD_RS2HAZ_2_port, Z(1) => 
                           sig_ADD_RS2HAZ_1_port, Z(0) => sig_ADD_RS2HAZ_0_port
                           );
   muxWR : mux21_NBIT5_1 port map( A(4) => sig_ADD_WR_4_port, A(3) => 
                           sig_ADD_WR_3_port, A(2) => sig_ADD_WR_2_port, A(1) 
                           => sig_ADD_WR_1_port, A(0) => sig_ADD_WR_0_port, 
                           B(4) => X_Logic0_port, B(3) => X_Logic0_port, B(2) 
                           => X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, S => n11, Z(4) => 
                           sig_ADD_WRHAZ_4_port, Z(3) => sig_ADD_WRHAZ_3_port, 
                           Z(2) => sig_ADD_WRHAZ_2_port, Z(1) => 
                           sig_ADD_WRHAZ_1_port, Z(0) => sig_ADD_WRHAZ_0_port);
   rf : register_file_NBIT_ADD5_NBIT_DATA32 port map( CLK => CLK, RST => RST, 
                           ENABLE => X_Logic1_port, RD1 => RD1, RD2 => RD2, WR 
                           => RF_WE, ADD_WR(4) => ADD_WR(4), ADD_WR(3) => 
                           ADD_WR(3), ADD_WR(2) => ADD_WR(2), ADD_WR(1) => 
                           ADD_WR(1), ADD_WR(0) => ADD_WR(0), ADD_RS1(4) => 
                           ADD_RS1_HDU_4_port, ADD_RS1(3) => n13, ADD_RS1(2) =>
                           n14, ADD_RS1(1) => n15, ADD_RS1(0) => 
                           ADD_RS1_HDU_0_port, ADD_RS2(4) => n16, ADD_RS2(3) =>
                           n17, ADD_RS2(2) => n18, ADD_RS2(1) => n19, 
                           ADD_RS2(0) => n20, DATAIN(31) => DATA_WR_IN(31), 
                           DATAIN(30) => DATA_WR_IN(30), DATAIN(29) => 
                           DATA_WR_IN(29), DATAIN(28) => DATA_WR_IN(28), 
                           DATAIN(27) => DATA_WR_IN(27), DATAIN(26) => 
                           DATA_WR_IN(26), DATAIN(25) => DATA_WR_IN(25), 
                           DATAIN(24) => DATA_WR_IN(24), DATAIN(23) => 
                           DATA_WR_IN(23), DATAIN(22) => DATA_WR_IN(22), 
                           DATAIN(21) => DATA_WR_IN(21), DATAIN(20) => 
                           DATA_WR_IN(20), DATAIN(19) => DATA_WR_IN(19), 
                           DATAIN(18) => DATA_WR_IN(18), DATAIN(17) => 
                           DATA_WR_IN(17), DATAIN(16) => DATA_WR_IN(16), 
                           DATAIN(15) => DATA_WR_IN(15), DATAIN(14) => 
                           DATA_WR_IN(14), DATAIN(13) => DATA_WR_IN(13), 
                           DATAIN(12) => DATA_WR_IN(12), DATAIN(11) => 
                           DATA_WR_IN(11), DATAIN(10) => DATA_WR_IN(10), 
                           DATAIN(9) => DATA_WR_IN(9), DATAIN(8) => 
                           DATA_WR_IN(8), DATAIN(7) => DATA_WR_IN(7), DATAIN(6)
                           => DATA_WR_IN(6), DATAIN(5) => DATA_WR_IN(5), 
                           DATAIN(4) => DATA_WR_IN(4), DATAIN(3) => 
                           DATA_WR_IN(3), DATAIN(2) => DATA_WR_IN(2), DATAIN(1)
                           => DATA_WR_IN(1), DATAIN(0) => DATA_WR_IN(0), 
                           OUT1(31) => A_OUT(31), OUT1(30) => A_OUT(30), 
                           OUT1(29) => A_OUT(29), OUT1(28) => A_OUT(28), 
                           OUT1(27) => A_OUT(27), OUT1(26) => A_OUT(26), 
                           OUT1(25) => A_OUT(25), OUT1(24) => A_OUT(24), 
                           OUT1(23) => A_OUT(23), OUT1(22) => A_OUT(22), 
                           OUT1(21) => A_OUT(21), OUT1(20) => A_OUT(20), 
                           OUT1(19) => A_OUT(19), OUT1(18) => A_OUT(18), 
                           OUT1(17) => A_OUT(17), OUT1(16) => A_OUT(16), 
                           OUT1(15) => A_OUT(15), OUT1(14) => A_OUT(14), 
                           OUT1(13) => A_OUT(13), OUT1(12) => A_OUT(12), 
                           OUT1(11) => A_OUT(11), OUT1(10) => A_OUT(10), 
                           OUT1(9) => A_OUT(9), OUT1(8) => A_OUT(8), OUT1(7) =>
                           A_OUT(7), OUT1(6) => A_OUT(6), OUT1(5) => A_OUT(5), 
                           OUT1(4) => A_OUT(4), OUT1(3) => A_OUT(3), OUT1(2) =>
                           A_OUT(2), OUT1(1) => A_OUT(1), OUT1(0) => A_OUT(0), 
                           OUT2(31) => B_OUT(31), OUT2(30) => B_OUT(30), 
                           OUT2(29) => B_OUT(29), OUT2(28) => B_OUT(28), 
                           OUT2(27) => B_OUT(27), OUT2(26) => B_OUT(26), 
                           OUT2(25) => B_OUT(25), OUT2(24) => B_OUT(24), 
                           OUT2(23) => B_OUT(23), OUT2(22) => B_OUT(22), 
                           OUT2(21) => B_OUT(21), OUT2(20) => B_OUT(20), 
                           OUT2(19) => B_OUT(19), OUT2(18) => B_OUT(18), 
                           OUT2(17) => B_OUT(17), OUT2(16) => B_OUT(16), 
                           OUT2(15) => B_OUT(15), OUT2(14) => B_OUT(14), 
                           OUT2(13) => B_OUT(13), OUT2(12) => B_OUT(12), 
                           OUT2(11) => B_OUT(11), OUT2(10) => B_OUT(10), 
                           OUT2(9) => B_OUT(9), OUT2(8) => B_OUT(8), OUT2(7) =>
                           B_OUT(7), OUT2(6) => B_OUT(6), OUT2(5) => B_OUT(5), 
                           OUT2(4) => B_OUT(4), OUT2(3) => B_OUT(3), OUT2(2) =>
                           B_OUT(2), OUT2(1) => B_OUT(1), OUT2(0) => B_OUT(0));
   U4 : BUF_X1 port map( A => Bubble, Z => n11);
   U5 : CLKBUF_X1 port map( A => n18, Z => ADD_RS2_HDU_2_port);
   U6 : CLKBUF_X1 port map( A => n14, Z => ADD_RS1_HDU_2_port);
   U7 : CLKBUF_X1 port map( A => n19, Z => ADD_RS2_HDU_1_port);
   U8 : CLKBUF_X1 port map( A => n15, Z => ADD_RS1_HDU_1_port);
   U9 : CLKBUF_X1 port map( A => n20, Z => ADD_RS2_HDU_0_port);
   U10 : CLKBUF_X1 port map( A => INS_IN(29), Z => n6);
   U11 : CLKBUF_X1 port map( A => INS_IN(30), Z => n7);
   U12 : CLKBUF_X1 port map( A => n16, Z => ADD_RS2_HDU_4_port);
   U13 : CLKBUF_X1 port map( A => n17, Z => ADD_RS2_HDU_3_port);
   U14 : CLKBUF_X1 port map( A => n13, Z => ADD_RS1_HDU_3_port);
   U15 : INV_X1 port map( A => RST, ZN => n12);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Fetch is

   port( CLK, RST, ZERO_FLAG : in std_logic;  PC_EXT, INS_IN : in 
         std_logic_vector (31 downto 0);  Bubble_in : in std_logic;  HDU_INS_IN
         , HDU_PC_IN, HDU_NPC_IN : in std_logic_vector (31 downto 0);  PC_OUT, 
         ADDR_OUT, NPC_OUT, INS_OUT : out std_logic_vector (31 downto 0));

end Fetch;

architecture SYN_struct of Fetch is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component Fetch_DW01_add_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component regn_N32_8
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_9
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component regn_N32_0
      port( DIN : in std_logic_vector (31 downto 0);  CLK, EN, RST : in 
            std_logic;  DOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_6
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Z : 
            out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, ADDR_OUT_31_port, ADDR_OUT_30_port, ADDR_OUT_29_port, 
      ADDR_OUT_28_port, ADDR_OUT_27_port, ADDR_OUT_26_port, ADDR_OUT_25_port, 
      ADDR_OUT_24_port, ADDR_OUT_23_port, ADDR_OUT_22_port, ADDR_OUT_21_port, 
      ADDR_OUT_20_port, ADDR_OUT_19_port, ADDR_OUT_18_port, ADDR_OUT_17_port, 
      ADDR_OUT_16_port, ADDR_OUT_15_port, ADDR_OUT_14_port, ADDR_OUT_13_port, 
      ADDR_OUT_12_port, ADDR_OUT_11_port, ADDR_OUT_10_port, ADDR_OUT_9_port, 
      ADDR_OUT_8_port, n6, ADDR_OUT_6_port, ADDR_OUT_5_port, ADDR_OUT_4_port, 
      ADDR_OUT_3_port, ADDR_OUT_2_port, ADDR_OUT_1_port, ADDR_OUT_0_port, 
      sig_RST, sig_NPC_31_port, sig_NPC_30_port, sig_NPC_29_port, 
      sig_NPC_28_port, sig_NPC_27_port, sig_NPC_26_port, sig_NPC_25_port, 
      sig_NPC_24_port, sig_NPC_23_port, sig_NPC_22_port, sig_NPC_21_port, 
      sig_NPC_20_port, sig_NPC_19_port, sig_NPC_18_port, sig_NPC_17_port, 
      sig_NPC_16_port, sig_NPC_15_port, sig_NPC_14_port, sig_NPC_13_port, 
      sig_NPC_12_port, sig_NPC_11_port, sig_NPC_10_port, sig_NPC_9_port, 
      sig_NPC_8_port, sig_NPC_7_port, sig_NPC_6_port, sig_NPC_5_port, 
      sig_NPC_4_port, sig_NPC_3_port, sig_NPC_2_port, sig_NPC_1_port, 
      sig_NPC_0_port, PC_MUX_OUT_31_port, PC_MUX_OUT_30_port, 
      PC_MUX_OUT_29_port, PC_MUX_OUT_28_port, PC_MUX_OUT_27_port, 
      PC_MUX_OUT_26_port, PC_MUX_OUT_25_port, PC_MUX_OUT_24_port, 
      PC_MUX_OUT_23_port, PC_MUX_OUT_22_port, PC_MUX_OUT_21_port, 
      PC_MUX_OUT_20_port, PC_MUX_OUT_19_port, PC_MUX_OUT_18_port, 
      PC_MUX_OUT_17_port, PC_MUX_OUT_16_port, PC_MUX_OUT_15_port, 
      PC_MUX_OUT_14_port, PC_MUX_OUT_13_port, PC_MUX_OUT_12_port, 
      PC_MUX_OUT_11_port, PC_MUX_OUT_10_port, PC_MUX_OUT_9_port, 
      PC_MUX_OUT_8_port, PC_MUX_OUT_7_port, PC_MUX_OUT_6_port, 
      PC_MUX_OUT_5_port, PC_MUX_OUT_4_port, PC_MUX_OUT_3_port, 
      PC_MUX_OUT_2_port, PC_MUX_OUT_1_port, PC_MUX_OUT_0_port, sig_INS_31_port,
      sig_INS_30_port, sig_INS_29_port, sig_INS_28_port, sig_INS_27_port, 
      sig_INS_26_port, sig_INS_25_port, sig_INS_24_port, sig_INS_23_port, 
      sig_INS_22_port, sig_INS_21_port, sig_INS_20_port, sig_INS_19_port, 
      sig_INS_18_port, sig_INS_17_port, sig_INS_16_port, sig_INS_15_port, 
      sig_INS_14_port, sig_INS_13_port, sig_INS_12_port, sig_INS_11_port, 
      sig_INS_10_port, sig_INS_9_port, sig_INS_8_port, sig_INS_7_port, 
      sig_INS_6_port, sig_INS_5_port, sig_INS_4_port, sig_INS_3_port, 
      sig_INS_2_port, sig_INS_1_port, sig_INS_0_port, n1, n2, n3, 
      ADDR_OUT_7_port, n5, n_1985 : std_logic;

begin
   ADDR_OUT <= ( ADDR_OUT_31_port, ADDR_OUT_30_port, ADDR_OUT_29_port, 
      ADDR_OUT_28_port, ADDR_OUT_27_port, ADDR_OUT_26_port, ADDR_OUT_25_port, 
      ADDR_OUT_24_port, ADDR_OUT_23_port, ADDR_OUT_22_port, ADDR_OUT_21_port, 
      ADDR_OUT_20_port, ADDR_OUT_19_port, ADDR_OUT_18_port, ADDR_OUT_17_port, 
      ADDR_OUT_16_port, ADDR_OUT_15_port, ADDR_OUT_14_port, ADDR_OUT_13_port, 
      ADDR_OUT_12_port, ADDR_OUT_11_port, ADDR_OUT_10_port, ADDR_OUT_9_port, 
      ADDR_OUT_8_port, ADDR_OUT_7_port, ADDR_OUT_6_port, ADDR_OUT_5_port, 
      ADDR_OUT_4_port, ADDR_OUT_3_port, ADDR_OUT_2_port, ADDR_OUT_1_port, 
      ADDR_OUT_0_port );
   
   X_Logic1_port <= '1';
   n1 <= '0';
   n2 <= '1';
   n3 <= '0';
   NPC_or_NPC_HDU : mux21_NBIT32_0 port map( A(31) => PC_EXT(31), A(30) => 
                           PC_EXT(30), A(29) => PC_EXT(29), A(28) => PC_EXT(28)
                           , A(27) => PC_EXT(27), A(26) => PC_EXT(26), A(25) =>
                           PC_EXT(25), A(24) => PC_EXT(24), A(23) => PC_EXT(23)
                           , A(22) => PC_EXT(22), A(21) => PC_EXT(21), A(20) =>
                           PC_EXT(20), A(19) => PC_EXT(19), A(18) => PC_EXT(18)
                           , A(17) => PC_EXT(17), A(16) => PC_EXT(16), A(15) =>
                           PC_EXT(15), A(14) => PC_EXT(14), A(13) => PC_EXT(13)
                           , A(12) => PC_EXT(12), A(11) => PC_EXT(11), A(10) =>
                           PC_EXT(10), A(9) => PC_EXT(9), A(8) => PC_EXT(8), 
                           A(7) => PC_EXT(7), A(6) => PC_EXT(6), A(5) => 
                           PC_EXT(5), A(4) => PC_EXT(4), A(3) => PC_EXT(3), 
                           A(2) => PC_EXT(2), A(1) => PC_EXT(1), A(0) => 
                           PC_EXT(0), B(31) => HDU_NPC_IN(31), B(30) => 
                           HDU_NPC_IN(30), B(29) => HDU_NPC_IN(29), B(28) => 
                           HDU_NPC_IN(28), B(27) => HDU_NPC_IN(27), B(26) => 
                           HDU_NPC_IN(26), B(25) => HDU_NPC_IN(25), B(24) => 
                           HDU_NPC_IN(24), B(23) => HDU_NPC_IN(23), B(22) => 
                           HDU_NPC_IN(22), B(21) => HDU_NPC_IN(21), B(20) => 
                           HDU_NPC_IN(20), B(19) => HDU_NPC_IN(19), B(18) => 
                           HDU_NPC_IN(18), B(17) => HDU_NPC_IN(17), B(16) => 
                           HDU_NPC_IN(16), B(15) => HDU_NPC_IN(15), B(14) => 
                           HDU_NPC_IN(14), B(13) => HDU_NPC_IN(13), B(12) => 
                           HDU_NPC_IN(12), B(11) => HDU_NPC_IN(11), B(10) => 
                           HDU_NPC_IN(10), B(9) => HDU_NPC_IN(9), B(8) => 
                           HDU_NPC_IN(8), B(7) => HDU_NPC_IN(7), B(6) => 
                           HDU_NPC_IN(6), B(5) => HDU_NPC_IN(5), B(4) => 
                           HDU_NPC_IN(4), B(3) => HDU_NPC_IN(3), B(2) => 
                           HDU_NPC_IN(2), B(1) => HDU_NPC_IN(1), B(0) => 
                           HDU_NPC_IN(0), S => Bubble_in, Z(31) => 
                           sig_NPC_31_port, Z(30) => sig_NPC_30_port, Z(29) => 
                           sig_NPC_29_port, Z(28) => sig_NPC_28_port, Z(27) => 
                           sig_NPC_27_port, Z(26) => sig_NPC_26_port, Z(25) => 
                           sig_NPC_25_port, Z(24) => sig_NPC_24_port, Z(23) => 
                           sig_NPC_23_port, Z(22) => sig_NPC_22_port, Z(21) => 
                           sig_NPC_21_port, Z(20) => sig_NPC_20_port, Z(19) => 
                           sig_NPC_19_port, Z(18) => sig_NPC_18_port, Z(17) => 
                           sig_NPC_17_port, Z(16) => sig_NPC_16_port, Z(15) => 
                           sig_NPC_15_port, Z(14) => sig_NPC_14_port, Z(13) => 
                           sig_NPC_13_port, Z(12) => sig_NPC_12_port, Z(11) => 
                           sig_NPC_11_port, Z(10) => sig_NPC_10_port, Z(9) => 
                           sig_NPC_9_port, Z(8) => sig_NPC_8_port, Z(7) => 
                           sig_NPC_7_port, Z(6) => sig_NPC_6_port, Z(5) => 
                           sig_NPC_5_port, Z(4) => sig_NPC_4_port, Z(3) => 
                           sig_NPC_3_port, Z(2) => sig_NPC_2_port, Z(1) => 
                           sig_NPC_1_port, Z(0) => sig_NPC_0_port);
   PC_or_PC_HDU : mux21_NBIT32_6 port map( A(31) => ADDR_OUT_31_port, A(30) => 
                           ADDR_OUT_30_port, A(29) => ADDR_OUT_29_port, A(28) 
                           => ADDR_OUT_28_port, A(27) => ADDR_OUT_27_port, 
                           A(26) => ADDR_OUT_26_port, A(25) => ADDR_OUT_25_port
                           , A(24) => ADDR_OUT_24_port, A(23) => 
                           ADDR_OUT_23_port, A(22) => ADDR_OUT_22_port, A(21) 
                           => ADDR_OUT_21_port, A(20) => ADDR_OUT_20_port, 
                           A(19) => ADDR_OUT_19_port, A(18) => ADDR_OUT_18_port
                           , A(17) => ADDR_OUT_17_port, A(16) => 
                           ADDR_OUT_16_port, A(15) => ADDR_OUT_15_port, A(14) 
                           => ADDR_OUT_14_port, A(13) => ADDR_OUT_13_port, 
                           A(12) => ADDR_OUT_12_port, A(11) => ADDR_OUT_11_port
                           , A(10) => ADDR_OUT_10_port, A(9) => ADDR_OUT_9_port
                           , A(8) => ADDR_OUT_8_port, A(7) => ADDR_OUT_7_port, 
                           A(6) => ADDR_OUT_6_port, A(5) => ADDR_OUT_5_port, 
                           A(4) => ADDR_OUT_4_port, A(3) => ADDR_OUT_3_port, 
                           A(2) => ADDR_OUT_2_port, A(1) => ADDR_OUT_1_port, 
                           A(0) => ADDR_OUT_0_port, B(31) => HDU_PC_IN(31), 
                           B(30) => HDU_PC_IN(30), B(29) => HDU_PC_IN(29), 
                           B(28) => HDU_PC_IN(28), B(27) => HDU_PC_IN(27), 
                           B(26) => HDU_PC_IN(26), B(25) => HDU_PC_IN(25), 
                           B(24) => HDU_PC_IN(24), B(23) => HDU_PC_IN(23), 
                           B(22) => HDU_PC_IN(22), B(21) => HDU_PC_IN(21), 
                           B(20) => HDU_PC_IN(20), B(19) => HDU_PC_IN(19), 
                           B(18) => HDU_PC_IN(18), B(17) => HDU_PC_IN(17), 
                           B(16) => HDU_PC_IN(16), B(15) => HDU_PC_IN(15), 
                           B(14) => HDU_PC_IN(14), B(13) => HDU_PC_IN(13), 
                           B(12) => HDU_PC_IN(12), B(11) => HDU_PC_IN(11), 
                           B(10) => HDU_PC_IN(10), B(9) => HDU_PC_IN(9), B(8) 
                           => HDU_PC_IN(8), B(7) => HDU_PC_IN(7), B(6) => 
                           HDU_PC_IN(6), B(5) => HDU_PC_IN(5), B(4) => 
                           HDU_PC_IN(4), B(3) => HDU_PC_IN(3), B(2) => 
                           HDU_PC_IN(2), B(1) => HDU_PC_IN(1), B(0) => 
                           HDU_PC_IN(0), S => Bubble_in, Z(31) => 
                           PC_MUX_OUT_31_port, Z(30) => PC_MUX_OUT_30_port, 
                           Z(29) => PC_MUX_OUT_29_port, Z(28) => 
                           PC_MUX_OUT_28_port, Z(27) => PC_MUX_OUT_27_port, 
                           Z(26) => PC_MUX_OUT_26_port, Z(25) => 
                           PC_MUX_OUT_25_port, Z(24) => PC_MUX_OUT_24_port, 
                           Z(23) => PC_MUX_OUT_23_port, Z(22) => 
                           PC_MUX_OUT_22_port, Z(21) => PC_MUX_OUT_21_port, 
                           Z(20) => PC_MUX_OUT_20_port, Z(19) => 
                           PC_MUX_OUT_19_port, Z(18) => PC_MUX_OUT_18_port, 
                           Z(17) => PC_MUX_OUT_17_port, Z(16) => 
                           PC_MUX_OUT_16_port, Z(15) => PC_MUX_OUT_15_port, 
                           Z(14) => PC_MUX_OUT_14_port, Z(13) => 
                           PC_MUX_OUT_13_port, Z(12) => PC_MUX_OUT_12_port, 
                           Z(11) => PC_MUX_OUT_11_port, Z(10) => 
                           PC_MUX_OUT_10_port, Z(9) => PC_MUX_OUT_9_port, Z(8) 
                           => PC_MUX_OUT_8_port, Z(7) => PC_MUX_OUT_7_port, 
                           Z(6) => PC_MUX_OUT_6_port, Z(5) => PC_MUX_OUT_5_port
                           , Z(4) => PC_MUX_OUT_4_port, Z(3) => 
                           PC_MUX_OUT_3_port, Z(2) => PC_MUX_OUT_2_port, Z(1) 
                           => PC_MUX_OUT_1_port, Z(0) => PC_MUX_OUT_0_port);
   INS_or_HDU_INS : mux21_NBIT32_5 port map( A(31) => INS_IN(31), A(30) => 
                           INS_IN(30), A(29) => INS_IN(29), A(28) => INS_IN(28)
                           , A(27) => INS_IN(27), A(26) => INS_IN(26), A(25) =>
                           INS_IN(25), A(24) => INS_IN(24), A(23) => INS_IN(23)
                           , A(22) => INS_IN(22), A(21) => INS_IN(21), A(20) =>
                           INS_IN(20), A(19) => INS_IN(19), A(18) => INS_IN(18)
                           , A(17) => INS_IN(17), A(16) => INS_IN(16), A(15) =>
                           INS_IN(15), A(14) => INS_IN(14), A(13) => INS_IN(13)
                           , A(12) => INS_IN(12), A(11) => INS_IN(11), A(10) =>
                           INS_IN(10), A(9) => INS_IN(9), A(8) => INS_IN(8), 
                           A(7) => INS_IN(7), A(6) => INS_IN(6), A(5) => 
                           INS_IN(5), A(4) => INS_IN(4), A(3) => INS_IN(3), 
                           A(2) => INS_IN(2), A(1) => INS_IN(1), A(0) => 
                           INS_IN(0), B(31) => HDU_INS_IN(31), B(30) => 
                           HDU_INS_IN(30), B(29) => HDU_INS_IN(29), B(28) => 
                           HDU_INS_IN(28), B(27) => HDU_INS_IN(27), B(26) => 
                           HDU_INS_IN(26), B(25) => HDU_INS_IN(25), B(24) => 
                           HDU_INS_IN(24), B(23) => HDU_INS_IN(23), B(22) => 
                           HDU_INS_IN(22), B(21) => HDU_INS_IN(21), B(20) => 
                           HDU_INS_IN(20), B(19) => HDU_INS_IN(19), B(18) => 
                           HDU_INS_IN(18), B(17) => HDU_INS_IN(17), B(16) => 
                           HDU_INS_IN(16), B(15) => HDU_INS_IN(15), B(14) => 
                           HDU_INS_IN(14), B(13) => HDU_INS_IN(13), B(12) => 
                           HDU_INS_IN(12), B(11) => HDU_INS_IN(11), B(10) => 
                           HDU_INS_IN(10), B(9) => HDU_INS_IN(9), B(8) => 
                           HDU_INS_IN(8), B(7) => HDU_INS_IN(7), B(6) => 
                           HDU_INS_IN(6), B(5) => HDU_INS_IN(5), B(4) => 
                           HDU_INS_IN(4), B(3) => HDU_INS_IN(3), B(2) => 
                           HDU_INS_IN(2), B(1) => HDU_INS_IN(1), B(0) => 
                           HDU_INS_IN(0), S => Bubble_in, Z(31) => 
                           sig_INS_31_port, Z(30) => sig_INS_30_port, Z(29) => 
                           sig_INS_29_port, Z(28) => sig_INS_28_port, Z(27) => 
                           sig_INS_27_port, Z(26) => sig_INS_26_port, Z(25) => 
                           sig_INS_25_port, Z(24) => sig_INS_24_port, Z(23) => 
                           sig_INS_23_port, Z(22) => sig_INS_22_port, Z(21) => 
                           sig_INS_21_port, Z(20) => sig_INS_20_port, Z(19) => 
                           sig_INS_19_port, Z(18) => sig_INS_18_port, Z(17) => 
                           sig_INS_17_port, Z(16) => sig_INS_16_port, Z(15) => 
                           sig_INS_15_port, Z(14) => sig_INS_14_port, Z(13) => 
                           sig_INS_13_port, Z(12) => sig_INS_12_port, Z(11) => 
                           sig_INS_11_port, Z(10) => sig_INS_10_port, Z(9) => 
                           sig_INS_9_port, Z(8) => sig_INS_8_port, Z(7) => 
                           sig_INS_7_port, Z(6) => sig_INS_6_port, Z(5) => 
                           sig_INS_5_port, Z(4) => sig_INS_4_port, Z(3) => 
                           sig_INS_3_port, Z(2) => sig_INS_2_port, Z(1) => 
                           sig_INS_1_port, Z(0) => sig_INS_0_port);
   PC : regn_N32_0 port map( DIN(31) => sig_NPC_31_port, DIN(30) => 
                           sig_NPC_30_port, DIN(29) => sig_NPC_29_port, DIN(28)
                           => sig_NPC_28_port, DIN(27) => sig_NPC_27_port, 
                           DIN(26) => sig_NPC_26_port, DIN(25) => 
                           sig_NPC_25_port, DIN(24) => sig_NPC_24_port, DIN(23)
                           => sig_NPC_23_port, DIN(22) => sig_NPC_22_port, 
                           DIN(21) => sig_NPC_21_port, DIN(20) => 
                           sig_NPC_20_port, DIN(19) => sig_NPC_19_port, DIN(18)
                           => sig_NPC_18_port, DIN(17) => sig_NPC_17_port, 
                           DIN(16) => sig_NPC_16_port, DIN(15) => 
                           sig_NPC_15_port, DIN(14) => sig_NPC_14_port, DIN(13)
                           => sig_NPC_13_port, DIN(12) => sig_NPC_12_port, 
                           DIN(11) => sig_NPC_11_port, DIN(10) => 
                           sig_NPC_10_port, DIN(9) => sig_NPC_9_port, DIN(8) =>
                           sig_NPC_8_port, DIN(7) => sig_NPC_7_port, DIN(6) => 
                           sig_NPC_6_port, DIN(5) => sig_NPC_5_port, DIN(4) => 
                           sig_NPC_4_port, DIN(3) => sig_NPC_3_port, DIN(2) => 
                           sig_NPC_2_port, DIN(1) => sig_NPC_1_port, DIN(0) => 
                           sig_NPC_0_port, CLK => CLK, EN => X_Logic1_port, RST
                           => RST, DOUT(31) => ADDR_OUT_31_port, DOUT(30) => 
                           ADDR_OUT_30_port, DOUT(29) => ADDR_OUT_29_port, 
                           DOUT(28) => ADDR_OUT_28_port, DOUT(27) => 
                           ADDR_OUT_27_port, DOUT(26) => ADDR_OUT_26_port, 
                           DOUT(25) => ADDR_OUT_25_port, DOUT(24) => 
                           ADDR_OUT_24_port, DOUT(23) => ADDR_OUT_23_port, 
                           DOUT(22) => ADDR_OUT_22_port, DOUT(21) => 
                           ADDR_OUT_21_port, DOUT(20) => ADDR_OUT_20_port, 
                           DOUT(19) => ADDR_OUT_19_port, DOUT(18) => 
                           ADDR_OUT_18_port, DOUT(17) => ADDR_OUT_17_port, 
                           DOUT(16) => ADDR_OUT_16_port, DOUT(15) => 
                           ADDR_OUT_15_port, DOUT(14) => ADDR_OUT_14_port, 
                           DOUT(13) => ADDR_OUT_13_port, DOUT(12) => 
                           ADDR_OUT_12_port, DOUT(11) => ADDR_OUT_11_port, 
                           DOUT(10) => ADDR_OUT_10_port, DOUT(9) => 
                           ADDR_OUT_9_port, DOUT(8) => ADDR_OUT_8_port, DOUT(7)
                           => n6, DOUT(6) => ADDR_OUT_6_port, DOUT(5) => 
                           ADDR_OUT_5_port, DOUT(4) => ADDR_OUT_4_port, DOUT(3)
                           => ADDR_OUT_3_port, DOUT(2) => ADDR_OUT_2_port, 
                           DOUT(1) => ADDR_OUT_1_port, DOUT(0) => 
                           ADDR_OUT_0_port);
   PC_reg : regn_N32_9 port map( DIN(31) => PC_MUX_OUT_31_port, DIN(30) => 
                           PC_MUX_OUT_30_port, DIN(29) => PC_MUX_OUT_29_port, 
                           DIN(28) => PC_MUX_OUT_28_port, DIN(27) => 
                           PC_MUX_OUT_27_port, DIN(26) => PC_MUX_OUT_26_port, 
                           DIN(25) => PC_MUX_OUT_25_port, DIN(24) => 
                           PC_MUX_OUT_24_port, DIN(23) => PC_MUX_OUT_23_port, 
                           DIN(22) => PC_MUX_OUT_22_port, DIN(21) => 
                           PC_MUX_OUT_21_port, DIN(20) => PC_MUX_OUT_20_port, 
                           DIN(19) => PC_MUX_OUT_19_port, DIN(18) => 
                           PC_MUX_OUT_18_port, DIN(17) => PC_MUX_OUT_17_port, 
                           DIN(16) => PC_MUX_OUT_16_port, DIN(15) => 
                           PC_MUX_OUT_15_port, DIN(14) => PC_MUX_OUT_14_port, 
                           DIN(13) => PC_MUX_OUT_13_port, DIN(12) => 
                           PC_MUX_OUT_12_port, DIN(11) => PC_MUX_OUT_11_port, 
                           DIN(10) => PC_MUX_OUT_10_port, DIN(9) => 
                           PC_MUX_OUT_9_port, DIN(8) => PC_MUX_OUT_8_port, 
                           DIN(7) => PC_MUX_OUT_7_port, DIN(6) => 
                           PC_MUX_OUT_6_port, DIN(5) => PC_MUX_OUT_5_port, 
                           DIN(4) => PC_MUX_OUT_4_port, DIN(3) => 
                           PC_MUX_OUT_3_port, DIN(2) => PC_MUX_OUT_2_port, 
                           DIN(1) => PC_MUX_OUT_1_port, DIN(0) => 
                           PC_MUX_OUT_0_port, CLK => CLK, EN => X_Logic1_port, 
                           RST => sig_RST, DOUT(31) => PC_OUT(31), DOUT(30) => 
                           PC_OUT(30), DOUT(29) => PC_OUT(29), DOUT(28) => 
                           PC_OUT(28), DOUT(27) => PC_OUT(27), DOUT(26) => 
                           PC_OUT(26), DOUT(25) => PC_OUT(25), DOUT(24) => 
                           PC_OUT(24), DOUT(23) => PC_OUT(23), DOUT(22) => 
                           PC_OUT(22), DOUT(21) => PC_OUT(21), DOUT(20) => 
                           PC_OUT(20), DOUT(19) => PC_OUT(19), DOUT(18) => 
                           PC_OUT(18), DOUT(17) => PC_OUT(17), DOUT(16) => 
                           PC_OUT(16), DOUT(15) => PC_OUT(15), DOUT(14) => 
                           PC_OUT(14), DOUT(13) => PC_OUT(13), DOUT(12) => 
                           PC_OUT(12), DOUT(11) => PC_OUT(11), DOUT(10) => 
                           PC_OUT(10), DOUT(9) => PC_OUT(9), DOUT(8) => 
                           PC_OUT(8), DOUT(7) => PC_OUT(7), DOUT(6) => 
                           PC_OUT(6), DOUT(5) => PC_OUT(5), DOUT(4) => 
                           PC_OUT(4), DOUT(3) => PC_OUT(3), DOUT(2) => 
                           PC_OUT(2), DOUT(1) => PC_OUT(1), DOUT(0) => 
                           PC_OUT(0));
   IR : regn_N32_8 port map( DIN(31) => sig_INS_31_port, DIN(30) => 
                           sig_INS_30_port, DIN(29) => sig_INS_29_port, DIN(28)
                           => sig_INS_28_port, DIN(27) => sig_INS_27_port, 
                           DIN(26) => sig_INS_26_port, DIN(25) => 
                           sig_INS_25_port, DIN(24) => sig_INS_24_port, DIN(23)
                           => sig_INS_23_port, DIN(22) => sig_INS_22_port, 
                           DIN(21) => sig_INS_21_port, DIN(20) => 
                           sig_INS_20_port, DIN(19) => sig_INS_19_port, DIN(18)
                           => sig_INS_18_port, DIN(17) => sig_INS_17_port, 
                           DIN(16) => sig_INS_16_port, DIN(15) => 
                           sig_INS_15_port, DIN(14) => sig_INS_14_port, DIN(13)
                           => sig_INS_13_port, DIN(12) => sig_INS_12_port, 
                           DIN(11) => sig_INS_11_port, DIN(10) => 
                           sig_INS_10_port, DIN(9) => sig_INS_9_port, DIN(8) =>
                           sig_INS_8_port, DIN(7) => sig_INS_7_port, DIN(6) => 
                           sig_INS_6_port, DIN(5) => sig_INS_5_port, DIN(4) => 
                           sig_INS_4_port, DIN(3) => sig_INS_3_port, DIN(2) => 
                           sig_INS_2_port, DIN(1) => sig_INS_1_port, DIN(0) => 
                           sig_INS_0_port, CLK => CLK, EN => X_Logic1_port, RST
                           => sig_RST, DOUT(31) => INS_OUT(31), DOUT(30) => 
                           INS_OUT(30), DOUT(29) => INS_OUT(29), DOUT(28) => 
                           INS_OUT(28), DOUT(27) => INS_OUT(27), DOUT(26) => 
                           INS_OUT(26), DOUT(25) => INS_OUT(25), DOUT(24) => 
                           INS_OUT(24), DOUT(23) => INS_OUT(23), DOUT(22) => 
                           INS_OUT(22), DOUT(21) => INS_OUT(21), DOUT(20) => 
                           INS_OUT(20), DOUT(19) => INS_OUT(19), DOUT(18) => 
                           INS_OUT(18), DOUT(17) => INS_OUT(17), DOUT(16) => 
                           INS_OUT(16), DOUT(15) => INS_OUT(15), DOUT(14) => 
                           INS_OUT(14), DOUT(13) => INS_OUT(13), DOUT(12) => 
                           INS_OUT(12), DOUT(11) => INS_OUT(11), DOUT(10) => 
                           INS_OUT(10), DOUT(9) => INS_OUT(9), DOUT(8) => 
                           INS_OUT(8), DOUT(7) => INS_OUT(7), DOUT(6) => 
                           INS_OUT(6), DOUT(5) => INS_OUT(5), DOUT(4) => 
                           INS_OUT(4), DOUT(3) => INS_OUT(3), DOUT(2) => 
                           INS_OUT(2), DOUT(1) => INS_OUT(1), DOUT(0) => 
                           INS_OUT(0));
   add_54 : Fetch_DW01_add_1 port map( A(31) => ADDR_OUT_31_port, A(30) => 
                           ADDR_OUT_30_port, A(29) => ADDR_OUT_29_port, A(28) 
                           => ADDR_OUT_28_port, A(27) => ADDR_OUT_27_port, 
                           A(26) => ADDR_OUT_26_port, A(25) => ADDR_OUT_25_port
                           , A(24) => ADDR_OUT_24_port, A(23) => 
                           ADDR_OUT_23_port, A(22) => ADDR_OUT_22_port, A(21) 
                           => ADDR_OUT_21_port, A(20) => ADDR_OUT_20_port, 
                           A(19) => ADDR_OUT_19_port, A(18) => ADDR_OUT_18_port
                           , A(17) => ADDR_OUT_17_port, A(16) => 
                           ADDR_OUT_16_port, A(15) => ADDR_OUT_15_port, A(14) 
                           => ADDR_OUT_14_port, A(13) => ADDR_OUT_13_port, 
                           A(12) => ADDR_OUT_12_port, A(11) => ADDR_OUT_11_port
                           , A(10) => ADDR_OUT_10_port, A(9) => ADDR_OUT_9_port
                           , A(8) => ADDR_OUT_8_port, A(7) => n6, A(6) => 
                           ADDR_OUT_6_port, A(5) => ADDR_OUT_5_port, A(4) => 
                           ADDR_OUT_4_port, A(3) => ADDR_OUT_3_port, A(2) => 
                           ADDR_OUT_2_port, A(1) => ADDR_OUT_1_port, A(0) => 
                           ADDR_OUT_0_port, B(31) => n1, B(30) => n1, B(29) => 
                           n1, B(28) => n1, B(27) => n1, B(26) => n1, B(25) => 
                           n1, B(24) => n1, B(23) => n1, B(22) => n1, B(21) => 
                           n1, B(20) => n1, B(19) => n1, B(18) => n1, B(17) => 
                           n1, B(16) => n1, B(15) => n1, B(14) => n1, B(13) => 
                           n1, B(12) => n1, B(11) => n1, B(10) => n1, B(9) => 
                           n1, B(8) => n1, B(7) => n1, B(6) => n1, B(5) => n1, 
                           B(4) => n1, B(3) => n1, B(2) => n2, B(1) => n1, B(0)
                           => n1, CI => n3, SUM(31) => NPC_OUT(31), SUM(30) => 
                           NPC_OUT(30), SUM(29) => NPC_OUT(29), SUM(28) => 
                           NPC_OUT(28), SUM(27) => NPC_OUT(27), SUM(26) => 
                           NPC_OUT(26), SUM(25) => NPC_OUT(25), SUM(24) => 
                           NPC_OUT(24), SUM(23) => NPC_OUT(23), SUM(22) => 
                           NPC_OUT(22), SUM(21) => NPC_OUT(21), SUM(20) => 
                           NPC_OUT(20), SUM(19) => NPC_OUT(19), SUM(18) => 
                           NPC_OUT(18), SUM(17) => NPC_OUT(17), SUM(16) => 
                           NPC_OUT(16), SUM(15) => NPC_OUT(15), SUM(14) => 
                           NPC_OUT(14), SUM(13) => NPC_OUT(13), SUM(12) => 
                           NPC_OUT(12), SUM(11) => NPC_OUT(11), SUM(10) => 
                           NPC_OUT(10), SUM(9) => NPC_OUT(9), SUM(8) => 
                           NPC_OUT(8), SUM(7) => NPC_OUT(7), SUM(6) => 
                           NPC_OUT(6), SUM(5) => NPC_OUT(5), SUM(4) => 
                           NPC_OUT(4), SUM(3) => NPC_OUT(3), SUM(2) => 
                           NPC_OUT(2), SUM(1) => NPC_OUT(1), SUM(0) => 
                           NPC_OUT(0), CO => n_1985);
   U6 : NOR2_X1 port map( A1 => ZERO_FLAG, A2 => n5, ZN => sig_RST);
   U7 : CLKBUF_X1 port map( A => n6, Z => ADDR_OUT_7_port);
   U8 : INV_X1 port map( A => RST, ZN => n5);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity hardwired_cu_NBIT32 is

   port( MUX_A_SEL : out std_logic;  MUX_B_SEL : out std_logic_vector (1 downto
         0);  ALU_OPC : out std_logic_vector (0 to 4);  ALU_OUTREG_EN, 
         DRAM_R_IN : out std_logic;  JUMP_TYPE : out std_logic_vector (1 downto
         0);  MEM_EN_IN, DRAM_W_IN, RF_WE : out std_logic;  LOAD_TYPE_IN : out 
         std_logic_vector (1 downto 0);  STORE_TYPE_IN, WB_MUX_SEL : out 
         std_logic;  INS_IN : in std_logic_vector (31 downto 0);  Bubble, Clk, 
         Rst : in std_logic);

end hardwired_cu_NBIT32;

architecture SYN_bhv of hardwired_cu_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal AluOP_E_4_port, AluOP_E_3_port, AluOP_E_2_port, AluOP_E_1_port, 
      AluOP_E_0_port, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, 
      n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n_1986, n_1987, n_1988, n_1989, n_1990 : std_logic;

begin
   
   ALU_OPC_reg_0_inst : DFFR_X1 port map( D => AluOP_E_0_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(4), QN => n_1986);
   WB_MUX_SEL <= '0';
   STORE_TYPE_IN <= '0';
   LOAD_TYPE_IN(0) <= '0';
   LOAD_TYPE_IN(1) <= '0';
   RF_WE <= '0';
   DRAM_W_IN <= '0';
   MEM_EN_IN <= '0';
   JUMP_TYPE(0) <= '0';
   JUMP_TYPE(1) <= '0';
   DRAM_R_IN <= '0';
   ALU_OUTREG_EN <= '0';
   MUX_B_SEL(0) <= '0';
   MUX_B_SEL(1) <= '0';
   MUX_A_SEL <= '0';
   U126 : NAND3_X1 port map( A1 => INS_IN(1), A2 => n25, A3 => INS_IN(0), ZN =>
                           n65);
   U127 : NAND3_X1 port map( A1 => n87, A2 => n64, A3 => n88, ZN => n51);
   U128 : XOR2_X1 port map( A => n28, B => INS_IN(1), Z => n91);
   U129 : NAND3_X1 port map( A1 => n92, A2 => n27, A3 => INS_IN(0), ZN => n37);
   U130 : NAND3_X1 port map( A1 => n10, A2 => n7, A3 => n33, ZN => n103);
   U131 : NAND3_X1 port map( A1 => n28, A2 => n27, A3 => n92, ZN => n39);
   U132 : NAND3_X1 port map( A1 => n110, A2 => n25, A3 => INS_IN(1), ZN => n38)
                           ;
   U133 : NAND3_X1 port map( A1 => n26, A2 => n27, A3 => n53, ZN => n106);
   U134 : NAND3_X1 port map( A1 => INS_IN(1), A2 => n28, A3 => n92, ZN => n43);
   U135 : NAND3_X1 port map( A1 => n23, A2 => n21, A3 => n113, ZN => n112);
   ALU_OPC_reg_3_inst : DFFR_X1 port map( D => AluOP_E_3_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(1), QN => n_1987);
   ALU_OPC_reg_1_inst : DFFR_X1 port map( D => AluOP_E_1_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(3), QN => n_1988);
   ALU_OPC_reg_4_inst : DFFR_X1 port map( D => AluOP_E_4_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(0), QN => n_1989);
   ALU_OPC_reg_2_inst : DFFR_X1 port map( D => AluOP_E_2_port, CK => Clk, RN =>
                           Rst, Q => ALU_OPC(2), QN => n_1990);
   U17 : INV_X1 port map( A => n79, ZN => n4);
   U18 : NAND2_X1 port map( A1 => n82, A2 => n66, ZN => n73);
   U19 : INV_X1 port map( A => n82, ZN => n5);
   U20 : INV_X1 port map( A => n66, ZN => n2);
   U21 : INV_X1 port map( A => n34, ZN => n13);
   U22 : NOR3_X1 port map( A1 => n33, A2 => n99, A3 => n11, ZN => n81);
   U23 : INV_X1 port map( A => n77, ZN => n11);
   U24 : NAND2_X1 port map( A1 => n70, A2 => n8, ZN => n79);
   U25 : NAND2_X1 port map( A1 => n70, A2 => n9, ZN => n82);
   U26 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => n54);
   U27 : OAI21_X1 port map( B1 => n100, B2 => n75, A => n101, ZN => n95);
   U28 : NOR3_X1 port map( A1 => n102, A2 => n4, A3 => n46, ZN => n100);
   U29 : OAI21_X1 port map( B1 => n14, B2 => n57, A => n73, ZN => n101);
   U30 : OAI21_X1 port map( B1 => n3, B2 => n60, A => n103, ZN => n102);
   U31 : AND4_X1 port map( A1 => n70, A2 => n57, A3 => n10, A4 => n7, ZN => n35
                           );
   U32 : NAND2_X1 port map( A1 => n75, A2 => n59, ZN => n34);
   U33 : NAND2_X1 port map( A1 => n9, A2 => n74, ZN => n66);
   U34 : INV_X1 port map( A => n60, ZN => n9);
   U35 : INV_X1 port map( A => n75, ZN => n12);
   U36 : INV_X1 port map( A => n59, ZN => n14);
   U37 : OAI221_X1 port map( B1 => n78, B2 => n79, C1 => n66, C2 => n11, A => 
                           n80, ZN => n67);
   U38 : NOR3_X1 port map( A1 => n77, A2 => n57, A3 => n12, ZN => n78);
   U39 : NOR2_X1 port map( A1 => n48, A2 => n81, ZN => n80);
   U40 : AND3_X1 port map( A1 => n8, A2 => n74, A3 => n57, ZN => n32);
   U41 : AND3_X1 port map( A1 => n8, A2 => n74, A3 => n77, ZN => n48);
   U42 : INV_X1 port map( A => n105, ZN => n1);
   U43 : AOI21_X1 port map( B1 => n57, B2 => n46, A => n81, ZN => n105);
   U44 : INV_X1 port map( A => n99, ZN => n8);
   U45 : INV_X1 port map( A => n51, ZN => n17);
   U46 : AOI21_X1 port map( B1 => n44, B2 => n45, A => Bubble, ZN => 
                           AluOP_E_3_port);
   U47 : AOI211_X1 port map( C1 => n14, C2 => n4, A => n54, B => n1, ZN => n44)
                           ;
   U48 : AOI221_X1 port map( B1 => n46, B2 => n34, C1 => n35, C2 => n47, A => 
                           n48, ZN => n45);
   U49 : OAI21_X1 port map( B1 => n49, B2 => n50, A => n17, ZN => n47);
   U50 : AOI21_X1 port map( B1 => n93, B2 => n94, A => Bubble, ZN => 
                           AluOP_E_0_port);
   U51 : NOR3_X1 port map( A1 => n95, A2 => n6, A3 => n96, ZN => n94);
   U52 : AOI221_X1 port map( B1 => n35, B2 => n104, C1 => n77, C2 => n4, A => 
                           n1, ZN => n93);
   U53 : INV_X1 port map( A => n68, ZN => n6);
   U54 : AOI22_X1 port map( A1 => n98, A2 => n77, B1 => n57, B2 => n99, ZN => 
                           n97);
   U55 : NAND2_X1 port map( A1 => n52, A2 => n89, ZN => n83);
   U56 : AOI21_X1 port map( B1 => n29, B2 => n30, A => Bubble, ZN => 
                           AluOP_E_4_port);
   U57 : AOI211_X1 port map( C1 => n31, C2 => n9, A => n2, B => n32, ZN => n30)
                           ;
   U58 : AOI22_X1 port map( A1 => n35, A2 => n36, B1 => n12, B2 => n4, ZN => 
                           n29);
   U59 : NOR2_X1 port map( A1 => n13, A2 => n33, ZN => n31);
   U60 : OAI21_X1 port map( B1 => n52, B2 => n41, A => n27, ZN => n90);
   U61 : NAND4_X1 port map( A1 => n37, A2 => n38, A3 => n39, A4 => n40, ZN => 
                           n36);
   U62 : AOI21_X1 port map( B1 => n41, B2 => n42, A => n20, ZN => n40);
   U63 : INV_X1 port map( A => n43, ZN => n20);
   U64 : AOI21_X1 port map( B1 => n55, B2 => n56, A => Bubble, ZN => 
                           AluOP_E_2_port);
   U65 : AOI211_X1 port map( C1 => n5, C2 => n12, A => n67, B => n54, ZN => n55
                           );
   U66 : AOI221_X1 port map( B1 => n2, B2 => n57, C1 => n35, C2 => n16, A => 
                           n58, ZN => n56);
   U67 : NOR3_X1 port map( A1 => n59, A2 => n33, A3 => n60, ZN => n58);
   U68 : NAND2_X1 port map( A1 => n89, A2 => n110, ZN => n87);
   U69 : NAND2_X1 port map( A1 => n89, A2 => n41, ZN => n64);
   U70 : AOI21_X1 port map( B1 => n71, B2 => n72, A => Bubble, ZN => 
                           AluOP_E_1_port);
   U71 : AOI221_X1 port map( B1 => n46, B2 => n34, C1 => n14, C2 => n73, A => 
                           n32, ZN => n72);
   U72 : AOI221_X1 port map( B1 => n35, B2 => n76, C1 => n5, C2 => n77, A => 
                           n67, ZN => n71);
   U73 : NAND4_X1 port map( A1 => n43, A2 => n37, A3 => n83, A4 => n84, ZN => 
                           n76);
   U74 : INV_X1 port map( A => n53, ZN => n19);
   U75 : INV_X1 port map( A => n38, ZN => n18);
   U76 : AND2_X1 port map( A1 => n41, A2 => n25, ZN => n92);
   U77 : INV_X1 port map( A => n50, ZN => n26);
   U78 : NOR3_X1 port map( A1 => n22, A2 => INS_IN(3), A3 => n112, ZN => n52);
   U79 : NOR3_X1 port map( A1 => n22, A2 => n24, A3 => n112, ZN => n41);
   U80 : INV_X1 port map( A => INS_IN(3), ZN => n24);
   U81 : NOR3_X1 port map( A1 => INS_IN(3), A2 => INS_IN(5), A3 => n112, ZN => 
                           n53);
   U82 : NOR3_X1 port map( A1 => n28, A2 => INS_IN(1), A3 => n25, ZN => n89);
   U83 : NOR4_X1 port map( A1 => INS_IN(7), A2 => INS_IN(10), A3 => INS_IN(9), 
                           A4 => INS_IN(8), ZN => n113);
   U84 : AOI221_X1 port map( B1 => n85, B2 => n52, C1 => n26, C2 => n86, A => 
                           n51, ZN => n84);
   U85 : NOR2_X1 port map( A1 => INS_IN(2), A2 => n91, ZN => n85);
   U86 : OAI21_X1 port map( B1 => n27, B2 => n19, A => n90, ZN => n86);
   U87 : NAND4_X1 port map( A1 => n88, A2 => n43, A3 => n106, A4 => n107, ZN =>
                           n104);
   U88 : AOI221_X1 port map( B1 => n108, B2 => n52, C1 => n18, C2 => INS_IN(0),
                           A => n62, ZN => n107);
   U89 : NOR2_X1 port map( A1 => INS_IN(2), A2 => INS_IN(0), ZN => n108);
   U90 : OAI21_X1 port map( B1 => INS_IN(1), B2 => n50, A => n65, ZN => n42);
   U91 : NAND4_X1 port map( A1 => n53, A2 => INS_IN(2), A3 => INS_IN(0), A4 => 
                           INS_IN(1), ZN => n88);
   U92 : NAND2_X1 port map( A1 => INS_IN(2), A2 => n28, ZN => n50);
   U93 : INV_X1 port map( A => INS_IN(1), ZN => n27);
   U94 : AOI21_X1 port map( B1 => n52, B2 => INS_IN(1), A => n53, ZN => n49);
   U95 : NAND4_X1 port map( A1 => n109, A2 => n83, A3 => n87, A4 => n39, ZN => 
                           n62);
   U96 : NAND4_X1 port map( A1 => INS_IN(3), A2 => n22, A3 => INS_IN(1), A4 => 
                           n111, ZN => n109);
   U97 : NOR2_X1 port map( A1 => n112, A2 => n50, ZN => n111);
   U98 : INV_X1 port map( A => INS_IN(0), ZN => n28);
   U99 : INV_X1 port map( A => INS_IN(5), ZN => n22);
   U100 : INV_X1 port map( A => INS_IN(2), ZN => n25);
   U101 : AND4_X1 port map( A1 => n113, A2 => n21, A3 => INS_IN(3), A4 => n114,
                           ZN => n110);
   U102 : NOR2_X1 port map( A1 => n23, A2 => n22, ZN => n114);
   U103 : INV_X1 port map( A => INS_IN(4), ZN => n23);
   U104 : INV_X1 port map( A => INS_IN(6), ZN => n21);
   U105 : INV_X1 port map( A => n61, ZN => n16);
   U106 : AOI211_X1 port map( C1 => n42, C2 => n52, A => n62, B => n63, ZN => 
                           n61);
   U107 : OAI211_X1 port map( C1 => n38, C2 => INS_IN(0), A => n37, B => n64, 
                           ZN => n63);
   U108 : NOR2_X1 port map( A1 => INS_IN(29), A2 => n10, ZN => n98);
   U109 : INV_X1 port map( A => INS_IN(29), ZN => n7);
   U110 : NAND2_X1 port map( A1 => INS_IN(29), A2 => n10, ZN => n60);
   U111 : INV_X1 port map( A => INS_IN(26), ZN => n15);
   U112 : NOR3_X1 port map( A1 => n3, A2 => INS_IN(30), A3 => n97, ZN => n96);
   U113 : AND2_X1 port map( A1 => INS_IN(30), A2 => n3, ZN => n74);
   U114 : NAND2_X1 port map( A1 => INS_IN(27), A2 => n15, ZN => n59);
   U115 : NAND2_X1 port map( A1 => INS_IN(26), A2 => INS_IN(27), ZN => n75);
   U116 : NOR2_X1 port map( A1 => n15, A2 => INS_IN(27), ZN => n77);
   U117 : NOR2_X1 port map( A1 => INS_IN(27), A2 => INS_IN(26), ZN => n57);
   U118 : NAND4_X1 port map( A1 => n70, A2 => n57, A3 => INS_IN(28), A4 => n7, 
                           ZN => n69);
   U119 : NAND4_X1 port map( A1 => n77, A2 => n70, A3 => INS_IN(28), A4 => n7, 
                           ZN => n68);
   U120 : AND3_X1 port map( A1 => INS_IN(28), A2 => n7, A3 => n74, ZN => n46);
   U121 : NAND2_X1 port map( A1 => INS_IN(29), A2 => INS_IN(28), ZN => n99);
   U122 : INV_X1 port map( A => INS_IN(28), ZN => n10);
   U123 : NAND2_X1 port map( A1 => INS_IN(31), A2 => INS_IN(30), ZN => n33);
   U124 : NOR2_X1 port map( A1 => INS_IN(31), A2 => INS_IN(30), ZN => n70);
   U125 : INV_X1 port map( A => INS_IN(31), ZN => n3);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity Datapath is

   port( CLK, RST : in std_logic;  INS_IN, DATA_IN : in std_logic_vector (31 
         downto 0);  MUX_A_SEL : in std_logic;  MUX_B_SEL : in std_logic_vector
         (1 downto 0);  ALU_OPC : in std_logic_vector (0 to 4);  ALU_OUTREG_EN 
         : in std_logic;  JUMP_TYPE : in std_logic_vector (1 downto 0);  
         DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, RF_WE : in std_logic;  LOAD_TYPE_IN :
         in std_logic_vector (1 downto 0);  STORE_TYPE_IN, WB_MUX_SEL : in 
         std_logic;  INS_OUT, IRAM_ADDR_OUT, DRAM_ADDR_OUT, DATA_OUT : out 
         std_logic_vector (31 downto 0);  DRAM_R_OUT, DRAM_W_OUT, Bubble_out : 
         out std_logic;  LOAD_TYPE_OUT : out std_logic_vector (1 downto 0);  
         STORE_TYPE_OUT : out std_logic);

end Datapath;

architecture SYN_struct of Datapath is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HazardDetection
      port( RST : in std_logic;  ADD_RS1, ADD_RS2, ADD_WR : in std_logic_vector
            (4 downto 0);  DRAM_R : in std_logic;  INS_IN, PC_IN : in 
            std_logic_vector (31 downto 0);  Bubble : out std_logic;  
            HDU_INS_OUT, HDU_PC_OUT, HDU_NPC_OUT : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Writeback
      port( WB_MUX_SEL : in std_logic;  DATA_IN, ALU_RES_IN : in 
            std_logic_vector (31 downto 0);  ADD_WR_IN : in std_logic_vector (4
            downto 0);  DATA_OUT : out std_logic_vector (31 downto 0);  
            ADD_WR_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component ff_2
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Memory
      port( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN : in std_logic;  PC_SEL :
            in std_logic_vector (1 downto 0);  NPC_IN, NPC_ABS, NPC_REL, 
            ALU_RES_IN, B_IN : in std_logic_vector (31 downto 0);  ADD_WR_IN : 
            in std_logic_vector (4 downto 0);  DRAM_DATA_IN : in 
            std_logic_vector (31 downto 0);  LOAD_TYPE_IN : in std_logic_vector
            (1 downto 0);  STORE_TYPE_IN : in std_logic;  PC_OUT : out 
            std_logic_vector (31 downto 0);  DRAM_R_OUT, DRAM_W_OUT : out 
            std_logic;  DRAM_ADDR_OUT, DRAM_DATA_OUT, DATA_OUT, ALU_RES_OUT, 
            OP_MEM : out std_logic_vector (31 downto 0);  ADD_WR_MEM, 
            ADD_WR_OUT : out std_logic_vector (4 downto 0);  LOAD_TYPE_OUT : 
            out std_logic_vector (1 downto 0);  STORE_TYPE_OUT : out std_logic
            );
   end component;
   
   component ff_0
      port( D, CLK, EN, RST : in std_logic;  Q : out std_logic);
   end component;
   
   component Execute
      port( CLK, RST, MUX_A_SEL : in std_logic;  MUX_B_SEL : in 
            std_logic_vector (1 downto 0);  ALU_OPC : in std_logic_vector (0 to
            4);  ALU_OUTREG_EN : in std_logic;  JUMP_TYPE : in std_logic_vector
            (1 downto 0);  PC_IN, A_IN, B_IN, IMM_IN : in std_logic_vector (31 
            downto 0);  ADD_WR_IN, ADD_RS1_IN, ADD_RS2_IN, ADD_WR_MEM, 
            ADD_WR_WB : in std_logic_vector (4 downto 0);  RF_WE_MEM, RF_WE_WB 
            : in std_logic;  OP_MEM, OP_WB : in std_logic_vector (31 downto 0);
            PC_SEL : out std_logic_vector (1 downto 0);  ZERO_FLAG : out 
            std_logic;  NPC_ABS, NPC_REL, ALU_RES, B_OUT : out std_logic_vector
            (31 downto 0);  ADD_WR_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component Decode
      port( CLK, RST, Bubble, RF_WE, ZERO_FLAG : in std_logic;  PC_IN, INS_IN :
            in std_logic_vector (31 downto 0);  ADD_WR : in std_logic_vector (4
            downto 0);  DATA_WR_IN : in std_logic_vector (31 downto 0);  PC_OUT
            , A_OUT, B_OUT, IMM_OUT : out std_logic_vector (31 downto 0);  
            ADD_RS1_HDU, ADD_RS2_HDU, ADD_WR_OUT, ADD_RS1_OUT, ADD_RS2_OUT : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component Fetch
      port( CLK, RST, ZERO_FLAG : in std_logic;  PC_EXT, INS_IN : in 
            std_logic_vector (31 downto 0);  Bubble_in : in std_logic;  
            HDU_INS_IN, HDU_PC_IN, HDU_NPC_IN : in std_logic_vector (31 downto 
            0);  PC_OUT, ADDR_OUT, NPC_OUT, INS_OUT : out std_logic_vector (31 
            downto 0));
   end component;
   
   signal X_Logic1_port, n8, n9, n10, n11, n12, n13, INS_OUT_25_port, 
      INS_OUT_24_port, INS_OUT_23_port, INS_OUT_22_port, INS_OUT_21_port, 
      INS_OUT_20_port, INS_OUT_19_port, INS_OUT_18_port, INS_OUT_17_port, 
      INS_OUT_16_port, INS_OUT_15_port, INS_OUT_14_port, INS_OUT_13_port, 
      INS_OUT_12_port, INS_OUT_11_port, INS_OUT_10_port, INS_OUT_9_port, 
      INS_OUT_8_port, INS_OUT_7_port, INS_OUT_6_port, INS_OUT_5_port, 
      INS_OUT_4_port, INS_OUT_3_port, INS_OUT_2_port, INS_OUT_1_port, 
      INS_OUT_0_port, n14, ZERO_FLAG_EX, PC_MEM_OUT_31_port, PC_MEM_OUT_30_port
      , PC_MEM_OUT_29_port, PC_MEM_OUT_28_port, PC_MEM_OUT_27_port, 
      PC_MEM_OUT_26_port, PC_MEM_OUT_25_port, PC_MEM_OUT_24_port, 
      PC_MEM_OUT_23_port, PC_MEM_OUT_22_port, PC_MEM_OUT_21_port, 
      PC_MEM_OUT_20_port, PC_MEM_OUT_19_port, PC_MEM_OUT_18_port, 
      PC_MEM_OUT_17_port, PC_MEM_OUT_16_port, PC_MEM_OUT_15_port, 
      PC_MEM_OUT_14_port, PC_MEM_OUT_13_port, PC_MEM_OUT_12_port, 
      PC_MEM_OUT_11_port, PC_MEM_OUT_10_port, PC_MEM_OUT_9_port, 
      PC_MEM_OUT_8_port, PC_MEM_OUT_7_port, PC_MEM_OUT_6_port, 
      PC_MEM_OUT_5_port, PC_MEM_OUT_4_port, PC_MEM_OUT_3_port, 
      PC_MEM_OUT_2_port, PC_MEM_OUT_1_port, PC_MEM_OUT_0_port, 
      sig_HDU_INS_OUT_31_port, sig_HDU_INS_OUT_30_port, sig_HDU_INS_OUT_29_port
      , sig_HDU_INS_OUT_28_port, sig_HDU_INS_OUT_27_port, 
      sig_HDU_INS_OUT_26_port, sig_HDU_INS_OUT_25_port, sig_HDU_INS_OUT_24_port
      , sig_HDU_INS_OUT_23_port, sig_HDU_INS_OUT_22_port, 
      sig_HDU_INS_OUT_21_port, sig_HDU_INS_OUT_20_port, sig_HDU_INS_OUT_19_port
      , sig_HDU_INS_OUT_18_port, sig_HDU_INS_OUT_17_port, 
      sig_HDU_INS_OUT_16_port, sig_HDU_INS_OUT_15_port, sig_HDU_INS_OUT_14_port
      , sig_HDU_INS_OUT_13_port, sig_HDU_INS_OUT_12_port, 
      sig_HDU_INS_OUT_11_port, sig_HDU_INS_OUT_10_port, sig_HDU_INS_OUT_9_port,
      sig_HDU_INS_OUT_8_port, sig_HDU_INS_OUT_7_port, sig_HDU_INS_OUT_6_port, 
      sig_HDU_INS_OUT_5_port, sig_HDU_INS_OUT_4_port, sig_HDU_INS_OUT_3_port, 
      sig_HDU_INS_OUT_2_port, sig_HDU_INS_OUT_1_port, sig_HDU_INS_OUT_0_port, 
      sig_HDU_PC_OUT_31_port, sig_HDU_PC_OUT_30_port, sig_HDU_PC_OUT_29_port, 
      sig_HDU_PC_OUT_28_port, sig_HDU_PC_OUT_27_port, sig_HDU_PC_OUT_26_port, 
      sig_HDU_PC_OUT_25_port, sig_HDU_PC_OUT_24_port, sig_HDU_PC_OUT_23_port, 
      sig_HDU_PC_OUT_22_port, sig_HDU_PC_OUT_21_port, sig_HDU_PC_OUT_20_port, 
      sig_HDU_PC_OUT_19_port, sig_HDU_PC_OUT_18_port, sig_HDU_PC_OUT_17_port, 
      sig_HDU_PC_OUT_16_port, sig_HDU_PC_OUT_15_port, sig_HDU_PC_OUT_14_port, 
      sig_HDU_PC_OUT_13_port, sig_HDU_PC_OUT_12_port, sig_HDU_PC_OUT_11_port, 
      sig_HDU_PC_OUT_10_port, sig_HDU_PC_OUT_9_port, sig_HDU_PC_OUT_8_port, 
      sig_HDU_PC_OUT_7_port, sig_HDU_PC_OUT_6_port, sig_HDU_PC_OUT_5_port, 
      sig_HDU_PC_OUT_4_port, sig_HDU_PC_OUT_3_port, sig_HDU_PC_OUT_2_port, 
      sig_HDU_PC_OUT_1_port, sig_HDU_PC_OUT_0_port, sig_HDU_NPC_OUT_31_port, 
      sig_HDU_NPC_OUT_30_port, sig_HDU_NPC_OUT_29_port, sig_HDU_NPC_OUT_28_port
      , sig_HDU_NPC_OUT_27_port, sig_HDU_NPC_OUT_26_port, 
      sig_HDU_NPC_OUT_25_port, sig_HDU_NPC_OUT_24_port, sig_HDU_NPC_OUT_23_port
      , sig_HDU_NPC_OUT_22_port, sig_HDU_NPC_OUT_21_port, 
      sig_HDU_NPC_OUT_20_port, sig_HDU_NPC_OUT_19_port, sig_HDU_NPC_OUT_18_port
      , sig_HDU_NPC_OUT_17_port, sig_HDU_NPC_OUT_16_port, 
      sig_HDU_NPC_OUT_15_port, sig_HDU_NPC_OUT_14_port, sig_HDU_NPC_OUT_13_port
      , sig_HDU_NPC_OUT_12_port, sig_HDU_NPC_OUT_11_port, 
      sig_HDU_NPC_OUT_10_port, sig_HDU_NPC_OUT_9_port, sig_HDU_NPC_OUT_8_port, 
      sig_HDU_NPC_OUT_7_port, sig_HDU_NPC_OUT_6_port, sig_HDU_NPC_OUT_5_port, 
      sig_HDU_NPC_OUT_4_port, sig_HDU_NPC_OUT_3_port, sig_HDU_NPC_OUT_2_port, 
      sig_HDU_NPC_OUT_1_port, sig_HDU_NPC_OUT_0_port, PC_FETCH_OUT_31_port, 
      PC_FETCH_OUT_30_port, PC_FETCH_OUT_29_port, PC_FETCH_OUT_28_port, 
      PC_FETCH_OUT_27_port, PC_FETCH_OUT_26_port, PC_FETCH_OUT_25_port, 
      PC_FETCH_OUT_24_port, PC_FETCH_OUT_23_port, PC_FETCH_OUT_22_port, 
      PC_FETCH_OUT_21_port, PC_FETCH_OUT_20_port, PC_FETCH_OUT_19_port, 
      PC_FETCH_OUT_18_port, PC_FETCH_OUT_17_port, PC_FETCH_OUT_16_port, 
      PC_FETCH_OUT_15_port, PC_FETCH_OUT_14_port, PC_FETCH_OUT_13_port, 
      PC_FETCH_OUT_12_port, PC_FETCH_OUT_11_port, PC_FETCH_OUT_10_port, 
      PC_FETCH_OUT_9_port, PC_FETCH_OUT_8_port, PC_FETCH_OUT_7_port, 
      PC_FETCH_OUT_6_port, PC_FETCH_OUT_5_port, PC_FETCH_OUT_4_port, 
      PC_FETCH_OUT_3_port, PC_FETCH_OUT_2_port, PC_FETCH_OUT_1_port, 
      PC_FETCH_OUT_0_port, NPC_FETCH_OUT_31_port, NPC_FETCH_OUT_30_port, 
      NPC_FETCH_OUT_29_port, NPC_FETCH_OUT_28_port, NPC_FETCH_OUT_27_port, 
      NPC_FETCH_OUT_26_port, NPC_FETCH_OUT_25_port, NPC_FETCH_OUT_24_port, 
      NPC_FETCH_OUT_23_port, NPC_FETCH_OUT_22_port, NPC_FETCH_OUT_21_port, 
      NPC_FETCH_OUT_20_port, NPC_FETCH_OUT_19_port, NPC_FETCH_OUT_18_port, 
      NPC_FETCH_OUT_17_port, NPC_FETCH_OUT_16_port, NPC_FETCH_OUT_15_port, 
      NPC_FETCH_OUT_14_port, NPC_FETCH_OUT_13_port, NPC_FETCH_OUT_12_port, 
      NPC_FETCH_OUT_11_port, NPC_FETCH_OUT_10_port, NPC_FETCH_OUT_9_port, 
      NPC_FETCH_OUT_8_port, NPC_FETCH_OUT_7_port, NPC_FETCH_OUT_6_port, 
      NPC_FETCH_OUT_5_port, NPC_FETCH_OUT_4_port, NPC_FETCH_OUT_3_port, 
      NPC_FETCH_OUT_2_port, NPC_FETCH_OUT_1_port, NPC_FETCH_OUT_0_port, 
      RF_WE_WB, ADD_WR_WB_4_port, ADD_WR_WB_3_port, ADD_WR_WB_2_port, 
      ADD_WR_WB_1_port, ADD_WR_WB_0_port, OP_WB_31_port, OP_WB_30_port, 
      OP_WB_29_port, OP_WB_28_port, OP_WB_27_port, OP_WB_26_port, OP_WB_25_port
      , OP_WB_24_port, OP_WB_23_port, OP_WB_22_port, OP_WB_21_port, 
      OP_WB_20_port, OP_WB_19_port, OP_WB_18_port, OP_WB_17_port, OP_WB_16_port
      , OP_WB_15_port, OP_WB_14_port, OP_WB_13_port, OP_WB_12_port, 
      OP_WB_11_port, OP_WB_10_port, OP_WB_9_port, OP_WB_8_port, OP_WB_7_port, 
      OP_WB_6_port, OP_WB_5_port, OP_WB_4_port, OP_WB_3_port, OP_WB_2_port, 
      OP_WB_1_port, OP_WB_0_port, PC_DECODE_OUT_31_port, PC_DECODE_OUT_30_port,
      PC_DECODE_OUT_29_port, PC_DECODE_OUT_28_port, PC_DECODE_OUT_27_port, 
      PC_DECODE_OUT_26_port, PC_DECODE_OUT_25_port, PC_DECODE_OUT_24_port, 
      PC_DECODE_OUT_23_port, PC_DECODE_OUT_22_port, PC_DECODE_OUT_21_port, 
      PC_DECODE_OUT_20_port, PC_DECODE_OUT_19_port, PC_DECODE_OUT_18_port, 
      PC_DECODE_OUT_17_port, PC_DECODE_OUT_16_port, PC_DECODE_OUT_15_port, 
      PC_DECODE_OUT_14_port, PC_DECODE_OUT_13_port, PC_DECODE_OUT_12_port, 
      PC_DECODE_OUT_11_port, PC_DECODE_OUT_10_port, PC_DECODE_OUT_9_port, 
      PC_DECODE_OUT_8_port, PC_DECODE_OUT_7_port, PC_DECODE_OUT_6_port, 
      PC_DECODE_OUT_5_port, PC_DECODE_OUT_4_port, PC_DECODE_OUT_3_port, 
      PC_DECODE_OUT_2_port, PC_DECODE_OUT_1_port, PC_DECODE_OUT_0_port, 
      A_DECODE_OUT_31_port, A_DECODE_OUT_30_port, A_DECODE_OUT_29_port, 
      A_DECODE_OUT_28_port, A_DECODE_OUT_27_port, A_DECODE_OUT_26_port, 
      A_DECODE_OUT_25_port, A_DECODE_OUT_24_port, A_DECODE_OUT_23_port, 
      A_DECODE_OUT_22_port, A_DECODE_OUT_21_port, A_DECODE_OUT_20_port, 
      A_DECODE_OUT_19_port, A_DECODE_OUT_18_port, A_DECODE_OUT_17_port, 
      A_DECODE_OUT_16_port, A_DECODE_OUT_15_port, A_DECODE_OUT_14_port, 
      A_DECODE_OUT_13_port, A_DECODE_OUT_12_port, A_DECODE_OUT_11_port, 
      A_DECODE_OUT_10_port, A_DECODE_OUT_9_port, A_DECODE_OUT_8_port, 
      A_DECODE_OUT_7_port, A_DECODE_OUT_6_port, A_DECODE_OUT_5_port, 
      A_DECODE_OUT_4_port, A_DECODE_OUT_3_port, A_DECODE_OUT_2_port, 
      A_DECODE_OUT_1_port, A_DECODE_OUT_0_port, B_DECODE_OUT_31_port, 
      B_DECODE_OUT_30_port, B_DECODE_OUT_29_port, B_DECODE_OUT_28_port, 
      B_DECODE_OUT_27_port, B_DECODE_OUT_26_port, B_DECODE_OUT_25_port, 
      B_DECODE_OUT_24_port, B_DECODE_OUT_23_port, B_DECODE_OUT_22_port, 
      B_DECODE_OUT_21_port, B_DECODE_OUT_20_port, B_DECODE_OUT_19_port, 
      B_DECODE_OUT_18_port, B_DECODE_OUT_17_port, B_DECODE_OUT_16_port, 
      B_DECODE_OUT_15_port, B_DECODE_OUT_14_port, B_DECODE_OUT_13_port, 
      B_DECODE_OUT_12_port, B_DECODE_OUT_11_port, B_DECODE_OUT_10_port, 
      B_DECODE_OUT_9_port, B_DECODE_OUT_8_port, B_DECODE_OUT_7_port, 
      B_DECODE_OUT_6_port, B_DECODE_OUT_5_port, B_DECODE_OUT_4_port, 
      B_DECODE_OUT_3_port, B_DECODE_OUT_2_port, B_DECODE_OUT_1_port, 
      B_DECODE_OUT_0_port, IMM_DECODE_OUT_31_port, IMM_DECODE_OUT_30_port, 
      IMM_DECODE_OUT_29_port, IMM_DECODE_OUT_28_port, IMM_DECODE_OUT_27_port, 
      IMM_DECODE_OUT_26_port, IMM_DECODE_OUT_25_port, IMM_DECODE_OUT_24_port, 
      IMM_DECODE_OUT_23_port, IMM_DECODE_OUT_22_port, IMM_DECODE_OUT_21_port, 
      IMM_DECODE_OUT_20_port, IMM_DECODE_OUT_19_port, IMM_DECODE_OUT_18_port, 
      IMM_DECODE_OUT_17_port, IMM_DECODE_OUT_16_port, IMM_DECODE_OUT_15_port, 
      IMM_DECODE_OUT_14_port, IMM_DECODE_OUT_13_port, IMM_DECODE_OUT_12_port, 
      IMM_DECODE_OUT_11_port, IMM_DECODE_OUT_10_port, IMM_DECODE_OUT_9_port, 
      IMM_DECODE_OUT_8_port, IMM_DECODE_OUT_7_port, IMM_DECODE_OUT_6_port, 
      IMM_DECODE_OUT_5_port, IMM_DECODE_OUT_4_port, IMM_DECODE_OUT_3_port, 
      IMM_DECODE_OUT_2_port, IMM_DECODE_OUT_1_port, IMM_DECODE_OUT_0_port, 
      ADD_RS1_HDU_4_port, ADD_RS1_HDU_3_port, ADD_RS1_HDU_2_port, 
      ADD_RS1_HDU_1_port, ADD_RS1_HDU_0_port, ADD_RS2_HDU_4_port, 
      ADD_RS2_HDU_3_port, ADD_RS2_HDU_2_port, ADD_RS2_HDU_1_port, 
      ADD_RS2_HDU_0_port, ADD_WR_DECODE_OUT_4_port, ADD_WR_DECODE_OUT_3_port, 
      ADD_WR_DECODE_OUT_2_port, ADD_WR_DECODE_OUT_1_port, 
      ADD_WR_DECODE_OUT_0_port, ADD_RS1_DECODE_OUT_4_port, 
      ADD_RS1_DECODE_OUT_3_port, ADD_RS1_DECODE_OUT_2_port, 
      ADD_RS1_DECODE_OUT_1_port, ADD_RS1_DECODE_OUT_0_port, 
      ADD_RS2_DECODE_OUT_4_port, ADD_RS2_DECODE_OUT_3_port, 
      ADD_RS2_DECODE_OUT_2_port, ADD_RS2_DECODE_OUT_1_port, 
      ADD_RS2_DECODE_OUT_0_port, ADD_WR_MEM_4_port, ADD_WR_MEM_3_port, 
      ADD_WR_MEM_2_port, ADD_WR_MEM_1_port, ADD_WR_MEM_0_port, OP_MEM_31_port, 
      OP_MEM_30_port, OP_MEM_29_port, OP_MEM_28_port, OP_MEM_27_port, 
      OP_MEM_26_port, OP_MEM_25_port, OP_MEM_24_port, OP_MEM_23_port, 
      OP_MEM_22_port, OP_MEM_21_port, OP_MEM_20_port, OP_MEM_19_port, 
      OP_MEM_18_port, OP_MEM_17_port, OP_MEM_16_port, OP_MEM_15_port, 
      OP_MEM_14_port, OP_MEM_13_port, OP_MEM_12_port, OP_MEM_11_port, 
      OP_MEM_10_port, OP_MEM_9_port, OP_MEM_8_port, OP_MEM_7_port, 
      OP_MEM_6_port, OP_MEM_5_port, OP_MEM_4_port, OP_MEM_3_port, OP_MEM_2_port
      , OP_MEM_1_port, OP_MEM_0_port, PC_SEL_EX_1_port, PC_SEL_EX_0_port, 
      NPC_ABS_EX_31_port, NPC_ABS_EX_30_port, NPC_ABS_EX_29_port, 
      NPC_ABS_EX_28_port, NPC_ABS_EX_27_port, NPC_ABS_EX_26_port, 
      NPC_ABS_EX_25_port, NPC_ABS_EX_24_port, NPC_ABS_EX_23_port, 
      NPC_ABS_EX_22_port, NPC_ABS_EX_21_port, NPC_ABS_EX_20_port, 
      NPC_ABS_EX_19_port, NPC_ABS_EX_18_port, NPC_ABS_EX_17_port, 
      NPC_ABS_EX_16_port, NPC_ABS_EX_15_port, NPC_ABS_EX_14_port, 
      NPC_ABS_EX_13_port, NPC_ABS_EX_12_port, NPC_ABS_EX_11_port, 
      NPC_ABS_EX_10_port, NPC_ABS_EX_9_port, NPC_ABS_EX_8_port, 
      NPC_ABS_EX_7_port, NPC_ABS_EX_6_port, NPC_ABS_EX_5_port, 
      NPC_ABS_EX_4_port, NPC_ABS_EX_3_port, NPC_ABS_EX_2_port, 
      NPC_ABS_EX_1_port, NPC_ABS_EX_0_port, NPC_REL_EX_31_port, 
      NPC_REL_EX_30_port, NPC_REL_EX_29_port, NPC_REL_EX_28_port, 
      NPC_REL_EX_27_port, NPC_REL_EX_26_port, NPC_REL_EX_25_port, 
      NPC_REL_EX_24_port, NPC_REL_EX_23_port, NPC_REL_EX_22_port, 
      NPC_REL_EX_21_port, NPC_REL_EX_20_port, NPC_REL_EX_19_port, 
      NPC_REL_EX_18_port, NPC_REL_EX_17_port, NPC_REL_EX_16_port, 
      NPC_REL_EX_15_port, NPC_REL_EX_14_port, NPC_REL_EX_13_port, 
      NPC_REL_EX_12_port, NPC_REL_EX_11_port, NPC_REL_EX_10_port, 
      NPC_REL_EX_9_port, NPC_REL_EX_8_port, NPC_REL_EX_7_port, 
      NPC_REL_EX_6_port, NPC_REL_EX_5_port, NPC_REL_EX_4_port, 
      NPC_REL_EX_3_port, NPC_REL_EX_2_port, NPC_REL_EX_1_port, 
      NPC_REL_EX_0_port, ALU_RES_EX_31_port, ALU_RES_EX_30_port, 
      ALU_RES_EX_29_port, ALU_RES_EX_28_port, ALU_RES_EX_27_port, 
      ALU_RES_EX_26_port, ALU_RES_EX_25_port, ALU_RES_EX_24_port, 
      ALU_RES_EX_23_port, ALU_RES_EX_22_port, ALU_RES_EX_21_port, 
      ALU_RES_EX_20_port, ALU_RES_EX_19_port, ALU_RES_EX_18_port, 
      ALU_RES_EX_17_port, ALU_RES_EX_16_port, ALU_RES_EX_15_port, 
      ALU_RES_EX_14_port, ALU_RES_EX_13_port, ALU_RES_EX_12_port, 
      ALU_RES_EX_11_port, ALU_RES_EX_10_port, ALU_RES_EX_9_port, 
      ALU_RES_EX_8_port, ALU_RES_EX_7_port, ALU_RES_EX_6_port, 
      ALU_RES_EX_5_port, ALU_RES_EX_4_port, ALU_RES_EX_3_port, 
      ALU_RES_EX_2_port, ALU_RES_EX_1_port, ALU_RES_EX_0_port, B_EX_OUT_31_port
      , B_EX_OUT_30_port, B_EX_OUT_29_port, B_EX_OUT_28_port, B_EX_OUT_27_port,
      B_EX_OUT_26_port, B_EX_OUT_25_port, B_EX_OUT_24_port, B_EX_OUT_23_port, 
      B_EX_OUT_22_port, B_EX_OUT_21_port, B_EX_OUT_20_port, B_EX_OUT_19_port, 
      B_EX_OUT_18_port, B_EX_OUT_17_port, B_EX_OUT_16_port, B_EX_OUT_15_port, 
      B_EX_OUT_14_port, B_EX_OUT_13_port, B_EX_OUT_12_port, B_EX_OUT_11_port, 
      B_EX_OUT_10_port, B_EX_OUT_9_port, B_EX_OUT_8_port, B_EX_OUT_7_port, 
      B_EX_OUT_6_port, B_EX_OUT_5_port, B_EX_OUT_4_port, B_EX_OUT_3_port, 
      B_EX_OUT_2_port, B_EX_OUT_1_port, B_EX_OUT_0_port, ADD_WR_EX_OUT_4_port, 
      ADD_WR_EX_OUT_3_port, ADD_WR_EX_OUT_2_port, ADD_WR_EX_OUT_1_port, 
      ADD_WR_EX_OUT_0_port, DRAM_R_MEM, DATA_MEM_OUT_31_port, 
      DATA_MEM_OUT_30_port, DATA_MEM_OUT_29_port, DATA_MEM_OUT_28_port, 
      DATA_MEM_OUT_27_port, DATA_MEM_OUT_26_port, DATA_MEM_OUT_25_port, 
      DATA_MEM_OUT_24_port, DATA_MEM_OUT_23_port, DATA_MEM_OUT_22_port, 
      DATA_MEM_OUT_21_port, DATA_MEM_OUT_20_port, DATA_MEM_OUT_19_port, 
      DATA_MEM_OUT_18_port, DATA_MEM_OUT_17_port, DATA_MEM_OUT_16_port, 
      DATA_MEM_OUT_15_port, DATA_MEM_OUT_14_port, DATA_MEM_OUT_13_port, 
      DATA_MEM_OUT_12_port, DATA_MEM_OUT_11_port, DATA_MEM_OUT_10_port, 
      DATA_MEM_OUT_9_port, DATA_MEM_OUT_8_port, DATA_MEM_OUT_7_port, 
      DATA_MEM_OUT_6_port, DATA_MEM_OUT_5_port, DATA_MEM_OUT_4_port, 
      DATA_MEM_OUT_3_port, DATA_MEM_OUT_2_port, DATA_MEM_OUT_1_port, 
      DATA_MEM_OUT_0_port, ALU_RES_MEM_31_port, ALU_RES_MEM_30_port, 
      ALU_RES_MEM_29_port, ALU_RES_MEM_28_port, ALU_RES_MEM_27_port, 
      ALU_RES_MEM_26_port, ALU_RES_MEM_25_port, ALU_RES_MEM_24_port, 
      ALU_RES_MEM_23_port, ALU_RES_MEM_22_port, ALU_RES_MEM_21_port, 
      ALU_RES_MEM_20_port, ALU_RES_MEM_19_port, ALU_RES_MEM_18_port, 
      ALU_RES_MEM_17_port, ALU_RES_MEM_16_port, ALU_RES_MEM_15_port, 
      ALU_RES_MEM_14_port, ALU_RES_MEM_13_port, ALU_RES_MEM_12_port, 
      ALU_RES_MEM_11_port, ALU_RES_MEM_10_port, ALU_RES_MEM_9_port, 
      ALU_RES_MEM_8_port, ALU_RES_MEM_7_port, ALU_RES_MEM_6_port, 
      ALU_RES_MEM_5_port, ALU_RES_MEM_4_port, ALU_RES_MEM_3_port, 
      ALU_RES_MEM_2_port, ALU_RES_MEM_1_port, ALU_RES_MEM_0_port, 
      ADD_WR_MEM_OUT_4_port, ADD_WR_MEM_OUT_3_port, ADD_WR_MEM_OUT_2_port, 
      ADD_WR_MEM_OUT_1_port, ADD_WR_MEM_OUT_0_port, INS_OUT_29_port, 
      INS_OUT_27_port, INS_OUT_26_port, INS_OUT_30_port, INS_OUT_28_port, 
      INS_OUT_31_port, Bubble_out_port : std_logic;

begin
   INS_OUT <= ( INS_OUT_31_port, INS_OUT_30_port, INS_OUT_29_port, 
      INS_OUT_28_port, INS_OUT_27_port, INS_OUT_26_port, INS_OUT_25_port, 
      INS_OUT_24_port, INS_OUT_23_port, INS_OUT_22_port, INS_OUT_21_port, 
      INS_OUT_20_port, INS_OUT_19_port, INS_OUT_18_port, INS_OUT_17_port, 
      INS_OUT_16_port, INS_OUT_15_port, INS_OUT_14_port, INS_OUT_13_port, 
      INS_OUT_12_port, INS_OUT_11_port, INS_OUT_10_port, INS_OUT_9_port, 
      INS_OUT_8_port, INS_OUT_7_port, INS_OUT_6_port, INS_OUT_5_port, 
      INS_OUT_4_port, INS_OUT_3_port, INS_OUT_2_port, INS_OUT_1_port, 
      INS_OUT_0_port );
   Bubble_out <= Bubble_out_port;
   
   X_Logic1_port <= '1';
   FetchStage : Fetch port map( CLK => CLK, RST => RST, ZERO_FLAG => 
                           ZERO_FLAG_EX, PC_EXT(31) => PC_MEM_OUT_31_port, 
                           PC_EXT(30) => PC_MEM_OUT_30_port, PC_EXT(29) => 
                           PC_MEM_OUT_29_port, PC_EXT(28) => PC_MEM_OUT_28_port
                           , PC_EXT(27) => PC_MEM_OUT_27_port, PC_EXT(26) => 
                           PC_MEM_OUT_26_port, PC_EXT(25) => PC_MEM_OUT_25_port
                           , PC_EXT(24) => PC_MEM_OUT_24_port, PC_EXT(23) => 
                           PC_MEM_OUT_23_port, PC_EXT(22) => PC_MEM_OUT_22_port
                           , PC_EXT(21) => PC_MEM_OUT_21_port, PC_EXT(20) => 
                           PC_MEM_OUT_20_port, PC_EXT(19) => PC_MEM_OUT_19_port
                           , PC_EXT(18) => PC_MEM_OUT_18_port, PC_EXT(17) => 
                           PC_MEM_OUT_17_port, PC_EXT(16) => PC_MEM_OUT_16_port
                           , PC_EXT(15) => PC_MEM_OUT_15_port, PC_EXT(14) => 
                           PC_MEM_OUT_14_port, PC_EXT(13) => PC_MEM_OUT_13_port
                           , PC_EXT(12) => PC_MEM_OUT_12_port, PC_EXT(11) => 
                           PC_MEM_OUT_11_port, PC_EXT(10) => PC_MEM_OUT_10_port
                           , PC_EXT(9) => PC_MEM_OUT_9_port, PC_EXT(8) => 
                           PC_MEM_OUT_8_port, PC_EXT(7) => PC_MEM_OUT_7_port, 
                           PC_EXT(6) => PC_MEM_OUT_6_port, PC_EXT(5) => 
                           PC_MEM_OUT_5_port, PC_EXT(4) => PC_MEM_OUT_4_port, 
                           PC_EXT(3) => PC_MEM_OUT_3_port, PC_EXT(2) => 
                           PC_MEM_OUT_2_port, PC_EXT(1) => PC_MEM_OUT_1_port, 
                           PC_EXT(0) => PC_MEM_OUT_0_port, INS_IN(31) => 
                           INS_IN(31), INS_IN(30) => INS_IN(30), INS_IN(29) => 
                           INS_IN(29), INS_IN(28) => INS_IN(28), INS_IN(27) => 
                           INS_IN(27), INS_IN(26) => INS_IN(26), INS_IN(25) => 
                           INS_IN(25), INS_IN(24) => INS_IN(24), INS_IN(23) => 
                           INS_IN(23), INS_IN(22) => INS_IN(22), INS_IN(21) => 
                           INS_IN(21), INS_IN(20) => INS_IN(20), INS_IN(19) => 
                           INS_IN(19), INS_IN(18) => INS_IN(18), INS_IN(17) => 
                           INS_IN(17), INS_IN(16) => INS_IN(16), INS_IN(15) => 
                           INS_IN(15), INS_IN(14) => INS_IN(14), INS_IN(13) => 
                           INS_IN(13), INS_IN(12) => INS_IN(12), INS_IN(11) => 
                           INS_IN(11), INS_IN(10) => INS_IN(10), INS_IN(9) => 
                           INS_IN(9), INS_IN(8) => INS_IN(8), INS_IN(7) => 
                           INS_IN(7), INS_IN(6) => INS_IN(6), INS_IN(5) => 
                           INS_IN(5), INS_IN(4) => INS_IN(4), INS_IN(3) => 
                           INS_IN(3), INS_IN(2) => INS_IN(2), INS_IN(1) => 
                           INS_IN(1), INS_IN(0) => INS_IN(0), Bubble_in => 
                           Bubble_out_port, HDU_INS_IN(31) => 
                           sig_HDU_INS_OUT_31_port, HDU_INS_IN(30) => 
                           sig_HDU_INS_OUT_30_port, HDU_INS_IN(29) => 
                           sig_HDU_INS_OUT_29_port, HDU_INS_IN(28) => 
                           sig_HDU_INS_OUT_28_port, HDU_INS_IN(27) => 
                           sig_HDU_INS_OUT_27_port, HDU_INS_IN(26) => 
                           sig_HDU_INS_OUT_26_port, HDU_INS_IN(25) => 
                           sig_HDU_INS_OUT_25_port, HDU_INS_IN(24) => 
                           sig_HDU_INS_OUT_24_port, HDU_INS_IN(23) => 
                           sig_HDU_INS_OUT_23_port, HDU_INS_IN(22) => 
                           sig_HDU_INS_OUT_22_port, HDU_INS_IN(21) => 
                           sig_HDU_INS_OUT_21_port, HDU_INS_IN(20) => 
                           sig_HDU_INS_OUT_20_port, HDU_INS_IN(19) => 
                           sig_HDU_INS_OUT_19_port, HDU_INS_IN(18) => 
                           sig_HDU_INS_OUT_18_port, HDU_INS_IN(17) => 
                           sig_HDU_INS_OUT_17_port, HDU_INS_IN(16) => 
                           sig_HDU_INS_OUT_16_port, HDU_INS_IN(15) => 
                           sig_HDU_INS_OUT_15_port, HDU_INS_IN(14) => 
                           sig_HDU_INS_OUT_14_port, HDU_INS_IN(13) => 
                           sig_HDU_INS_OUT_13_port, HDU_INS_IN(12) => 
                           sig_HDU_INS_OUT_12_port, HDU_INS_IN(11) => 
                           sig_HDU_INS_OUT_11_port, HDU_INS_IN(10) => 
                           sig_HDU_INS_OUT_10_port, HDU_INS_IN(9) => 
                           sig_HDU_INS_OUT_9_port, HDU_INS_IN(8) => 
                           sig_HDU_INS_OUT_8_port, HDU_INS_IN(7) => 
                           sig_HDU_INS_OUT_7_port, HDU_INS_IN(6) => 
                           sig_HDU_INS_OUT_6_port, HDU_INS_IN(5) => 
                           sig_HDU_INS_OUT_5_port, HDU_INS_IN(4) => 
                           sig_HDU_INS_OUT_4_port, HDU_INS_IN(3) => 
                           sig_HDU_INS_OUT_3_port, HDU_INS_IN(2) => 
                           sig_HDU_INS_OUT_2_port, HDU_INS_IN(1) => 
                           sig_HDU_INS_OUT_1_port, HDU_INS_IN(0) => 
                           sig_HDU_INS_OUT_0_port, HDU_PC_IN(31) => 
                           sig_HDU_PC_OUT_31_port, HDU_PC_IN(30) => 
                           sig_HDU_PC_OUT_30_port, HDU_PC_IN(29) => 
                           sig_HDU_PC_OUT_29_port, HDU_PC_IN(28) => 
                           sig_HDU_PC_OUT_28_port, HDU_PC_IN(27) => 
                           sig_HDU_PC_OUT_27_port, HDU_PC_IN(26) => 
                           sig_HDU_PC_OUT_26_port, HDU_PC_IN(25) => 
                           sig_HDU_PC_OUT_25_port, HDU_PC_IN(24) => 
                           sig_HDU_PC_OUT_24_port, HDU_PC_IN(23) => 
                           sig_HDU_PC_OUT_23_port, HDU_PC_IN(22) => 
                           sig_HDU_PC_OUT_22_port, HDU_PC_IN(21) => 
                           sig_HDU_PC_OUT_21_port, HDU_PC_IN(20) => 
                           sig_HDU_PC_OUT_20_port, HDU_PC_IN(19) => 
                           sig_HDU_PC_OUT_19_port, HDU_PC_IN(18) => 
                           sig_HDU_PC_OUT_18_port, HDU_PC_IN(17) => 
                           sig_HDU_PC_OUT_17_port, HDU_PC_IN(16) => 
                           sig_HDU_PC_OUT_16_port, HDU_PC_IN(15) => 
                           sig_HDU_PC_OUT_15_port, HDU_PC_IN(14) => 
                           sig_HDU_PC_OUT_14_port, HDU_PC_IN(13) => 
                           sig_HDU_PC_OUT_13_port, HDU_PC_IN(12) => 
                           sig_HDU_PC_OUT_12_port, HDU_PC_IN(11) => 
                           sig_HDU_PC_OUT_11_port, HDU_PC_IN(10) => 
                           sig_HDU_PC_OUT_10_port, HDU_PC_IN(9) => 
                           sig_HDU_PC_OUT_9_port, HDU_PC_IN(8) => 
                           sig_HDU_PC_OUT_8_port, HDU_PC_IN(7) => 
                           sig_HDU_PC_OUT_7_port, HDU_PC_IN(6) => 
                           sig_HDU_PC_OUT_6_port, HDU_PC_IN(5) => 
                           sig_HDU_PC_OUT_5_port, HDU_PC_IN(4) => 
                           sig_HDU_PC_OUT_4_port, HDU_PC_IN(3) => 
                           sig_HDU_PC_OUT_3_port, HDU_PC_IN(2) => 
                           sig_HDU_PC_OUT_2_port, HDU_PC_IN(1) => 
                           sig_HDU_PC_OUT_1_port, HDU_PC_IN(0) => 
                           sig_HDU_PC_OUT_0_port, HDU_NPC_IN(31) => 
                           sig_HDU_NPC_OUT_31_port, HDU_NPC_IN(30) => 
                           sig_HDU_NPC_OUT_30_port, HDU_NPC_IN(29) => 
                           sig_HDU_NPC_OUT_29_port, HDU_NPC_IN(28) => 
                           sig_HDU_NPC_OUT_28_port, HDU_NPC_IN(27) => 
                           sig_HDU_NPC_OUT_27_port, HDU_NPC_IN(26) => 
                           sig_HDU_NPC_OUT_26_port, HDU_NPC_IN(25) => 
                           sig_HDU_NPC_OUT_25_port, HDU_NPC_IN(24) => 
                           sig_HDU_NPC_OUT_24_port, HDU_NPC_IN(23) => 
                           sig_HDU_NPC_OUT_23_port, HDU_NPC_IN(22) => 
                           sig_HDU_NPC_OUT_22_port, HDU_NPC_IN(21) => 
                           sig_HDU_NPC_OUT_21_port, HDU_NPC_IN(20) => 
                           sig_HDU_NPC_OUT_20_port, HDU_NPC_IN(19) => 
                           sig_HDU_NPC_OUT_19_port, HDU_NPC_IN(18) => 
                           sig_HDU_NPC_OUT_18_port, HDU_NPC_IN(17) => 
                           sig_HDU_NPC_OUT_17_port, HDU_NPC_IN(16) => 
                           sig_HDU_NPC_OUT_16_port, HDU_NPC_IN(15) => 
                           sig_HDU_NPC_OUT_15_port, HDU_NPC_IN(14) => 
                           sig_HDU_NPC_OUT_14_port, HDU_NPC_IN(13) => 
                           sig_HDU_NPC_OUT_13_port, HDU_NPC_IN(12) => 
                           sig_HDU_NPC_OUT_12_port, HDU_NPC_IN(11) => 
                           sig_HDU_NPC_OUT_11_port, HDU_NPC_IN(10) => 
                           sig_HDU_NPC_OUT_10_port, HDU_NPC_IN(9) => 
                           sig_HDU_NPC_OUT_9_port, HDU_NPC_IN(8) => 
                           sig_HDU_NPC_OUT_8_port, HDU_NPC_IN(7) => 
                           sig_HDU_NPC_OUT_7_port, HDU_NPC_IN(6) => 
                           sig_HDU_NPC_OUT_6_port, HDU_NPC_IN(5) => 
                           sig_HDU_NPC_OUT_5_port, HDU_NPC_IN(4) => 
                           sig_HDU_NPC_OUT_4_port, HDU_NPC_IN(3) => 
                           sig_HDU_NPC_OUT_3_port, HDU_NPC_IN(2) => 
                           sig_HDU_NPC_OUT_2_port, HDU_NPC_IN(1) => 
                           sig_HDU_NPC_OUT_1_port, HDU_NPC_IN(0) => 
                           sig_HDU_NPC_OUT_0_port, PC_OUT(31) => 
                           PC_FETCH_OUT_31_port, PC_OUT(30) => 
                           PC_FETCH_OUT_30_port, PC_OUT(29) => 
                           PC_FETCH_OUT_29_port, PC_OUT(28) => 
                           PC_FETCH_OUT_28_port, PC_OUT(27) => 
                           PC_FETCH_OUT_27_port, PC_OUT(26) => 
                           PC_FETCH_OUT_26_port, PC_OUT(25) => 
                           PC_FETCH_OUT_25_port, PC_OUT(24) => 
                           PC_FETCH_OUT_24_port, PC_OUT(23) => 
                           PC_FETCH_OUT_23_port, PC_OUT(22) => 
                           PC_FETCH_OUT_22_port, PC_OUT(21) => 
                           PC_FETCH_OUT_21_port, PC_OUT(20) => 
                           PC_FETCH_OUT_20_port, PC_OUT(19) => 
                           PC_FETCH_OUT_19_port, PC_OUT(18) => 
                           PC_FETCH_OUT_18_port, PC_OUT(17) => 
                           PC_FETCH_OUT_17_port, PC_OUT(16) => 
                           PC_FETCH_OUT_16_port, PC_OUT(15) => 
                           PC_FETCH_OUT_15_port, PC_OUT(14) => 
                           PC_FETCH_OUT_14_port, PC_OUT(13) => 
                           PC_FETCH_OUT_13_port, PC_OUT(12) => 
                           PC_FETCH_OUT_12_port, PC_OUT(11) => 
                           PC_FETCH_OUT_11_port, PC_OUT(10) => 
                           PC_FETCH_OUT_10_port, PC_OUT(9) => 
                           PC_FETCH_OUT_9_port, PC_OUT(8) => 
                           PC_FETCH_OUT_8_port, PC_OUT(7) => 
                           PC_FETCH_OUT_7_port, PC_OUT(6) => 
                           PC_FETCH_OUT_6_port, PC_OUT(5) => 
                           PC_FETCH_OUT_5_port, PC_OUT(4) => 
                           PC_FETCH_OUT_4_port, PC_OUT(3) => 
                           PC_FETCH_OUT_3_port, PC_OUT(2) => 
                           PC_FETCH_OUT_2_port, PC_OUT(1) => 
                           PC_FETCH_OUT_1_port, PC_OUT(0) => 
                           PC_FETCH_OUT_0_port, ADDR_OUT(31) => 
                           IRAM_ADDR_OUT(31), ADDR_OUT(30) => IRAM_ADDR_OUT(30)
                           , ADDR_OUT(29) => IRAM_ADDR_OUT(29), ADDR_OUT(28) =>
                           IRAM_ADDR_OUT(28), ADDR_OUT(27) => IRAM_ADDR_OUT(27)
                           , ADDR_OUT(26) => IRAM_ADDR_OUT(26), ADDR_OUT(25) =>
                           IRAM_ADDR_OUT(25), ADDR_OUT(24) => IRAM_ADDR_OUT(24)
                           , ADDR_OUT(23) => IRAM_ADDR_OUT(23), ADDR_OUT(22) =>
                           IRAM_ADDR_OUT(22), ADDR_OUT(21) => IRAM_ADDR_OUT(21)
                           , ADDR_OUT(20) => IRAM_ADDR_OUT(20), ADDR_OUT(19) =>
                           IRAM_ADDR_OUT(19), ADDR_OUT(18) => IRAM_ADDR_OUT(18)
                           , ADDR_OUT(17) => IRAM_ADDR_OUT(17), ADDR_OUT(16) =>
                           IRAM_ADDR_OUT(16), ADDR_OUT(15) => IRAM_ADDR_OUT(15)
                           , ADDR_OUT(14) => IRAM_ADDR_OUT(14), ADDR_OUT(13) =>
                           IRAM_ADDR_OUT(13), ADDR_OUT(12) => IRAM_ADDR_OUT(12)
                           , ADDR_OUT(11) => IRAM_ADDR_OUT(11), ADDR_OUT(10) =>
                           IRAM_ADDR_OUT(10), ADDR_OUT(9) => IRAM_ADDR_OUT(9), 
                           ADDR_OUT(8) => IRAM_ADDR_OUT(8), ADDR_OUT(7) => 
                           IRAM_ADDR_OUT(7), ADDR_OUT(6) => IRAM_ADDR_OUT(6), 
                           ADDR_OUT(5) => IRAM_ADDR_OUT(5), ADDR_OUT(4) => 
                           IRAM_ADDR_OUT(4), ADDR_OUT(3) => IRAM_ADDR_OUT(3), 
                           ADDR_OUT(2) => IRAM_ADDR_OUT(2), ADDR_OUT(1) => 
                           IRAM_ADDR_OUT(1), ADDR_OUT(0) => IRAM_ADDR_OUT(0), 
                           NPC_OUT(31) => NPC_FETCH_OUT_31_port, NPC_OUT(30) =>
                           NPC_FETCH_OUT_30_port, NPC_OUT(29) => 
                           NPC_FETCH_OUT_29_port, NPC_OUT(28) => 
                           NPC_FETCH_OUT_28_port, NPC_OUT(27) => 
                           NPC_FETCH_OUT_27_port, NPC_OUT(26) => 
                           NPC_FETCH_OUT_26_port, NPC_OUT(25) => 
                           NPC_FETCH_OUT_25_port, NPC_OUT(24) => 
                           NPC_FETCH_OUT_24_port, NPC_OUT(23) => 
                           NPC_FETCH_OUT_23_port, NPC_OUT(22) => 
                           NPC_FETCH_OUT_22_port, NPC_OUT(21) => 
                           NPC_FETCH_OUT_21_port, NPC_OUT(20) => 
                           NPC_FETCH_OUT_20_port, NPC_OUT(19) => 
                           NPC_FETCH_OUT_19_port, NPC_OUT(18) => 
                           NPC_FETCH_OUT_18_port, NPC_OUT(17) => 
                           NPC_FETCH_OUT_17_port, NPC_OUT(16) => 
                           NPC_FETCH_OUT_16_port, NPC_OUT(15) => 
                           NPC_FETCH_OUT_15_port, NPC_OUT(14) => 
                           NPC_FETCH_OUT_14_port, NPC_OUT(13) => 
                           NPC_FETCH_OUT_13_port, NPC_OUT(12) => 
                           NPC_FETCH_OUT_12_port, NPC_OUT(11) => 
                           NPC_FETCH_OUT_11_port, NPC_OUT(10) => 
                           NPC_FETCH_OUT_10_port, NPC_OUT(9) => 
                           NPC_FETCH_OUT_9_port, NPC_OUT(8) => 
                           NPC_FETCH_OUT_8_port, NPC_OUT(7) => 
                           NPC_FETCH_OUT_7_port, NPC_OUT(6) => 
                           NPC_FETCH_OUT_6_port, NPC_OUT(5) => 
                           NPC_FETCH_OUT_5_port, NPC_OUT(4) => 
                           NPC_FETCH_OUT_4_port, NPC_OUT(3) => 
                           NPC_FETCH_OUT_3_port, NPC_OUT(2) => 
                           NPC_FETCH_OUT_2_port, NPC_OUT(1) => 
                           NPC_FETCH_OUT_1_port, NPC_OUT(0) => 
                           NPC_FETCH_OUT_0_port, INS_OUT(31) => n8, INS_OUT(30)
                           => n9, INS_OUT(29) => n10, INS_OUT(28) => n11, 
                           INS_OUT(27) => n12, INS_OUT(26) => n13, INS_OUT(25) 
                           => INS_OUT_25_port, INS_OUT(24) => INS_OUT_24_port, 
                           INS_OUT(23) => INS_OUT_23_port, INS_OUT(22) => 
                           INS_OUT_22_port, INS_OUT(21) => INS_OUT_21_port, 
                           INS_OUT(20) => INS_OUT_20_port, INS_OUT(19) => 
                           INS_OUT_19_port, INS_OUT(18) => INS_OUT_18_port, 
                           INS_OUT(17) => INS_OUT_17_port, INS_OUT(16) => 
                           INS_OUT_16_port, INS_OUT(15) => INS_OUT_15_port, 
                           INS_OUT(14) => INS_OUT_14_port, INS_OUT(13) => 
                           INS_OUT_13_port, INS_OUT(12) => INS_OUT_12_port, 
                           INS_OUT(11) => INS_OUT_11_port, INS_OUT(10) => 
                           INS_OUT_10_port, INS_OUT(9) => INS_OUT_9_port, 
                           INS_OUT(8) => INS_OUT_8_port, INS_OUT(7) => 
                           INS_OUT_7_port, INS_OUT(6) => INS_OUT_6_port, 
                           INS_OUT(5) => INS_OUT_5_port, INS_OUT(4) => 
                           INS_OUT_4_port, INS_OUT(3) => INS_OUT_3_port, 
                           INS_OUT(2) => INS_OUT_2_port, INS_OUT(1) => 
                           INS_OUT_1_port, INS_OUT(0) => INS_OUT_0_port);
   DecodeStage : Decode port map( CLK => CLK, RST => RST, Bubble => 
                           Bubble_out_port, RF_WE => RF_WE_WB, ZERO_FLAG => 
                           ZERO_FLAG_EX, PC_IN(31) => PC_FETCH_OUT_31_port, 
                           PC_IN(30) => PC_FETCH_OUT_30_port, PC_IN(29) => 
                           PC_FETCH_OUT_29_port, PC_IN(28) => 
                           PC_FETCH_OUT_28_port, PC_IN(27) => 
                           PC_FETCH_OUT_27_port, PC_IN(26) => 
                           PC_FETCH_OUT_26_port, PC_IN(25) => 
                           PC_FETCH_OUT_25_port, PC_IN(24) => 
                           PC_FETCH_OUT_24_port, PC_IN(23) => 
                           PC_FETCH_OUT_23_port, PC_IN(22) => 
                           PC_FETCH_OUT_22_port, PC_IN(21) => 
                           PC_FETCH_OUT_21_port, PC_IN(20) => 
                           PC_FETCH_OUT_20_port, PC_IN(19) => 
                           PC_FETCH_OUT_19_port, PC_IN(18) => 
                           PC_FETCH_OUT_18_port, PC_IN(17) => 
                           PC_FETCH_OUT_17_port, PC_IN(16) => 
                           PC_FETCH_OUT_16_port, PC_IN(15) => 
                           PC_FETCH_OUT_15_port, PC_IN(14) => 
                           PC_FETCH_OUT_14_port, PC_IN(13) => 
                           PC_FETCH_OUT_13_port, PC_IN(12) => 
                           PC_FETCH_OUT_12_port, PC_IN(11) => 
                           PC_FETCH_OUT_11_port, PC_IN(10) => 
                           PC_FETCH_OUT_10_port, PC_IN(9) => 
                           PC_FETCH_OUT_9_port, PC_IN(8) => PC_FETCH_OUT_8_port
                           , PC_IN(7) => PC_FETCH_OUT_7_port, PC_IN(6) => 
                           PC_FETCH_OUT_6_port, PC_IN(5) => PC_FETCH_OUT_5_port
                           , PC_IN(4) => PC_FETCH_OUT_4_port, PC_IN(3) => 
                           PC_FETCH_OUT_3_port, PC_IN(2) => PC_FETCH_OUT_2_port
                           , PC_IN(1) => PC_FETCH_OUT_1_port, PC_IN(0) => 
                           PC_FETCH_OUT_0_port, INS_IN(31) => n8, INS_IN(30) =>
                           n9, INS_IN(29) => n10, INS_IN(28) => n11, INS_IN(27)
                           => n12, INS_IN(26) => n13, INS_IN(25) => 
                           INS_OUT_25_port, INS_IN(24) => INS_OUT_24_port, 
                           INS_IN(23) => INS_OUT_23_port, INS_IN(22) => 
                           INS_OUT_22_port, INS_IN(21) => INS_OUT_21_port, 
                           INS_IN(20) => INS_OUT_20_port, INS_IN(19) => 
                           INS_OUT_19_port, INS_IN(18) => INS_OUT_18_port, 
                           INS_IN(17) => INS_OUT_17_port, INS_IN(16) => 
                           INS_OUT_16_port, INS_IN(15) => INS_OUT_15_port, 
                           INS_IN(14) => INS_OUT_14_port, INS_IN(13) => 
                           INS_OUT_13_port, INS_IN(12) => INS_OUT_12_port, 
                           INS_IN(11) => INS_OUT_11_port, INS_IN(10) => 
                           INS_OUT_10_port, INS_IN(9) => INS_OUT_9_port, 
                           INS_IN(8) => INS_OUT_8_port, INS_IN(7) => 
                           INS_OUT_7_port, INS_IN(6) => INS_OUT_6_port, 
                           INS_IN(5) => INS_OUT_5_port, INS_IN(4) => 
                           INS_OUT_4_port, INS_IN(3) => INS_OUT_3_port, 
                           INS_IN(2) => INS_OUT_2_port, INS_IN(1) => 
                           INS_OUT_1_port, INS_IN(0) => INS_OUT_0_port, 
                           ADD_WR(4) => ADD_WR_WB_4_port, ADD_WR(3) => 
                           ADD_WR_WB_3_port, ADD_WR(2) => ADD_WR_WB_2_port, 
                           ADD_WR(1) => ADD_WR_WB_1_port, ADD_WR(0) => 
                           ADD_WR_WB_0_port, DATA_WR_IN(31) => OP_WB_31_port, 
                           DATA_WR_IN(30) => OP_WB_30_port, DATA_WR_IN(29) => 
                           OP_WB_29_port, DATA_WR_IN(28) => OP_WB_28_port, 
                           DATA_WR_IN(27) => OP_WB_27_port, DATA_WR_IN(26) => 
                           OP_WB_26_port, DATA_WR_IN(25) => OP_WB_25_port, 
                           DATA_WR_IN(24) => OP_WB_24_port, DATA_WR_IN(23) => 
                           OP_WB_23_port, DATA_WR_IN(22) => OP_WB_22_port, 
                           DATA_WR_IN(21) => OP_WB_21_port, DATA_WR_IN(20) => 
                           OP_WB_20_port, DATA_WR_IN(19) => OP_WB_19_port, 
                           DATA_WR_IN(18) => OP_WB_18_port, DATA_WR_IN(17) => 
                           OP_WB_17_port, DATA_WR_IN(16) => OP_WB_16_port, 
                           DATA_WR_IN(15) => OP_WB_15_port, DATA_WR_IN(14) => 
                           OP_WB_14_port, DATA_WR_IN(13) => OP_WB_13_port, 
                           DATA_WR_IN(12) => OP_WB_12_port, DATA_WR_IN(11) => 
                           OP_WB_11_port, DATA_WR_IN(10) => OP_WB_10_port, 
                           DATA_WR_IN(9) => OP_WB_9_port, DATA_WR_IN(8) => 
                           OP_WB_8_port, DATA_WR_IN(7) => OP_WB_7_port, 
                           DATA_WR_IN(6) => OP_WB_6_port, DATA_WR_IN(5) => 
                           OP_WB_5_port, DATA_WR_IN(4) => OP_WB_4_port, 
                           DATA_WR_IN(3) => OP_WB_3_port, DATA_WR_IN(2) => 
                           OP_WB_2_port, DATA_WR_IN(1) => OP_WB_1_port, 
                           DATA_WR_IN(0) => OP_WB_0_port, PC_OUT(31) => 
                           PC_DECODE_OUT_31_port, PC_OUT(30) => 
                           PC_DECODE_OUT_30_port, PC_OUT(29) => 
                           PC_DECODE_OUT_29_port, PC_OUT(28) => 
                           PC_DECODE_OUT_28_port, PC_OUT(27) => 
                           PC_DECODE_OUT_27_port, PC_OUT(26) => 
                           PC_DECODE_OUT_26_port, PC_OUT(25) => 
                           PC_DECODE_OUT_25_port, PC_OUT(24) => 
                           PC_DECODE_OUT_24_port, PC_OUT(23) => 
                           PC_DECODE_OUT_23_port, PC_OUT(22) => 
                           PC_DECODE_OUT_22_port, PC_OUT(21) => 
                           PC_DECODE_OUT_21_port, PC_OUT(20) => 
                           PC_DECODE_OUT_20_port, PC_OUT(19) => 
                           PC_DECODE_OUT_19_port, PC_OUT(18) => 
                           PC_DECODE_OUT_18_port, PC_OUT(17) => 
                           PC_DECODE_OUT_17_port, PC_OUT(16) => 
                           PC_DECODE_OUT_16_port, PC_OUT(15) => 
                           PC_DECODE_OUT_15_port, PC_OUT(14) => 
                           PC_DECODE_OUT_14_port, PC_OUT(13) => 
                           PC_DECODE_OUT_13_port, PC_OUT(12) => 
                           PC_DECODE_OUT_12_port, PC_OUT(11) => 
                           PC_DECODE_OUT_11_port, PC_OUT(10) => 
                           PC_DECODE_OUT_10_port, PC_OUT(9) => 
                           PC_DECODE_OUT_9_port, PC_OUT(8) => 
                           PC_DECODE_OUT_8_port, PC_OUT(7) => 
                           PC_DECODE_OUT_7_port, PC_OUT(6) => 
                           PC_DECODE_OUT_6_port, PC_OUT(5) => 
                           PC_DECODE_OUT_5_port, PC_OUT(4) => 
                           PC_DECODE_OUT_4_port, PC_OUT(3) => 
                           PC_DECODE_OUT_3_port, PC_OUT(2) => 
                           PC_DECODE_OUT_2_port, PC_OUT(1) => 
                           PC_DECODE_OUT_1_port, PC_OUT(0) => 
                           PC_DECODE_OUT_0_port, A_OUT(31) => 
                           A_DECODE_OUT_31_port, A_OUT(30) => 
                           A_DECODE_OUT_30_port, A_OUT(29) => 
                           A_DECODE_OUT_29_port, A_OUT(28) => 
                           A_DECODE_OUT_28_port, A_OUT(27) => 
                           A_DECODE_OUT_27_port, A_OUT(26) => 
                           A_DECODE_OUT_26_port, A_OUT(25) => 
                           A_DECODE_OUT_25_port, A_OUT(24) => 
                           A_DECODE_OUT_24_port, A_OUT(23) => 
                           A_DECODE_OUT_23_port, A_OUT(22) => 
                           A_DECODE_OUT_22_port, A_OUT(21) => 
                           A_DECODE_OUT_21_port, A_OUT(20) => 
                           A_DECODE_OUT_20_port, A_OUT(19) => 
                           A_DECODE_OUT_19_port, A_OUT(18) => 
                           A_DECODE_OUT_18_port, A_OUT(17) => 
                           A_DECODE_OUT_17_port, A_OUT(16) => 
                           A_DECODE_OUT_16_port, A_OUT(15) => 
                           A_DECODE_OUT_15_port, A_OUT(14) => 
                           A_DECODE_OUT_14_port, A_OUT(13) => 
                           A_DECODE_OUT_13_port, A_OUT(12) => 
                           A_DECODE_OUT_12_port, A_OUT(11) => 
                           A_DECODE_OUT_11_port, A_OUT(10) => 
                           A_DECODE_OUT_10_port, A_OUT(9) => 
                           A_DECODE_OUT_9_port, A_OUT(8) => A_DECODE_OUT_8_port
                           , A_OUT(7) => A_DECODE_OUT_7_port, A_OUT(6) => 
                           A_DECODE_OUT_6_port, A_OUT(5) => A_DECODE_OUT_5_port
                           , A_OUT(4) => A_DECODE_OUT_4_port, A_OUT(3) => 
                           A_DECODE_OUT_3_port, A_OUT(2) => A_DECODE_OUT_2_port
                           , A_OUT(1) => A_DECODE_OUT_1_port, A_OUT(0) => 
                           A_DECODE_OUT_0_port, B_OUT(31) => 
                           B_DECODE_OUT_31_port, B_OUT(30) => 
                           B_DECODE_OUT_30_port, B_OUT(29) => 
                           B_DECODE_OUT_29_port, B_OUT(28) => 
                           B_DECODE_OUT_28_port, B_OUT(27) => 
                           B_DECODE_OUT_27_port, B_OUT(26) => 
                           B_DECODE_OUT_26_port, B_OUT(25) => 
                           B_DECODE_OUT_25_port, B_OUT(24) => 
                           B_DECODE_OUT_24_port, B_OUT(23) => 
                           B_DECODE_OUT_23_port, B_OUT(22) => 
                           B_DECODE_OUT_22_port, B_OUT(21) => 
                           B_DECODE_OUT_21_port, B_OUT(20) => 
                           B_DECODE_OUT_20_port, B_OUT(19) => 
                           B_DECODE_OUT_19_port, B_OUT(18) => 
                           B_DECODE_OUT_18_port, B_OUT(17) => 
                           B_DECODE_OUT_17_port, B_OUT(16) => 
                           B_DECODE_OUT_16_port, B_OUT(15) => 
                           B_DECODE_OUT_15_port, B_OUT(14) => 
                           B_DECODE_OUT_14_port, B_OUT(13) => 
                           B_DECODE_OUT_13_port, B_OUT(12) => 
                           B_DECODE_OUT_12_port, B_OUT(11) => 
                           B_DECODE_OUT_11_port, B_OUT(10) => 
                           B_DECODE_OUT_10_port, B_OUT(9) => 
                           B_DECODE_OUT_9_port, B_OUT(8) => B_DECODE_OUT_8_port
                           , B_OUT(7) => B_DECODE_OUT_7_port, B_OUT(6) => 
                           B_DECODE_OUT_6_port, B_OUT(5) => B_DECODE_OUT_5_port
                           , B_OUT(4) => B_DECODE_OUT_4_port, B_OUT(3) => 
                           B_DECODE_OUT_3_port, B_OUT(2) => B_DECODE_OUT_2_port
                           , B_OUT(1) => B_DECODE_OUT_1_port, B_OUT(0) => 
                           B_DECODE_OUT_0_port, IMM_OUT(31) => 
                           IMM_DECODE_OUT_31_port, IMM_OUT(30) => 
                           IMM_DECODE_OUT_30_port, IMM_OUT(29) => 
                           IMM_DECODE_OUT_29_port, IMM_OUT(28) => 
                           IMM_DECODE_OUT_28_port, IMM_OUT(27) => 
                           IMM_DECODE_OUT_27_port, IMM_OUT(26) => 
                           IMM_DECODE_OUT_26_port, IMM_OUT(25) => 
                           IMM_DECODE_OUT_25_port, IMM_OUT(24) => 
                           IMM_DECODE_OUT_24_port, IMM_OUT(23) => 
                           IMM_DECODE_OUT_23_port, IMM_OUT(22) => 
                           IMM_DECODE_OUT_22_port, IMM_OUT(21) => 
                           IMM_DECODE_OUT_21_port, IMM_OUT(20) => 
                           IMM_DECODE_OUT_20_port, IMM_OUT(19) => 
                           IMM_DECODE_OUT_19_port, IMM_OUT(18) => 
                           IMM_DECODE_OUT_18_port, IMM_OUT(17) => 
                           IMM_DECODE_OUT_17_port, IMM_OUT(16) => 
                           IMM_DECODE_OUT_16_port, IMM_OUT(15) => 
                           IMM_DECODE_OUT_15_port, IMM_OUT(14) => 
                           IMM_DECODE_OUT_14_port, IMM_OUT(13) => 
                           IMM_DECODE_OUT_13_port, IMM_OUT(12) => 
                           IMM_DECODE_OUT_12_port, IMM_OUT(11) => 
                           IMM_DECODE_OUT_11_port, IMM_OUT(10) => 
                           IMM_DECODE_OUT_10_port, IMM_OUT(9) => 
                           IMM_DECODE_OUT_9_port, IMM_OUT(8) => 
                           IMM_DECODE_OUT_8_port, IMM_OUT(7) => 
                           IMM_DECODE_OUT_7_port, IMM_OUT(6) => 
                           IMM_DECODE_OUT_6_port, IMM_OUT(5) => 
                           IMM_DECODE_OUT_5_port, IMM_OUT(4) => 
                           IMM_DECODE_OUT_4_port, IMM_OUT(3) => 
                           IMM_DECODE_OUT_3_port, IMM_OUT(2) => 
                           IMM_DECODE_OUT_2_port, IMM_OUT(1) => 
                           IMM_DECODE_OUT_1_port, IMM_OUT(0) => 
                           IMM_DECODE_OUT_0_port, ADD_RS1_HDU(4) => 
                           ADD_RS1_HDU_4_port, ADD_RS1_HDU(3) => 
                           ADD_RS1_HDU_3_port, ADD_RS1_HDU(2) => 
                           ADD_RS1_HDU_2_port, ADD_RS1_HDU(1) => 
                           ADD_RS1_HDU_1_port, ADD_RS1_HDU(0) => 
                           ADD_RS1_HDU_0_port, ADD_RS2_HDU(4) => 
                           ADD_RS2_HDU_4_port, ADD_RS2_HDU(3) => 
                           ADD_RS2_HDU_3_port, ADD_RS2_HDU(2) => 
                           ADD_RS2_HDU_2_port, ADD_RS2_HDU(1) => 
                           ADD_RS2_HDU_1_port, ADD_RS2_HDU(0) => 
                           ADD_RS2_HDU_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_DECODE_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_DECODE_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_DECODE_OUT_0_port, ADD_RS1_OUT(4) => 
                           ADD_RS1_DECODE_OUT_4_port, ADD_RS1_OUT(3) => 
                           ADD_RS1_DECODE_OUT_3_port, ADD_RS1_OUT(2) => 
                           ADD_RS1_DECODE_OUT_2_port, ADD_RS1_OUT(1) => 
                           ADD_RS1_DECODE_OUT_1_port, ADD_RS1_OUT(0) => 
                           ADD_RS1_DECODE_OUT_0_port, ADD_RS2_OUT(4) => 
                           ADD_RS2_DECODE_OUT_4_port, ADD_RS2_OUT(3) => 
                           ADD_RS2_DECODE_OUT_3_port, ADD_RS2_OUT(2) => 
                           ADD_RS2_DECODE_OUT_2_port, ADD_RS2_OUT(1) => 
                           ADD_RS2_DECODE_OUT_1_port, ADD_RS2_OUT(0) => 
                           ADD_RS2_DECODE_OUT_0_port);
   ExecuteStage : Execute port map( CLK => CLK, RST => RST, MUX_A_SEL => 
                           MUX_A_SEL, MUX_B_SEL(1) => MUX_B_SEL(1), 
                           MUX_B_SEL(0) => MUX_B_SEL(0), ALU_OPC(0) => 
                           ALU_OPC(0), ALU_OPC(1) => ALU_OPC(1), ALU_OPC(2) => 
                           ALU_OPC(2), ALU_OPC(3) => ALU_OPC(3), ALU_OPC(4) => 
                           ALU_OPC(4), ALU_OUTREG_EN => ALU_OUTREG_EN, 
                           JUMP_TYPE(1) => JUMP_TYPE(1), JUMP_TYPE(0) => 
                           JUMP_TYPE(0), PC_IN(31) => PC_DECODE_OUT_31_port, 
                           PC_IN(30) => PC_DECODE_OUT_30_port, PC_IN(29) => 
                           PC_DECODE_OUT_29_port, PC_IN(28) => 
                           PC_DECODE_OUT_28_port, PC_IN(27) => 
                           PC_DECODE_OUT_27_port, PC_IN(26) => 
                           PC_DECODE_OUT_26_port, PC_IN(25) => 
                           PC_DECODE_OUT_25_port, PC_IN(24) => 
                           PC_DECODE_OUT_24_port, PC_IN(23) => 
                           PC_DECODE_OUT_23_port, PC_IN(22) => 
                           PC_DECODE_OUT_22_port, PC_IN(21) => 
                           PC_DECODE_OUT_21_port, PC_IN(20) => 
                           PC_DECODE_OUT_20_port, PC_IN(19) => 
                           PC_DECODE_OUT_19_port, PC_IN(18) => 
                           PC_DECODE_OUT_18_port, PC_IN(17) => 
                           PC_DECODE_OUT_17_port, PC_IN(16) => 
                           PC_DECODE_OUT_16_port, PC_IN(15) => 
                           PC_DECODE_OUT_15_port, PC_IN(14) => 
                           PC_DECODE_OUT_14_port, PC_IN(13) => 
                           PC_DECODE_OUT_13_port, PC_IN(12) => 
                           PC_DECODE_OUT_12_port, PC_IN(11) => 
                           PC_DECODE_OUT_11_port, PC_IN(10) => 
                           PC_DECODE_OUT_10_port, PC_IN(9) => 
                           PC_DECODE_OUT_9_port, PC_IN(8) => 
                           PC_DECODE_OUT_8_port, PC_IN(7) => 
                           PC_DECODE_OUT_7_port, PC_IN(6) => 
                           PC_DECODE_OUT_6_port, PC_IN(5) => 
                           PC_DECODE_OUT_5_port, PC_IN(4) => 
                           PC_DECODE_OUT_4_port, PC_IN(3) => 
                           PC_DECODE_OUT_3_port, PC_IN(2) => 
                           PC_DECODE_OUT_2_port, PC_IN(1) => 
                           PC_DECODE_OUT_1_port, PC_IN(0) => 
                           PC_DECODE_OUT_0_port, A_IN(31) => 
                           A_DECODE_OUT_31_port, A_IN(30) => 
                           A_DECODE_OUT_30_port, A_IN(29) => 
                           A_DECODE_OUT_29_port, A_IN(28) => 
                           A_DECODE_OUT_28_port, A_IN(27) => 
                           A_DECODE_OUT_27_port, A_IN(26) => 
                           A_DECODE_OUT_26_port, A_IN(25) => 
                           A_DECODE_OUT_25_port, A_IN(24) => 
                           A_DECODE_OUT_24_port, A_IN(23) => 
                           A_DECODE_OUT_23_port, A_IN(22) => 
                           A_DECODE_OUT_22_port, A_IN(21) => 
                           A_DECODE_OUT_21_port, A_IN(20) => 
                           A_DECODE_OUT_20_port, A_IN(19) => 
                           A_DECODE_OUT_19_port, A_IN(18) => 
                           A_DECODE_OUT_18_port, A_IN(17) => 
                           A_DECODE_OUT_17_port, A_IN(16) => 
                           A_DECODE_OUT_16_port, A_IN(15) => 
                           A_DECODE_OUT_15_port, A_IN(14) => 
                           A_DECODE_OUT_14_port, A_IN(13) => 
                           A_DECODE_OUT_13_port, A_IN(12) => 
                           A_DECODE_OUT_12_port, A_IN(11) => 
                           A_DECODE_OUT_11_port, A_IN(10) => 
                           A_DECODE_OUT_10_port, A_IN(9) => A_DECODE_OUT_9_port
                           , A_IN(8) => A_DECODE_OUT_8_port, A_IN(7) => 
                           A_DECODE_OUT_7_port, A_IN(6) => A_DECODE_OUT_6_port,
                           A_IN(5) => A_DECODE_OUT_5_port, A_IN(4) => 
                           A_DECODE_OUT_4_port, A_IN(3) => A_DECODE_OUT_3_port,
                           A_IN(2) => A_DECODE_OUT_2_port, A_IN(1) => 
                           A_DECODE_OUT_1_port, A_IN(0) => A_DECODE_OUT_0_port,
                           B_IN(31) => B_DECODE_OUT_31_port, B_IN(30) => 
                           B_DECODE_OUT_30_port, B_IN(29) => 
                           B_DECODE_OUT_29_port, B_IN(28) => 
                           B_DECODE_OUT_28_port, B_IN(27) => 
                           B_DECODE_OUT_27_port, B_IN(26) => 
                           B_DECODE_OUT_26_port, B_IN(25) => 
                           B_DECODE_OUT_25_port, B_IN(24) => 
                           B_DECODE_OUT_24_port, B_IN(23) => 
                           B_DECODE_OUT_23_port, B_IN(22) => 
                           B_DECODE_OUT_22_port, B_IN(21) => 
                           B_DECODE_OUT_21_port, B_IN(20) => 
                           B_DECODE_OUT_20_port, B_IN(19) => 
                           B_DECODE_OUT_19_port, B_IN(18) => 
                           B_DECODE_OUT_18_port, B_IN(17) => 
                           B_DECODE_OUT_17_port, B_IN(16) => 
                           B_DECODE_OUT_16_port, B_IN(15) => 
                           B_DECODE_OUT_15_port, B_IN(14) => 
                           B_DECODE_OUT_14_port, B_IN(13) => 
                           B_DECODE_OUT_13_port, B_IN(12) => 
                           B_DECODE_OUT_12_port, B_IN(11) => 
                           B_DECODE_OUT_11_port, B_IN(10) => 
                           B_DECODE_OUT_10_port, B_IN(9) => B_DECODE_OUT_9_port
                           , B_IN(8) => B_DECODE_OUT_8_port, B_IN(7) => 
                           B_DECODE_OUT_7_port, B_IN(6) => B_DECODE_OUT_6_port,
                           B_IN(5) => B_DECODE_OUT_5_port, B_IN(4) => 
                           B_DECODE_OUT_4_port, B_IN(3) => B_DECODE_OUT_3_port,
                           B_IN(2) => B_DECODE_OUT_2_port, B_IN(1) => 
                           B_DECODE_OUT_1_port, B_IN(0) => B_DECODE_OUT_0_port,
                           IMM_IN(31) => IMM_DECODE_OUT_31_port, IMM_IN(30) => 
                           IMM_DECODE_OUT_30_port, IMM_IN(29) => 
                           IMM_DECODE_OUT_29_port, IMM_IN(28) => 
                           IMM_DECODE_OUT_28_port, IMM_IN(27) => 
                           IMM_DECODE_OUT_27_port, IMM_IN(26) => 
                           IMM_DECODE_OUT_26_port, IMM_IN(25) => 
                           IMM_DECODE_OUT_25_port, IMM_IN(24) => 
                           IMM_DECODE_OUT_24_port, IMM_IN(23) => 
                           IMM_DECODE_OUT_23_port, IMM_IN(22) => 
                           IMM_DECODE_OUT_22_port, IMM_IN(21) => 
                           IMM_DECODE_OUT_21_port, IMM_IN(20) => 
                           IMM_DECODE_OUT_20_port, IMM_IN(19) => 
                           IMM_DECODE_OUT_19_port, IMM_IN(18) => 
                           IMM_DECODE_OUT_18_port, IMM_IN(17) => 
                           IMM_DECODE_OUT_17_port, IMM_IN(16) => 
                           IMM_DECODE_OUT_16_port, IMM_IN(15) => 
                           IMM_DECODE_OUT_15_port, IMM_IN(14) => 
                           IMM_DECODE_OUT_14_port, IMM_IN(13) => 
                           IMM_DECODE_OUT_13_port, IMM_IN(12) => 
                           IMM_DECODE_OUT_12_port, IMM_IN(11) => 
                           IMM_DECODE_OUT_11_port, IMM_IN(10) => 
                           IMM_DECODE_OUT_10_port, IMM_IN(9) => 
                           IMM_DECODE_OUT_9_port, IMM_IN(8) => 
                           IMM_DECODE_OUT_8_port, IMM_IN(7) => 
                           IMM_DECODE_OUT_7_port, IMM_IN(6) => 
                           IMM_DECODE_OUT_6_port, IMM_IN(5) => 
                           IMM_DECODE_OUT_5_port, IMM_IN(4) => 
                           IMM_DECODE_OUT_4_port, IMM_IN(3) => 
                           IMM_DECODE_OUT_3_port, IMM_IN(2) => 
                           IMM_DECODE_OUT_2_port, IMM_IN(1) => 
                           IMM_DECODE_OUT_1_port, IMM_IN(0) => 
                           IMM_DECODE_OUT_0_port, ADD_WR_IN(4) => 
                           ADD_WR_DECODE_OUT_4_port, ADD_WR_IN(3) => 
                           ADD_WR_DECODE_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_DECODE_OUT_0_port, ADD_RS1_IN(4) => 
                           ADD_RS1_DECODE_OUT_4_port, ADD_RS1_IN(3) => 
                           ADD_RS1_DECODE_OUT_3_port, ADD_RS1_IN(2) => 
                           ADD_RS1_DECODE_OUT_2_port, ADD_RS1_IN(1) => 
                           ADD_RS1_DECODE_OUT_1_port, ADD_RS1_IN(0) => 
                           ADD_RS1_DECODE_OUT_0_port, ADD_RS2_IN(4) => 
                           ADD_RS2_DECODE_OUT_4_port, ADD_RS2_IN(3) => 
                           ADD_RS2_DECODE_OUT_3_port, ADD_RS2_IN(2) => 
                           ADD_RS2_DECODE_OUT_2_port, ADD_RS2_IN(1) => 
                           ADD_RS2_DECODE_OUT_1_port, ADD_RS2_IN(0) => 
                           ADD_RS2_DECODE_OUT_0_port, ADD_WR_MEM(4) => 
                           ADD_WR_MEM_4_port, ADD_WR_MEM(3) => 
                           ADD_WR_MEM_3_port, ADD_WR_MEM(2) => 
                           ADD_WR_MEM_2_port, ADD_WR_MEM(1) => 
                           ADD_WR_MEM_1_port, ADD_WR_MEM(0) => 
                           ADD_WR_MEM_0_port, ADD_WR_WB(4) => ADD_WR_WB_4_port,
                           ADD_WR_WB(3) => ADD_WR_WB_3_port, ADD_WR_WB(2) => 
                           ADD_WR_WB_2_port, ADD_WR_WB(1) => ADD_WR_WB_1_port, 
                           ADD_WR_WB(0) => ADD_WR_WB_0_port, RF_WE_MEM => RF_WE
                           , RF_WE_WB => RF_WE_WB, OP_MEM(31) => OP_MEM_31_port
                           , OP_MEM(30) => OP_MEM_30_port, OP_MEM(29) => 
                           OP_MEM_29_port, OP_MEM(28) => OP_MEM_28_port, 
                           OP_MEM(27) => OP_MEM_27_port, OP_MEM(26) => 
                           OP_MEM_26_port, OP_MEM(25) => OP_MEM_25_port, 
                           OP_MEM(24) => OP_MEM_24_port, OP_MEM(23) => 
                           OP_MEM_23_port, OP_MEM(22) => OP_MEM_22_port, 
                           OP_MEM(21) => OP_MEM_21_port, OP_MEM(20) => 
                           OP_MEM_20_port, OP_MEM(19) => OP_MEM_19_port, 
                           OP_MEM(18) => OP_MEM_18_port, OP_MEM(17) => 
                           OP_MEM_17_port, OP_MEM(16) => OP_MEM_16_port, 
                           OP_MEM(15) => OP_MEM_15_port, OP_MEM(14) => 
                           OP_MEM_14_port, OP_MEM(13) => OP_MEM_13_port, 
                           OP_MEM(12) => OP_MEM_12_port, OP_MEM(11) => 
                           OP_MEM_11_port, OP_MEM(10) => OP_MEM_10_port, 
                           OP_MEM(9) => OP_MEM_9_port, OP_MEM(8) => 
                           OP_MEM_8_port, OP_MEM(7) => OP_MEM_7_port, OP_MEM(6)
                           => OP_MEM_6_port, OP_MEM(5) => OP_MEM_5_port, 
                           OP_MEM(4) => OP_MEM_4_port, OP_MEM(3) => 
                           OP_MEM_3_port, OP_MEM(2) => OP_MEM_2_port, OP_MEM(1)
                           => OP_MEM_1_port, OP_MEM(0) => OP_MEM_0_port, 
                           OP_WB(31) => OP_WB_31_port, OP_WB(30) => 
                           OP_WB_30_port, OP_WB(29) => OP_WB_29_port, OP_WB(28)
                           => OP_WB_28_port, OP_WB(27) => OP_WB_27_port, 
                           OP_WB(26) => OP_WB_26_port, OP_WB(25) => 
                           OP_WB_25_port, OP_WB(24) => OP_WB_24_port, OP_WB(23)
                           => OP_WB_23_port, OP_WB(22) => OP_WB_22_port, 
                           OP_WB(21) => OP_WB_21_port, OP_WB(20) => 
                           OP_WB_20_port, OP_WB(19) => OP_WB_19_port, OP_WB(18)
                           => OP_WB_18_port, OP_WB(17) => OP_WB_17_port, 
                           OP_WB(16) => OP_WB_16_port, OP_WB(15) => 
                           OP_WB_15_port, OP_WB(14) => OP_WB_14_port, OP_WB(13)
                           => OP_WB_13_port, OP_WB(12) => OP_WB_12_port, 
                           OP_WB(11) => OP_WB_11_port, OP_WB(10) => 
                           OP_WB_10_port, OP_WB(9) => OP_WB_9_port, OP_WB(8) =>
                           OP_WB_8_port, OP_WB(7) => OP_WB_7_port, OP_WB(6) => 
                           OP_WB_6_port, OP_WB(5) => OP_WB_5_port, OP_WB(4) => 
                           OP_WB_4_port, OP_WB(3) => OP_WB_3_port, OP_WB(2) => 
                           OP_WB_2_port, OP_WB(1) => OP_WB_1_port, OP_WB(0) => 
                           OP_WB_0_port, PC_SEL(1) => PC_SEL_EX_1_port, 
                           PC_SEL(0) => PC_SEL_EX_0_port, ZERO_FLAG => 
                           ZERO_FLAG_EX, NPC_ABS(31) => NPC_ABS_EX_31_port, 
                           NPC_ABS(30) => NPC_ABS_EX_30_port, NPC_ABS(29) => 
                           NPC_ABS_EX_29_port, NPC_ABS(28) => 
                           NPC_ABS_EX_28_port, NPC_ABS(27) => 
                           NPC_ABS_EX_27_port, NPC_ABS(26) => 
                           NPC_ABS_EX_26_port, NPC_ABS(25) => 
                           NPC_ABS_EX_25_port, NPC_ABS(24) => 
                           NPC_ABS_EX_24_port, NPC_ABS(23) => 
                           NPC_ABS_EX_23_port, NPC_ABS(22) => 
                           NPC_ABS_EX_22_port, NPC_ABS(21) => 
                           NPC_ABS_EX_21_port, NPC_ABS(20) => 
                           NPC_ABS_EX_20_port, NPC_ABS(19) => 
                           NPC_ABS_EX_19_port, NPC_ABS(18) => 
                           NPC_ABS_EX_18_port, NPC_ABS(17) => 
                           NPC_ABS_EX_17_port, NPC_ABS(16) => 
                           NPC_ABS_EX_16_port, NPC_ABS(15) => 
                           NPC_ABS_EX_15_port, NPC_ABS(14) => 
                           NPC_ABS_EX_14_port, NPC_ABS(13) => 
                           NPC_ABS_EX_13_port, NPC_ABS(12) => 
                           NPC_ABS_EX_12_port, NPC_ABS(11) => 
                           NPC_ABS_EX_11_port, NPC_ABS(10) => 
                           NPC_ABS_EX_10_port, NPC_ABS(9) => NPC_ABS_EX_9_port,
                           NPC_ABS(8) => NPC_ABS_EX_8_port, NPC_ABS(7) => 
                           NPC_ABS_EX_7_port, NPC_ABS(6) => NPC_ABS_EX_6_port, 
                           NPC_ABS(5) => NPC_ABS_EX_5_port, NPC_ABS(4) => 
                           NPC_ABS_EX_4_port, NPC_ABS(3) => NPC_ABS_EX_3_port, 
                           NPC_ABS(2) => NPC_ABS_EX_2_port, NPC_ABS(1) => 
                           NPC_ABS_EX_1_port, NPC_ABS(0) => NPC_ABS_EX_0_port, 
                           NPC_REL(31) => NPC_REL_EX_31_port, NPC_REL(30) => 
                           NPC_REL_EX_30_port, NPC_REL(29) => 
                           NPC_REL_EX_29_port, NPC_REL(28) => 
                           NPC_REL_EX_28_port, NPC_REL(27) => 
                           NPC_REL_EX_27_port, NPC_REL(26) => 
                           NPC_REL_EX_26_port, NPC_REL(25) => 
                           NPC_REL_EX_25_port, NPC_REL(24) => 
                           NPC_REL_EX_24_port, NPC_REL(23) => 
                           NPC_REL_EX_23_port, NPC_REL(22) => 
                           NPC_REL_EX_22_port, NPC_REL(21) => 
                           NPC_REL_EX_21_port, NPC_REL(20) => 
                           NPC_REL_EX_20_port, NPC_REL(19) => 
                           NPC_REL_EX_19_port, NPC_REL(18) => 
                           NPC_REL_EX_18_port, NPC_REL(17) => 
                           NPC_REL_EX_17_port, NPC_REL(16) => 
                           NPC_REL_EX_16_port, NPC_REL(15) => 
                           NPC_REL_EX_15_port, NPC_REL(14) => 
                           NPC_REL_EX_14_port, NPC_REL(13) => 
                           NPC_REL_EX_13_port, NPC_REL(12) => 
                           NPC_REL_EX_12_port, NPC_REL(11) => 
                           NPC_REL_EX_11_port, NPC_REL(10) => 
                           NPC_REL_EX_10_port, NPC_REL(9) => NPC_REL_EX_9_port,
                           NPC_REL(8) => NPC_REL_EX_8_port, NPC_REL(7) => 
                           NPC_REL_EX_7_port, NPC_REL(6) => NPC_REL_EX_6_port, 
                           NPC_REL(5) => NPC_REL_EX_5_port, NPC_REL(4) => 
                           NPC_REL_EX_4_port, NPC_REL(3) => NPC_REL_EX_3_port, 
                           NPC_REL(2) => NPC_REL_EX_2_port, NPC_REL(1) => 
                           NPC_REL_EX_1_port, NPC_REL(0) => NPC_REL_EX_0_port, 
                           ALU_RES(31) => ALU_RES_EX_31_port, ALU_RES(30) => 
                           ALU_RES_EX_30_port, ALU_RES(29) => 
                           ALU_RES_EX_29_port, ALU_RES(28) => 
                           ALU_RES_EX_28_port, ALU_RES(27) => 
                           ALU_RES_EX_27_port, ALU_RES(26) => 
                           ALU_RES_EX_26_port, ALU_RES(25) => 
                           ALU_RES_EX_25_port, ALU_RES(24) => 
                           ALU_RES_EX_24_port, ALU_RES(23) => 
                           ALU_RES_EX_23_port, ALU_RES(22) => 
                           ALU_RES_EX_22_port, ALU_RES(21) => 
                           ALU_RES_EX_21_port, ALU_RES(20) => 
                           ALU_RES_EX_20_port, ALU_RES(19) => 
                           ALU_RES_EX_19_port, ALU_RES(18) => 
                           ALU_RES_EX_18_port, ALU_RES(17) => 
                           ALU_RES_EX_17_port, ALU_RES(16) => 
                           ALU_RES_EX_16_port, ALU_RES(15) => 
                           ALU_RES_EX_15_port, ALU_RES(14) => 
                           ALU_RES_EX_14_port, ALU_RES(13) => 
                           ALU_RES_EX_13_port, ALU_RES(12) => 
                           ALU_RES_EX_12_port, ALU_RES(11) => 
                           ALU_RES_EX_11_port, ALU_RES(10) => 
                           ALU_RES_EX_10_port, ALU_RES(9) => ALU_RES_EX_9_port,
                           ALU_RES(8) => ALU_RES_EX_8_port, ALU_RES(7) => 
                           ALU_RES_EX_7_port, ALU_RES(6) => ALU_RES_EX_6_port, 
                           ALU_RES(5) => ALU_RES_EX_5_port, ALU_RES(4) => 
                           ALU_RES_EX_4_port, ALU_RES(3) => ALU_RES_EX_3_port, 
                           ALU_RES(2) => ALU_RES_EX_2_port, ALU_RES(1) => 
                           ALU_RES_EX_1_port, ALU_RES(0) => ALU_RES_EX_0_port, 
                           B_OUT(31) => B_EX_OUT_31_port, B_OUT(30) => 
                           B_EX_OUT_30_port, B_OUT(29) => B_EX_OUT_29_port, 
                           B_OUT(28) => B_EX_OUT_28_port, B_OUT(27) => 
                           B_EX_OUT_27_port, B_OUT(26) => B_EX_OUT_26_port, 
                           B_OUT(25) => B_EX_OUT_25_port, B_OUT(24) => 
                           B_EX_OUT_24_port, B_OUT(23) => B_EX_OUT_23_port, 
                           B_OUT(22) => B_EX_OUT_22_port, B_OUT(21) => 
                           B_EX_OUT_21_port, B_OUT(20) => B_EX_OUT_20_port, 
                           B_OUT(19) => B_EX_OUT_19_port, B_OUT(18) => 
                           B_EX_OUT_18_port, B_OUT(17) => B_EX_OUT_17_port, 
                           B_OUT(16) => B_EX_OUT_16_port, B_OUT(15) => 
                           B_EX_OUT_15_port, B_OUT(14) => B_EX_OUT_14_port, 
                           B_OUT(13) => B_EX_OUT_13_port, B_OUT(12) => 
                           B_EX_OUT_12_port, B_OUT(11) => B_EX_OUT_11_port, 
                           B_OUT(10) => B_EX_OUT_10_port, B_OUT(9) => 
                           B_EX_OUT_9_port, B_OUT(8) => B_EX_OUT_8_port, 
                           B_OUT(7) => B_EX_OUT_7_port, B_OUT(6) => 
                           B_EX_OUT_6_port, B_OUT(5) => B_EX_OUT_5_port, 
                           B_OUT(4) => B_EX_OUT_4_port, B_OUT(3) => 
                           B_EX_OUT_3_port, B_OUT(2) => B_EX_OUT_2_port, 
                           B_OUT(1) => B_EX_OUT_1_port, B_OUT(0) => 
                           B_EX_OUT_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_EX_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_EX_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_EX_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_EX_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_EX_OUT_0_port);
   DRAM_R_ff : ff_0 port map( D => DRAM_R_IN, CLK => CLK, EN => X_Logic1_port, 
                           RST => RST, Q => DRAM_R_MEM);
   MemoryStage : Memory port map( CLK => CLK, RST => RST, MEM_EN_IN => 
                           MEM_EN_IN, DRAM_R_IN => DRAM_R_MEM, DRAM_W_IN => 
                           DRAM_W_IN, PC_SEL(1) => PC_SEL_EX_1_port, PC_SEL(0) 
                           => PC_SEL_EX_0_port, NPC_IN(31) => 
                           NPC_FETCH_OUT_31_port, NPC_IN(30) => 
                           NPC_FETCH_OUT_30_port, NPC_IN(29) => 
                           NPC_FETCH_OUT_29_port, NPC_IN(28) => 
                           NPC_FETCH_OUT_28_port, NPC_IN(27) => 
                           NPC_FETCH_OUT_27_port, NPC_IN(26) => 
                           NPC_FETCH_OUT_26_port, NPC_IN(25) => 
                           NPC_FETCH_OUT_25_port, NPC_IN(24) => 
                           NPC_FETCH_OUT_24_port, NPC_IN(23) => 
                           NPC_FETCH_OUT_23_port, NPC_IN(22) => 
                           NPC_FETCH_OUT_22_port, NPC_IN(21) => 
                           NPC_FETCH_OUT_21_port, NPC_IN(20) => 
                           NPC_FETCH_OUT_20_port, NPC_IN(19) => 
                           NPC_FETCH_OUT_19_port, NPC_IN(18) => 
                           NPC_FETCH_OUT_18_port, NPC_IN(17) => 
                           NPC_FETCH_OUT_17_port, NPC_IN(16) => 
                           NPC_FETCH_OUT_16_port, NPC_IN(15) => 
                           NPC_FETCH_OUT_15_port, NPC_IN(14) => 
                           NPC_FETCH_OUT_14_port, NPC_IN(13) => 
                           NPC_FETCH_OUT_13_port, NPC_IN(12) => 
                           NPC_FETCH_OUT_12_port, NPC_IN(11) => 
                           NPC_FETCH_OUT_11_port, NPC_IN(10) => 
                           NPC_FETCH_OUT_10_port, NPC_IN(9) => 
                           NPC_FETCH_OUT_9_port, NPC_IN(8) => 
                           NPC_FETCH_OUT_8_port, NPC_IN(7) => 
                           NPC_FETCH_OUT_7_port, NPC_IN(6) => 
                           NPC_FETCH_OUT_6_port, NPC_IN(5) => 
                           NPC_FETCH_OUT_5_port, NPC_IN(4) => 
                           NPC_FETCH_OUT_4_port, NPC_IN(3) => 
                           NPC_FETCH_OUT_3_port, NPC_IN(2) => 
                           NPC_FETCH_OUT_2_port, NPC_IN(1) => 
                           NPC_FETCH_OUT_1_port, NPC_IN(0) => 
                           NPC_FETCH_OUT_0_port, NPC_ABS(31) => 
                           NPC_ABS_EX_31_port, NPC_ABS(30) => 
                           NPC_ABS_EX_30_port, NPC_ABS(29) => 
                           NPC_ABS_EX_29_port, NPC_ABS(28) => 
                           NPC_ABS_EX_28_port, NPC_ABS(27) => 
                           NPC_ABS_EX_27_port, NPC_ABS(26) => 
                           NPC_ABS_EX_26_port, NPC_ABS(25) => 
                           NPC_ABS_EX_25_port, NPC_ABS(24) => 
                           NPC_ABS_EX_24_port, NPC_ABS(23) => 
                           NPC_ABS_EX_23_port, NPC_ABS(22) => 
                           NPC_ABS_EX_22_port, NPC_ABS(21) => 
                           NPC_ABS_EX_21_port, NPC_ABS(20) => 
                           NPC_ABS_EX_20_port, NPC_ABS(19) => 
                           NPC_ABS_EX_19_port, NPC_ABS(18) => 
                           NPC_ABS_EX_18_port, NPC_ABS(17) => 
                           NPC_ABS_EX_17_port, NPC_ABS(16) => 
                           NPC_ABS_EX_16_port, NPC_ABS(15) => 
                           NPC_ABS_EX_15_port, NPC_ABS(14) => 
                           NPC_ABS_EX_14_port, NPC_ABS(13) => 
                           NPC_ABS_EX_13_port, NPC_ABS(12) => 
                           NPC_ABS_EX_12_port, NPC_ABS(11) => 
                           NPC_ABS_EX_11_port, NPC_ABS(10) => 
                           NPC_ABS_EX_10_port, NPC_ABS(9) => NPC_ABS_EX_9_port,
                           NPC_ABS(8) => NPC_ABS_EX_8_port, NPC_ABS(7) => 
                           NPC_ABS_EX_7_port, NPC_ABS(6) => NPC_ABS_EX_6_port, 
                           NPC_ABS(5) => NPC_ABS_EX_5_port, NPC_ABS(4) => 
                           NPC_ABS_EX_4_port, NPC_ABS(3) => NPC_ABS_EX_3_port, 
                           NPC_ABS(2) => NPC_ABS_EX_2_port, NPC_ABS(1) => 
                           NPC_ABS_EX_1_port, NPC_ABS(0) => NPC_ABS_EX_0_port, 
                           NPC_REL(31) => NPC_REL_EX_31_port, NPC_REL(30) => 
                           NPC_REL_EX_30_port, NPC_REL(29) => 
                           NPC_REL_EX_29_port, NPC_REL(28) => 
                           NPC_REL_EX_28_port, NPC_REL(27) => 
                           NPC_REL_EX_27_port, NPC_REL(26) => 
                           NPC_REL_EX_26_port, NPC_REL(25) => 
                           NPC_REL_EX_25_port, NPC_REL(24) => 
                           NPC_REL_EX_24_port, NPC_REL(23) => 
                           NPC_REL_EX_23_port, NPC_REL(22) => 
                           NPC_REL_EX_22_port, NPC_REL(21) => 
                           NPC_REL_EX_21_port, NPC_REL(20) => 
                           NPC_REL_EX_20_port, NPC_REL(19) => 
                           NPC_REL_EX_19_port, NPC_REL(18) => 
                           NPC_REL_EX_18_port, NPC_REL(17) => 
                           NPC_REL_EX_17_port, NPC_REL(16) => 
                           NPC_REL_EX_16_port, NPC_REL(15) => 
                           NPC_REL_EX_15_port, NPC_REL(14) => 
                           NPC_REL_EX_14_port, NPC_REL(13) => 
                           NPC_REL_EX_13_port, NPC_REL(12) => 
                           NPC_REL_EX_12_port, NPC_REL(11) => 
                           NPC_REL_EX_11_port, NPC_REL(10) => 
                           NPC_REL_EX_10_port, NPC_REL(9) => NPC_REL_EX_9_port,
                           NPC_REL(8) => NPC_REL_EX_8_port, NPC_REL(7) => 
                           NPC_REL_EX_7_port, NPC_REL(6) => NPC_REL_EX_6_port, 
                           NPC_REL(5) => NPC_REL_EX_5_port, NPC_REL(4) => 
                           NPC_REL_EX_4_port, NPC_REL(3) => NPC_REL_EX_3_port, 
                           NPC_REL(2) => NPC_REL_EX_2_port, NPC_REL(1) => 
                           NPC_REL_EX_1_port, NPC_REL(0) => NPC_REL_EX_0_port, 
                           ALU_RES_IN(31) => ALU_RES_EX_31_port, ALU_RES_IN(30)
                           => ALU_RES_EX_30_port, ALU_RES_IN(29) => 
                           ALU_RES_EX_29_port, ALU_RES_IN(28) => 
                           ALU_RES_EX_28_port, ALU_RES_IN(27) => 
                           ALU_RES_EX_27_port, ALU_RES_IN(26) => 
                           ALU_RES_EX_26_port, ALU_RES_IN(25) => 
                           ALU_RES_EX_25_port, ALU_RES_IN(24) => 
                           ALU_RES_EX_24_port, ALU_RES_IN(23) => 
                           ALU_RES_EX_23_port, ALU_RES_IN(22) => 
                           ALU_RES_EX_22_port, ALU_RES_IN(21) => 
                           ALU_RES_EX_21_port, ALU_RES_IN(20) => 
                           ALU_RES_EX_20_port, ALU_RES_IN(19) => 
                           ALU_RES_EX_19_port, ALU_RES_IN(18) => 
                           ALU_RES_EX_18_port, ALU_RES_IN(17) => 
                           ALU_RES_EX_17_port, ALU_RES_IN(16) => 
                           ALU_RES_EX_16_port, ALU_RES_IN(15) => 
                           ALU_RES_EX_15_port, ALU_RES_IN(14) => 
                           ALU_RES_EX_14_port, ALU_RES_IN(13) => 
                           ALU_RES_EX_13_port, ALU_RES_IN(12) => 
                           ALU_RES_EX_12_port, ALU_RES_IN(11) => 
                           ALU_RES_EX_11_port, ALU_RES_IN(10) => 
                           ALU_RES_EX_10_port, ALU_RES_IN(9) => 
                           ALU_RES_EX_9_port, ALU_RES_IN(8) => 
                           ALU_RES_EX_8_port, ALU_RES_IN(7) => 
                           ALU_RES_EX_7_port, ALU_RES_IN(6) => 
                           ALU_RES_EX_6_port, ALU_RES_IN(5) => 
                           ALU_RES_EX_5_port, ALU_RES_IN(4) => 
                           ALU_RES_EX_4_port, ALU_RES_IN(3) => 
                           ALU_RES_EX_3_port, ALU_RES_IN(2) => 
                           ALU_RES_EX_2_port, ALU_RES_IN(1) => 
                           ALU_RES_EX_1_port, ALU_RES_IN(0) => 
                           ALU_RES_EX_0_port, B_IN(31) => B_EX_OUT_31_port, 
                           B_IN(30) => B_EX_OUT_30_port, B_IN(29) => 
                           B_EX_OUT_29_port, B_IN(28) => B_EX_OUT_28_port, 
                           B_IN(27) => B_EX_OUT_27_port, B_IN(26) => 
                           B_EX_OUT_26_port, B_IN(25) => B_EX_OUT_25_port, 
                           B_IN(24) => B_EX_OUT_24_port, B_IN(23) => 
                           B_EX_OUT_23_port, B_IN(22) => B_EX_OUT_22_port, 
                           B_IN(21) => B_EX_OUT_21_port, B_IN(20) => 
                           B_EX_OUT_20_port, B_IN(19) => B_EX_OUT_19_port, 
                           B_IN(18) => B_EX_OUT_18_port, B_IN(17) => 
                           B_EX_OUT_17_port, B_IN(16) => B_EX_OUT_16_port, 
                           B_IN(15) => B_EX_OUT_15_port, B_IN(14) => 
                           B_EX_OUT_14_port, B_IN(13) => B_EX_OUT_13_port, 
                           B_IN(12) => B_EX_OUT_12_port, B_IN(11) => 
                           B_EX_OUT_11_port, B_IN(10) => B_EX_OUT_10_port, 
                           B_IN(9) => B_EX_OUT_9_port, B_IN(8) => 
                           B_EX_OUT_8_port, B_IN(7) => B_EX_OUT_7_port, B_IN(6)
                           => B_EX_OUT_6_port, B_IN(5) => B_EX_OUT_5_port, 
                           B_IN(4) => B_EX_OUT_4_port, B_IN(3) => 
                           B_EX_OUT_3_port, B_IN(2) => B_EX_OUT_2_port, B_IN(1)
                           => B_EX_OUT_1_port, B_IN(0) => B_EX_OUT_0_port, 
                           ADD_WR_IN(4) => ADD_WR_EX_OUT_4_port, ADD_WR_IN(3) 
                           => ADD_WR_EX_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_EX_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_EX_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_EX_OUT_0_port, DRAM_DATA_IN(31) => 
                           DATA_IN(31), DRAM_DATA_IN(30) => DATA_IN(30), 
                           DRAM_DATA_IN(29) => DATA_IN(29), DRAM_DATA_IN(28) =>
                           DATA_IN(28), DRAM_DATA_IN(27) => DATA_IN(27), 
                           DRAM_DATA_IN(26) => DATA_IN(26), DRAM_DATA_IN(25) =>
                           DATA_IN(25), DRAM_DATA_IN(24) => DATA_IN(24), 
                           DRAM_DATA_IN(23) => DATA_IN(23), DRAM_DATA_IN(22) =>
                           DATA_IN(22), DRAM_DATA_IN(21) => DATA_IN(21), 
                           DRAM_DATA_IN(20) => DATA_IN(20), DRAM_DATA_IN(19) =>
                           DATA_IN(19), DRAM_DATA_IN(18) => DATA_IN(18), 
                           DRAM_DATA_IN(17) => DATA_IN(17), DRAM_DATA_IN(16) =>
                           DATA_IN(16), DRAM_DATA_IN(15) => DATA_IN(15), 
                           DRAM_DATA_IN(14) => DATA_IN(14), DRAM_DATA_IN(13) =>
                           DATA_IN(13), DRAM_DATA_IN(12) => DATA_IN(12), 
                           DRAM_DATA_IN(11) => DATA_IN(11), DRAM_DATA_IN(10) =>
                           DATA_IN(10), DRAM_DATA_IN(9) => DATA_IN(9), 
                           DRAM_DATA_IN(8) => DATA_IN(8), DRAM_DATA_IN(7) => 
                           DATA_IN(7), DRAM_DATA_IN(6) => DATA_IN(6), 
                           DRAM_DATA_IN(5) => DATA_IN(5), DRAM_DATA_IN(4) => 
                           DATA_IN(4), DRAM_DATA_IN(3) => DATA_IN(3), 
                           DRAM_DATA_IN(2) => DATA_IN(2), DRAM_DATA_IN(1) => 
                           DATA_IN(1), DRAM_DATA_IN(0) => DATA_IN(0), 
                           LOAD_TYPE_IN(1) => LOAD_TYPE_IN(1), LOAD_TYPE_IN(0) 
                           => LOAD_TYPE_IN(0), STORE_TYPE_IN => STORE_TYPE_IN, 
                           PC_OUT(31) => PC_MEM_OUT_31_port, PC_OUT(30) => 
                           PC_MEM_OUT_30_port, PC_OUT(29) => PC_MEM_OUT_29_port
                           , PC_OUT(28) => PC_MEM_OUT_28_port, PC_OUT(27) => 
                           PC_MEM_OUT_27_port, PC_OUT(26) => PC_MEM_OUT_26_port
                           , PC_OUT(25) => PC_MEM_OUT_25_port, PC_OUT(24) => 
                           PC_MEM_OUT_24_port, PC_OUT(23) => PC_MEM_OUT_23_port
                           , PC_OUT(22) => PC_MEM_OUT_22_port, PC_OUT(21) => 
                           PC_MEM_OUT_21_port, PC_OUT(20) => PC_MEM_OUT_20_port
                           , PC_OUT(19) => PC_MEM_OUT_19_port, PC_OUT(18) => 
                           PC_MEM_OUT_18_port, PC_OUT(17) => PC_MEM_OUT_17_port
                           , PC_OUT(16) => PC_MEM_OUT_16_port, PC_OUT(15) => 
                           PC_MEM_OUT_15_port, PC_OUT(14) => PC_MEM_OUT_14_port
                           , PC_OUT(13) => PC_MEM_OUT_13_port, PC_OUT(12) => 
                           PC_MEM_OUT_12_port, PC_OUT(11) => PC_MEM_OUT_11_port
                           , PC_OUT(10) => PC_MEM_OUT_10_port, PC_OUT(9) => 
                           PC_MEM_OUT_9_port, PC_OUT(8) => PC_MEM_OUT_8_port, 
                           PC_OUT(7) => PC_MEM_OUT_7_port, PC_OUT(6) => 
                           PC_MEM_OUT_6_port, PC_OUT(5) => PC_MEM_OUT_5_port, 
                           PC_OUT(4) => PC_MEM_OUT_4_port, PC_OUT(3) => 
                           PC_MEM_OUT_3_port, PC_OUT(2) => PC_MEM_OUT_2_port, 
                           PC_OUT(1) => PC_MEM_OUT_1_port, PC_OUT(0) => 
                           PC_MEM_OUT_0_port, DRAM_R_OUT => DRAM_R_OUT, 
                           DRAM_W_OUT => DRAM_W_OUT, DRAM_ADDR_OUT(31) => 
                           DRAM_ADDR_OUT(31), DRAM_ADDR_OUT(30) => 
                           DRAM_ADDR_OUT(30), DRAM_ADDR_OUT(29) => 
                           DRAM_ADDR_OUT(29), DRAM_ADDR_OUT(28) => 
                           DRAM_ADDR_OUT(28), DRAM_ADDR_OUT(27) => 
                           DRAM_ADDR_OUT(27), DRAM_ADDR_OUT(26) => 
                           DRAM_ADDR_OUT(26), DRAM_ADDR_OUT(25) => 
                           DRAM_ADDR_OUT(25), DRAM_ADDR_OUT(24) => 
                           DRAM_ADDR_OUT(24), DRAM_ADDR_OUT(23) => 
                           DRAM_ADDR_OUT(23), DRAM_ADDR_OUT(22) => 
                           DRAM_ADDR_OUT(22), DRAM_ADDR_OUT(21) => 
                           DRAM_ADDR_OUT(21), DRAM_ADDR_OUT(20) => 
                           DRAM_ADDR_OUT(20), DRAM_ADDR_OUT(19) => 
                           DRAM_ADDR_OUT(19), DRAM_ADDR_OUT(18) => 
                           DRAM_ADDR_OUT(18), DRAM_ADDR_OUT(17) => 
                           DRAM_ADDR_OUT(17), DRAM_ADDR_OUT(16) => 
                           DRAM_ADDR_OUT(16), DRAM_ADDR_OUT(15) => 
                           DRAM_ADDR_OUT(15), DRAM_ADDR_OUT(14) => 
                           DRAM_ADDR_OUT(14), DRAM_ADDR_OUT(13) => 
                           DRAM_ADDR_OUT(13), DRAM_ADDR_OUT(12) => 
                           DRAM_ADDR_OUT(12), DRAM_ADDR_OUT(11) => 
                           DRAM_ADDR_OUT(11), DRAM_ADDR_OUT(10) => 
                           DRAM_ADDR_OUT(10), DRAM_ADDR_OUT(9) => 
                           DRAM_ADDR_OUT(9), DRAM_ADDR_OUT(8) => 
                           DRAM_ADDR_OUT(8), DRAM_ADDR_OUT(7) => 
                           DRAM_ADDR_OUT(7), DRAM_ADDR_OUT(6) => 
                           DRAM_ADDR_OUT(6), DRAM_ADDR_OUT(5) => 
                           DRAM_ADDR_OUT(5), DRAM_ADDR_OUT(4) => 
                           DRAM_ADDR_OUT(4), DRAM_ADDR_OUT(3) => 
                           DRAM_ADDR_OUT(3), DRAM_ADDR_OUT(2) => 
                           DRAM_ADDR_OUT(2), DRAM_ADDR_OUT(1) => 
                           DRAM_ADDR_OUT(1), DRAM_ADDR_OUT(0) => 
                           DRAM_ADDR_OUT(0), DRAM_DATA_OUT(31) => DATA_OUT(31),
                           DRAM_DATA_OUT(30) => DATA_OUT(30), DRAM_DATA_OUT(29)
                           => DATA_OUT(29), DRAM_DATA_OUT(28) => DATA_OUT(28), 
                           DRAM_DATA_OUT(27) => DATA_OUT(27), DRAM_DATA_OUT(26)
                           => DATA_OUT(26), DRAM_DATA_OUT(25) => DATA_OUT(25), 
                           DRAM_DATA_OUT(24) => DATA_OUT(24), DRAM_DATA_OUT(23)
                           => DATA_OUT(23), DRAM_DATA_OUT(22) => DATA_OUT(22), 
                           DRAM_DATA_OUT(21) => DATA_OUT(21), DRAM_DATA_OUT(20)
                           => DATA_OUT(20), DRAM_DATA_OUT(19) => DATA_OUT(19), 
                           DRAM_DATA_OUT(18) => DATA_OUT(18), DRAM_DATA_OUT(17)
                           => DATA_OUT(17), DRAM_DATA_OUT(16) => DATA_OUT(16), 
                           DRAM_DATA_OUT(15) => DATA_OUT(15), DRAM_DATA_OUT(14)
                           => DATA_OUT(14), DRAM_DATA_OUT(13) => DATA_OUT(13), 
                           DRAM_DATA_OUT(12) => DATA_OUT(12), DRAM_DATA_OUT(11)
                           => DATA_OUT(11), DRAM_DATA_OUT(10) => DATA_OUT(10), 
                           DRAM_DATA_OUT(9) => DATA_OUT(9), DRAM_DATA_OUT(8) =>
                           DATA_OUT(8), DRAM_DATA_OUT(7) => DATA_OUT(7), 
                           DRAM_DATA_OUT(6) => DATA_OUT(6), DRAM_DATA_OUT(5) =>
                           DATA_OUT(5), DRAM_DATA_OUT(4) => DATA_OUT(4), 
                           DRAM_DATA_OUT(3) => DATA_OUT(3), DRAM_DATA_OUT(2) =>
                           DATA_OUT(2), DRAM_DATA_OUT(1) => DATA_OUT(1), 
                           DRAM_DATA_OUT(0) => DATA_OUT(0), DATA_OUT(31) => 
                           DATA_MEM_OUT_31_port, DATA_OUT(30) => 
                           DATA_MEM_OUT_30_port, DATA_OUT(29) => 
                           DATA_MEM_OUT_29_port, DATA_OUT(28) => 
                           DATA_MEM_OUT_28_port, DATA_OUT(27) => 
                           DATA_MEM_OUT_27_port, DATA_OUT(26) => 
                           DATA_MEM_OUT_26_port, DATA_OUT(25) => 
                           DATA_MEM_OUT_25_port, DATA_OUT(24) => 
                           DATA_MEM_OUT_24_port, DATA_OUT(23) => 
                           DATA_MEM_OUT_23_port, DATA_OUT(22) => 
                           DATA_MEM_OUT_22_port, DATA_OUT(21) => 
                           DATA_MEM_OUT_21_port, DATA_OUT(20) => 
                           DATA_MEM_OUT_20_port, DATA_OUT(19) => 
                           DATA_MEM_OUT_19_port, DATA_OUT(18) => 
                           DATA_MEM_OUT_18_port, DATA_OUT(17) => 
                           DATA_MEM_OUT_17_port, DATA_OUT(16) => 
                           DATA_MEM_OUT_16_port, DATA_OUT(15) => 
                           DATA_MEM_OUT_15_port, DATA_OUT(14) => 
                           DATA_MEM_OUT_14_port, DATA_OUT(13) => 
                           DATA_MEM_OUT_13_port, DATA_OUT(12) => 
                           DATA_MEM_OUT_12_port, DATA_OUT(11) => 
                           DATA_MEM_OUT_11_port, DATA_OUT(10) => 
                           DATA_MEM_OUT_10_port, DATA_OUT(9) => 
                           DATA_MEM_OUT_9_port, DATA_OUT(8) => 
                           DATA_MEM_OUT_8_port, DATA_OUT(7) => 
                           DATA_MEM_OUT_7_port, DATA_OUT(6) => 
                           DATA_MEM_OUT_6_port, DATA_OUT(5) => 
                           DATA_MEM_OUT_5_port, DATA_OUT(4) => 
                           DATA_MEM_OUT_4_port, DATA_OUT(3) => 
                           DATA_MEM_OUT_3_port, DATA_OUT(2) => 
                           DATA_MEM_OUT_2_port, DATA_OUT(1) => 
                           DATA_MEM_OUT_1_port, DATA_OUT(0) => 
                           DATA_MEM_OUT_0_port, ALU_RES_OUT(31) => 
                           ALU_RES_MEM_31_port, ALU_RES_OUT(30) => 
                           ALU_RES_MEM_30_port, ALU_RES_OUT(29) => 
                           ALU_RES_MEM_29_port, ALU_RES_OUT(28) => 
                           ALU_RES_MEM_28_port, ALU_RES_OUT(27) => 
                           ALU_RES_MEM_27_port, ALU_RES_OUT(26) => 
                           ALU_RES_MEM_26_port, ALU_RES_OUT(25) => 
                           ALU_RES_MEM_25_port, ALU_RES_OUT(24) => 
                           ALU_RES_MEM_24_port, ALU_RES_OUT(23) => 
                           ALU_RES_MEM_23_port, ALU_RES_OUT(22) => 
                           ALU_RES_MEM_22_port, ALU_RES_OUT(21) => 
                           ALU_RES_MEM_21_port, ALU_RES_OUT(20) => 
                           ALU_RES_MEM_20_port, ALU_RES_OUT(19) => 
                           ALU_RES_MEM_19_port, ALU_RES_OUT(18) => 
                           ALU_RES_MEM_18_port, ALU_RES_OUT(17) => 
                           ALU_RES_MEM_17_port, ALU_RES_OUT(16) => 
                           ALU_RES_MEM_16_port, ALU_RES_OUT(15) => 
                           ALU_RES_MEM_15_port, ALU_RES_OUT(14) => 
                           ALU_RES_MEM_14_port, ALU_RES_OUT(13) => 
                           ALU_RES_MEM_13_port, ALU_RES_OUT(12) => 
                           ALU_RES_MEM_12_port, ALU_RES_OUT(11) => 
                           ALU_RES_MEM_11_port, ALU_RES_OUT(10) => 
                           ALU_RES_MEM_10_port, ALU_RES_OUT(9) => 
                           ALU_RES_MEM_9_port, ALU_RES_OUT(8) => 
                           ALU_RES_MEM_8_port, ALU_RES_OUT(7) => 
                           ALU_RES_MEM_7_port, ALU_RES_OUT(6) => 
                           ALU_RES_MEM_6_port, ALU_RES_OUT(5) => 
                           ALU_RES_MEM_5_port, ALU_RES_OUT(4) => 
                           ALU_RES_MEM_4_port, ALU_RES_OUT(3) => 
                           ALU_RES_MEM_3_port, ALU_RES_OUT(2) => 
                           ALU_RES_MEM_2_port, ALU_RES_OUT(1) => 
                           ALU_RES_MEM_1_port, ALU_RES_OUT(0) => 
                           ALU_RES_MEM_0_port, OP_MEM(31) => OP_MEM_31_port, 
                           OP_MEM(30) => OP_MEM_30_port, OP_MEM(29) => 
                           OP_MEM_29_port, OP_MEM(28) => OP_MEM_28_port, 
                           OP_MEM(27) => OP_MEM_27_port, OP_MEM(26) => 
                           OP_MEM_26_port, OP_MEM(25) => OP_MEM_25_port, 
                           OP_MEM(24) => OP_MEM_24_port, OP_MEM(23) => 
                           OP_MEM_23_port, OP_MEM(22) => OP_MEM_22_port, 
                           OP_MEM(21) => OP_MEM_21_port, OP_MEM(20) => 
                           OP_MEM_20_port, OP_MEM(19) => OP_MEM_19_port, 
                           OP_MEM(18) => OP_MEM_18_port, OP_MEM(17) => 
                           OP_MEM_17_port, OP_MEM(16) => OP_MEM_16_port, 
                           OP_MEM(15) => OP_MEM_15_port, OP_MEM(14) => 
                           OP_MEM_14_port, OP_MEM(13) => OP_MEM_13_port, 
                           OP_MEM(12) => OP_MEM_12_port, OP_MEM(11) => 
                           OP_MEM_11_port, OP_MEM(10) => OP_MEM_10_port, 
                           OP_MEM(9) => OP_MEM_9_port, OP_MEM(8) => 
                           OP_MEM_8_port, OP_MEM(7) => OP_MEM_7_port, OP_MEM(6)
                           => OP_MEM_6_port, OP_MEM(5) => OP_MEM_5_port, 
                           OP_MEM(4) => OP_MEM_4_port, OP_MEM(3) => 
                           OP_MEM_3_port, OP_MEM(2) => OP_MEM_2_port, OP_MEM(1)
                           => OP_MEM_1_port, OP_MEM(0) => OP_MEM_0_port, 
                           ADD_WR_MEM(4) => ADD_WR_MEM_4_port, ADD_WR_MEM(3) =>
                           ADD_WR_MEM_3_port, ADD_WR_MEM(2) => 
                           ADD_WR_MEM_2_port, ADD_WR_MEM(1) => 
                           ADD_WR_MEM_1_port, ADD_WR_MEM(0) => 
                           ADD_WR_MEM_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_MEM_OUT_4_port, ADD_WR_OUT(3) => 
                           ADD_WR_MEM_OUT_3_port, ADD_WR_OUT(2) => 
                           ADD_WR_MEM_OUT_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_MEM_OUT_1_port, ADD_WR_OUT(0) => 
                           ADD_WR_MEM_OUT_0_port, LOAD_TYPE_OUT(1) => 
                           LOAD_TYPE_OUT(1), LOAD_TYPE_OUT(0) => 
                           LOAD_TYPE_OUT(0), STORE_TYPE_OUT => STORE_TYPE_OUT);
   RF_WE_ff : ff_2 port map( D => RF_WE, CLK => CLK, EN => X_Logic1_port, RST 
                           => RST, Q => RF_WE_WB);
   WritebackStage : Writeback port map( WB_MUX_SEL => WB_MUX_SEL, DATA_IN(31) 
                           => DATA_MEM_OUT_31_port, DATA_IN(30) => 
                           DATA_MEM_OUT_30_port, DATA_IN(29) => 
                           DATA_MEM_OUT_29_port, DATA_IN(28) => 
                           DATA_MEM_OUT_28_port, DATA_IN(27) => 
                           DATA_MEM_OUT_27_port, DATA_IN(26) => 
                           DATA_MEM_OUT_26_port, DATA_IN(25) => 
                           DATA_MEM_OUT_25_port, DATA_IN(24) => 
                           DATA_MEM_OUT_24_port, DATA_IN(23) => 
                           DATA_MEM_OUT_23_port, DATA_IN(22) => 
                           DATA_MEM_OUT_22_port, DATA_IN(21) => 
                           DATA_MEM_OUT_21_port, DATA_IN(20) => 
                           DATA_MEM_OUT_20_port, DATA_IN(19) => 
                           DATA_MEM_OUT_19_port, DATA_IN(18) => 
                           DATA_MEM_OUT_18_port, DATA_IN(17) => 
                           DATA_MEM_OUT_17_port, DATA_IN(16) => 
                           DATA_MEM_OUT_16_port, DATA_IN(15) => 
                           DATA_MEM_OUT_15_port, DATA_IN(14) => 
                           DATA_MEM_OUT_14_port, DATA_IN(13) => 
                           DATA_MEM_OUT_13_port, DATA_IN(12) => 
                           DATA_MEM_OUT_12_port, DATA_IN(11) => 
                           DATA_MEM_OUT_11_port, DATA_IN(10) => 
                           DATA_MEM_OUT_10_port, DATA_IN(9) => 
                           DATA_MEM_OUT_9_port, DATA_IN(8) => 
                           DATA_MEM_OUT_8_port, DATA_IN(7) => 
                           DATA_MEM_OUT_7_port, DATA_IN(6) => 
                           DATA_MEM_OUT_6_port, DATA_IN(5) => 
                           DATA_MEM_OUT_5_port, DATA_IN(4) => 
                           DATA_MEM_OUT_4_port, DATA_IN(3) => 
                           DATA_MEM_OUT_3_port, DATA_IN(2) => 
                           DATA_MEM_OUT_2_port, DATA_IN(1) => 
                           DATA_MEM_OUT_1_port, DATA_IN(0) => 
                           DATA_MEM_OUT_0_port, ALU_RES_IN(31) => 
                           ALU_RES_MEM_31_port, ALU_RES_IN(30) => 
                           ALU_RES_MEM_30_port, ALU_RES_IN(29) => 
                           ALU_RES_MEM_29_port, ALU_RES_IN(28) => 
                           ALU_RES_MEM_28_port, ALU_RES_IN(27) => 
                           ALU_RES_MEM_27_port, ALU_RES_IN(26) => 
                           ALU_RES_MEM_26_port, ALU_RES_IN(25) => 
                           ALU_RES_MEM_25_port, ALU_RES_IN(24) => 
                           ALU_RES_MEM_24_port, ALU_RES_IN(23) => 
                           ALU_RES_MEM_23_port, ALU_RES_IN(22) => 
                           ALU_RES_MEM_22_port, ALU_RES_IN(21) => 
                           ALU_RES_MEM_21_port, ALU_RES_IN(20) => 
                           ALU_RES_MEM_20_port, ALU_RES_IN(19) => 
                           ALU_RES_MEM_19_port, ALU_RES_IN(18) => 
                           ALU_RES_MEM_18_port, ALU_RES_IN(17) => 
                           ALU_RES_MEM_17_port, ALU_RES_IN(16) => 
                           ALU_RES_MEM_16_port, ALU_RES_IN(15) => 
                           ALU_RES_MEM_15_port, ALU_RES_IN(14) => 
                           ALU_RES_MEM_14_port, ALU_RES_IN(13) => 
                           ALU_RES_MEM_13_port, ALU_RES_IN(12) => 
                           ALU_RES_MEM_12_port, ALU_RES_IN(11) => 
                           ALU_RES_MEM_11_port, ALU_RES_IN(10) => 
                           ALU_RES_MEM_10_port, ALU_RES_IN(9) => 
                           ALU_RES_MEM_9_port, ALU_RES_IN(8) => 
                           ALU_RES_MEM_8_port, ALU_RES_IN(7) => 
                           ALU_RES_MEM_7_port, ALU_RES_IN(6) => 
                           ALU_RES_MEM_6_port, ALU_RES_IN(5) => 
                           ALU_RES_MEM_5_port, ALU_RES_IN(4) => 
                           ALU_RES_MEM_4_port, ALU_RES_IN(3) => 
                           ALU_RES_MEM_3_port, ALU_RES_IN(2) => 
                           ALU_RES_MEM_2_port, ALU_RES_IN(1) => 
                           ALU_RES_MEM_1_port, ALU_RES_IN(0) => 
                           ALU_RES_MEM_0_port, ADD_WR_IN(4) => 
                           ADD_WR_MEM_OUT_4_port, ADD_WR_IN(3) => 
                           ADD_WR_MEM_OUT_3_port, ADD_WR_IN(2) => 
                           ADD_WR_MEM_OUT_2_port, ADD_WR_IN(1) => 
                           ADD_WR_MEM_OUT_1_port, ADD_WR_IN(0) => 
                           ADD_WR_MEM_OUT_0_port, DATA_OUT(31) => OP_WB_31_port
                           , DATA_OUT(30) => OP_WB_30_port, DATA_OUT(29) => 
                           OP_WB_29_port, DATA_OUT(28) => OP_WB_28_port, 
                           DATA_OUT(27) => OP_WB_27_port, DATA_OUT(26) => 
                           OP_WB_26_port, DATA_OUT(25) => OP_WB_25_port, 
                           DATA_OUT(24) => OP_WB_24_port, DATA_OUT(23) => 
                           OP_WB_23_port, DATA_OUT(22) => OP_WB_22_port, 
                           DATA_OUT(21) => OP_WB_21_port, DATA_OUT(20) => 
                           OP_WB_20_port, DATA_OUT(19) => OP_WB_19_port, 
                           DATA_OUT(18) => OP_WB_18_port, DATA_OUT(17) => 
                           OP_WB_17_port, DATA_OUT(16) => OP_WB_16_port, 
                           DATA_OUT(15) => OP_WB_15_port, DATA_OUT(14) => 
                           OP_WB_14_port, DATA_OUT(13) => OP_WB_13_port, 
                           DATA_OUT(12) => OP_WB_12_port, DATA_OUT(11) => 
                           OP_WB_11_port, DATA_OUT(10) => OP_WB_10_port, 
                           DATA_OUT(9) => OP_WB_9_port, DATA_OUT(8) => 
                           OP_WB_8_port, DATA_OUT(7) => OP_WB_7_port, 
                           DATA_OUT(6) => OP_WB_6_port, DATA_OUT(5) => 
                           OP_WB_5_port, DATA_OUT(4) => OP_WB_4_port, 
                           DATA_OUT(3) => OP_WB_3_port, DATA_OUT(2) => 
                           OP_WB_2_port, DATA_OUT(1) => OP_WB_1_port, 
                           DATA_OUT(0) => OP_WB_0_port, ADD_WR_OUT(4) => 
                           ADD_WR_WB_4_port, ADD_WR_OUT(3) => ADD_WR_WB_3_port,
                           ADD_WR_OUT(2) => ADD_WR_WB_2_port, ADD_WR_OUT(1) => 
                           ADD_WR_WB_1_port, ADD_WR_OUT(0) => ADD_WR_WB_0_port)
                           ;
   HDU : HazardDetection port map( RST => RST, ADD_RS1(4) => ADD_RS1_HDU_4_port
                           , ADD_RS1(3) => ADD_RS1_HDU_3_port, ADD_RS1(2) => 
                           ADD_RS1_HDU_2_port, ADD_RS1(1) => ADD_RS1_HDU_1_port
                           , ADD_RS1(0) => ADD_RS1_HDU_0_port, ADD_RS2(4) => 
                           ADD_RS2_HDU_4_port, ADD_RS2(3) => ADD_RS2_HDU_3_port
                           , ADD_RS2(2) => ADD_RS2_HDU_2_port, ADD_RS2(1) => 
                           ADD_RS2_HDU_1_port, ADD_RS2(0) => ADD_RS2_HDU_0_port
                           , ADD_WR(4) => ADD_WR_DECODE_OUT_4_port, ADD_WR(3) 
                           => ADD_WR_DECODE_OUT_3_port, ADD_WR(2) => 
                           ADD_WR_DECODE_OUT_2_port, ADD_WR(1) => 
                           ADD_WR_DECODE_OUT_1_port, ADD_WR(0) => 
                           ADD_WR_DECODE_OUT_0_port, DRAM_R => DRAM_R_IN, 
                           INS_IN(31) => INS_OUT_31_port, INS_IN(30) => 
                           INS_OUT_30_port, INS_IN(29) => INS_OUT_29_port, 
                           INS_IN(28) => INS_OUT_28_port, INS_IN(27) => 
                           INS_OUT_27_port, INS_IN(26) => INS_OUT_26_port, 
                           INS_IN(25) => INS_OUT_25_port, INS_IN(24) => 
                           INS_OUT_24_port, INS_IN(23) => INS_OUT_23_port, 
                           INS_IN(22) => INS_OUT_22_port, INS_IN(21) => 
                           INS_OUT_21_port, INS_IN(20) => INS_OUT_20_port, 
                           INS_IN(19) => INS_OUT_19_port, INS_IN(18) => 
                           INS_OUT_18_port, INS_IN(17) => INS_OUT_17_port, 
                           INS_IN(16) => INS_OUT_16_port, INS_IN(15) => 
                           INS_OUT_15_port, INS_IN(14) => INS_OUT_14_port, 
                           INS_IN(13) => INS_OUT_13_port, INS_IN(12) => 
                           INS_OUT_12_port, INS_IN(11) => INS_OUT_11_port, 
                           INS_IN(10) => INS_OUT_10_port, INS_IN(9) => 
                           INS_OUT_9_port, INS_IN(8) => INS_OUT_8_port, 
                           INS_IN(7) => INS_OUT_7_port, INS_IN(6) => 
                           INS_OUT_6_port, INS_IN(5) => INS_OUT_5_port, 
                           INS_IN(4) => INS_OUT_4_port, INS_IN(3) => 
                           INS_OUT_3_port, INS_IN(2) => INS_OUT_2_port, 
                           INS_IN(1) => INS_OUT_1_port, INS_IN(0) => 
                           INS_OUT_0_port, PC_IN(31) => PC_FETCH_OUT_31_port, 
                           PC_IN(30) => PC_FETCH_OUT_30_port, PC_IN(29) => 
                           PC_FETCH_OUT_29_port, PC_IN(28) => 
                           PC_FETCH_OUT_28_port, PC_IN(27) => 
                           PC_FETCH_OUT_27_port, PC_IN(26) => 
                           PC_FETCH_OUT_26_port, PC_IN(25) => 
                           PC_FETCH_OUT_25_port, PC_IN(24) => 
                           PC_FETCH_OUT_24_port, PC_IN(23) => 
                           PC_FETCH_OUT_23_port, PC_IN(22) => 
                           PC_FETCH_OUT_22_port, PC_IN(21) => 
                           PC_FETCH_OUT_21_port, PC_IN(20) => 
                           PC_FETCH_OUT_20_port, PC_IN(19) => 
                           PC_FETCH_OUT_19_port, PC_IN(18) => 
                           PC_FETCH_OUT_18_port, PC_IN(17) => 
                           PC_FETCH_OUT_17_port, PC_IN(16) => 
                           PC_FETCH_OUT_16_port, PC_IN(15) => 
                           PC_FETCH_OUT_15_port, PC_IN(14) => 
                           PC_FETCH_OUT_14_port, PC_IN(13) => 
                           PC_FETCH_OUT_13_port, PC_IN(12) => 
                           PC_FETCH_OUT_12_port, PC_IN(11) => 
                           PC_FETCH_OUT_11_port, PC_IN(10) => 
                           PC_FETCH_OUT_10_port, PC_IN(9) => 
                           PC_FETCH_OUT_9_port, PC_IN(8) => PC_FETCH_OUT_8_port
                           , PC_IN(7) => PC_FETCH_OUT_7_port, PC_IN(6) => 
                           PC_FETCH_OUT_6_port, PC_IN(5) => PC_FETCH_OUT_5_port
                           , PC_IN(4) => PC_FETCH_OUT_4_port, PC_IN(3) => 
                           PC_FETCH_OUT_3_port, PC_IN(2) => PC_FETCH_OUT_2_port
                           , PC_IN(1) => PC_FETCH_OUT_1_port, PC_IN(0) => 
                           PC_FETCH_OUT_0_port, Bubble => n14, HDU_INS_OUT(31) 
                           => sig_HDU_INS_OUT_31_port, HDU_INS_OUT(30) => 
                           sig_HDU_INS_OUT_30_port, HDU_INS_OUT(29) => 
                           sig_HDU_INS_OUT_29_port, HDU_INS_OUT(28) => 
                           sig_HDU_INS_OUT_28_port, HDU_INS_OUT(27) => 
                           sig_HDU_INS_OUT_27_port, HDU_INS_OUT(26) => 
                           sig_HDU_INS_OUT_26_port, HDU_INS_OUT(25) => 
                           sig_HDU_INS_OUT_25_port, HDU_INS_OUT(24) => 
                           sig_HDU_INS_OUT_24_port, HDU_INS_OUT(23) => 
                           sig_HDU_INS_OUT_23_port, HDU_INS_OUT(22) => 
                           sig_HDU_INS_OUT_22_port, HDU_INS_OUT(21) => 
                           sig_HDU_INS_OUT_21_port, HDU_INS_OUT(20) => 
                           sig_HDU_INS_OUT_20_port, HDU_INS_OUT(19) => 
                           sig_HDU_INS_OUT_19_port, HDU_INS_OUT(18) => 
                           sig_HDU_INS_OUT_18_port, HDU_INS_OUT(17) => 
                           sig_HDU_INS_OUT_17_port, HDU_INS_OUT(16) => 
                           sig_HDU_INS_OUT_16_port, HDU_INS_OUT(15) => 
                           sig_HDU_INS_OUT_15_port, HDU_INS_OUT(14) => 
                           sig_HDU_INS_OUT_14_port, HDU_INS_OUT(13) => 
                           sig_HDU_INS_OUT_13_port, HDU_INS_OUT(12) => 
                           sig_HDU_INS_OUT_12_port, HDU_INS_OUT(11) => 
                           sig_HDU_INS_OUT_11_port, HDU_INS_OUT(10) => 
                           sig_HDU_INS_OUT_10_port, HDU_INS_OUT(9) => 
                           sig_HDU_INS_OUT_9_port, HDU_INS_OUT(8) => 
                           sig_HDU_INS_OUT_8_port, HDU_INS_OUT(7) => 
                           sig_HDU_INS_OUT_7_port, HDU_INS_OUT(6) => 
                           sig_HDU_INS_OUT_6_port, HDU_INS_OUT(5) => 
                           sig_HDU_INS_OUT_5_port, HDU_INS_OUT(4) => 
                           sig_HDU_INS_OUT_4_port, HDU_INS_OUT(3) => 
                           sig_HDU_INS_OUT_3_port, HDU_INS_OUT(2) => 
                           sig_HDU_INS_OUT_2_port, HDU_INS_OUT(1) => 
                           sig_HDU_INS_OUT_1_port, HDU_INS_OUT(0) => 
                           sig_HDU_INS_OUT_0_port, HDU_PC_OUT(31) => 
                           sig_HDU_PC_OUT_31_port, HDU_PC_OUT(30) => 
                           sig_HDU_PC_OUT_30_port, HDU_PC_OUT(29) => 
                           sig_HDU_PC_OUT_29_port, HDU_PC_OUT(28) => 
                           sig_HDU_PC_OUT_28_port, HDU_PC_OUT(27) => 
                           sig_HDU_PC_OUT_27_port, HDU_PC_OUT(26) => 
                           sig_HDU_PC_OUT_26_port, HDU_PC_OUT(25) => 
                           sig_HDU_PC_OUT_25_port, HDU_PC_OUT(24) => 
                           sig_HDU_PC_OUT_24_port, HDU_PC_OUT(23) => 
                           sig_HDU_PC_OUT_23_port, HDU_PC_OUT(22) => 
                           sig_HDU_PC_OUT_22_port, HDU_PC_OUT(21) => 
                           sig_HDU_PC_OUT_21_port, HDU_PC_OUT(20) => 
                           sig_HDU_PC_OUT_20_port, HDU_PC_OUT(19) => 
                           sig_HDU_PC_OUT_19_port, HDU_PC_OUT(18) => 
                           sig_HDU_PC_OUT_18_port, HDU_PC_OUT(17) => 
                           sig_HDU_PC_OUT_17_port, HDU_PC_OUT(16) => 
                           sig_HDU_PC_OUT_16_port, HDU_PC_OUT(15) => 
                           sig_HDU_PC_OUT_15_port, HDU_PC_OUT(14) => 
                           sig_HDU_PC_OUT_14_port, HDU_PC_OUT(13) => 
                           sig_HDU_PC_OUT_13_port, HDU_PC_OUT(12) => 
                           sig_HDU_PC_OUT_12_port, HDU_PC_OUT(11) => 
                           sig_HDU_PC_OUT_11_port, HDU_PC_OUT(10) => 
                           sig_HDU_PC_OUT_10_port, HDU_PC_OUT(9) => 
                           sig_HDU_PC_OUT_9_port, HDU_PC_OUT(8) => 
                           sig_HDU_PC_OUT_8_port, HDU_PC_OUT(7) => 
                           sig_HDU_PC_OUT_7_port, HDU_PC_OUT(6) => 
                           sig_HDU_PC_OUT_6_port, HDU_PC_OUT(5) => 
                           sig_HDU_PC_OUT_5_port, HDU_PC_OUT(4) => 
                           sig_HDU_PC_OUT_4_port, HDU_PC_OUT(3) => 
                           sig_HDU_PC_OUT_3_port, HDU_PC_OUT(2) => 
                           sig_HDU_PC_OUT_2_port, HDU_PC_OUT(1) => 
                           sig_HDU_PC_OUT_1_port, HDU_PC_OUT(0) => 
                           sig_HDU_PC_OUT_0_port, HDU_NPC_OUT(31) => 
                           sig_HDU_NPC_OUT_31_port, HDU_NPC_OUT(30) => 
                           sig_HDU_NPC_OUT_30_port, HDU_NPC_OUT(29) => 
                           sig_HDU_NPC_OUT_29_port, HDU_NPC_OUT(28) => 
                           sig_HDU_NPC_OUT_28_port, HDU_NPC_OUT(27) => 
                           sig_HDU_NPC_OUT_27_port, HDU_NPC_OUT(26) => 
                           sig_HDU_NPC_OUT_26_port, HDU_NPC_OUT(25) => 
                           sig_HDU_NPC_OUT_25_port, HDU_NPC_OUT(24) => 
                           sig_HDU_NPC_OUT_24_port, HDU_NPC_OUT(23) => 
                           sig_HDU_NPC_OUT_23_port, HDU_NPC_OUT(22) => 
                           sig_HDU_NPC_OUT_22_port, HDU_NPC_OUT(21) => 
                           sig_HDU_NPC_OUT_21_port, HDU_NPC_OUT(20) => 
                           sig_HDU_NPC_OUT_20_port, HDU_NPC_OUT(19) => 
                           sig_HDU_NPC_OUT_19_port, HDU_NPC_OUT(18) => 
                           sig_HDU_NPC_OUT_18_port, HDU_NPC_OUT(17) => 
                           sig_HDU_NPC_OUT_17_port, HDU_NPC_OUT(16) => 
                           sig_HDU_NPC_OUT_16_port, HDU_NPC_OUT(15) => 
                           sig_HDU_NPC_OUT_15_port, HDU_NPC_OUT(14) => 
                           sig_HDU_NPC_OUT_14_port, HDU_NPC_OUT(13) => 
                           sig_HDU_NPC_OUT_13_port, HDU_NPC_OUT(12) => 
                           sig_HDU_NPC_OUT_12_port, HDU_NPC_OUT(11) => 
                           sig_HDU_NPC_OUT_11_port, HDU_NPC_OUT(10) => 
                           sig_HDU_NPC_OUT_10_port, HDU_NPC_OUT(9) => 
                           sig_HDU_NPC_OUT_9_port, HDU_NPC_OUT(8) => 
                           sig_HDU_NPC_OUT_8_port, HDU_NPC_OUT(7) => 
                           sig_HDU_NPC_OUT_7_port, HDU_NPC_OUT(6) => 
                           sig_HDU_NPC_OUT_6_port, HDU_NPC_OUT(5) => 
                           sig_HDU_NPC_OUT_5_port, HDU_NPC_OUT(4) => 
                           sig_HDU_NPC_OUT_4_port, HDU_NPC_OUT(3) => 
                           sig_HDU_NPC_OUT_3_port, HDU_NPC_OUT(2) => 
                           sig_HDU_NPC_OUT_2_port, HDU_NPC_OUT(1) => 
                           sig_HDU_NPC_OUT_1_port, HDU_NPC_OUT(0) => 
                           sig_HDU_NPC_OUT_0_port);
   U2 : BUF_X1 port map( A => n14, Z => Bubble_out_port);
   U3 : CLKBUF_X1 port map( A => n10, Z => INS_OUT_29_port);
   U4 : CLKBUF_X1 port map( A => n12, Z => INS_OUT_27_port);
   U5 : CLKBUF_X1 port map( A => n13, Z => INS_OUT_26_port);
   U6 : CLKBUF_X1 port map( A => n9, Z => INS_OUT_30_port);
   U7 : CLKBUF_X1 port map( A => n11, Z => INS_OUT_28_port);
   U8 : CLKBUF_X1 port map( A => n8, Z => INS_OUT_31_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( Clk, Rst : in std_logic);

end DLX;

architecture SYN_dlx_rtl of DLX is

   component DRAM
      port( Clk, Rst : in std_logic;  ADDR_IN, DATA_IN : in std_logic_vector 
            (31 downto 0);  LOAD_TYPE : in std_logic_vector (1 downto 0);  
            STORE_TYPE, DRAM_W, DRAM_R : in std_logic;  DATA_OUT : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component IRAM
      port( Rst : in std_logic;  Addr : in std_logic_vector (31 downto 0);  
            Iout : out std_logic_vector (31 downto 0));
   end component;
   
   component hardwired_cu_NBIT32
      port( MUX_A_SEL : out std_logic;  MUX_B_SEL : out std_logic_vector (1 
            downto 0);  ALU_OPC : out std_logic_vector (0 to 4);  ALU_OUTREG_EN
            , DRAM_R_IN : out std_logic;  JUMP_TYPE : out std_logic_vector (1 
            downto 0);  MEM_EN_IN, DRAM_W_IN, RF_WE : out std_logic;  
            LOAD_TYPE_IN : out std_logic_vector (1 downto 0);  STORE_TYPE_IN, 
            WB_MUX_SEL : out std_logic;  INS_IN : in std_logic_vector (31 
            downto 0);  Bubble, Clk, Rst : in std_logic);
   end component;
   
   component Datapath
      port( CLK, RST : in std_logic;  INS_IN, DATA_IN : in std_logic_vector (31
            downto 0);  MUX_A_SEL : in std_logic;  MUX_B_SEL : in 
            std_logic_vector (1 downto 0);  ALU_OPC : in std_logic_vector (0 to
            4);  ALU_OUTREG_EN : in std_logic;  JUMP_TYPE : in std_logic_vector
            (1 downto 0);  DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, RF_WE : in 
            std_logic;  LOAD_TYPE_IN : in std_logic_vector (1 downto 0);  
            STORE_TYPE_IN, WB_MUX_SEL : in std_logic;  INS_OUT, IRAM_ADDR_OUT, 
            DRAM_ADDR_OUT, DATA_OUT : out std_logic_vector (31 downto 0);  
            DRAM_R_OUT, DRAM_W_OUT, Bubble_out : out std_logic;  LOAD_TYPE_OUT 
            : out std_logic_vector (1 downto 0);  STORE_TYPE_OUT : out 
            std_logic);
   end component;
   
   signal INS_IN_31_port, INS_IN_30_port, INS_IN_29_port, INS_IN_28_port, 
      INS_IN_27_port, INS_IN_26_port, INS_IN_25_port, INS_IN_24_port, 
      INS_IN_23_port, INS_IN_22_port, INS_IN_21_port, INS_IN_20_port, 
      INS_IN_19_port, INS_IN_18_port, INS_IN_17_port, INS_IN_16_port, 
      INS_IN_15_port, INS_IN_14_port, INS_IN_13_port, INS_IN_12_port, 
      INS_IN_11_port, INS_IN_10_port, INS_IN_9_port, INS_IN_8_port, 
      INS_IN_7_port, INS_IN_6_port, INS_IN_5_port, INS_IN_4_port, INS_IN_3_port
      , INS_IN_2_port, INS_IN_1_port, INS_IN_0_port, DATA_IN_31_port, 
      DATA_IN_30_port, DATA_IN_29_port, DATA_IN_28_port, DATA_IN_27_port, 
      DATA_IN_26_port, DATA_IN_25_port, DATA_IN_24_port, DATA_IN_23_port, 
      DATA_IN_22_port, DATA_IN_21_port, DATA_IN_20_port, DATA_IN_19_port, 
      DATA_IN_18_port, DATA_IN_17_port, DATA_IN_16_port, DATA_IN_15_port, 
      DATA_IN_14_port, DATA_IN_13_port, DATA_IN_12_port, DATA_IN_11_port, 
      DATA_IN_10_port, DATA_IN_9_port, DATA_IN_8_port, DATA_IN_7_port, 
      DATA_IN_6_port, DATA_IN_5_port, DATA_IN_4_port, DATA_IN_3_port, 
      DATA_IN_2_port, DATA_IN_1_port, DATA_IN_0_port, MUX_A_SEL, 
      MUX_B_SEL_1_port, MUX_B_SEL_0_port, ALU_OPC_4_port, ALU_OPC_3_port, 
      ALU_OPC_2_port, ALU_OPC_1_port, ALU_OPC_0_port, ALU_OUTREG_EN, 
      JUMP_TYPE_1_port, JUMP_TYPE_0_port, DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, 
      RF_WE, LOAD_TYPE_IN_1_port, LOAD_TYPE_IN_0_port, STORE_TYPE_IN, 
      WB_MUX_SEL, INST_31_port, INST_30_port, INST_29_port, INST_28_port, 
      INST_27_port, INST_26_port, INST_25_port, INST_24_port, INST_23_port, 
      INST_22_port, INST_21_port, INST_20_port, INST_19_port, INST_18_port, 
      INST_17_port, INST_16_port, INST_15_port, INST_14_port, INST_13_port, 
      INST_12_port, INST_11_port, INST_10_port, INST_9_port, INST_8_port, 
      INST_7_port, INST_6_port, INST_5_port, INST_4_port, INST_3_port, 
      INST_2_port, INST_1_port, INST_0_port, IRAM_ADDR_OUT_31_port, 
      IRAM_ADDR_OUT_30_port, IRAM_ADDR_OUT_29_port, IRAM_ADDR_OUT_28_port, 
      IRAM_ADDR_OUT_27_port, IRAM_ADDR_OUT_26_port, IRAM_ADDR_OUT_25_port, 
      IRAM_ADDR_OUT_24_port, IRAM_ADDR_OUT_23_port, IRAM_ADDR_OUT_22_port, 
      IRAM_ADDR_OUT_21_port, IRAM_ADDR_OUT_20_port, IRAM_ADDR_OUT_19_port, 
      IRAM_ADDR_OUT_18_port, IRAM_ADDR_OUT_17_port, IRAM_ADDR_OUT_16_port, 
      IRAM_ADDR_OUT_15_port, IRAM_ADDR_OUT_14_port, IRAM_ADDR_OUT_13_port, 
      IRAM_ADDR_OUT_12_port, IRAM_ADDR_OUT_11_port, IRAM_ADDR_OUT_10_port, 
      IRAM_ADDR_OUT_9_port, IRAM_ADDR_OUT_8_port, IRAM_ADDR_OUT_7_port, 
      IRAM_ADDR_OUT_6_port, IRAM_ADDR_OUT_5_port, IRAM_ADDR_OUT_4_port, 
      IRAM_ADDR_OUT_3_port, IRAM_ADDR_OUT_2_port, IRAM_ADDR_OUT_1_port, 
      IRAM_ADDR_OUT_0_port, DRAM_ADDR_OUT_31_port, DRAM_ADDR_OUT_30_port, 
      DRAM_ADDR_OUT_29_port, DRAM_ADDR_OUT_28_port, DRAM_ADDR_OUT_27_port, 
      DRAM_ADDR_OUT_26_port, DRAM_ADDR_OUT_25_port, DRAM_ADDR_OUT_24_port, 
      DRAM_ADDR_OUT_23_port, DRAM_ADDR_OUT_22_port, DRAM_ADDR_OUT_21_port, 
      DRAM_ADDR_OUT_20_port, DRAM_ADDR_OUT_19_port, DRAM_ADDR_OUT_18_port, 
      DRAM_ADDR_OUT_17_port, DRAM_ADDR_OUT_16_port, DRAM_ADDR_OUT_15_port, 
      DRAM_ADDR_OUT_14_port, DRAM_ADDR_OUT_13_port, DRAM_ADDR_OUT_12_port, 
      DRAM_ADDR_OUT_11_port, DRAM_ADDR_OUT_10_port, DRAM_ADDR_OUT_9_port, 
      DRAM_ADDR_OUT_8_port, DRAM_ADDR_OUT_7_port, DRAM_ADDR_OUT_6_port, 
      DRAM_ADDR_OUT_5_port, DRAM_ADDR_OUT_4_port, DRAM_ADDR_OUT_3_port, 
      DRAM_ADDR_OUT_2_port, DRAM_ADDR_OUT_1_port, DRAM_ADDR_OUT_0_port, 
      DATA_OUT_31_port, DATA_OUT_30_port, DATA_OUT_29_port, DATA_OUT_28_port, 
      DATA_OUT_27_port, DATA_OUT_26_port, DATA_OUT_25_port, DATA_OUT_24_port, 
      DATA_OUT_23_port, DATA_OUT_22_port, DATA_OUT_21_port, DATA_OUT_20_port, 
      DATA_OUT_19_port, DATA_OUT_18_port, DATA_OUT_17_port, DATA_OUT_16_port, 
      DATA_OUT_15_port, DATA_OUT_14_port, DATA_OUT_13_port, DATA_OUT_12_port, 
      DATA_OUT_11_port, DATA_OUT_10_port, DATA_OUT_9_port, DATA_OUT_8_port, 
      DATA_OUT_7_port, DATA_OUT_6_port, DATA_OUT_5_port, DATA_OUT_4_port, 
      DATA_OUT_3_port, DATA_OUT_2_port, DATA_OUT_1_port, DATA_OUT_0_port, 
      DRAM_R_OUT, DRAM_W_OUT, Bubble, LOAD_TYPE_OUT_1_port, 
      LOAD_TYPE_OUT_0_port, STORE_TYPE_OUT, n_1991, n_1992, n_1993, n_1994, 
      n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, 
      n_2004 : std_logic;

begin
   
   DP : Datapath port map( CLK => Clk, RST => Rst, INS_IN(31) => INS_IN_31_port
                           , INS_IN(30) => INS_IN_30_port, INS_IN(29) => 
                           INS_IN_29_port, INS_IN(28) => INS_IN_28_port, 
                           INS_IN(27) => INS_IN_27_port, INS_IN(26) => 
                           INS_IN_26_port, INS_IN(25) => INS_IN_25_port, 
                           INS_IN(24) => INS_IN_24_port, INS_IN(23) => 
                           INS_IN_23_port, INS_IN(22) => INS_IN_22_port, 
                           INS_IN(21) => INS_IN_21_port, INS_IN(20) => 
                           INS_IN_20_port, INS_IN(19) => INS_IN_19_port, 
                           INS_IN(18) => INS_IN_18_port, INS_IN(17) => 
                           INS_IN_17_port, INS_IN(16) => INS_IN_16_port, 
                           INS_IN(15) => INS_IN_15_port, INS_IN(14) => 
                           INS_IN_14_port, INS_IN(13) => INS_IN_13_port, 
                           INS_IN(12) => INS_IN_12_port, INS_IN(11) => 
                           INS_IN_11_port, INS_IN(10) => INS_IN_10_port, 
                           INS_IN(9) => INS_IN_9_port, INS_IN(8) => 
                           INS_IN_8_port, INS_IN(7) => INS_IN_7_port, INS_IN(6)
                           => INS_IN_6_port, INS_IN(5) => INS_IN_5_port, 
                           INS_IN(4) => INS_IN_4_port, INS_IN(3) => 
                           INS_IN_3_port, INS_IN(2) => INS_IN_2_port, INS_IN(1)
                           => INS_IN_1_port, INS_IN(0) => INS_IN_0_port, 
                           DATA_IN(31) => DATA_IN_31_port, DATA_IN(30) => 
                           DATA_IN_30_port, DATA_IN(29) => DATA_IN_29_port, 
                           DATA_IN(28) => DATA_IN_28_port, DATA_IN(27) => 
                           DATA_IN_27_port, DATA_IN(26) => DATA_IN_26_port, 
                           DATA_IN(25) => DATA_IN_25_port, DATA_IN(24) => 
                           DATA_IN_24_port, DATA_IN(23) => DATA_IN_23_port, 
                           DATA_IN(22) => DATA_IN_22_port, DATA_IN(21) => 
                           DATA_IN_21_port, DATA_IN(20) => DATA_IN_20_port, 
                           DATA_IN(19) => DATA_IN_19_port, DATA_IN(18) => 
                           DATA_IN_18_port, DATA_IN(17) => DATA_IN_17_port, 
                           DATA_IN(16) => DATA_IN_16_port, DATA_IN(15) => 
                           DATA_IN_15_port, DATA_IN(14) => DATA_IN_14_port, 
                           DATA_IN(13) => DATA_IN_13_port, DATA_IN(12) => 
                           DATA_IN_12_port, DATA_IN(11) => DATA_IN_11_port, 
                           DATA_IN(10) => DATA_IN_10_port, DATA_IN(9) => 
                           DATA_IN_9_port, DATA_IN(8) => DATA_IN_8_port, 
                           DATA_IN(7) => DATA_IN_7_port, DATA_IN(6) => 
                           DATA_IN_6_port, DATA_IN(5) => DATA_IN_5_port, 
                           DATA_IN(4) => DATA_IN_4_port, DATA_IN(3) => 
                           DATA_IN_3_port, DATA_IN(2) => DATA_IN_2_port, 
                           DATA_IN(1) => DATA_IN_1_port, DATA_IN(0) => 
                           DATA_IN_0_port, MUX_A_SEL => MUX_A_SEL, MUX_B_SEL(1)
                           => MUX_B_SEL_1_port, MUX_B_SEL(0) => 
                           MUX_B_SEL_0_port, ALU_OPC(0) => ALU_OPC_4_port, 
                           ALU_OPC(1) => ALU_OPC_3_port, ALU_OPC(2) => 
                           ALU_OPC_2_port, ALU_OPC(3) => ALU_OPC_1_port, 
                           ALU_OPC(4) => ALU_OPC_0_port, ALU_OUTREG_EN => 
                           ALU_OUTREG_EN, JUMP_TYPE(1) => JUMP_TYPE_1_port, 
                           JUMP_TYPE(0) => JUMP_TYPE_0_port, DRAM_R_IN => 
                           DRAM_R_IN, MEM_EN_IN => MEM_EN_IN, DRAM_W_IN => 
                           DRAM_W_IN, RF_WE => RF_WE, LOAD_TYPE_IN(1) => 
                           LOAD_TYPE_IN_1_port, LOAD_TYPE_IN(0) => 
                           LOAD_TYPE_IN_0_port, STORE_TYPE_IN => STORE_TYPE_IN,
                           WB_MUX_SEL => WB_MUX_SEL, INS_OUT(31) => 
                           INST_31_port, INS_OUT(30) => INST_30_port, 
                           INS_OUT(29) => INST_29_port, INS_OUT(28) => 
                           INST_28_port, INS_OUT(27) => INST_27_port, 
                           INS_OUT(26) => INST_26_port, INS_OUT(25) => 
                           INST_25_port, INS_OUT(24) => INST_24_port, 
                           INS_OUT(23) => INST_23_port, INS_OUT(22) => 
                           INST_22_port, INS_OUT(21) => INST_21_port, 
                           INS_OUT(20) => INST_20_port, INS_OUT(19) => 
                           INST_19_port, INS_OUT(18) => INST_18_port, 
                           INS_OUT(17) => INST_17_port, INS_OUT(16) => 
                           INST_16_port, INS_OUT(15) => INST_15_port, 
                           INS_OUT(14) => INST_14_port, INS_OUT(13) => 
                           INST_13_port, INS_OUT(12) => INST_12_port, 
                           INS_OUT(11) => INST_11_port, INS_OUT(10) => 
                           INST_10_port, INS_OUT(9) => INST_9_port, INS_OUT(8) 
                           => INST_8_port, INS_OUT(7) => INST_7_port, 
                           INS_OUT(6) => INST_6_port, INS_OUT(5) => INST_5_port
                           , INS_OUT(4) => INST_4_port, INS_OUT(3) => 
                           INST_3_port, INS_OUT(2) => INST_2_port, INS_OUT(1) 
                           => INST_1_port, INS_OUT(0) => INST_0_port, 
                           IRAM_ADDR_OUT(31) => IRAM_ADDR_OUT_31_port, 
                           IRAM_ADDR_OUT(30) => IRAM_ADDR_OUT_30_port, 
                           IRAM_ADDR_OUT(29) => IRAM_ADDR_OUT_29_port, 
                           IRAM_ADDR_OUT(28) => IRAM_ADDR_OUT_28_port, 
                           IRAM_ADDR_OUT(27) => IRAM_ADDR_OUT_27_port, 
                           IRAM_ADDR_OUT(26) => IRAM_ADDR_OUT_26_port, 
                           IRAM_ADDR_OUT(25) => IRAM_ADDR_OUT_25_port, 
                           IRAM_ADDR_OUT(24) => IRAM_ADDR_OUT_24_port, 
                           IRAM_ADDR_OUT(23) => IRAM_ADDR_OUT_23_port, 
                           IRAM_ADDR_OUT(22) => IRAM_ADDR_OUT_22_port, 
                           IRAM_ADDR_OUT(21) => IRAM_ADDR_OUT_21_port, 
                           IRAM_ADDR_OUT(20) => IRAM_ADDR_OUT_20_port, 
                           IRAM_ADDR_OUT(19) => IRAM_ADDR_OUT_19_port, 
                           IRAM_ADDR_OUT(18) => IRAM_ADDR_OUT_18_port, 
                           IRAM_ADDR_OUT(17) => IRAM_ADDR_OUT_17_port, 
                           IRAM_ADDR_OUT(16) => IRAM_ADDR_OUT_16_port, 
                           IRAM_ADDR_OUT(15) => IRAM_ADDR_OUT_15_port, 
                           IRAM_ADDR_OUT(14) => IRAM_ADDR_OUT_14_port, 
                           IRAM_ADDR_OUT(13) => IRAM_ADDR_OUT_13_port, 
                           IRAM_ADDR_OUT(12) => IRAM_ADDR_OUT_12_port, 
                           IRAM_ADDR_OUT(11) => IRAM_ADDR_OUT_11_port, 
                           IRAM_ADDR_OUT(10) => IRAM_ADDR_OUT_10_port, 
                           IRAM_ADDR_OUT(9) => IRAM_ADDR_OUT_9_port, 
                           IRAM_ADDR_OUT(8) => IRAM_ADDR_OUT_8_port, 
                           IRAM_ADDR_OUT(7) => IRAM_ADDR_OUT_7_port, 
                           IRAM_ADDR_OUT(6) => IRAM_ADDR_OUT_6_port, 
                           IRAM_ADDR_OUT(5) => IRAM_ADDR_OUT_5_port, 
                           IRAM_ADDR_OUT(4) => IRAM_ADDR_OUT_4_port, 
                           IRAM_ADDR_OUT(3) => IRAM_ADDR_OUT_3_port, 
                           IRAM_ADDR_OUT(2) => IRAM_ADDR_OUT_2_port, 
                           IRAM_ADDR_OUT(1) => IRAM_ADDR_OUT_1_port, 
                           IRAM_ADDR_OUT(0) => IRAM_ADDR_OUT_0_port, 
                           DRAM_ADDR_OUT(31) => DRAM_ADDR_OUT_31_port, 
                           DRAM_ADDR_OUT(30) => DRAM_ADDR_OUT_30_port, 
                           DRAM_ADDR_OUT(29) => DRAM_ADDR_OUT_29_port, 
                           DRAM_ADDR_OUT(28) => DRAM_ADDR_OUT_28_port, 
                           DRAM_ADDR_OUT(27) => DRAM_ADDR_OUT_27_port, 
                           DRAM_ADDR_OUT(26) => DRAM_ADDR_OUT_26_port, 
                           DRAM_ADDR_OUT(25) => DRAM_ADDR_OUT_25_port, 
                           DRAM_ADDR_OUT(24) => DRAM_ADDR_OUT_24_port, 
                           DRAM_ADDR_OUT(23) => DRAM_ADDR_OUT_23_port, 
                           DRAM_ADDR_OUT(22) => DRAM_ADDR_OUT_22_port, 
                           DRAM_ADDR_OUT(21) => DRAM_ADDR_OUT_21_port, 
                           DRAM_ADDR_OUT(20) => DRAM_ADDR_OUT_20_port, 
                           DRAM_ADDR_OUT(19) => DRAM_ADDR_OUT_19_port, 
                           DRAM_ADDR_OUT(18) => DRAM_ADDR_OUT_18_port, 
                           DRAM_ADDR_OUT(17) => DRAM_ADDR_OUT_17_port, 
                           DRAM_ADDR_OUT(16) => DRAM_ADDR_OUT_16_port, 
                           DRAM_ADDR_OUT(15) => DRAM_ADDR_OUT_15_port, 
                           DRAM_ADDR_OUT(14) => DRAM_ADDR_OUT_14_port, 
                           DRAM_ADDR_OUT(13) => DRAM_ADDR_OUT_13_port, 
                           DRAM_ADDR_OUT(12) => DRAM_ADDR_OUT_12_port, 
                           DRAM_ADDR_OUT(11) => DRAM_ADDR_OUT_11_port, 
                           DRAM_ADDR_OUT(10) => DRAM_ADDR_OUT_10_port, 
                           DRAM_ADDR_OUT(9) => DRAM_ADDR_OUT_9_port, 
                           DRAM_ADDR_OUT(8) => DRAM_ADDR_OUT_8_port, 
                           DRAM_ADDR_OUT(7) => DRAM_ADDR_OUT_7_port, 
                           DRAM_ADDR_OUT(6) => DRAM_ADDR_OUT_6_port, 
                           DRAM_ADDR_OUT(5) => DRAM_ADDR_OUT_5_port, 
                           DRAM_ADDR_OUT(4) => DRAM_ADDR_OUT_4_port, 
                           DRAM_ADDR_OUT(3) => DRAM_ADDR_OUT_3_port, 
                           DRAM_ADDR_OUT(2) => DRAM_ADDR_OUT_2_port, 
                           DRAM_ADDR_OUT(1) => DRAM_ADDR_OUT_1_port, 
                           DRAM_ADDR_OUT(0) => DRAM_ADDR_OUT_0_port, 
                           DATA_OUT(31) => DATA_OUT_31_port, DATA_OUT(30) => 
                           DATA_OUT_30_port, DATA_OUT(29) => DATA_OUT_29_port, 
                           DATA_OUT(28) => DATA_OUT_28_port, DATA_OUT(27) => 
                           DATA_OUT_27_port, DATA_OUT(26) => DATA_OUT_26_port, 
                           DATA_OUT(25) => DATA_OUT_25_port, DATA_OUT(24) => 
                           DATA_OUT_24_port, DATA_OUT(23) => DATA_OUT_23_port, 
                           DATA_OUT(22) => DATA_OUT_22_port, DATA_OUT(21) => 
                           DATA_OUT_21_port, DATA_OUT(20) => DATA_OUT_20_port, 
                           DATA_OUT(19) => DATA_OUT_19_port, DATA_OUT(18) => 
                           DATA_OUT_18_port, DATA_OUT(17) => DATA_OUT_17_port, 
                           DATA_OUT(16) => DATA_OUT_16_port, DATA_OUT(15) => 
                           DATA_OUT_15_port, DATA_OUT(14) => DATA_OUT_14_port, 
                           DATA_OUT(13) => DATA_OUT_13_port, DATA_OUT(12) => 
                           DATA_OUT_12_port, DATA_OUT(11) => DATA_OUT_11_port, 
                           DATA_OUT(10) => DATA_OUT_10_port, DATA_OUT(9) => 
                           DATA_OUT_9_port, DATA_OUT(8) => DATA_OUT_8_port, 
                           DATA_OUT(7) => DATA_OUT_7_port, DATA_OUT(6) => 
                           DATA_OUT_6_port, DATA_OUT(5) => DATA_OUT_5_port, 
                           DATA_OUT(4) => DATA_OUT_4_port, DATA_OUT(3) => 
                           DATA_OUT_3_port, DATA_OUT(2) => DATA_OUT_2_port, 
                           DATA_OUT(1) => DATA_OUT_1_port, DATA_OUT(0) => 
                           DATA_OUT_0_port, DRAM_R_OUT => DRAM_R_OUT, 
                           DRAM_W_OUT => DRAM_W_OUT, Bubble_out => Bubble, 
                           LOAD_TYPE_OUT(1) => LOAD_TYPE_OUT_1_port, 
                           LOAD_TYPE_OUT(0) => LOAD_TYPE_OUT_0_port, 
                           STORE_TYPE_OUT => STORE_TYPE_OUT);
   CU : hardwired_cu_NBIT32 port map( MUX_A_SEL => n_1991, MUX_B_SEL(1) => 
                           n_1992, MUX_B_SEL(0) => n_1993, ALU_OPC(0) => 
                           ALU_OPC_4_port, ALU_OPC(1) => ALU_OPC_3_port, 
                           ALU_OPC(2) => ALU_OPC_2_port, ALU_OPC(3) => 
                           ALU_OPC_1_port, ALU_OPC(4) => ALU_OPC_0_port, 
                           ALU_OUTREG_EN => n_1994, DRAM_R_IN => n_1995, 
                           JUMP_TYPE(1) => n_1996, JUMP_TYPE(0) => n_1997, 
                           MEM_EN_IN => n_1998, DRAM_W_IN => n_1999, RF_WE => 
                           n_2000, LOAD_TYPE_IN(1) => n_2001, LOAD_TYPE_IN(0) 
                           => n_2002, STORE_TYPE_IN => n_2003, WB_MUX_SEL => 
                           n_2004, INS_IN(31) => INST_31_port, INS_IN(30) => 
                           INST_30_port, INS_IN(29) => INST_29_port, INS_IN(28)
                           => INST_28_port, INS_IN(27) => INST_27_port, 
                           INS_IN(26) => INST_26_port, INS_IN(25) => 
                           INST_25_port, INS_IN(24) => INST_24_port, INS_IN(23)
                           => INST_23_port, INS_IN(22) => INST_22_port, 
                           INS_IN(21) => INST_21_port, INS_IN(20) => 
                           INST_20_port, INS_IN(19) => INST_19_port, INS_IN(18)
                           => INST_18_port, INS_IN(17) => INST_17_port, 
                           INS_IN(16) => INST_16_port, INS_IN(15) => 
                           INST_15_port, INS_IN(14) => INST_14_port, INS_IN(13)
                           => INST_13_port, INS_IN(12) => INST_12_port, 
                           INS_IN(11) => INST_11_port, INS_IN(10) => 
                           INST_10_port, INS_IN(9) => INST_9_port, INS_IN(8) =>
                           INST_8_port, INS_IN(7) => INST_7_port, INS_IN(6) => 
                           INST_6_port, INS_IN(5) => INST_5_port, INS_IN(4) => 
                           INST_4_port, INS_IN(3) => INST_3_port, INS_IN(2) => 
                           INST_2_port, INS_IN(1) => INST_1_port, INS_IN(0) => 
                           INST_0_port, Bubble => Bubble, Clk => Clk, Rst => 
                           Rst);
   IRAM_I : IRAM port map( Rst => Rst, Addr(31) => IRAM_ADDR_OUT_31_port, 
                           Addr(30) => IRAM_ADDR_OUT_30_port, Addr(29) => 
                           IRAM_ADDR_OUT_29_port, Addr(28) => 
                           IRAM_ADDR_OUT_28_port, Addr(27) => 
                           IRAM_ADDR_OUT_27_port, Addr(26) => 
                           IRAM_ADDR_OUT_26_port, Addr(25) => 
                           IRAM_ADDR_OUT_25_port, Addr(24) => 
                           IRAM_ADDR_OUT_24_port, Addr(23) => 
                           IRAM_ADDR_OUT_23_port, Addr(22) => 
                           IRAM_ADDR_OUT_22_port, Addr(21) => 
                           IRAM_ADDR_OUT_21_port, Addr(20) => 
                           IRAM_ADDR_OUT_20_port, Addr(19) => 
                           IRAM_ADDR_OUT_19_port, Addr(18) => 
                           IRAM_ADDR_OUT_18_port, Addr(17) => 
                           IRAM_ADDR_OUT_17_port, Addr(16) => 
                           IRAM_ADDR_OUT_16_port, Addr(15) => 
                           IRAM_ADDR_OUT_15_port, Addr(14) => 
                           IRAM_ADDR_OUT_14_port, Addr(13) => 
                           IRAM_ADDR_OUT_13_port, Addr(12) => 
                           IRAM_ADDR_OUT_12_port, Addr(11) => 
                           IRAM_ADDR_OUT_11_port, Addr(10) => 
                           IRAM_ADDR_OUT_10_port, Addr(9) => 
                           IRAM_ADDR_OUT_9_port, Addr(8) => 
                           IRAM_ADDR_OUT_8_port, Addr(7) => 
                           IRAM_ADDR_OUT_7_port, Addr(6) => 
                           IRAM_ADDR_OUT_6_port, Addr(5) => 
                           IRAM_ADDR_OUT_5_port, Addr(4) => 
                           IRAM_ADDR_OUT_4_port, Addr(3) => 
                           IRAM_ADDR_OUT_3_port, Addr(2) => 
                           IRAM_ADDR_OUT_2_port, Addr(1) => 
                           IRAM_ADDR_OUT_1_port, Addr(0) => 
                           IRAM_ADDR_OUT_0_port, Iout(31) => INS_IN_31_port, 
                           Iout(30) => INS_IN_30_port, Iout(29) => 
                           INS_IN_29_port, Iout(28) => INS_IN_28_port, Iout(27)
                           => INS_IN_27_port, Iout(26) => INS_IN_26_port, 
                           Iout(25) => INS_IN_25_port, Iout(24) => 
                           INS_IN_24_port, Iout(23) => INS_IN_23_port, Iout(22)
                           => INS_IN_22_port, Iout(21) => INS_IN_21_port, 
                           Iout(20) => INS_IN_20_port, Iout(19) => 
                           INS_IN_19_port, Iout(18) => INS_IN_18_port, Iout(17)
                           => INS_IN_17_port, Iout(16) => INS_IN_16_port, 
                           Iout(15) => INS_IN_15_port, Iout(14) => 
                           INS_IN_14_port, Iout(13) => INS_IN_13_port, Iout(12)
                           => INS_IN_12_port, Iout(11) => INS_IN_11_port, 
                           Iout(10) => INS_IN_10_port, Iout(9) => INS_IN_9_port
                           , Iout(8) => INS_IN_8_port, Iout(7) => INS_IN_7_port
                           , Iout(6) => INS_IN_6_port, Iout(5) => INS_IN_5_port
                           , Iout(4) => INS_IN_4_port, Iout(3) => INS_IN_3_port
                           , Iout(2) => INS_IN_2_port, Iout(1) => INS_IN_1_port
                           , Iout(0) => INS_IN_0_port);
   DRAM_I : DRAM port map( Clk => Clk, Rst => Rst, ADDR_IN(31) => 
                           DRAM_ADDR_OUT_31_port, ADDR_IN(30) => 
                           DRAM_ADDR_OUT_30_port, ADDR_IN(29) => 
                           DRAM_ADDR_OUT_29_port, ADDR_IN(28) => 
                           DRAM_ADDR_OUT_28_port, ADDR_IN(27) => 
                           DRAM_ADDR_OUT_27_port, ADDR_IN(26) => 
                           DRAM_ADDR_OUT_26_port, ADDR_IN(25) => 
                           DRAM_ADDR_OUT_25_port, ADDR_IN(24) => 
                           DRAM_ADDR_OUT_24_port, ADDR_IN(23) => 
                           DRAM_ADDR_OUT_23_port, ADDR_IN(22) => 
                           DRAM_ADDR_OUT_22_port, ADDR_IN(21) => 
                           DRAM_ADDR_OUT_21_port, ADDR_IN(20) => 
                           DRAM_ADDR_OUT_20_port, ADDR_IN(19) => 
                           DRAM_ADDR_OUT_19_port, ADDR_IN(18) => 
                           DRAM_ADDR_OUT_18_port, ADDR_IN(17) => 
                           DRAM_ADDR_OUT_17_port, ADDR_IN(16) => 
                           DRAM_ADDR_OUT_16_port, ADDR_IN(15) => 
                           DRAM_ADDR_OUT_15_port, ADDR_IN(14) => 
                           DRAM_ADDR_OUT_14_port, ADDR_IN(13) => 
                           DRAM_ADDR_OUT_13_port, ADDR_IN(12) => 
                           DRAM_ADDR_OUT_12_port, ADDR_IN(11) => 
                           DRAM_ADDR_OUT_11_port, ADDR_IN(10) => 
                           DRAM_ADDR_OUT_10_port, ADDR_IN(9) => 
                           DRAM_ADDR_OUT_9_port, ADDR_IN(8) => 
                           DRAM_ADDR_OUT_8_port, ADDR_IN(7) => 
                           DRAM_ADDR_OUT_7_port, ADDR_IN(6) => 
                           DRAM_ADDR_OUT_6_port, ADDR_IN(5) => 
                           DRAM_ADDR_OUT_5_port, ADDR_IN(4) => 
                           DRAM_ADDR_OUT_4_port, ADDR_IN(3) => 
                           DRAM_ADDR_OUT_3_port, ADDR_IN(2) => 
                           DRAM_ADDR_OUT_2_port, ADDR_IN(1) => 
                           DRAM_ADDR_OUT_1_port, ADDR_IN(0) => 
                           DRAM_ADDR_OUT_0_port, DATA_IN(31) => 
                           DATA_OUT_31_port, DATA_IN(30) => DATA_OUT_30_port, 
                           DATA_IN(29) => DATA_OUT_29_port, DATA_IN(28) => 
                           DATA_OUT_28_port, DATA_IN(27) => DATA_OUT_27_port, 
                           DATA_IN(26) => DATA_OUT_26_port, DATA_IN(25) => 
                           DATA_OUT_25_port, DATA_IN(24) => DATA_OUT_24_port, 
                           DATA_IN(23) => DATA_OUT_23_port, DATA_IN(22) => 
                           DATA_OUT_22_port, DATA_IN(21) => DATA_OUT_21_port, 
                           DATA_IN(20) => DATA_OUT_20_port, DATA_IN(19) => 
                           DATA_OUT_19_port, DATA_IN(18) => DATA_OUT_18_port, 
                           DATA_IN(17) => DATA_OUT_17_port, DATA_IN(16) => 
                           DATA_OUT_16_port, DATA_IN(15) => DATA_OUT_15_port, 
                           DATA_IN(14) => DATA_OUT_14_port, DATA_IN(13) => 
                           DATA_OUT_13_port, DATA_IN(12) => DATA_OUT_12_port, 
                           DATA_IN(11) => DATA_OUT_11_port, DATA_IN(10) => 
                           DATA_OUT_10_port, DATA_IN(9) => DATA_OUT_9_port, 
                           DATA_IN(8) => DATA_OUT_8_port, DATA_IN(7) => 
                           DATA_OUT_7_port, DATA_IN(6) => DATA_OUT_6_port, 
                           DATA_IN(5) => DATA_OUT_5_port, DATA_IN(4) => 
                           DATA_OUT_4_port, DATA_IN(3) => DATA_OUT_3_port, 
                           DATA_IN(2) => DATA_OUT_2_port, DATA_IN(1) => 
                           DATA_OUT_1_port, DATA_IN(0) => DATA_OUT_0_port, 
                           LOAD_TYPE(1) => LOAD_TYPE_OUT_1_port, LOAD_TYPE(0) 
                           => LOAD_TYPE_OUT_0_port, STORE_TYPE => 
                           STORE_TYPE_OUT, DRAM_W => DRAM_W_OUT, DRAM_R => 
                           DRAM_R_OUT, DATA_OUT(31) => DATA_IN_31_port, 
                           DATA_OUT(30) => DATA_IN_30_port, DATA_OUT(29) => 
                           DATA_IN_29_port, DATA_OUT(28) => DATA_IN_28_port, 
                           DATA_OUT(27) => DATA_IN_27_port, DATA_OUT(26) => 
                           DATA_IN_26_port, DATA_OUT(25) => DATA_IN_25_port, 
                           DATA_OUT(24) => DATA_IN_24_port, DATA_OUT(23) => 
                           DATA_IN_23_port, DATA_OUT(22) => DATA_IN_22_port, 
                           DATA_OUT(21) => DATA_IN_21_port, DATA_OUT(20) => 
                           DATA_IN_20_port, DATA_OUT(19) => DATA_IN_19_port, 
                           DATA_OUT(18) => DATA_IN_18_port, DATA_OUT(17) => 
                           DATA_IN_17_port, DATA_OUT(16) => DATA_IN_16_port, 
                           DATA_OUT(15) => DATA_IN_15_port, DATA_OUT(14) => 
                           DATA_IN_14_port, DATA_OUT(13) => DATA_IN_13_port, 
                           DATA_OUT(12) => DATA_IN_12_port, DATA_OUT(11) => 
                           DATA_IN_11_port, DATA_OUT(10) => DATA_IN_10_port, 
                           DATA_OUT(9) => DATA_IN_9_port, DATA_OUT(8) => 
                           DATA_IN_8_port, DATA_OUT(7) => DATA_IN_7_port, 
                           DATA_OUT(6) => DATA_IN_6_port, DATA_OUT(5) => 
                           DATA_IN_5_port, DATA_OUT(4) => DATA_IN_4_port, 
                           DATA_OUT(3) => DATA_IN_3_port, DATA_OUT(2) => 
                           DATA_IN_2_port, DATA_OUT(1) => DATA_IN_1_port, 
                           DATA_OUT(0) => DATA_IN_0_port);
   WB_MUX_SEL <= '0';
   STORE_TYPE_IN <= '0';
   LOAD_TYPE_IN_0_port <= '0';
   LOAD_TYPE_IN_1_port <= '0';
   RF_WE <= '0';
   DRAM_W_IN <= '0';
   MEM_EN_IN <= '0';
   JUMP_TYPE_0_port <= '0';
   JUMP_TYPE_1_port <= '0';
   DRAM_R_IN <= '0';
   ALU_OUTREG_EN <= '0';
   MUX_B_SEL_0_port <= '0';
   MUX_B_SEL_1_port <= '0';
   MUX_A_SEL <= '0';

end SYN_dlx_rtl;
