library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;
use work.constants.all;

entity tb_shifter is
end entity;

architecture test of tb_shifter is

  component shifter is
	generic(NBIT : integer);
	port( A           : in std_logic_vector(NBIT-1 downto 0); -- Operand to shift
	      B           : in std_logic_vector(NBIT-1 downto 0); -- Shift amount
	      LOGIC_ARITH : in std_logic;	-- 1 = logic, 0 = arith
	      LEFT_RIGHT  : in std_logic;	-- 1 = left, 0 = right
	      RES         : out std_logic_vector(NBIT-1 downto 0)
	);
 end component;

  constant tb_period : time := 10ns;
  signal A : std_logic_vector(NBIT-1 downto 0);
  signal B : std_logic_vector(NBIT-1 downto 0);
  signal LOGIC_ARITH : std_logic;
  signal LEFT_RIGHT: std_logic;
  signal RES : std_logic_vector(NBIT-1 downto 0);

begin
    
  dut_shifter : shifter
  generic map (NBIT => 32)
  port map (A => A,
            B => B,
            LOGIC_ARITH => LOGIC_ARITH,
            LEFT_RIGHT => LEFT_RIGHT,
            RES => RES);

  stimuli : process
                procedure apply_stimuli (
                        constant A_val : in std_logic_vector(NBIT-1 downto 0);
                        constant B_val : in integer;
                        constant LOGIC_ARITH_val : in std_logic;
                        constant LEFT_RIGHT_val: in std_logic;
                        signal A : out std_logic_vector(NBIT-1 downto 0);
                        signal B : out std_logic_vector(NBIT-1 downto 0);
                        signal LOGIC_ARITH : out std_logic;
                        signal LEFT_RIGHT: out std_logic ) is
                begin
                        A <= A_val;
                        B <= std_logic_vector(to_signed(B_val, NBIT));
                        LOGIC_ARITH <= LOGIC_ARITH_val;
                        LEFT_RIGHT <= LEFT_RIGHT_val;
                        wait for tb_period;
                end apply_stimuli;
  begin

   --apply_stimuli( , , '', '', A, B, LOGIC_ARITH, LEFT_RIGHT);
   
   -- x"F003_00F0" => 4,026,728,688
  
  for i in 0 to 4 loop
     apply_stimuli(x"0000_001A", i*2, '1', '0', A, B, LOGIC_ARITH, LEFT_RIGHT);
     apply_stimuli(x"0000_001A", i*2, '0', '0', A, B, LOGIC_ARITH, LEFT_RIGHT);
     apply_stimuli(x"0000_001A", i*2, '1', '1', A, B, LOGIC_ARITH, LEFT_RIGHT);
     apply_stimuli(x"0000_001A", i*2, '0', '1', A, B, LOGIC_ARITH, LEFT_RIGHT);
    
  
	   apply_stimuli(x"F003_8830", i*2, '1', '0', A, B, LOGIC_ARITH, LEFT_RIGHT);
   	  apply_stimuli(x"F003_8830", i*2, '0', '0', A, B, LOGIC_ARITH, LEFT_RIGHT);
   	  apply_stimuli(x"F003_8830", i*2, '1', '1', A, B, LOGIC_ARITH, LEFT_RIGHT);
   	  apply_stimuli(x"F003_8830", i*2, '0', '1', A, B, LOGIC_ARITH, LEFT_RIGHT);
--( -268238608)
  end loop;
 
  end process;
  
  

end test;
