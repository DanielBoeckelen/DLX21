
module mux21_NBIT32_0 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;

  MUX2_X1 U1 ( .A(B[29]), .B(A[29]), .S(n1), .Z(Z[29]) );
  INV_X32 U2 ( .A(n12), .ZN(n1) );
  NAND2_X1 U3 ( .A1(B[26]), .A2(n12), .ZN(n9) );
  INV_X1 U4 ( .A(n13), .ZN(n11) );
  INV_X1 U5 ( .A(n13), .ZN(n12) );
  MUX2_X1 U6 ( .A(A[19]), .B(B[19]), .S(S), .Z(Z[19]) );
  MUX2_X1 U7 ( .A(A[15]), .B(B[15]), .S(S), .Z(Z[15]) );
  NAND2_X1 U8 ( .A1(A[17]), .A2(n14), .ZN(n2) );
  NAND2_X1 U9 ( .A1(B[17]), .A2(n11), .ZN(n3) );
  NAND2_X1 U10 ( .A1(n2), .A2(n3), .ZN(Z[17]) );
  NAND2_X1 U11 ( .A1(A[28]), .A2(n14), .ZN(n4) );
  NAND2_X1 U12 ( .A1(B[28]), .A2(n11), .ZN(n5) );
  NAND2_X1 U13 ( .A1(n4), .A2(n5), .ZN(Z[28]) );
  NAND2_X1 U14 ( .A1(A[30]), .A2(n13), .ZN(n6) );
  NAND2_X1 U15 ( .A1(B[30]), .A2(n11), .ZN(n7) );
  NAND2_X1 U16 ( .A1(n6), .A2(n7), .ZN(Z[30]) );
  NAND2_X1 U17 ( .A1(A[26]), .A2(n14), .ZN(n8) );
  NAND2_X1 U18 ( .A1(n8), .A2(n9), .ZN(Z[26]) );
  INV_X1 U19 ( .A(n14), .ZN(n10) );
  INV_X1 U20 ( .A(S), .ZN(n13) );
  INV_X1 U21 ( .A(S), .ZN(n14) );
  MUX2_X1 U22 ( .A(A[0]), .B(B[0]), .S(n10), .Z(Z[0]) );
  MUX2_X1 U23 ( .A(A[1]), .B(B[1]), .S(n10), .Z(Z[1]) );
  MUX2_X1 U24 ( .A(A[2]), .B(B[2]), .S(n10), .Z(Z[2]) );
  MUX2_X1 U25 ( .A(A[3]), .B(B[3]), .S(n10), .Z(Z[3]) );
  MUX2_X1 U26 ( .A(A[4]), .B(B[4]), .S(n10), .Z(Z[4]) );
  MUX2_X1 U27 ( .A(A[5]), .B(B[5]), .S(n10), .Z(Z[5]) );
  MUX2_X1 U28 ( .A(A[6]), .B(B[6]), .S(n10), .Z(Z[6]) );
  MUX2_X1 U29 ( .A(A[7]), .B(B[7]), .S(n10), .Z(Z[7]) );
  MUX2_X1 U30 ( .A(A[8]), .B(B[8]), .S(n10), .Z(Z[8]) );
  MUX2_X1 U31 ( .A(A[9]), .B(B[9]), .S(n10), .Z(Z[9]) );
  MUX2_X1 U32 ( .A(A[10]), .B(B[10]), .S(n10), .Z(Z[10]) );
  MUX2_X1 U33 ( .A(A[11]), .B(B[11]), .S(n10), .Z(Z[11]) );
  MUX2_X1 U34 ( .A(A[12]), .B(B[12]), .S(n11), .Z(Z[12]) );
  MUX2_X1 U35 ( .A(A[13]), .B(B[13]), .S(n11), .Z(Z[13]) );
  MUX2_X1 U36 ( .A(A[14]), .B(B[14]), .S(n11), .Z(Z[14]) );
  MUX2_X1 U37 ( .A(A[16]), .B(B[16]), .S(n11), .Z(Z[16]) );
  MUX2_X1 U38 ( .A(A[18]), .B(B[18]), .S(n11), .Z(Z[18]) );
  MUX2_X1 U39 ( .A(A[20]), .B(B[20]), .S(n11), .Z(Z[20]) );
  MUX2_X1 U40 ( .A(A[21]), .B(B[21]), .S(n11), .Z(Z[21]) );
  MUX2_X1 U41 ( .A(A[22]), .B(B[22]), .S(n11), .Z(Z[22]) );
  AOI22_X1 U42 ( .A1(B[23]), .A2(n12), .B1(A[23]), .B2(n14), .ZN(n15) );
  INV_X1 U43 ( .A(n15), .ZN(Z[23]) );
  MUX2_X1 U44 ( .A(A[24]), .B(B[24]), .S(n11), .Z(Z[24]) );
  MUX2_X1 U45 ( .A(A[25]), .B(B[25]), .S(n12), .Z(Z[25]) );
  AOI22_X1 U46 ( .A1(A[27]), .A2(n13), .B1(B[27]), .B2(n12), .ZN(n16) );
  INV_X1 U47 ( .A(n16), .ZN(Z[27]) );
  AOI22_X1 U48 ( .A1(A[31]), .A2(n13), .B1(B[31]), .B2(n12), .ZN(n17) );
  INV_X1 U49 ( .A(n17), .ZN(Z[31]) );
endmodule


module mux21_NBIT32_5 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3;

  BUF_X1 U1 ( .A(S), .Z(n1) );
  BUF_X1 U2 ( .A(S), .Z(n2) );
  BUF_X1 U3 ( .A(S), .Z(n3) );
  MUX2_X1 U4 ( .A(A[0]), .B(B[0]), .S(n1), .Z(Z[0]) );
  MUX2_X1 U5 ( .A(A[1]), .B(B[1]), .S(n1), .Z(Z[1]) );
  MUX2_X1 U6 ( .A(A[2]), .B(B[2]), .S(n1), .Z(Z[2]) );
  MUX2_X1 U7 ( .A(A[3]), .B(B[3]), .S(n1), .Z(Z[3]) );
  MUX2_X1 U8 ( .A(A[4]), .B(B[4]), .S(n1), .Z(Z[4]) );
  MUX2_X1 U9 ( .A(A[5]), .B(B[5]), .S(n1), .Z(Z[5]) );
  MUX2_X1 U10 ( .A(A[6]), .B(B[6]), .S(n1), .Z(Z[6]) );
  MUX2_X1 U11 ( .A(A[7]), .B(B[7]), .S(n1), .Z(Z[7]) );
  MUX2_X1 U12 ( .A(A[8]), .B(B[8]), .S(n1), .Z(Z[8]) );
  MUX2_X1 U13 ( .A(A[9]), .B(B[9]), .S(n1), .Z(Z[9]) );
  MUX2_X1 U14 ( .A(A[10]), .B(B[10]), .S(n1), .Z(Z[10]) );
  MUX2_X1 U15 ( .A(A[11]), .B(B[11]), .S(n1), .Z(Z[11]) );
  MUX2_X1 U16 ( .A(A[12]), .B(B[12]), .S(n2), .Z(Z[12]) );
  MUX2_X1 U17 ( .A(A[13]), .B(B[13]), .S(n2), .Z(Z[13]) );
  MUX2_X1 U18 ( .A(A[14]), .B(B[14]), .S(n2), .Z(Z[14]) );
  MUX2_X1 U19 ( .A(A[15]), .B(B[15]), .S(n2), .Z(Z[15]) );
  MUX2_X1 U20 ( .A(A[16]), .B(B[16]), .S(n2), .Z(Z[16]) );
  MUX2_X1 U21 ( .A(A[17]), .B(B[17]), .S(n2), .Z(Z[17]) );
  MUX2_X1 U22 ( .A(A[18]), .B(B[18]), .S(n2), .Z(Z[18]) );
  MUX2_X1 U23 ( .A(A[19]), .B(B[19]), .S(n2), .Z(Z[19]) );
  MUX2_X1 U24 ( .A(A[20]), .B(B[20]), .S(n2), .Z(Z[20]) );
  MUX2_X1 U25 ( .A(A[21]), .B(B[21]), .S(n2), .Z(Z[21]) );
  MUX2_X1 U26 ( .A(A[22]), .B(B[22]), .S(n2), .Z(Z[22]) );
  MUX2_X1 U27 ( .A(A[23]), .B(B[23]), .S(n2), .Z(Z[23]) );
  MUX2_X1 U28 ( .A(A[24]), .B(B[24]), .S(n3), .Z(Z[24]) );
  MUX2_X1 U29 ( .A(A[25]), .B(B[25]), .S(n3), .Z(Z[25]) );
  MUX2_X1 U30 ( .A(A[26]), .B(B[26]), .S(n3), .Z(Z[26]) );
  MUX2_X1 U31 ( .A(A[27]), .B(B[27]), .S(n3), .Z(Z[27]) );
  MUX2_X1 U32 ( .A(A[28]), .B(B[28]), .S(n3), .Z(Z[28]) );
  MUX2_X1 U33 ( .A(A[29]), .B(B[29]), .S(n3), .Z(Z[29]) );
  MUX2_X1 U34 ( .A(A[30]), .B(B[30]), .S(n3), .Z(Z[30]) );
  MUX2_X1 U35 ( .A(A[31]), .B(B[31]), .S(n3), .Z(Z[31]) );
endmodule


module mux21_NBIT32_4 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111;

  INV_X1 U1 ( .A(n15), .ZN(n4) );
  INV_X1 U2 ( .A(n15), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n7) );
  BUF_X1 U4 ( .A(n3), .Z(n13) );
  BUF_X1 U5 ( .A(n2), .Z(n12) );
  BUF_X1 U6 ( .A(n2), .Z(n10) );
  BUF_X1 U7 ( .A(n1), .Z(n9) );
  BUF_X1 U8 ( .A(n2), .Z(n11) );
  BUF_X1 U9 ( .A(n1), .Z(n8) );
  BUF_X1 U10 ( .A(n3), .Z(n15) );
  BUF_X1 U11 ( .A(n3), .Z(n14) );
  BUF_X1 U12 ( .A(S), .Z(n3) );
  BUF_X1 U13 ( .A(S), .Z(n2) );
  BUF_X1 U14 ( .A(S), .Z(n1) );
  INV_X1 U15 ( .A(n91), .ZN(Z[1]) );
  AOI22_X1 U16 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(n11), .ZN(n91) );
  INV_X1 U17 ( .A(n102), .ZN(Z[2]) );
  AOI22_X1 U18 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n8), .ZN(n102) );
  INV_X1 U19 ( .A(n105), .ZN(Z[3]) );
  AOI22_X1 U20 ( .A1(A[3]), .A2(n6), .B1(B[3]), .B2(n8), .ZN(n105) );
  INV_X1 U21 ( .A(n106), .ZN(Z[4]) );
  AOI22_X1 U22 ( .A1(A[4]), .A2(n6), .B1(B[4]), .B2(n8), .ZN(n106) );
  INV_X1 U23 ( .A(n107), .ZN(Z[5]) );
  AOI22_X1 U24 ( .A1(A[5]), .A2(n6), .B1(B[5]), .B2(n7), .ZN(n107) );
  INV_X1 U25 ( .A(n108), .ZN(Z[6]) );
  AOI22_X1 U26 ( .A1(A[6]), .A2(n6), .B1(B[6]), .B2(n7), .ZN(n108) );
  INV_X1 U27 ( .A(n109), .ZN(Z[7]) );
  AOI22_X1 U28 ( .A1(A[7]), .A2(n6), .B1(B[7]), .B2(n7), .ZN(n109) );
  INV_X1 U29 ( .A(n110), .ZN(Z[8]) );
  AOI22_X1 U30 ( .A1(A[8]), .A2(n6), .B1(B[8]), .B2(n7), .ZN(n110) );
  INV_X1 U31 ( .A(n81), .ZN(Z[10]) );
  AOI22_X1 U32 ( .A1(A[10]), .A2(n4), .B1(B[10]), .B2(n14), .ZN(n81) );
  INV_X1 U33 ( .A(n82), .ZN(Z[11]) );
  AOI22_X1 U34 ( .A1(A[11]), .A2(n4), .B1(B[11]), .B2(n14), .ZN(n82) );
  INV_X1 U35 ( .A(n83), .ZN(Z[12]) );
  AOI22_X1 U36 ( .A1(A[12]), .A2(n4), .B1(B[12]), .B2(n13), .ZN(n83) );
  INV_X1 U37 ( .A(n84), .ZN(Z[13]) );
  AOI22_X1 U38 ( .A1(A[13]), .A2(n4), .B1(B[13]), .B2(n13), .ZN(n84) );
  INV_X1 U39 ( .A(n85), .ZN(Z[14]) );
  AOI22_X1 U40 ( .A1(A[14]), .A2(n4), .B1(B[14]), .B2(n13), .ZN(n85) );
  INV_X1 U41 ( .A(n86), .ZN(Z[15]) );
  AOI22_X1 U42 ( .A1(A[15]), .A2(n4), .B1(B[15]), .B2(n13), .ZN(n86) );
  INV_X1 U43 ( .A(n87), .ZN(Z[16]) );
  AOI22_X1 U44 ( .A1(A[16]), .A2(n4), .B1(B[16]), .B2(n12), .ZN(n87) );
  INV_X1 U45 ( .A(n88), .ZN(Z[17]) );
  AOI22_X1 U46 ( .A1(A[17]), .A2(n4), .B1(B[17]), .B2(n12), .ZN(n88) );
  INV_X1 U47 ( .A(n89), .ZN(Z[18]) );
  AOI22_X1 U48 ( .A1(A[18]), .A2(n4), .B1(B[18]), .B2(n12), .ZN(n89) );
  INV_X1 U49 ( .A(n90), .ZN(Z[19]) );
  AOI22_X1 U50 ( .A1(A[19]), .A2(n4), .B1(B[19]), .B2(n12), .ZN(n90) );
  INV_X1 U51 ( .A(n92), .ZN(Z[20]) );
  AOI22_X1 U52 ( .A1(A[20]), .A2(n5), .B1(B[20]), .B2(n11), .ZN(n92) );
  INV_X1 U53 ( .A(n93), .ZN(Z[21]) );
  AOI22_X1 U54 ( .A1(A[21]), .A2(n5), .B1(B[21]), .B2(n11), .ZN(n93) );
  INV_X1 U55 ( .A(n94), .ZN(Z[22]) );
  AOI22_X1 U56 ( .A1(A[22]), .A2(n5), .B1(B[22]), .B2(n10), .ZN(n94) );
  INV_X1 U57 ( .A(n95), .ZN(Z[23]) );
  AOI22_X1 U58 ( .A1(A[23]), .A2(n5), .B1(B[23]), .B2(n10), .ZN(n95) );
  INV_X1 U59 ( .A(n96), .ZN(Z[24]) );
  AOI22_X1 U60 ( .A1(A[24]), .A2(n5), .B1(B[24]), .B2(n10), .ZN(n96) );
  INV_X1 U61 ( .A(n97), .ZN(Z[25]) );
  AOI22_X1 U62 ( .A1(A[25]), .A2(n5), .B1(B[25]), .B2(n10), .ZN(n97) );
  INV_X1 U63 ( .A(n98), .ZN(Z[26]) );
  AOI22_X1 U64 ( .A1(A[26]), .A2(n5), .B1(B[26]), .B2(n9), .ZN(n98) );
  INV_X1 U65 ( .A(n99), .ZN(Z[27]) );
  AOI22_X1 U66 ( .A1(A[27]), .A2(n5), .B1(B[27]), .B2(n9), .ZN(n99) );
  INV_X1 U67 ( .A(n100), .ZN(Z[28]) );
  AOI22_X1 U68 ( .A1(A[28]), .A2(n5), .B1(B[28]), .B2(n9), .ZN(n100) );
  INV_X1 U69 ( .A(n101), .ZN(Z[29]) );
  AOI22_X1 U70 ( .A1(A[29]), .A2(n5), .B1(B[29]), .B2(n9), .ZN(n101) );
  INV_X1 U71 ( .A(n103), .ZN(Z[30]) );
  AOI22_X1 U72 ( .A1(A[30]), .A2(n5), .B1(B[30]), .B2(n11), .ZN(n103) );
  INV_X1 U73 ( .A(n104), .ZN(Z[31]) );
  AOI22_X1 U74 ( .A1(A[31]), .A2(n6), .B1(B[31]), .B2(n8), .ZN(n104) );
  INV_X1 U75 ( .A(n111), .ZN(Z[9]) );
  AOI22_X1 U76 ( .A1(A[9]), .A2(n6), .B1(n14), .B2(B[9]), .ZN(n111) );
  INV_X1 U77 ( .A(n80), .ZN(Z[0]) );
  AOI22_X1 U78 ( .A1(A[0]), .A2(n4), .B1(B[0]), .B2(n14), .ZN(n80) );
  INV_X1 U79 ( .A(n15), .ZN(n6) );
endmodule


module regn_N32_0 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n31, n99, n101, n102, n103, n104, n105, n106, n107, n108,
         n110, n111, n112, n113, n114, n115, n116;

  DFFR_X1 \DOUT_reg[31]  ( .D(n96), .CK(CLK), .RN(n19), .Q(DOUT[31]), .QN(n64)
         );
  DFFR_X1 \DOUT_reg[30]  ( .D(n95), .CK(CLK), .RN(n19), .Q(DOUT[30]), .QN(n63)
         );
  DFFR_X1 \DOUT_reg[28]  ( .D(n93), .CK(CLK), .RN(n19), .Q(DOUT[28]), .QN(n61)
         );
  DFFR_X1 \DOUT_reg[26]  ( .D(n91), .CK(CLK), .RN(n19), .Q(DOUT[26]), .QN(n59)
         );
  DFFR_X1 \DOUT_reg[25]  ( .D(n90), .CK(CLK), .RN(n19), .Q(DOUT[25]), .QN(n58)
         );
  DFFR_X1 \DOUT_reg[24]  ( .D(n89), .CK(CLK), .RN(n19), .Q(n117), .QN(n57) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n88), .CK(CLK), .RN(n18), .Q(DOUT[23]), .QN(n56)
         );
  DFFR_X1 \DOUT_reg[22]  ( .D(n87), .CK(CLK), .RN(n18), .Q(DOUT[22]), .QN(n55)
         );
  DFFR_X1 \DOUT_reg[21]  ( .D(n86), .CK(CLK), .RN(n18), .Q(DOUT[21]), .QN(n54)
         );
  DFFR_X1 \DOUT_reg[20]  ( .D(n85), .CK(CLK), .RN(n18), .Q(DOUT[20]), .QN(n53)
         );
  DFFR_X1 \DOUT_reg[19]  ( .D(n84), .CK(CLK), .RN(n18), .Q(DOUT[19]), .QN(n52)
         );
  DFFR_X1 \DOUT_reg[18]  ( .D(n83), .CK(CLK), .RN(n18), .Q(DOUT[18]), .QN(n51)
         );
  DFFR_X1 \DOUT_reg[17]  ( .D(n82), .CK(CLK), .RN(n18), .Q(DOUT[17]), .QN(n50)
         );
  DFFR_X1 \DOUT_reg[16]  ( .D(n81), .CK(CLK), .RN(n18), .Q(n118), .QN(n49) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n80), .CK(CLK), .RN(n18), .Q(DOUT[15]), .QN(n48)
         );
  DFFR_X1 \DOUT_reg[14]  ( .D(n79), .CK(CLK), .RN(n18), .QN(n47) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n78), .CK(CLK), .RN(n18), .Q(n119), .QN(n46) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n77), .CK(CLK), .RN(n18), .Q(n120), .QN(n45) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n76), .CK(CLK), .RN(n17), .Q(DOUT[11]), .QN(n44)
         );
  DFFR_X1 \DOUT_reg[10]  ( .D(n75), .CK(CLK), .RN(n17), .Q(n121), .QN(n43) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n74), .CK(CLK), .RN(n17), .Q(n122), .QN(n42) );
  DFFR_X1 \DOUT_reg[8]  ( .D(n73), .CK(CLK), .RN(n17), .Q(n123), .QN(n41) );
  DFFR_X1 \DOUT_reg[7]  ( .D(n72), .CK(CLK), .RN(n17), .Q(n124), .QN(n40) );
  DFFR_X1 \DOUT_reg[6]  ( .D(n71), .CK(CLK), .RN(n17), .Q(n125), .QN(n39) );
  DFFR_X1 \DOUT_reg[5]  ( .D(n70), .CK(CLK), .RN(n17), .Q(n126), .QN(n38) );
  DFFR_X1 \DOUT_reg[4]  ( .D(n69), .CK(CLK), .RN(n17), .Q(n127), .QN(n37) );
  DFFR_X1 \DOUT_reg[3]  ( .D(n68), .CK(CLK), .RN(n17), .Q(n128), .QN(n36) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n67), .CK(CLK), .RN(n17), .Q(n129), .QN(n35) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n66), .CK(CLK), .RN(n17), .Q(DOUT[1]), .QN(n34)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n65), .CK(CLK), .RN(n17), .Q(DOUT[0]), .QN(n33)
         );
  DFFR_X1 \DOUT_reg[27]  ( .D(n92), .CK(CLK), .RN(n19), .Q(DOUT[27]), .QN(n60)
         );
  DFFR_X2 \DOUT_reg[29]  ( .D(n94), .CK(CLK), .RN(n19), .Q(DOUT[29]), .QN(n62)
         );
  INV_X1 U2 ( .A(EN), .ZN(n5) );
  INV_X1 U3 ( .A(EN), .ZN(n4) );
  INV_X1 U4 ( .A(EN), .ZN(n6) );
  INV_X1 U5 ( .A(EN), .ZN(n7) );
  INV_X1 U6 ( .A(EN), .ZN(n3) );
  INV_X1 U7 ( .A(EN), .ZN(n2) );
  INV_X1 U8 ( .A(EN), .ZN(n1) );
  MUX2_X1 U9 ( .A(DIN[0]), .B(n20), .S(n1), .Z(n65) );
  MUX2_X1 U10 ( .A(DIN[4]), .B(n127), .S(n2), .Z(n69) );
  MUX2_X1 U11 ( .A(DIN[3]), .B(n128), .S(n3), .Z(n68) );
  MUX2_X1 U12 ( .A(DIN[5]), .B(n126), .S(n4), .Z(n70) );
  MUX2_X1 U13 ( .A(DIN[1]), .B(n21), .S(n5), .Z(n66) );
  MUX2_X1 U14 ( .A(DIN[6]), .B(n125), .S(n5), .Z(n71) );
  MUX2_X1 U15 ( .A(DIN[10]), .B(n121), .S(n6), .Z(n75) );
  MUX2_X1 U16 ( .A(DIN[16]), .B(n118), .S(n7), .Z(n81) );
  INV_X1 U17 ( .A(n49), .ZN(DOUT[16]) );
  MUX2_X1 U18 ( .A(DIN[24]), .B(n117), .S(n3), .Z(n89) );
  MUX2_X1 U19 ( .A(DIN[8]), .B(n123), .S(n2), .Z(n73) );
  MUX2_X1 U20 ( .A(DIN[12]), .B(n120), .S(n1), .Z(n77) );
  NAND2_X1 U21 ( .A1(DIN[7]), .A2(EN), .ZN(n8) );
  NAND2_X1 U22 ( .A1(n124), .A2(n108), .ZN(n9) );
  NAND2_X1 U23 ( .A1(n8), .A2(n9), .ZN(n72) );
  OR2_X1 U24 ( .A1(n58), .A2(EN), .ZN(n10) );
  NAND2_X1 U25 ( .A1(n110), .A2(n10), .ZN(n90) );
  OR2_X2 U26 ( .A1(n62), .A2(EN), .ZN(n11) );
  NAND2_X1 U27 ( .A1(n114), .A2(n11), .ZN(n94) );
  OR2_X1 U28 ( .A1(n61), .A2(EN), .ZN(n12) );
  NAND2_X1 U29 ( .A1(n113), .A2(n12), .ZN(n93) );
  OR2_X1 U30 ( .A1(n63), .A2(EN), .ZN(n13) );
  NAND2_X1 U31 ( .A1(n115), .A2(n13), .ZN(n95) );
  OR2_X2 U32 ( .A1(n50), .A2(EN), .ZN(n14) );
  NAND2_X1 U33 ( .A1(n101), .A2(n14), .ZN(n82) );
  OR2_X2 U34 ( .A1(n44), .A2(EN), .ZN(n15) );
  NAND2_X1 U35 ( .A1(n31), .A2(n15), .ZN(n76) );
  OR2_X2 U36 ( .A1(n59), .A2(EN), .ZN(n16) );
  NAND2_X1 U37 ( .A1(n111), .A2(n16), .ZN(n91) );
  BUF_X1 U38 ( .A(RST), .Z(n17) );
  BUF_X1 U39 ( .A(RST), .Z(n18) );
  BUF_X1 U40 ( .A(RST), .Z(n19) );
  INV_X1 U41 ( .A(EN), .ZN(n108) );
  OAI22_X1 U42 ( .A1(n107), .A2(n108), .B1(n56), .B2(EN), .ZN(n88) );
  INV_X1 U43 ( .A(DIN[23]), .ZN(n107) );
  INV_X1 U44 ( .A(n33), .ZN(n20) );
  INV_X1 U45 ( .A(n34), .ZN(n21) );
  INV_X1 U46 ( .A(n35), .ZN(DOUT[2]) );
  MUX2_X1 U47 ( .A(n129), .B(DIN[2]), .S(EN), .Z(n67) );
  INV_X1 U48 ( .A(n36), .ZN(DOUT[3]) );
  INV_X1 U49 ( .A(n37), .ZN(DOUT[4]) );
  INV_X1 U50 ( .A(n38), .ZN(DOUT[5]) );
  INV_X1 U51 ( .A(n39), .ZN(DOUT[6]) );
  INV_X1 U52 ( .A(n40), .ZN(DOUT[7]) );
  INV_X1 U53 ( .A(n41), .ZN(DOUT[8]) );
  INV_X1 U54 ( .A(n42), .ZN(DOUT[9]) );
  MUX2_X1 U55 ( .A(n122), .B(DIN[9]), .S(EN), .Z(n74) );
  INV_X1 U56 ( .A(n43), .ZN(DOUT[10]) );
  NAND2_X1 U57 ( .A1(DIN[11]), .A2(EN), .ZN(n31) );
  INV_X1 U58 ( .A(n45), .ZN(DOUT[12]) );
  INV_X1 U59 ( .A(n46), .ZN(DOUT[13]) );
  MUX2_X1 U60 ( .A(n119), .B(DIN[13]), .S(EN), .Z(n78) );
  INV_X1 U61 ( .A(n47), .ZN(DOUT[14]) );
  MUX2_X1 U62 ( .A(DOUT[14]), .B(DIN[14]), .S(EN), .Z(n79) );
  NAND2_X1 U63 ( .A1(DIN[15]), .A2(EN), .ZN(n99) );
  OAI21_X1 U64 ( .B1(n48), .B2(EN), .A(n99), .ZN(n80) );
  NAND2_X1 U65 ( .A1(DIN[17]), .A2(EN), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[18]), .A2(EN), .ZN(n102) );
  OAI21_X1 U67 ( .B1(n51), .B2(EN), .A(n102), .ZN(n83) );
  NAND2_X1 U68 ( .A1(DIN[19]), .A2(EN), .ZN(n103) );
  OAI21_X1 U69 ( .B1(n52), .B2(EN), .A(n103), .ZN(n84) );
  NAND2_X1 U70 ( .A1(DIN[20]), .A2(EN), .ZN(n104) );
  OAI21_X1 U71 ( .B1(n53), .B2(EN), .A(n104), .ZN(n85) );
  NAND2_X1 U72 ( .A1(DIN[21]), .A2(EN), .ZN(n105) );
  OAI21_X1 U73 ( .B1(n54), .B2(EN), .A(n105), .ZN(n86) );
  NAND2_X1 U74 ( .A1(DIN[22]), .A2(EN), .ZN(n106) );
  OAI21_X1 U75 ( .B1(n55), .B2(EN), .A(n106), .ZN(n87) );
  INV_X1 U76 ( .A(n57), .ZN(DOUT[24]) );
  NAND2_X1 U77 ( .A1(DIN[25]), .A2(EN), .ZN(n110) );
  NAND2_X1 U78 ( .A1(DIN[26]), .A2(EN), .ZN(n111) );
  NAND2_X1 U79 ( .A1(DIN[27]), .A2(EN), .ZN(n112) );
  OAI21_X1 U80 ( .B1(n60), .B2(EN), .A(n112), .ZN(n92) );
  NAND2_X1 U81 ( .A1(DIN[28]), .A2(EN), .ZN(n113) );
  NAND2_X1 U82 ( .A1(DIN[29]), .A2(EN), .ZN(n114) );
  NAND2_X1 U83 ( .A1(DIN[30]), .A2(EN), .ZN(n115) );
  NAND2_X1 U84 ( .A1(DIN[31]), .A2(EN), .ZN(n116) );
  OAI21_X1 U85 ( .B1(n64), .B2(EN), .A(n116), .ZN(n96) );
endmodule


module regn_N32_10 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n68, n69, n70;

  DFFR_X1 \DOUT_reg[31]  ( .D(n36), .CK(CLK), .RN(n3), .Q(DOUT[31]) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n37), .CK(CLK), .RN(n3), .Q(DOUT[30]) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n38), .CK(CLK), .RN(n3), .Q(DOUT[29]) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n39), .CK(CLK), .RN(n3), .Q(DOUT[28]) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n40), .CK(CLK), .RN(n3), .Q(DOUT[27]) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n41), .CK(CLK), .RN(n3), .Q(DOUT[26]) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n42), .CK(CLK), .RN(n3), .Q(DOUT[25]) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n43), .CK(CLK), .RN(n3), .Q(DOUT[24]) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n44), .CK(CLK), .RN(n2), .Q(DOUT[23]) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n45), .CK(CLK), .RN(n2), .Q(DOUT[22]) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n46), .CK(CLK), .RN(n2), .Q(DOUT[21]) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n47), .CK(CLK), .RN(n2), .Q(DOUT[20]) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n48), .CK(CLK), .RN(n2), .Q(DOUT[19]) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n49), .CK(CLK), .RN(n2), .Q(DOUT[18]) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n50), .CK(CLK), .RN(n2), .Q(DOUT[17]) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n51), .CK(CLK), .RN(n2), .Q(DOUT[16]) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n52), .CK(CLK), .RN(n2), .Q(DOUT[15]) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n53), .CK(CLK), .RN(n2), .Q(DOUT[14]) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n54), .CK(CLK), .RN(n2), .Q(DOUT[13]) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n55), .CK(CLK), .RN(n2), .Q(DOUT[12]) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n56), .CK(CLK), .RN(n1), .Q(DOUT[11]) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n57), .CK(CLK), .RN(n1), .Q(DOUT[10]) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n58), .CK(CLK), .RN(n1), .Q(DOUT[9]) );
  DFFR_X1 \DOUT_reg[8]  ( .D(n59), .CK(CLK), .RN(n1), .Q(DOUT[8]) );
  DFFR_X1 \DOUT_reg[7]  ( .D(n60), .CK(CLK), .RN(n1), .Q(DOUT[7]) );
  DFFR_X1 \DOUT_reg[6]  ( .D(n61), .CK(CLK), .RN(n1), .Q(DOUT[6]) );
  DFFR_X1 \DOUT_reg[5]  ( .D(n62), .CK(CLK), .RN(n1), .Q(DOUT[5]) );
  DFFR_X1 \DOUT_reg[4]  ( .D(n63), .CK(CLK), .RN(n1), .Q(DOUT[4]) );
  DFFR_X1 \DOUT_reg[3]  ( .D(n64), .CK(CLK), .RN(n1), .Q(DOUT[3]) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n68), .CK(CLK), .RN(n1), .Q(DOUT[2]) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n69), .CK(CLK), .RN(n1), .Q(DOUT[1]) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n70), .CK(CLK), .RN(n1), .Q(DOUT[0]) );
  BUF_X1 U2 ( .A(RST), .Z(n1) );
  BUF_X1 U3 ( .A(RST), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n3) );
  MUX2_X1 U5 ( .A(DOUT[0]), .B(DIN[0]), .S(EN), .Z(n70) );
  MUX2_X1 U6 ( .A(DOUT[1]), .B(DIN[1]), .S(EN), .Z(n69) );
  MUX2_X1 U7 ( .A(DOUT[2]), .B(DIN[2]), .S(EN), .Z(n68) );
  MUX2_X1 U8 ( .A(DOUT[3]), .B(DIN[3]), .S(EN), .Z(n64) );
  MUX2_X1 U9 ( .A(DOUT[4]), .B(DIN[4]), .S(EN), .Z(n63) );
  MUX2_X1 U10 ( .A(DOUT[5]), .B(DIN[5]), .S(EN), .Z(n62) );
  MUX2_X1 U11 ( .A(DOUT[6]), .B(DIN[6]), .S(EN), .Z(n61) );
  MUX2_X1 U12 ( .A(DOUT[7]), .B(DIN[7]), .S(EN), .Z(n60) );
  MUX2_X1 U13 ( .A(DOUT[8]), .B(DIN[8]), .S(EN), .Z(n59) );
  MUX2_X1 U14 ( .A(DOUT[9]), .B(DIN[9]), .S(EN), .Z(n58) );
  MUX2_X1 U15 ( .A(DOUT[10]), .B(DIN[10]), .S(EN), .Z(n57) );
  MUX2_X1 U16 ( .A(DOUT[11]), .B(DIN[11]), .S(EN), .Z(n56) );
  MUX2_X1 U17 ( .A(DOUT[12]), .B(DIN[12]), .S(EN), .Z(n55) );
  MUX2_X1 U18 ( .A(DOUT[13]), .B(DIN[13]), .S(EN), .Z(n54) );
  MUX2_X1 U19 ( .A(DOUT[14]), .B(DIN[14]), .S(EN), .Z(n53) );
  MUX2_X1 U20 ( .A(DOUT[15]), .B(DIN[15]), .S(EN), .Z(n52) );
  MUX2_X1 U21 ( .A(DOUT[16]), .B(DIN[16]), .S(EN), .Z(n51) );
  MUX2_X1 U22 ( .A(DOUT[17]), .B(DIN[17]), .S(EN), .Z(n50) );
  MUX2_X1 U23 ( .A(DOUT[18]), .B(DIN[18]), .S(EN), .Z(n49) );
  MUX2_X1 U24 ( .A(DOUT[19]), .B(DIN[19]), .S(EN), .Z(n48) );
  MUX2_X1 U25 ( .A(DOUT[20]), .B(DIN[20]), .S(EN), .Z(n47) );
  MUX2_X1 U26 ( .A(DOUT[21]), .B(DIN[21]), .S(EN), .Z(n46) );
  MUX2_X1 U27 ( .A(DOUT[22]), .B(DIN[22]), .S(EN), .Z(n45) );
  MUX2_X1 U28 ( .A(DOUT[23]), .B(DIN[23]), .S(EN), .Z(n44) );
  MUX2_X1 U29 ( .A(DOUT[24]), .B(DIN[24]), .S(EN), .Z(n43) );
  MUX2_X1 U30 ( .A(DOUT[25]), .B(DIN[25]), .S(EN), .Z(n42) );
  MUX2_X1 U31 ( .A(DOUT[26]), .B(DIN[26]), .S(EN), .Z(n41) );
  MUX2_X1 U32 ( .A(DOUT[27]), .B(DIN[27]), .S(EN), .Z(n40) );
  MUX2_X1 U33 ( .A(DOUT[28]), .B(DIN[28]), .S(EN), .Z(n39) );
  MUX2_X1 U34 ( .A(DOUT[29]), .B(DIN[29]), .S(EN), .Z(n38) );
  MUX2_X1 U35 ( .A(DOUT[30]), .B(DIN[30]), .S(EN), .Z(n37) );
  MUX2_X1 U36 ( .A(DOUT[31]), .B(DIN[31]), .S(EN), .Z(n36) );
endmodule


module regn_N32_9 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(
        n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(
        n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(
        n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(
        n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(
        n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(
        n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(
        n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(
        n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(
        n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(
        n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(
        n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(
        n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(
        n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(
        n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(
        n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(
        n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(
        n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(
        n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(
        n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(
        n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(
        n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(
        n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U6 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U7 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U8 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U9 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U10 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U11 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U12 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U13 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U14 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U15 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U16 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U17 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U18 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U19 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U20 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U21 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U22 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U23 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U24 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U25 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U26 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U27 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U28 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U29 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U30 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U31 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U32 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U33 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U34 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U35 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U36 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U37 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U38 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U39 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U40 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U41 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U42 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U43 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U44 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U45 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U46 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U47 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U48 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U49 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U50 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U51 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U52 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U53 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U54 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U55 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U56 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U57 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U58 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U59 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U60 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U61 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U62 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U63 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U64 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
  OAI21_X1 U65 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U66 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U67 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U68 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
endmodule


module Fetch_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XNOR2_X1 U2 ( .A(n116), .B(n69), .ZN(SUM[5]) );
  XOR2_X1 U3 ( .A(n1), .B(n3), .Z(SUM[14]) );
  AND2_X1 U4 ( .A1(n109), .A2(n59), .ZN(n1) );
  AND2_X1 U5 ( .A1(n2), .A2(n109), .ZN(n107) );
  AND2_X1 U6 ( .A1(n59), .A2(n3), .ZN(n2) );
  INV_X1 U7 ( .A(n108), .ZN(n3) );
  BUF_X1 U8 ( .A(n58), .Z(n26) );
  AND2_X1 U9 ( .A1(A[24]), .A2(A[25]), .ZN(n4) );
  AND2_X1 U10 ( .A1(n70), .A2(n31), .ZN(n5) );
  BUF_X1 U11 ( .A(A[4]), .Z(n20) );
  INV_X1 U12 ( .A(n10), .ZN(n6) );
  XOR2_X1 U13 ( .A(n7), .B(n35), .Z(SUM[9]) );
  NOR2_X1 U14 ( .A1(n76), .A2(n22), .ZN(n7) );
  CLKBUF_X1 U15 ( .A(A[16]), .Z(n8) );
  AND2_X1 U16 ( .A1(n57), .A2(n41), .ZN(n9) );
  INV_X1 U17 ( .A(n53), .ZN(n10) );
  AND2_X1 U18 ( .A1(n69), .A2(n11), .ZN(n13) );
  NOR2_X1 U19 ( .A1(n116), .A2(n10), .ZN(n11) );
  XOR2_X1 U20 ( .A(n12), .B(n72), .Z(SUM[8]) );
  NOR2_X1 U21 ( .A1(n76), .A2(n75), .ZN(n12) );
  NOR2_X1 U22 ( .A1(n78), .A2(n116), .ZN(n77) );
  XOR2_X1 U23 ( .A(n13), .B(n36), .Z(SUM[7]) );
  XOR2_X1 U24 ( .A(A[12]), .B(n14), .Z(SUM[12]) );
  NOR2_X1 U25 ( .A1(n62), .A2(n19), .ZN(n14) );
  XNOR2_X1 U26 ( .A(n15), .B(n111), .ZN(SUM[13]) );
  AND2_X1 U27 ( .A1(n23), .A2(n12), .ZN(n15) );
  BUF_X1 U28 ( .A(n113), .Z(n16) );
  NOR2_X1 U29 ( .A1(n76), .A2(n17), .ZN(n59) );
  NAND2_X1 U30 ( .A1(n18), .A2(n60), .ZN(n17) );
  AND2_X1 U31 ( .A1(A[3]), .A2(A[2]), .ZN(n18) );
  AND2_X1 U32 ( .A1(A[2]), .A2(A[3]), .ZN(n79) );
  NAND4_X1 U33 ( .A1(n112), .A2(n46), .A3(n31), .A4(n35), .ZN(n19) );
  XOR2_X1 U34 ( .A(n21), .B(n43), .Z(SUM[21]) );
  AND2_X1 U35 ( .A1(n26), .A2(n9), .ZN(n21) );
  NAND2_X1 U36 ( .A1(n18), .A2(A[8]), .ZN(n22) );
  NOR2_X1 U37 ( .A1(n19), .A2(n105), .ZN(n23) );
  NAND2_X1 U38 ( .A1(A[16]), .A2(A[17]), .ZN(n24) );
  CLKBUF_X1 U39 ( .A(A[2]), .Z(n25) );
  XOR2_X1 U40 ( .A(n54), .B(A[31]), .Z(SUM[31]) );
  CLKBUF_X1 U41 ( .A(n57), .Z(n27) );
  XNOR2_X1 U42 ( .A(n28), .B(n88), .ZN(SUM[29]) );
  NOR2_X1 U43 ( .A1(n71), .A2(n86), .ZN(n28) );
  XOR2_X1 U44 ( .A(n48), .B(n29), .Z(SUM[17]) );
  AND2_X1 U45 ( .A1(n26), .A2(n8), .ZN(n29) );
  NAND2_X1 U46 ( .A1(n114), .A2(n115), .ZN(n30) );
  BUF_X1 U47 ( .A(A[10]), .Z(n31) );
  AND2_X1 U48 ( .A1(n45), .A2(n85), .ZN(n89) );
  AND2_X1 U49 ( .A1(n61), .A2(n4), .ZN(n92) );
  NOR3_X1 U50 ( .A1(n83), .A2(n82), .A3(n81), .ZN(n54) );
  CLKBUF_X1 U51 ( .A(A[3]), .Z(n32) );
  CLKBUF_X1 U52 ( .A(A[15]), .Z(n33) );
  CLKBUF_X1 U53 ( .A(A[23]), .Z(n34) );
  BUF_X1 U54 ( .A(A[9]), .Z(n35) );
  CLKBUF_X1 U55 ( .A(A[7]), .Z(n36) );
  CLKBUF_X1 U56 ( .A(A[22]), .Z(n37) );
  XNOR2_X1 U57 ( .A(n38), .B(n90), .ZN(SUM[28]) );
  NOR2_X1 U58 ( .A1(n71), .A2(n44), .ZN(n38) );
  AND2_X1 U59 ( .A1(n4), .A2(A[26]), .ZN(n39) );
  AND2_X1 U60 ( .A1(n61), .A2(n39), .ZN(n66) );
  XOR2_X1 U61 ( .A(n40), .B(n41), .Z(SUM[20]) );
  AND2_X1 U62 ( .A1(n27), .A2(n58), .ZN(n40) );
  AND2_X1 U63 ( .A1(n101), .A2(n102), .ZN(n45) );
  BUF_X1 U64 ( .A(A[20]), .Z(n41) );
  NOR2_X1 U65 ( .A1(n87), .A2(n90), .ZN(n42) );
  CLKBUF_X1 U66 ( .A(A[21]), .Z(n43) );
  CLKBUF_X1 U67 ( .A(n87), .Z(n44) );
  INV_X1 U68 ( .A(n113), .ZN(n46) );
  AND3_X1 U69 ( .A1(A[22]), .A2(A[21]), .A3(A[23]), .ZN(n47) );
  AND2_X1 U70 ( .A1(n47), .A2(n41), .ZN(n63) );
  CLKBUF_X1 U71 ( .A(A[17]), .Z(n48) );
  NAND2_X1 U72 ( .A1(A[19]), .A2(A[18]), .ZN(n96) );
  AND2_X1 U73 ( .A1(A[5]), .A2(A[4]), .ZN(n114) );
  CLKBUF_X1 U74 ( .A(A[6]), .Z(n53) );
  AND2_X1 U75 ( .A1(n63), .A2(n94), .ZN(n49) );
  OR2_X1 U76 ( .A1(n87), .A2(n90), .ZN(n86) );
  AND2_X1 U77 ( .A1(A[16]), .A2(A[17]), .ZN(n50) );
  AND2_X1 U78 ( .A1(n45), .A2(n50), .ZN(n64) );
  XNOR2_X1 U79 ( .A(n92), .B(n93), .ZN(SUM[26]) );
  AND3_X1 U80 ( .A1(n45), .A2(n9), .A3(n43), .ZN(n51) );
  AND3_X1 U81 ( .A1(n9), .A2(n45), .A3(n43), .ZN(n65) );
  XOR2_X1 U82 ( .A(n52), .B(A[25]), .Z(SUM[25]) );
  AND2_X1 U83 ( .A1(A[24]), .A2(n89), .ZN(n52) );
  NOR2_X1 U84 ( .A1(n55), .A2(n56), .ZN(n102) );
  NAND4_X1 U85 ( .A1(A[3]), .A2(A[5]), .A3(A[6]), .A4(A[7]), .ZN(n55) );
  NAND3_X1 U86 ( .A1(A[4]), .A2(A[2]), .A3(A[9]), .ZN(n56) );
  NOR2_X1 U87 ( .A1(n96), .A2(n97), .ZN(n57) );
  AND2_X1 U88 ( .A1(A[7]), .A2(A[6]), .ZN(n115) );
  AND2_X1 U89 ( .A1(n101), .A2(n102), .ZN(n58) );
  INV_X1 U90 ( .A(n111), .ZN(n60) );
  AND2_X1 U91 ( .A1(n45), .A2(n85), .ZN(n61) );
  OR2_X1 U92 ( .A1(n30), .A2(n75), .ZN(n62) );
  NOR2_X1 U93 ( .A1(n110), .A2(n105), .ZN(n109) );
  AND2_X1 U94 ( .A1(n63), .A2(n94), .ZN(n85) );
  XNOR2_X1 U95 ( .A(n95), .B(n34), .ZN(SUM[23]) );
  NOR2_X1 U96 ( .A1(n30), .A2(n75), .ZN(n73) );
  NOR2_X1 U97 ( .A1(n24), .A2(n96), .ZN(n94) );
  INV_X1 U98 ( .A(n74), .ZN(n72) );
  AND2_X1 U99 ( .A1(n64), .A2(n98), .ZN(n67) );
  INV_X1 U100 ( .A(A[27]), .ZN(n91) );
  INV_X1 U101 ( .A(n33), .ZN(n106) );
  INV_X1 U102 ( .A(n74), .ZN(n112) );
  XNOR2_X1 U103 ( .A(n68), .B(n80), .ZN(SUM[30]) );
  OR2_X1 U104 ( .A1(n83), .A2(n82), .ZN(n68) );
  XOR2_X1 U105 ( .A(n64), .B(n98), .Z(SUM[18]) );
  XOR2_X1 U106 ( .A(n26), .B(n8), .Z(SUM[16]) );
  XOR2_X1 U107 ( .A(n77), .B(n6), .Z(SUM[6]) );
  XOR2_X1 U108 ( .A(n25), .B(n32), .Z(SUM[3]) );
  XOR2_X1 U109 ( .A(n18), .B(n20), .Z(SUM[4]) );
  XOR2_X1 U110 ( .A(n70), .B(n31), .Z(SUM[10]) );
  XOR2_X1 U111 ( .A(n89), .B(A[24]), .Z(SUM[24]) );
  XOR2_X1 U112 ( .A(n51), .B(n37), .Z(SUM[22]) );
  INV_X1 U113 ( .A(n100), .ZN(n98) );
  AND2_X1 U114 ( .A1(n79), .A2(n20), .ZN(n69) );
  INV_X1 U115 ( .A(A[26]), .ZN(n93) );
  INV_X1 U116 ( .A(A[28]), .ZN(n90) );
  INV_X1 U117 ( .A(n81), .ZN(n80) );
  INV_X1 U118 ( .A(A[30]), .ZN(n81) );
  AND3_X1 U119 ( .A1(n73), .A2(n35), .A3(A[8]), .ZN(n70) );
  INV_X1 U120 ( .A(n88), .ZN(n84) );
  INV_X1 U121 ( .A(A[29]), .ZN(n88) );
  INV_X1 U122 ( .A(A[11]), .ZN(n113) );
  INV_X1 U123 ( .A(A[8]), .ZN(n74) );
  INV_X1 U124 ( .A(n25), .ZN(SUM[2]) );
  NAND4_X1 U125 ( .A1(A[24]), .A2(A[25]), .A3(A[26]), .A4(A[27]), .ZN(n87) );
  INV_X1 U126 ( .A(A[19]), .ZN(n99) );
  INV_X1 U127 ( .A(A[18]), .ZN(n100) );
  NAND2_X1 U128 ( .A1(A[16]), .A2(A[17]), .ZN(n97) );
  XNOR2_X1 U129 ( .A(n66), .B(n91), .ZN(SUM[27]) );
  INV_X1 U130 ( .A(A[13]), .ZN(n111) );
  NAND2_X1 U131 ( .A1(n65), .A2(n37), .ZN(n95) );
  INV_X1 U132 ( .A(A[5]), .ZN(n116) );
  XNOR2_X1 U133 ( .A(n67), .B(n99), .ZN(SUM[19]) );
  NAND2_X1 U134 ( .A1(n114), .A2(n115), .ZN(n76) );
  NAND2_X1 U135 ( .A1(n58), .A2(n85), .ZN(n71) );
  NOR2_X1 U136 ( .A1(n103), .A2(n104), .ZN(n101) );
  INV_X1 U137 ( .A(A[12]), .ZN(n105) );
  NAND4_X1 U138 ( .A1(n112), .A2(n46), .A3(n31), .A4(n35), .ZN(n110) );
  NAND4_X1 U139 ( .A1(A[14]), .A2(A[15]), .A3(A[13]), .A4(A[10]), .ZN(n103) );
  XNOR2_X1 U140 ( .A(n5), .B(n16), .ZN(SUM[11]) );
  INV_X1 U141 ( .A(n69), .ZN(n78) );
  INV_X1 U142 ( .A(n58), .ZN(n83) );
  NAND3_X1 U143 ( .A1(n49), .A2(n42), .A3(n84), .ZN(n82) );
  NAND3_X1 U144 ( .A1(A[8]), .A2(A[11]), .A3(A[12]), .ZN(n104) );
  XNOR2_X1 U145 ( .A(n107), .B(n106), .ZN(SUM[15]) );
  INV_X1 U146 ( .A(A[14]), .ZN(n108) );
  INV_X1 U147 ( .A(n79), .ZN(n75) );
endmodule


module Fetch ( CLK, RST, ZERO_FLAG, PC_EXT, INS_IN, Bubble_in, HDU_INS_IN, 
        HDU_PC_IN, HDU_NPC_IN, PC_OUT, ADDR_OUT, NPC_OUT, INS_OUT );
  input [31:0] PC_EXT;
  input [31:0] INS_IN;
  input [31:0] HDU_INS_IN;
  input [31:0] HDU_PC_IN;
  input [31:0] HDU_NPC_IN;
  output [31:0] PC_OUT;
  output [31:0] ADDR_OUT;
  output [31:0] NPC_OUT;
  output [31:0] INS_OUT;
  input CLK, RST, ZERO_FLAG, Bubble_in;
  wire   n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, sig_RST, n26;
  wire   [31:0] sig_NPC;
  wire   [31:0] PC_MUX_OUT;
  wire   [31:0] sig_INS;

  mux21_NBIT32_0 NPC_or_NPC_HDU ( .A(PC_EXT), .B(HDU_NPC_IN), .S(Bubble_in), 
        .Z(sig_NPC) );
  mux21_NBIT32_5 PC_or_PC_HDU ( .A(ADDR_OUT), .B(HDU_PC_IN), .S(Bubble_in), 
        .Z(PC_MUX_OUT) );
  mux21_NBIT32_4 INS_or_HDU_INS ( .A(INS_IN), .B(HDU_INS_IN), .S(Bubble_in), 
        .Z(sig_INS) );
  regn_N32_0 PC ( .DIN(sig_NPC), .CLK(CLK), .EN(1'b1), .RST(RST), .DOUT({
        ADDR_OUT[31:28], n27, n28, ADDR_OUT[25:24], n29, n30, n31, 
        ADDR_OUT[20], n32, n33, n34, n35, n36, n37, n38, ADDR_OUT[12], n39, 
        n40, n41, n42, n43, n44, n45, n46, n47, n48, ADDR_OUT[1:0]}) );
  regn_N32_10 PC_reg ( .DIN(PC_MUX_OUT), .CLK(CLK), .EN(1'b1), .RST(sig_RST), 
        .DOUT(PC_OUT) );
  regn_N32_9 IR ( .DIN(sig_INS), .CLK(CLK), .EN(1'b1), .RST(sig_RST), .DOUT(
        INS_OUT) );
  Fetch_DW01_add_3 add_54 ( .A({ADDR_OUT[31:28], n27, n28, ADDR_OUT[25:24], 
        n29, n30, n31, ADDR_OUT[20], n32, n33, n34, n35, n36, n37, n38, 
        ADDR_OUT[12], n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
        ADDR_OUT[1:0]}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(NPC_OUT) );
  BUF_X1 U6 ( .A(n46), .Z(ADDR_OUT[4]) );
  CLKBUF_X1 U7 ( .A(n29), .Z(ADDR_OUT[23]) );
  CLKBUF_X1 U8 ( .A(n30), .Z(ADDR_OUT[22]) );
  CLKBUF_X1 U9 ( .A(n28), .Z(ADDR_OUT[26]) );
  CLKBUF_X1 U10 ( .A(n41), .Z(ADDR_OUT[9]) );
  CLKBUF_X1 U11 ( .A(n42), .Z(ADDR_OUT[8]) );
  CLKBUF_X1 U12 ( .A(n48), .Z(ADDR_OUT[2]) );
  CLKBUF_X1 U13 ( .A(n47), .Z(ADDR_OUT[3]) );
  CLKBUF_X1 U14 ( .A(n31), .Z(ADDR_OUT[21]) );
  CLKBUF_X1 U15 ( .A(n32), .Z(ADDR_OUT[19]) );
  CLKBUF_X1 U16 ( .A(n33), .Z(ADDR_OUT[18]) );
  CLKBUF_X1 U17 ( .A(n35), .Z(ADDR_OUT[16]) );
  CLKBUF_X1 U18 ( .A(n27), .Z(ADDR_OUT[27]) );
  CLKBUF_X1 U19 ( .A(n43), .Z(ADDR_OUT[7]) );
  NOR2_X1 U20 ( .A1(ZERO_FLAG), .A2(n26), .ZN(sig_RST) );
  CLKBUF_X1 U21 ( .A(n36), .Z(ADDR_OUT[15]) );
  CLKBUF_X1 U22 ( .A(n37), .Z(ADDR_OUT[14]) );
  CLKBUF_X1 U23 ( .A(n45), .Z(ADDR_OUT[5]) );
  CLKBUF_X1 U24 ( .A(n40), .Z(ADDR_OUT[10]) );
  CLKBUF_X1 U25 ( .A(n34), .Z(ADDR_OUT[17]) );
  CLKBUF_X1 U26 ( .A(n39), .Z(ADDR_OUT[11]) );
  CLKBUF_X1 U27 ( .A(n38), .Z(ADDR_OUT[13]) );
  CLKBUF_X1 U28 ( .A(n44), .Z(ADDR_OUT[6]) );
  INV_X1 U29 ( .A(RST), .ZN(n26) );
endmodule


module instruction_type ( INST_IN, Rtype, Itype, Jtype );
  input [31:0] INST_IN;
  output Rtype, Itype, Jtype;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n1, n2, n3, n4, n5,
         n6, n7, n8;

  OAI33_X1 U21 ( .A1(n5), .A2(INST_IN[29]), .A3(n2), .B1(n4), .B2(INST_IN[30]), 
        .B3(INST_IN[26]), .ZN(n17) );
  NOR2_X1 U1 ( .A1(n9), .A2(n10), .ZN(Rtype) );
  OAI22_X1 U2 ( .A1(n10), .A2(n5), .B1(n7), .B2(n4), .ZN(n16) );
  NOR2_X1 U3 ( .A1(n9), .A2(n6), .ZN(Jtype) );
  NAND4_X1 U4 ( .A1(n5), .A2(n4), .A3(n3), .A4(n1), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n6), .A2(n8), .ZN(n10) );
  INV_X1 U6 ( .A(n14), .ZN(n7) );
  INV_X1 U7 ( .A(n18), .ZN(n2) );
  OAI221_X1 U8 ( .B1(n7), .B2(INST_IN[30]), .C1(n3), .C2(INST_IN[26]), .A(n10), 
        .ZN(n18) );
  OAI211_X1 U9 ( .C1(INST_IN[31]), .C2(n11), .A(n12), .B(n13), .ZN(Itype) );
  NAND4_X1 U10 ( .A1(INST_IN[29]), .A2(INST_IN[28]), .A3(n14), .A4(n1), .ZN(
        n13) );
  NAND4_X1 U11 ( .A1(INST_IN[31]), .A2(INST_IN[27]), .A3(n15), .A4(INST_IN[26]), .ZN(n12) );
  AOI21_X1 U12 ( .B1(INST_IN[30]), .B2(n16), .A(n17), .ZN(n11) );
  NOR2_X1 U13 ( .A1(n8), .A2(INST_IN[27]), .ZN(n14) );
  NOR2_X1 U14 ( .A1(INST_IN[30]), .A2(INST_IN[28]), .ZN(n15) );
  INV_X1 U15 ( .A(INST_IN[30]), .ZN(n3) );
  INV_X1 U16 ( .A(INST_IN[28]), .ZN(n5) );
  INV_X1 U17 ( .A(INST_IN[29]), .ZN(n4) );
  INV_X1 U18 ( .A(INST_IN[26]), .ZN(n8) );
  INV_X1 U19 ( .A(INST_IN[31]), .ZN(n1) );
  INV_X1 U20 ( .A(INST_IN[27]), .ZN(n6) );
endmodule


module instruction_decomposition ( INST_IN, Rtype, Itype, Jtype, ADD_RS1, 
        ADD_RS2, ADD_WR, IMM );
  input [31:0] INST_IN;
  output [4:0] ADD_RS1;
  output [4:0] ADD_RS2;
  output [4:0] ADD_WR;
  output [31:0] IMM;
  input Rtype, Itype, Jtype;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n1, n2,
         \IMM[31] , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20;
  assign IMM[25] = \IMM[31] ;
  assign IMM[26] = \IMM[31] ;
  assign IMM[27] = \IMM[31] ;
  assign IMM[28] = \IMM[31] ;
  assign IMM[29] = \IMM[31] ;
  assign IMM[30] = \IMM[31] ;
  assign IMM[31] = \IMM[31] ;

  NAND3_X1 U72 ( .A1(INST_IN[29]), .A2(INST_IN[27]), .A3(INST_IN[31]), .ZN(n31) );
  NAND3_X1 U73 ( .A1(INST_IN[26]), .A2(Itype), .A3(n32), .ZN(n30) );
  INV_X1 U2 ( .A(Rtype), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n28), .A2(Jtype), .ZN(n24) );
  INV_X1 U4 ( .A(n27), .ZN(n2) );
  OAI21_X1 U5 ( .B1(Itype), .B2(Jtype), .A(n4), .ZN(n27) );
  NOR2_X1 U6 ( .A1(Rtype), .A2(Itype), .ZN(n28) );
  NOR2_X1 U7 ( .A1(n28), .A2(n7), .ZN(ADD_RS1[3]) );
  NOR2_X1 U8 ( .A1(n1), .A2(n12), .ZN(ADD_RS2[3]) );
  NOR2_X1 U9 ( .A1(n28), .A2(n10), .ZN(ADD_RS1[0]) );
  NOR2_X1 U10 ( .A1(n1), .A2(n15), .ZN(ADD_RS2[0]) );
  NOR2_X1 U11 ( .A1(n1), .A2(n11), .ZN(ADD_RS2[4]) );
  OR2_X1 U12 ( .A1(n26), .A2(n16), .ZN(n25) );
  NOR2_X1 U13 ( .A1(n28), .A2(n8), .ZN(ADD_RS1[2]) );
  NOR2_X1 U14 ( .A1(n1), .A2(n13), .ZN(ADD_RS2[2]) );
  NOR2_X1 U15 ( .A1(n28), .A2(n9), .ZN(ADD_RS1[1]) );
  NOR2_X1 U16 ( .A1(n1), .A2(n14), .ZN(ADD_RS2[1]) );
  NAND2_X1 U17 ( .A1(Itype), .A2(n4), .ZN(n26) );
  INV_X1 U18 ( .A(Itype), .ZN(n5) );
  AND2_X1 U19 ( .A1(INST_IN[0]), .A2(n2), .ZN(IMM[0]) );
  AND2_X1 U20 ( .A1(INST_IN[1]), .A2(n2), .ZN(IMM[1]) );
  AND2_X1 U21 ( .A1(INST_IN[2]), .A2(n2), .ZN(IMM[2]) );
  AND2_X1 U22 ( .A1(INST_IN[3]), .A2(n2), .ZN(IMM[3]) );
  AND2_X1 U23 ( .A1(INST_IN[4]), .A2(n2), .ZN(IMM[4]) );
  AND2_X1 U24 ( .A1(INST_IN[5]), .A2(n2), .ZN(IMM[5]) );
  AND2_X1 U25 ( .A1(INST_IN[6]), .A2(n2), .ZN(IMM[6]) );
  AND2_X1 U26 ( .A1(INST_IN[7]), .A2(n2), .ZN(IMM[7]) );
  AND2_X1 U27 ( .A1(INST_IN[8]), .A2(n2), .ZN(IMM[8]) );
  AND2_X1 U28 ( .A1(INST_IN[9]), .A2(n2), .ZN(IMM[9]) );
  AND2_X1 U29 ( .A1(INST_IN[10]), .A2(n2), .ZN(IMM[10]) );
  NOR2_X1 U30 ( .A1(n27), .A2(n20), .ZN(IMM[11]) );
  NOR2_X1 U31 ( .A1(n27), .A2(n19), .ZN(IMM[12]) );
  NOR2_X1 U32 ( .A1(n27), .A2(n18), .ZN(IMM[13]) );
  NOR2_X1 U33 ( .A1(n27), .A2(n17), .ZN(IMM[14]) );
  NOR2_X1 U34 ( .A1(n27), .A2(n16), .ZN(IMM[15]) );
  OAI21_X1 U35 ( .B1(n24), .B2(n15), .A(n25), .ZN(IMM[16]) );
  OAI21_X1 U36 ( .B1(n24), .B2(n14), .A(n25), .ZN(IMM[17]) );
  OAI21_X1 U37 ( .B1(n24), .B2(n13), .A(n25), .ZN(IMM[18]) );
  OAI21_X1 U38 ( .B1(n24), .B2(n12), .A(n25), .ZN(IMM[19]) );
  OAI21_X1 U39 ( .B1(n24), .B2(n11), .A(n25), .ZN(IMM[20]) );
  OAI21_X1 U40 ( .B1(n24), .B2(n10), .A(n25), .ZN(IMM[21]) );
  OAI21_X1 U41 ( .B1(n24), .B2(n9), .A(n25), .ZN(IMM[22]) );
  OAI21_X1 U42 ( .B1(n24), .B2(n8), .A(n25), .ZN(IMM[23]) );
  OAI21_X1 U43 ( .B1(n24), .B2(n7), .A(n25), .ZN(IMM[24]) );
  OAI221_X1 U44 ( .B1(n26), .B2(n15), .C1(n20), .C2(n4), .A(n24), .ZN(
        ADD_WR[0]) );
  OAI221_X1 U45 ( .B1(n26), .B2(n14), .C1(n19), .C2(n4), .A(n24), .ZN(
        ADD_WR[1]) );
  OAI221_X1 U46 ( .B1(n26), .B2(n13), .C1(n18), .C2(n4), .A(n24), .ZN(
        ADD_WR[2]) );
  OAI221_X1 U47 ( .B1(n26), .B2(n12), .C1(n17), .C2(n4), .A(n24), .ZN(
        ADD_WR[3]) );
  OAI221_X1 U48 ( .B1(n26), .B2(n11), .C1(n16), .C2(n4), .A(n24), .ZN(
        ADD_WR[4]) );
  NOR2_X1 U49 ( .A1(n28), .A2(n6), .ZN(ADD_RS1[4]) );
  INV_X1 U50 ( .A(INST_IN[25]), .ZN(n6) );
  INV_X1 U51 ( .A(n29), .ZN(n1) );
  OAI21_X1 U52 ( .B1(n30), .B2(n31), .A(n4), .ZN(n29) );
  INV_X1 U53 ( .A(INST_IN[15]), .ZN(n16) );
  INV_X1 U54 ( .A(INST_IN[16]), .ZN(n15) );
  INV_X1 U55 ( .A(INST_IN[17]), .ZN(n14) );
  INV_X1 U56 ( .A(INST_IN[19]), .ZN(n12) );
  INV_X1 U57 ( .A(INST_IN[18]), .ZN(n13) );
  INV_X1 U58 ( .A(INST_IN[20]), .ZN(n11) );
  NOR2_X1 U59 ( .A1(INST_IN[30]), .A2(INST_IN[28]), .ZN(n32) );
  INV_X1 U60 ( .A(n21), .ZN(\IMM[31] ) );
  OAI21_X1 U61 ( .B1(n22), .B2(n23), .A(n4), .ZN(n21) );
  AND3_X1 U62 ( .A1(Jtype), .A2(n5), .A3(INST_IN[25]), .ZN(n22) );
  NOR2_X1 U63 ( .A1(n16), .A2(n5), .ZN(n23) );
  INV_X1 U64 ( .A(INST_IN[21]), .ZN(n10) );
  INV_X1 U65 ( .A(INST_IN[24]), .ZN(n7) );
  INV_X1 U66 ( .A(INST_IN[22]), .ZN(n9) );
  INV_X1 U67 ( .A(INST_IN[23]), .ZN(n8) );
  INV_X1 U68 ( .A(INST_IN[11]), .ZN(n20) );
  INV_X1 U69 ( .A(INST_IN[12]), .ZN(n19) );
  INV_X1 U70 ( .A(INST_IN[13]), .ZN(n18) );
  INV_X1 U71 ( .A(INST_IN[14]), .ZN(n17) );
endmodule


module regn_N32_8 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n68, n69, n70;

  DFFR_X1 \DOUT_reg[31]  ( .D(n36), .CK(CLK), .RN(n3), .Q(DOUT[31]) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n37), .CK(CLK), .RN(n3), .Q(DOUT[30]) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n38), .CK(CLK), .RN(n3), .Q(DOUT[29]) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n39), .CK(CLK), .RN(n3), .Q(DOUT[28]) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n40), .CK(CLK), .RN(n3), .Q(DOUT[27]) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n41), .CK(CLK), .RN(n3), .Q(DOUT[26]) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n42), .CK(CLK), .RN(n3), .Q(DOUT[25]) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n43), .CK(CLK), .RN(n3), .Q(DOUT[24]) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n44), .CK(CLK), .RN(n2), .Q(DOUT[23]) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n45), .CK(CLK), .RN(n2), .Q(DOUT[22]) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n46), .CK(CLK), .RN(n2), .Q(DOUT[21]) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n47), .CK(CLK), .RN(n2), .Q(DOUT[20]) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n48), .CK(CLK), .RN(n2), .Q(DOUT[19]) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n49), .CK(CLK), .RN(n2), .Q(DOUT[18]) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n50), .CK(CLK), .RN(n2), .Q(DOUT[17]) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n51), .CK(CLK), .RN(n2), .Q(DOUT[16]) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n52), .CK(CLK), .RN(n2), .Q(DOUT[15]) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n53), .CK(CLK), .RN(n2), .Q(DOUT[14]) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n54), .CK(CLK), .RN(n2), .Q(DOUT[13]) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n55), .CK(CLK), .RN(n2), .Q(DOUT[12]) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n56), .CK(CLK), .RN(n1), .Q(DOUT[11]) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n57), .CK(CLK), .RN(n1), .Q(DOUT[10]) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n58), .CK(CLK), .RN(n1), .Q(DOUT[9]) );
  DFFR_X1 \DOUT_reg[8]  ( .D(n59), .CK(CLK), .RN(n1), .Q(DOUT[8]) );
  DFFR_X1 \DOUT_reg[7]  ( .D(n60), .CK(CLK), .RN(n1), .Q(DOUT[7]) );
  DFFR_X1 \DOUT_reg[6]  ( .D(n61), .CK(CLK), .RN(n1), .Q(DOUT[6]) );
  DFFR_X1 \DOUT_reg[5]  ( .D(n62), .CK(CLK), .RN(n1), .Q(DOUT[5]) );
  DFFR_X1 \DOUT_reg[4]  ( .D(n63), .CK(CLK), .RN(n1), .Q(DOUT[4]) );
  DFFR_X1 \DOUT_reg[3]  ( .D(n64), .CK(CLK), .RN(n1), .Q(DOUT[3]) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n68), .CK(CLK), .RN(n1), .Q(DOUT[2]) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n69), .CK(CLK), .RN(n1), .Q(DOUT[1]) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n70), .CK(CLK), .RN(n1), .Q(DOUT[0]) );
  BUF_X1 U2 ( .A(RST), .Z(n1) );
  BUF_X1 U3 ( .A(RST), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n3) );
  MUX2_X1 U5 ( .A(DOUT[0]), .B(DIN[0]), .S(EN), .Z(n70) );
  MUX2_X1 U6 ( .A(DOUT[1]), .B(DIN[1]), .S(EN), .Z(n69) );
  MUX2_X1 U7 ( .A(DOUT[2]), .B(DIN[2]), .S(EN), .Z(n68) );
  MUX2_X1 U8 ( .A(DOUT[3]), .B(DIN[3]), .S(EN), .Z(n64) );
  MUX2_X1 U9 ( .A(DOUT[4]), .B(DIN[4]), .S(EN), .Z(n63) );
  MUX2_X1 U10 ( .A(DOUT[5]), .B(DIN[5]), .S(EN), .Z(n62) );
  MUX2_X1 U11 ( .A(DOUT[6]), .B(DIN[6]), .S(EN), .Z(n61) );
  MUX2_X1 U12 ( .A(DOUT[7]), .B(DIN[7]), .S(EN), .Z(n60) );
  MUX2_X1 U13 ( .A(DOUT[8]), .B(DIN[8]), .S(EN), .Z(n59) );
  MUX2_X1 U14 ( .A(DOUT[9]), .B(DIN[9]), .S(EN), .Z(n58) );
  MUX2_X1 U15 ( .A(DOUT[10]), .B(DIN[10]), .S(EN), .Z(n57) );
  MUX2_X1 U16 ( .A(DOUT[11]), .B(DIN[11]), .S(EN), .Z(n56) );
  MUX2_X1 U17 ( .A(DOUT[12]), .B(DIN[12]), .S(EN), .Z(n55) );
  MUX2_X1 U18 ( .A(DOUT[13]), .B(DIN[13]), .S(EN), .Z(n54) );
  MUX2_X1 U19 ( .A(DOUT[14]), .B(DIN[14]), .S(EN), .Z(n53) );
  MUX2_X1 U20 ( .A(DOUT[15]), .B(DIN[15]), .S(EN), .Z(n52) );
  MUX2_X1 U21 ( .A(DOUT[16]), .B(DIN[16]), .S(EN), .Z(n51) );
  MUX2_X1 U22 ( .A(DOUT[17]), .B(DIN[17]), .S(EN), .Z(n50) );
  MUX2_X1 U23 ( .A(DOUT[18]), .B(DIN[18]), .S(EN), .Z(n49) );
  MUX2_X1 U24 ( .A(DOUT[19]), .B(DIN[19]), .S(EN), .Z(n48) );
  MUX2_X1 U25 ( .A(DOUT[20]), .B(DIN[20]), .S(EN), .Z(n47) );
  MUX2_X1 U26 ( .A(DOUT[21]), .B(DIN[21]), .S(EN), .Z(n46) );
  MUX2_X1 U27 ( .A(DOUT[22]), .B(DIN[22]), .S(EN), .Z(n45) );
  MUX2_X1 U28 ( .A(DOUT[23]), .B(DIN[23]), .S(EN), .Z(n44) );
  MUX2_X1 U29 ( .A(DOUT[24]), .B(DIN[24]), .S(EN), .Z(n43) );
  MUX2_X1 U30 ( .A(DOUT[25]), .B(DIN[25]), .S(EN), .Z(n42) );
  MUX2_X1 U31 ( .A(DOUT[26]), .B(DIN[26]), .S(EN), .Z(n41) );
  MUX2_X1 U32 ( .A(DOUT[27]), .B(DIN[27]), .S(EN), .Z(n40) );
  MUX2_X1 U33 ( .A(DOUT[28]), .B(DIN[28]), .S(EN), .Z(n39) );
  MUX2_X1 U34 ( .A(DOUT[29]), .B(DIN[29]), .S(EN), .Z(n38) );
  MUX2_X1 U35 ( .A(DOUT[30]), .B(DIN[30]), .S(EN), .Z(n37) );
  MUX2_X1 U36 ( .A(DOUT[31]), .B(DIN[31]), .S(EN), .Z(n36) );
endmodule


module regn_N32_7 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n68, n69, n70;

  DFFR_X1 \DOUT_reg[31]  ( .D(n36), .CK(CLK), .RN(n3), .Q(DOUT[31]) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n37), .CK(CLK), .RN(n3), .Q(DOUT[30]) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n38), .CK(CLK), .RN(n3), .Q(DOUT[29]) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n39), .CK(CLK), .RN(n3), .Q(DOUT[28]) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n40), .CK(CLK), .RN(n3), .Q(DOUT[27]) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n41), .CK(CLK), .RN(n3), .Q(DOUT[26]) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n42), .CK(CLK), .RN(n3), .Q(DOUT[25]) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n43), .CK(CLK), .RN(n3), .Q(DOUT[24]) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n44), .CK(CLK), .RN(n2), .Q(DOUT[23]) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n45), .CK(CLK), .RN(n2), .Q(DOUT[22]) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n46), .CK(CLK), .RN(n2), .Q(DOUT[21]) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n47), .CK(CLK), .RN(n2), .Q(DOUT[20]) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n48), .CK(CLK), .RN(n2), .Q(DOUT[19]) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n49), .CK(CLK), .RN(n2), .Q(DOUT[18]) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n50), .CK(CLK), .RN(n2), .Q(DOUT[17]) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n51), .CK(CLK), .RN(n2), .Q(DOUT[16]) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n52), .CK(CLK), .RN(n2), .Q(DOUT[15]) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n53), .CK(CLK), .RN(n2), .Q(DOUT[14]) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n54), .CK(CLK), .RN(n2), .Q(DOUT[13]) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n55), .CK(CLK), .RN(n2), .Q(DOUT[12]) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n56), .CK(CLK), .RN(n1), .Q(DOUT[11]) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n57), .CK(CLK), .RN(n1), .Q(DOUT[10]) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n58), .CK(CLK), .RN(n1), .Q(DOUT[9]) );
  DFFR_X1 \DOUT_reg[8]  ( .D(n59), .CK(CLK), .RN(n1), .Q(DOUT[8]) );
  DFFR_X1 \DOUT_reg[7]  ( .D(n60), .CK(CLK), .RN(n1), .Q(DOUT[7]) );
  DFFR_X1 \DOUT_reg[6]  ( .D(n61), .CK(CLK), .RN(n1), .Q(DOUT[6]) );
  DFFR_X1 \DOUT_reg[5]  ( .D(n62), .CK(CLK), .RN(n1), .Q(DOUT[5]) );
  DFFR_X1 \DOUT_reg[4]  ( .D(n63), .CK(CLK), .RN(n1), .Q(DOUT[4]) );
  DFFR_X1 \DOUT_reg[3]  ( .D(n64), .CK(CLK), .RN(n1), .Q(DOUT[3]) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n68), .CK(CLK), .RN(n1), .Q(DOUT[2]) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n69), .CK(CLK), .RN(n1), .Q(DOUT[1]) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n70), .CK(CLK), .RN(n1), .Q(DOUT[0]) );
  BUF_X1 U2 ( .A(RST), .Z(n1) );
  BUF_X1 U3 ( .A(RST), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n3) );
  MUX2_X1 U5 ( .A(DOUT[0]), .B(DIN[0]), .S(EN), .Z(n70) );
  MUX2_X1 U6 ( .A(DOUT[1]), .B(DIN[1]), .S(EN), .Z(n69) );
  MUX2_X1 U7 ( .A(DOUT[2]), .B(DIN[2]), .S(EN), .Z(n68) );
  MUX2_X1 U8 ( .A(DOUT[3]), .B(DIN[3]), .S(EN), .Z(n64) );
  MUX2_X1 U9 ( .A(DOUT[4]), .B(DIN[4]), .S(EN), .Z(n63) );
  MUX2_X1 U10 ( .A(DOUT[5]), .B(DIN[5]), .S(EN), .Z(n62) );
  MUX2_X1 U11 ( .A(DOUT[6]), .B(DIN[6]), .S(EN), .Z(n61) );
  MUX2_X1 U12 ( .A(DOUT[7]), .B(DIN[7]), .S(EN), .Z(n60) );
  MUX2_X1 U13 ( .A(DOUT[8]), .B(DIN[8]), .S(EN), .Z(n59) );
  MUX2_X1 U14 ( .A(DOUT[9]), .B(DIN[9]), .S(EN), .Z(n58) );
  MUX2_X1 U15 ( .A(DOUT[10]), .B(DIN[10]), .S(EN), .Z(n57) );
  MUX2_X1 U16 ( .A(DOUT[11]), .B(DIN[11]), .S(EN), .Z(n56) );
  MUX2_X1 U17 ( .A(DOUT[12]), .B(DIN[12]), .S(EN), .Z(n55) );
  MUX2_X1 U18 ( .A(DOUT[13]), .B(DIN[13]), .S(EN), .Z(n54) );
  MUX2_X1 U19 ( .A(DOUT[14]), .B(DIN[14]), .S(EN), .Z(n53) );
  MUX2_X1 U20 ( .A(DOUT[15]), .B(DIN[15]), .S(EN), .Z(n52) );
  MUX2_X1 U21 ( .A(DOUT[16]), .B(DIN[16]), .S(EN), .Z(n51) );
  MUX2_X1 U22 ( .A(DOUT[17]), .B(DIN[17]), .S(EN), .Z(n50) );
  MUX2_X1 U23 ( .A(DOUT[18]), .B(DIN[18]), .S(EN), .Z(n49) );
  MUX2_X1 U24 ( .A(DOUT[19]), .B(DIN[19]), .S(EN), .Z(n48) );
  MUX2_X1 U25 ( .A(DOUT[20]), .B(DIN[20]), .S(EN), .Z(n47) );
  MUX2_X1 U26 ( .A(DOUT[21]), .B(DIN[21]), .S(EN), .Z(n46) );
  MUX2_X1 U27 ( .A(DOUT[22]), .B(DIN[22]), .S(EN), .Z(n45) );
  MUX2_X1 U28 ( .A(DOUT[23]), .B(DIN[23]), .S(EN), .Z(n44) );
  MUX2_X1 U29 ( .A(DOUT[24]), .B(DIN[24]), .S(EN), .Z(n43) );
  MUX2_X1 U30 ( .A(DOUT[25]), .B(DIN[25]), .S(EN), .Z(n42) );
  MUX2_X1 U31 ( .A(DOUT[26]), .B(DIN[26]), .S(EN), .Z(n41) );
  MUX2_X1 U32 ( .A(DOUT[27]), .B(DIN[27]), .S(EN), .Z(n40) );
  MUX2_X1 U33 ( .A(DOUT[28]), .B(DIN[28]), .S(EN), .Z(n39) );
  MUX2_X1 U34 ( .A(DOUT[29]), .B(DIN[29]), .S(EN), .Z(n38) );
  MUX2_X1 U35 ( .A(DOUT[30]), .B(DIN[30]), .S(EN), .Z(n37) );
  MUX2_X1 U36 ( .A(DOUT[31]), .B(DIN[31]), .S(EN), .Z(n36) );
endmodule


module regn_N5_0 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n11, n12, n13, n14, n15;

  DFFR_X1 \DOUT_reg[4]  ( .D(n15), .CK(CLK), .RN(RST), .Q(DOUT[4]) );
  DFFR_X1 \DOUT_reg[3]  ( .D(n14), .CK(CLK), .RN(RST), .Q(DOUT[3]) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n13), .CK(CLK), .RN(RST), .Q(DOUT[2]) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n12), .CK(CLK), .RN(RST), .Q(DOUT[1]) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n11), .CK(CLK), .RN(RST), .Q(DOUT[0]) );
  MUX2_X1 U2 ( .A(DOUT[0]), .B(DIN[0]), .S(EN), .Z(n11) );
  MUX2_X1 U3 ( .A(DOUT[1]), .B(DIN[1]), .S(EN), .Z(n12) );
  MUX2_X1 U4 ( .A(DOUT[2]), .B(DIN[2]), .S(EN), .Z(n13) );
  MUX2_X1 U5 ( .A(DOUT[3]), .B(DIN[3]), .S(EN), .Z(n14) );
  MUX2_X1 U6 ( .A(DOUT[4]), .B(DIN[4]), .S(EN), .Z(n15) );
endmodule


module regn_N5_4 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n6, n7, n8, n9, n10;

  DFFR_X1 \DOUT_reg[4]  ( .D(n6), .CK(CLK), .RN(RST), .Q(DOUT[4]) );
  DFFR_X1 \DOUT_reg[3]  ( .D(n7), .CK(CLK), .RN(RST), .Q(DOUT[3]) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n8), .CK(CLK), .RN(RST), .Q(DOUT[2]) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n9), .CK(CLK), .RN(RST), .Q(DOUT[1]) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n10), .CK(CLK), .RN(RST), .Q(DOUT[0]) );
  MUX2_X1 U2 ( .A(DOUT[0]), .B(DIN[0]), .S(EN), .Z(n10) );
  MUX2_X1 U3 ( .A(DOUT[1]), .B(DIN[1]), .S(EN), .Z(n9) );
  MUX2_X1 U4 ( .A(DOUT[2]), .B(DIN[2]), .S(EN), .Z(n8) );
  MUX2_X1 U5 ( .A(DOUT[3]), .B(DIN[3]), .S(EN), .Z(n7) );
  MUX2_X1 U6 ( .A(DOUT[4]), .B(DIN[4]), .S(EN), .Z(n6) );
endmodule


module regn_N5_3 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n6, n7, n8, n9, n10;

  DFFR_X1 \DOUT_reg[4]  ( .D(n6), .CK(CLK), .RN(RST), .Q(DOUT[4]) );
  DFFR_X1 \DOUT_reg[3]  ( .D(n7), .CK(CLK), .RN(RST), .Q(DOUT[3]) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n8), .CK(CLK), .RN(RST), .Q(DOUT[2]) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n9), .CK(CLK), .RN(RST), .Q(DOUT[1]) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n10), .CK(CLK), .RN(RST), .Q(DOUT[0]) );
  MUX2_X1 U2 ( .A(DOUT[0]), .B(DIN[0]), .S(EN), .Z(n10) );
  MUX2_X1 U3 ( .A(DOUT[1]), .B(DIN[1]), .S(EN), .Z(n9) );
  MUX2_X1 U4 ( .A(DOUT[2]), .B(DIN[2]), .S(EN), .Z(n8) );
  MUX2_X1 U5 ( .A(DOUT[3]), .B(DIN[3]), .S(EN), .Z(n7) );
  MUX2_X1 U6 ( .A(DOUT[4]), .B(DIN[4]), .S(EN), .Z(n6) );
endmodule


module register_file_NBIT_ADD5_NBIT_DATA32 ( CLK, RST, ENABLE, RD1, RD2, WR, 
        ADD_WR, ADD_RS1, ADD_RS2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RST, ENABLE, RD1, RD2, WR;
  wire   n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605;

  DFFR_X1 \REGISTERS_reg[10][31]  ( .D(n3430), .CK(CLK), .RN(n434), .Q(n3869)
         );
  DFFR_X1 \REGISTERS_reg[10][30]  ( .D(n3429), .CK(CLK), .RN(n434), .Q(n3868)
         );
  DFFR_X1 \REGISTERS_reg[10][29]  ( .D(n3428), .CK(CLK), .RN(n434), .Q(n3867)
         );
  DFFR_X1 \REGISTERS_reg[10][28]  ( .D(n3427), .CK(CLK), .RN(n434), .Q(n3866)
         );
  DFFR_X1 \REGISTERS_reg[10][27]  ( .D(n3426), .CK(CLK), .RN(n434), .Q(n3865)
         );
  DFFR_X1 \REGISTERS_reg[10][26]  ( .D(n3425), .CK(CLK), .RN(n434), .Q(n3864)
         );
  DFFR_X1 \REGISTERS_reg[10][25]  ( .D(n3424), .CK(CLK), .RN(n434), .Q(n3863)
         );
  DFFR_X1 \REGISTERS_reg[10][24]  ( .D(n3423), .CK(CLK), .RN(n434), .Q(n3862)
         );
  DFFR_X1 \REGISTERS_reg[10][23]  ( .D(n3422), .CK(CLK), .RN(n434), .Q(n3861)
         );
  DFFR_X1 \REGISTERS_reg[10][22]  ( .D(n3421), .CK(CLK), .RN(n434), .Q(n3860)
         );
  DFFR_X1 \REGISTERS_reg[10][21]  ( .D(n3420), .CK(CLK), .RN(n434), .Q(n3859)
         );
  DFFR_X1 \REGISTERS_reg[10][20]  ( .D(n3419), .CK(CLK), .RN(n434), .Q(n3858)
         );
  DFFR_X1 \REGISTERS_reg[10][19]  ( .D(n3418), .CK(CLK), .RN(n435), .Q(n3857)
         );
  DFFR_X1 \REGISTERS_reg[10][18]  ( .D(n3417), .CK(CLK), .RN(n435), .Q(n3856)
         );
  DFFR_X1 \REGISTERS_reg[10][17]  ( .D(n3416), .CK(CLK), .RN(n435), .Q(n3855)
         );
  DFFR_X1 \REGISTERS_reg[10][16]  ( .D(n3415), .CK(CLK), .RN(n435), .Q(n3854)
         );
  DFFR_X1 \REGISTERS_reg[10][15]  ( .D(n3414), .CK(CLK), .RN(n435), .Q(n3853)
         );
  DFFR_X1 \REGISTERS_reg[10][14]  ( .D(n3413), .CK(CLK), .RN(n435), .Q(n3852)
         );
  DFFR_X1 \REGISTERS_reg[10][13]  ( .D(n3412), .CK(CLK), .RN(n435), .Q(n3851)
         );
  DFFR_X1 \REGISTERS_reg[10][12]  ( .D(n3411), .CK(CLK), .RN(n435), .Q(n3850)
         );
  DFFR_X1 \REGISTERS_reg[10][11]  ( .D(n3410), .CK(CLK), .RN(n435), .Q(n3849)
         );
  DFFR_X1 \REGISTERS_reg[10][10]  ( .D(n3409), .CK(CLK), .RN(n435), .Q(n3848)
         );
  DFFR_X1 \REGISTERS_reg[10][9]  ( .D(n3408), .CK(CLK), .RN(n435), .Q(n3847)
         );
  DFFR_X1 \REGISTERS_reg[10][8]  ( .D(n3407), .CK(CLK), .RN(n435), .Q(n3846)
         );
  DFFR_X1 \REGISTERS_reg[10][7]  ( .D(n3406), .CK(CLK), .RN(n436), .Q(n3845)
         );
  DFFR_X1 \REGISTERS_reg[10][6]  ( .D(n3405), .CK(CLK), .RN(n436), .Q(n3844)
         );
  DFFR_X1 \REGISTERS_reg[10][5]  ( .D(n3404), .CK(CLK), .RN(n436), .Q(n3843)
         );
  DFFR_X1 \REGISTERS_reg[10][4]  ( .D(n3403), .CK(CLK), .RN(n436), .Q(n3842)
         );
  DFFR_X1 \REGISTERS_reg[10][3]  ( .D(n3402), .CK(CLK), .RN(n436), .Q(n3841)
         );
  DFFR_X1 \REGISTERS_reg[10][2]  ( .D(n3401), .CK(CLK), .RN(n436), .Q(n3840)
         );
  DFFR_X1 \REGISTERS_reg[10][1]  ( .D(n3400), .CK(CLK), .RN(n436), .Q(n3839)
         );
  DFFR_X1 \REGISTERS_reg[10][0]  ( .D(n3399), .CK(CLK), .RN(n436), .Q(n3838)
         );
  DFFR_X1 \REGISTERS_reg[11][31]  ( .D(n3398), .CK(CLK), .RN(n436), .Q(n3837)
         );
  DFFR_X1 \REGISTERS_reg[11][30]  ( .D(n3397), .CK(CLK), .RN(n436), .Q(n3836)
         );
  DFFR_X1 \REGISTERS_reg[11][29]  ( .D(n3396), .CK(CLK), .RN(n436), .Q(n3835)
         );
  DFFR_X1 \REGISTERS_reg[11][28]  ( .D(n3395), .CK(CLK), .RN(n436), .Q(n3834)
         );
  DFFR_X1 \REGISTERS_reg[11][27]  ( .D(n3394), .CK(CLK), .RN(n437), .Q(n3833)
         );
  DFFR_X1 \REGISTERS_reg[11][26]  ( .D(n3393), .CK(CLK), .RN(n437), .Q(n3832)
         );
  DFFR_X1 \REGISTERS_reg[11][25]  ( .D(n3392), .CK(CLK), .RN(n437), .Q(n3831)
         );
  DFFR_X1 \REGISTERS_reg[11][24]  ( .D(n3391), .CK(CLK), .RN(n437), .Q(n3830)
         );
  DFFR_X1 \REGISTERS_reg[11][23]  ( .D(n3390), .CK(CLK), .RN(n437), .Q(n3829)
         );
  DFFR_X1 \REGISTERS_reg[11][22]  ( .D(n3389), .CK(CLK), .RN(n437), .Q(n3828)
         );
  DFFR_X1 \REGISTERS_reg[11][21]  ( .D(n3388), .CK(CLK), .RN(n437), .Q(n3827)
         );
  DFFR_X1 \REGISTERS_reg[11][20]  ( .D(n3387), .CK(CLK), .RN(n437), .Q(n3826)
         );
  DFFR_X1 \REGISTERS_reg[11][19]  ( .D(n3386), .CK(CLK), .RN(n437), .Q(n3825)
         );
  DFFR_X1 \REGISTERS_reg[11][18]  ( .D(n3385), .CK(CLK), .RN(n437), .Q(n3824)
         );
  DFFR_X1 \REGISTERS_reg[11][17]  ( .D(n3384), .CK(CLK), .RN(n437), .Q(n3823)
         );
  DFFR_X1 \REGISTERS_reg[11][16]  ( .D(n3383), .CK(CLK), .RN(n437), .Q(n3822)
         );
  DFFR_X1 \REGISTERS_reg[11][15]  ( .D(n3382), .CK(CLK), .RN(n438), .Q(n3821)
         );
  DFFR_X1 \REGISTERS_reg[11][14]  ( .D(n3381), .CK(CLK), .RN(n438), .Q(n3820)
         );
  DFFR_X1 \REGISTERS_reg[11][13]  ( .D(n3380), .CK(CLK), .RN(n438), .Q(n3819)
         );
  DFFR_X1 \REGISTERS_reg[11][12]  ( .D(n3379), .CK(CLK), .RN(n438), .Q(n3818)
         );
  DFFR_X1 \REGISTERS_reg[11][11]  ( .D(n3378), .CK(CLK), .RN(n438), .Q(n3817)
         );
  DFFR_X1 \REGISTERS_reg[11][10]  ( .D(n3377), .CK(CLK), .RN(n438), .Q(n3816)
         );
  DFFR_X1 \REGISTERS_reg[11][9]  ( .D(n3376), .CK(CLK), .RN(n438), .Q(n3815)
         );
  DFFR_X1 \REGISTERS_reg[11][8]  ( .D(n3375), .CK(CLK), .RN(n438), .Q(n3814)
         );
  DFFR_X1 \REGISTERS_reg[11][7]  ( .D(n3374), .CK(CLK), .RN(n438), .Q(n3813)
         );
  DFFR_X1 \REGISTERS_reg[11][6]  ( .D(n3373), .CK(CLK), .RN(n438), .Q(n3812)
         );
  DFFR_X1 \REGISTERS_reg[11][5]  ( .D(n3372), .CK(CLK), .RN(n438), .Q(n3811)
         );
  DFFR_X1 \REGISTERS_reg[11][4]  ( .D(n3371), .CK(CLK), .RN(n438), .Q(n3810)
         );
  DFFR_X1 \REGISTERS_reg[11][3]  ( .D(n3370), .CK(CLK), .RN(n439), .Q(n3809)
         );
  DFFR_X1 \REGISTERS_reg[11][2]  ( .D(n3369), .CK(CLK), .RN(n439), .Q(n3808)
         );
  DFFR_X1 \REGISTERS_reg[11][1]  ( .D(n3368), .CK(CLK), .RN(n439), .Q(n3807)
         );
  DFFR_X1 \REGISTERS_reg[11][0]  ( .D(n3367), .CK(CLK), .RN(n439), .Q(n3806)
         );
  DFFR_X1 \REGISTERS_reg[14][31]  ( .D(n3366), .CK(CLK), .RN(n444), .Q(n3741)
         );
  DFFR_X1 \REGISTERS_reg[14][30]  ( .D(n3365), .CK(CLK), .RN(n444), .Q(n3740)
         );
  DFFR_X1 \REGISTERS_reg[14][29]  ( .D(n3364), .CK(CLK), .RN(n444), .Q(n3739)
         );
  DFFR_X1 \REGISTERS_reg[14][28]  ( .D(n3363), .CK(CLK), .RN(n444), .Q(n3738)
         );
  DFFR_X1 \REGISTERS_reg[14][27]  ( .D(n3362), .CK(CLK), .RN(n445), .Q(n3737)
         );
  DFFR_X1 \REGISTERS_reg[14][26]  ( .D(n3361), .CK(CLK), .RN(n445), .Q(n3736)
         );
  DFFR_X1 \REGISTERS_reg[14][25]  ( .D(n3360), .CK(CLK), .RN(n445), .Q(n3735)
         );
  DFFR_X1 \REGISTERS_reg[14][24]  ( .D(n3359), .CK(CLK), .RN(n445), .Q(n3734)
         );
  DFFR_X1 \REGISTERS_reg[14][23]  ( .D(n3358), .CK(CLK), .RN(n445), .Q(n3733)
         );
  DFFR_X1 \REGISTERS_reg[14][22]  ( .D(n3357), .CK(CLK), .RN(n445), .Q(n3732)
         );
  DFFR_X1 \REGISTERS_reg[14][21]  ( .D(n3356), .CK(CLK), .RN(n445), .Q(n3731)
         );
  DFFR_X1 \REGISTERS_reg[14][20]  ( .D(n3355), .CK(CLK), .RN(n445), .Q(n3730)
         );
  DFFR_X1 \REGISTERS_reg[14][19]  ( .D(n3354), .CK(CLK), .RN(n445), .Q(n3729)
         );
  DFFR_X1 \REGISTERS_reg[14][18]  ( .D(n3353), .CK(CLK), .RN(n445), .Q(n3728)
         );
  DFFR_X1 \REGISTERS_reg[14][17]  ( .D(n3352), .CK(CLK), .RN(n445), .Q(n3727)
         );
  DFFR_X1 \REGISTERS_reg[14][16]  ( .D(n3351), .CK(CLK), .RN(n445), .Q(n3726)
         );
  DFFR_X1 \REGISTERS_reg[14][15]  ( .D(n3350), .CK(CLK), .RN(n446), .Q(n3725)
         );
  DFFR_X1 \REGISTERS_reg[14][14]  ( .D(n3349), .CK(CLK), .RN(n446), .Q(n3724)
         );
  DFFR_X1 \REGISTERS_reg[14][13]  ( .D(n3348), .CK(CLK), .RN(n446), .Q(n3723)
         );
  DFFR_X1 \REGISTERS_reg[14][12]  ( .D(n3347), .CK(CLK), .RN(n446), .Q(n3722)
         );
  DFFR_X1 \REGISTERS_reg[14][11]  ( .D(n3346), .CK(CLK), .RN(n446), .Q(n3721)
         );
  DFFR_X1 \REGISTERS_reg[14][10]  ( .D(n3345), .CK(CLK), .RN(n446), .Q(n3720)
         );
  DFFR_X1 \REGISTERS_reg[14][9]  ( .D(n3344), .CK(CLK), .RN(n446), .Q(n3719)
         );
  DFFR_X1 \REGISTERS_reg[14][8]  ( .D(n3343), .CK(CLK), .RN(n446), .Q(n3718)
         );
  DFFR_X1 \REGISTERS_reg[14][7]  ( .D(n3342), .CK(CLK), .RN(n446), .Q(n3717)
         );
  DFFR_X1 \REGISTERS_reg[14][6]  ( .D(n3341), .CK(CLK), .RN(n446), .Q(n3716)
         );
  DFFR_X1 \REGISTERS_reg[14][5]  ( .D(n3340), .CK(CLK), .RN(n446), .Q(n3715)
         );
  DFFR_X1 \REGISTERS_reg[14][4]  ( .D(n3339), .CK(CLK), .RN(n446), .Q(n3714)
         );
  DFFR_X1 \REGISTERS_reg[14][3]  ( .D(n3338), .CK(CLK), .RN(n447), .Q(n3713)
         );
  DFFR_X1 \REGISTERS_reg[14][2]  ( .D(n3337), .CK(CLK), .RN(n447), .Q(n3712)
         );
  DFFR_X1 \REGISTERS_reg[14][1]  ( .D(n3336), .CK(CLK), .RN(n447), .Q(n3711)
         );
  DFFR_X1 \REGISTERS_reg[14][0]  ( .D(n3335), .CK(CLK), .RN(n447), .Q(n3710)
         );
  DFFR_X1 \REGISTERS_reg[15][31]  ( .D(n3334), .CK(CLK), .RN(n447), .Q(n3709)
         );
  DFFR_X1 \REGISTERS_reg[15][30]  ( .D(n3333), .CK(CLK), .RN(n447), .Q(n3708)
         );
  DFFR_X1 \REGISTERS_reg[15][29]  ( .D(n3332), .CK(CLK), .RN(n447), .Q(n3707)
         );
  DFFR_X1 \REGISTERS_reg[15][28]  ( .D(n3331), .CK(CLK), .RN(n447), .Q(n3706)
         );
  DFFR_X1 \REGISTERS_reg[15][27]  ( .D(n3330), .CK(CLK), .RN(n447), .Q(n3705)
         );
  DFFR_X1 \REGISTERS_reg[15][26]  ( .D(n3329), .CK(CLK), .RN(n447), .Q(n3704)
         );
  DFFR_X1 \REGISTERS_reg[15][25]  ( .D(n3328), .CK(CLK), .RN(n447), .Q(n3703)
         );
  DFFR_X1 \REGISTERS_reg[15][24]  ( .D(n3327), .CK(CLK), .RN(n447), .Q(n3702)
         );
  DFFR_X1 \REGISTERS_reg[15][23]  ( .D(n3326), .CK(CLK), .RN(n448), .Q(n3701)
         );
  DFFR_X1 \REGISTERS_reg[15][22]  ( .D(n3325), .CK(CLK), .RN(n448), .Q(n3700)
         );
  DFFR_X1 \REGISTERS_reg[15][21]  ( .D(n3324), .CK(CLK), .RN(n448), .Q(n3699)
         );
  DFFR_X1 \REGISTERS_reg[15][20]  ( .D(n3323), .CK(CLK), .RN(n448), .Q(n3698)
         );
  DFFR_X1 \REGISTERS_reg[15][19]  ( .D(n3322), .CK(CLK), .RN(n448), .Q(n3697)
         );
  DFFR_X1 \REGISTERS_reg[15][18]  ( .D(n3321), .CK(CLK), .RN(n448), .Q(n3696)
         );
  DFFR_X1 \REGISTERS_reg[15][17]  ( .D(n3320), .CK(CLK), .RN(n448), .Q(n3695)
         );
  DFFR_X1 \REGISTERS_reg[15][16]  ( .D(n3319), .CK(CLK), .RN(n448), .Q(n3694)
         );
  DFFR_X1 \REGISTERS_reg[15][15]  ( .D(n3318), .CK(CLK), .RN(n448), .Q(n3693)
         );
  DFFR_X1 \REGISTERS_reg[15][14]  ( .D(n3317), .CK(CLK), .RN(n448), .Q(n3692)
         );
  DFFR_X1 \REGISTERS_reg[15][13]  ( .D(n3316), .CK(CLK), .RN(n448), .Q(n3691)
         );
  DFFR_X1 \REGISTERS_reg[15][12]  ( .D(n3315), .CK(CLK), .RN(n448), .Q(n3690)
         );
  DFFR_X1 \REGISTERS_reg[15][11]  ( .D(n3314), .CK(CLK), .RN(n449), .Q(n3689)
         );
  DFFR_X1 \REGISTERS_reg[15][10]  ( .D(n3313), .CK(CLK), .RN(n449), .Q(n3688)
         );
  DFFR_X1 \REGISTERS_reg[15][9]  ( .D(n3312), .CK(CLK), .RN(n449), .Q(n3687)
         );
  DFFR_X1 \REGISTERS_reg[15][8]  ( .D(n3311), .CK(CLK), .RN(n449), .Q(n3686)
         );
  DFFR_X1 \REGISTERS_reg[15][7]  ( .D(n3310), .CK(CLK), .RN(n449), .Q(n3685)
         );
  DFFR_X1 \REGISTERS_reg[15][6]  ( .D(n3309), .CK(CLK), .RN(n449), .Q(n3684)
         );
  DFFR_X1 \REGISTERS_reg[15][5]  ( .D(n3308), .CK(CLK), .RN(n449), .Q(n3683)
         );
  DFFR_X1 \REGISTERS_reg[15][4]  ( .D(n3307), .CK(CLK), .RN(n449), .Q(n3682)
         );
  DFFR_X1 \REGISTERS_reg[15][3]  ( .D(n3306), .CK(CLK), .RN(n449), .Q(n3681)
         );
  DFFR_X1 \REGISTERS_reg[15][2]  ( .D(n3305), .CK(CLK), .RN(n449), .Q(n3680)
         );
  DFFR_X1 \REGISTERS_reg[15][1]  ( .D(n3304), .CK(CLK), .RN(n449), .Q(n3679)
         );
  DFFR_X1 \REGISTERS_reg[15][0]  ( .D(n3303), .CK(CLK), .RN(n449), .Q(n3678)
         );
  DFFR_X1 \REGISTERS_reg[18][30]  ( .D(n3301), .CK(CLK), .RN(n455), .Q(n3644)
         );
  DFFR_X1 \REGISTERS_reg[18][29]  ( .D(n3300), .CK(CLK), .RN(n455), .Q(n3643)
         );
  DFFR_X1 \REGISTERS_reg[18][28]  ( .D(n3299), .CK(CLK), .RN(n455), .Q(n3642)
         );
  DFFR_X1 \REGISTERS_reg[18][27]  ( .D(n3298), .CK(CLK), .RN(n455), .Q(n3641)
         );
  DFFR_X1 \REGISTERS_reg[18][26]  ( .D(n3297), .CK(CLK), .RN(n455), .Q(n3640)
         );
  DFFR_X1 \REGISTERS_reg[18][25]  ( .D(n3296), .CK(CLK), .RN(n455), .Q(n3639)
         );
  DFFR_X1 \REGISTERS_reg[18][24]  ( .D(n3295), .CK(CLK), .RN(n455), .Q(n3638)
         );
  DFFR_X1 \REGISTERS_reg[18][23]  ( .D(n3294), .CK(CLK), .RN(n456), .Q(n3637)
         );
  DFFR_X1 \REGISTERS_reg[18][22]  ( .D(n3293), .CK(CLK), .RN(n456), .Q(n3636)
         );
  DFFR_X1 \REGISTERS_reg[18][21]  ( .D(n3292), .CK(CLK), .RN(n456), .Q(n3635)
         );
  DFFR_X1 \REGISTERS_reg[18][20]  ( .D(n3291), .CK(CLK), .RN(n456), .Q(n3634)
         );
  DFFR_X1 \REGISTERS_reg[18][19]  ( .D(n3290), .CK(CLK), .RN(n456), .Q(n3633)
         );
  DFFR_X1 \REGISTERS_reg[18][18]  ( .D(n3289), .CK(CLK), .RN(n456), .Q(n3632)
         );
  DFFR_X1 \REGISTERS_reg[18][17]  ( .D(n3288), .CK(CLK), .RN(n456), .Q(n3631)
         );
  DFFR_X1 \REGISTERS_reg[18][16]  ( .D(n3287), .CK(CLK), .RN(n456), .Q(n3630)
         );
  DFFR_X1 \REGISTERS_reg[18][15]  ( .D(n3286), .CK(CLK), .RN(n456), .Q(n3629)
         );
  DFFR_X1 \REGISTERS_reg[18][14]  ( .D(n3285), .CK(CLK), .RN(n456), .Q(n3628)
         );
  DFFR_X1 \REGISTERS_reg[18][13]  ( .D(n3284), .CK(CLK), .RN(n456), .Q(n3627)
         );
  DFFR_X1 \REGISTERS_reg[18][12]  ( .D(n3283), .CK(CLK), .RN(n456), .Q(n3626)
         );
  DFFR_X1 \REGISTERS_reg[18][11]  ( .D(n3282), .CK(CLK), .RN(n457), .Q(n3625)
         );
  DFFR_X1 \REGISTERS_reg[18][10]  ( .D(n3281), .CK(CLK), .RN(n457), .Q(n3624)
         );
  DFFR_X1 \REGISTERS_reg[18][9]  ( .D(n3280), .CK(CLK), .RN(n457), .Q(n3623)
         );
  DFFR_X1 \REGISTERS_reg[18][8]  ( .D(n3279), .CK(CLK), .RN(n457), .Q(n3622)
         );
  DFFR_X1 \REGISTERS_reg[18][7]  ( .D(n3278), .CK(CLK), .RN(n457), .Q(n3621)
         );
  DFFR_X1 \REGISTERS_reg[18][6]  ( .D(n3277), .CK(CLK), .RN(n457), .Q(n3620)
         );
  DFFR_X1 \REGISTERS_reg[18][5]  ( .D(n3276), .CK(CLK), .RN(n457), .Q(n3619)
         );
  DFFR_X1 \REGISTERS_reg[18][4]  ( .D(n3275), .CK(CLK), .RN(n457), .Q(n3618)
         );
  DFFR_X1 \REGISTERS_reg[18][3]  ( .D(n3274), .CK(CLK), .RN(n457), .Q(n3617)
         );
  DFFR_X1 \REGISTERS_reg[18][2]  ( .D(n3273), .CK(CLK), .RN(n457), .Q(n3616)
         );
  DFFR_X1 \REGISTERS_reg[18][1]  ( .D(n3272), .CK(CLK), .RN(n457), .Q(n3615)
         );
  DFFR_X1 \REGISTERS_reg[18][0]  ( .D(n3271), .CK(CLK), .RN(n457), .Q(n3614)
         );
  DFFR_X1 \REGISTERS_reg[19][31]  ( .D(n3270), .CK(CLK), .RN(n458), .Q(n3613)
         );
  DFFR_X1 \REGISTERS_reg[19][30]  ( .D(n3269), .CK(CLK), .RN(n458), .Q(n3612)
         );
  DFFR_X1 \REGISTERS_reg[19][29]  ( .D(n3268), .CK(CLK), .RN(n458), .Q(n3611)
         );
  DFFR_X1 \REGISTERS_reg[19][28]  ( .D(n3267), .CK(CLK), .RN(n458), .Q(n3610)
         );
  DFFR_X1 \REGISTERS_reg[19][27]  ( .D(n3266), .CK(CLK), .RN(n458), .Q(n3609)
         );
  DFFR_X1 \REGISTERS_reg[19][26]  ( .D(n3265), .CK(CLK), .RN(n458), .Q(n3608)
         );
  DFFR_X1 \REGISTERS_reg[19][25]  ( .D(n3264), .CK(CLK), .RN(n458), .Q(n3607)
         );
  DFFR_X1 \REGISTERS_reg[19][24]  ( .D(n3263), .CK(CLK), .RN(n458), .Q(n3606)
         );
  DFFR_X1 \REGISTERS_reg[19][23]  ( .D(n3262), .CK(CLK), .RN(n458), .Q(n3605)
         );
  DFFR_X1 \REGISTERS_reg[19][22]  ( .D(n3261), .CK(CLK), .RN(n458), .Q(n3604)
         );
  DFFR_X1 \REGISTERS_reg[19][21]  ( .D(n3260), .CK(CLK), .RN(n458), .Q(n3603)
         );
  DFFR_X1 \REGISTERS_reg[19][20]  ( .D(n3259), .CK(CLK), .RN(n458), .Q(n3602)
         );
  DFFR_X1 \REGISTERS_reg[19][19]  ( .D(n3258), .CK(CLK), .RN(n459), .Q(n3601)
         );
  DFFR_X1 \REGISTERS_reg[19][18]  ( .D(n3257), .CK(CLK), .RN(n459), .Q(n3600)
         );
  DFFR_X1 \REGISTERS_reg[19][17]  ( .D(n3256), .CK(CLK), .RN(n459), .Q(n3599)
         );
  DFFR_X1 \REGISTERS_reg[19][16]  ( .D(n3255), .CK(CLK), .RN(n459), .Q(n3598)
         );
  DFFR_X1 \REGISTERS_reg[19][15]  ( .D(n3254), .CK(CLK), .RN(n459), .Q(n3597)
         );
  DFFR_X1 \REGISTERS_reg[19][14]  ( .D(n3253), .CK(CLK), .RN(n459), .Q(n3596)
         );
  DFFR_X1 \REGISTERS_reg[19][13]  ( .D(n3252), .CK(CLK), .RN(n459), .Q(n3595)
         );
  DFFR_X1 \REGISTERS_reg[19][12]  ( .D(n3251), .CK(CLK), .RN(n459), .Q(n3594)
         );
  DFFR_X1 \REGISTERS_reg[19][11]  ( .D(n3250), .CK(CLK), .RN(n459), .Q(n3593)
         );
  DFFR_X1 \REGISTERS_reg[19][10]  ( .D(n3249), .CK(CLK), .RN(n459), .Q(n3592)
         );
  DFFR_X1 \REGISTERS_reg[19][9]  ( .D(n3248), .CK(CLK), .RN(n459), .Q(n3591)
         );
  DFFR_X1 \REGISTERS_reg[19][8]  ( .D(n3247), .CK(CLK), .RN(n459), .Q(n3590)
         );
  DFFR_X1 \REGISTERS_reg[19][7]  ( .D(n3246), .CK(CLK), .RN(n460), .Q(n3589)
         );
  DFFR_X1 \REGISTERS_reg[19][6]  ( .D(n3245), .CK(CLK), .RN(n460), .Q(n3588)
         );
  DFFR_X1 \REGISTERS_reg[19][5]  ( .D(n3244), .CK(CLK), .RN(n460), .Q(n3587)
         );
  DFFR_X1 \REGISTERS_reg[19][4]  ( .D(n3243), .CK(CLK), .RN(n460), .Q(n3586)
         );
  DFFR_X1 \REGISTERS_reg[19][3]  ( .D(n3242), .CK(CLK), .RN(n460), .Q(n3585)
         );
  DFFR_X1 \REGISTERS_reg[19][2]  ( .D(n3241), .CK(CLK), .RN(n460), .Q(n3584)
         );
  DFFR_X1 \REGISTERS_reg[19][1]  ( .D(n3240), .CK(CLK), .RN(n460), .Q(n3583)
         );
  DFFR_X1 \REGISTERS_reg[19][0]  ( .D(n3239), .CK(CLK), .RN(n460), .Q(n3582)
         );
  DFFR_X1 \REGISTERS_reg[25][31]  ( .D(n3142), .CK(CLK), .RN(n474), .Q(n2845)
         );
  DFFR_X1 \REGISTERS_reg[25][30]  ( .D(n3141), .CK(CLK), .RN(n474), .Q(n2844)
         );
  DFFR_X1 \REGISTERS_reg[25][29]  ( .D(n3140), .CK(CLK), .RN(n474), .Q(n2843)
         );
  DFFR_X1 \REGISTERS_reg[25][28]  ( .D(n3139), .CK(CLK), .RN(n474), .Q(n2842)
         );
  DFFR_X1 \REGISTERS_reg[25][27]  ( .D(n3138), .CK(CLK), .RN(n474), .Q(n2841)
         );
  DFFR_X1 \REGISTERS_reg[25][26]  ( .D(n3137), .CK(CLK), .RN(n474), .Q(n2840)
         );
  DFFR_X1 \REGISTERS_reg[25][25]  ( .D(n3136), .CK(CLK), .RN(n474), .Q(n2839)
         );
  DFFR_X1 \REGISTERS_reg[25][24]  ( .D(n3135), .CK(CLK), .RN(n474), .Q(n2838)
         );
  DFFR_X1 \REGISTERS_reg[25][23]  ( .D(n3134), .CK(CLK), .RN(n474), .Q(n2837)
         );
  DFFR_X1 \REGISTERS_reg[25][22]  ( .D(n3133), .CK(CLK), .RN(n474), .Q(n2836)
         );
  DFFR_X1 \REGISTERS_reg[25][21]  ( .D(n3132), .CK(CLK), .RN(n474), .Q(n2835)
         );
  DFFR_X1 \REGISTERS_reg[25][20]  ( .D(n3131), .CK(CLK), .RN(n474), .Q(n2834)
         );
  DFFR_X1 \REGISTERS_reg[25][19]  ( .D(n3130), .CK(CLK), .RN(n475), .Q(n2833)
         );
  DFFR_X1 \REGISTERS_reg[25][18]  ( .D(n3129), .CK(CLK), .RN(n475), .Q(n2832)
         );
  DFFR_X1 \REGISTERS_reg[25][17]  ( .D(n3128), .CK(CLK), .RN(n475), .Q(n2831)
         );
  DFFR_X1 \REGISTERS_reg[25][16]  ( .D(n3127), .CK(CLK), .RN(n475), .Q(n2830)
         );
  DFFR_X1 \REGISTERS_reg[25][15]  ( .D(n3126), .CK(CLK), .RN(n475), .Q(n2829)
         );
  DFFR_X1 \REGISTERS_reg[25][14]  ( .D(n3125), .CK(CLK), .RN(n475), .Q(n2828)
         );
  DFFR_X1 \REGISTERS_reg[25][13]  ( .D(n3124), .CK(CLK), .RN(n475), .Q(n2827)
         );
  DFFR_X1 \REGISTERS_reg[25][12]  ( .D(n3123), .CK(CLK), .RN(n475), .Q(n2826)
         );
  DFFR_X1 \REGISTERS_reg[25][11]  ( .D(n3122), .CK(CLK), .RN(n475), .Q(n2825)
         );
  DFFR_X1 \REGISTERS_reg[25][10]  ( .D(n3121), .CK(CLK), .RN(n475), .Q(n2824)
         );
  DFFR_X1 \REGISTERS_reg[25][9]  ( .D(n3120), .CK(CLK), .RN(n475), .Q(n2823)
         );
  DFFR_X1 \REGISTERS_reg[25][8]  ( .D(n3119), .CK(CLK), .RN(n475), .Q(n2822)
         );
  DFFR_X1 \REGISTERS_reg[25][7]  ( .D(n3118), .CK(CLK), .RN(n476), .Q(n2821)
         );
  DFFR_X1 \REGISTERS_reg[25][6]  ( .D(n3117), .CK(CLK), .RN(n476), .Q(n2820)
         );
  DFFR_X1 \REGISTERS_reg[25][5]  ( .D(n3116), .CK(CLK), .RN(n476), .Q(n2819)
         );
  DFFR_X1 \REGISTERS_reg[25][4]  ( .D(n3115), .CK(CLK), .RN(n476), .Q(n2818)
         );
  DFFR_X1 \REGISTERS_reg[25][3]  ( .D(n3114), .CK(CLK), .RN(n476), .Q(n2817)
         );
  DFFR_X1 \REGISTERS_reg[25][2]  ( .D(n3113), .CK(CLK), .RN(n476), .Q(n2816)
         );
  DFFR_X1 \REGISTERS_reg[25][1]  ( .D(n3112), .CK(CLK), .RN(n476), .Q(n2815)
         );
  DFFR_X1 \REGISTERS_reg[25][0]  ( .D(n3111), .CK(CLK), .RN(n476), .Q(n2814)
         );
  DFFR_X1 \REGISTERS_reg[29][31]  ( .D(n3078), .CK(CLK), .RN(n484), .Q(n2781)
         );
  DFFR_X1 \REGISTERS_reg[29][30]  ( .D(n3077), .CK(CLK), .RN(n484), .Q(n2780)
         );
  DFFR_X1 \REGISTERS_reg[29][29]  ( .D(n3076), .CK(CLK), .RN(n484), .Q(n2779)
         );
  DFFR_X1 \REGISTERS_reg[29][28]  ( .D(n3075), .CK(CLK), .RN(n484), .Q(n2778)
         );
  DFFR_X1 \REGISTERS_reg[29][27]  ( .D(n3074), .CK(CLK), .RN(n485), .Q(n2777)
         );
  DFFR_X1 \REGISTERS_reg[29][26]  ( .D(n3073), .CK(CLK), .RN(n485), .Q(n2776)
         );
  DFFR_X1 \REGISTERS_reg[29][25]  ( .D(n3072), .CK(CLK), .RN(n485), .Q(n2775)
         );
  DFFR_X1 \REGISTERS_reg[29][24]  ( .D(n3071), .CK(CLK), .RN(n485), .Q(n2774)
         );
  DFFR_X1 \REGISTERS_reg[29][23]  ( .D(n3070), .CK(CLK), .RN(n485), .Q(n2773)
         );
  DFFR_X1 \REGISTERS_reg[29][22]  ( .D(n3069), .CK(CLK), .RN(n485), .Q(n2772)
         );
  DFFR_X1 \REGISTERS_reg[29][21]  ( .D(n3068), .CK(CLK), .RN(n485), .Q(n2771)
         );
  DFFR_X1 \REGISTERS_reg[29][20]  ( .D(n3067), .CK(CLK), .RN(n485), .Q(n2770)
         );
  DFFR_X1 \REGISTERS_reg[29][19]  ( .D(n3066), .CK(CLK), .RN(n485), .Q(n2769)
         );
  DFFR_X1 \REGISTERS_reg[29][18]  ( .D(n3065), .CK(CLK), .RN(n485), .Q(n2768)
         );
  DFFR_X1 \REGISTERS_reg[29][17]  ( .D(n3064), .CK(CLK), .RN(n485), .Q(n2767)
         );
  DFFR_X1 \REGISTERS_reg[29][16]  ( .D(n3063), .CK(CLK), .RN(n485), .Q(n2766)
         );
  DFFR_X1 \REGISTERS_reg[29][15]  ( .D(n3062), .CK(CLK), .RN(n486), .Q(n2765)
         );
  DFFR_X1 \REGISTERS_reg[29][14]  ( .D(n3061), .CK(CLK), .RN(n486), .Q(n2764)
         );
  DFFR_X1 \REGISTERS_reg[29][13]  ( .D(n3060), .CK(CLK), .RN(n486), .Q(n2763)
         );
  DFFR_X1 \REGISTERS_reg[29][12]  ( .D(n3059), .CK(CLK), .RN(n486), .Q(n2762)
         );
  DFFR_X1 \REGISTERS_reg[29][11]  ( .D(n3058), .CK(CLK), .RN(n486), .Q(n2761)
         );
  DFFR_X1 \REGISTERS_reg[29][10]  ( .D(n3057), .CK(CLK), .RN(n486), .Q(n2760)
         );
  DFFR_X1 \REGISTERS_reg[29][9]  ( .D(n3056), .CK(CLK), .RN(n486), .Q(n2759)
         );
  DFFR_X1 \REGISTERS_reg[29][8]  ( .D(n3055), .CK(CLK), .RN(n486), .Q(n2758)
         );
  DFFR_X1 \REGISTERS_reg[29][7]  ( .D(n3054), .CK(CLK), .RN(n486), .Q(n2757)
         );
  DFFR_X1 \REGISTERS_reg[29][6]  ( .D(n3053), .CK(CLK), .RN(n486), .Q(n2756)
         );
  DFFR_X1 \REGISTERS_reg[29][5]  ( .D(n3052), .CK(CLK), .RN(n486), .Q(n2755)
         );
  DFFR_X1 \REGISTERS_reg[29][4]  ( .D(n3051), .CK(CLK), .RN(n486), .Q(n2754)
         );
  DFFR_X1 \REGISTERS_reg[29][3]  ( .D(n3050), .CK(CLK), .RN(n487), .Q(n2753)
         );
  DFFR_X1 \REGISTERS_reg[29][2]  ( .D(n3049), .CK(CLK), .RN(n487), .Q(n2752)
         );
  DFFR_X1 \REGISTERS_reg[29][1]  ( .D(n3048), .CK(CLK), .RN(n487), .Q(n2751)
         );
  DFFR_X1 \REGISTERS_reg[29][0]  ( .D(n3047), .CK(CLK), .RN(n487), .Q(n2750)
         );
  DFF_X1 \OUT2_reg[31]  ( .D(n3015), .CK(CLK), .Q(OUT2[31]), .QN(n2654) );
  DFF_X1 \OUT2_reg[30]  ( .D(n3016), .CK(CLK), .Q(OUT2[30]), .QN(n2655) );
  DFF_X1 \OUT2_reg[29]  ( .D(n3017), .CK(CLK), .Q(OUT2[29]), .QN(n2656) );
  DFF_X1 \OUT2_reg[28]  ( .D(n3018), .CK(CLK), .Q(OUT2[28]), .QN(n2657) );
  DFF_X1 \OUT2_reg[27]  ( .D(n3019), .CK(CLK), .Q(OUT2[27]), .QN(n2658) );
  DFF_X1 \OUT2_reg[26]  ( .D(n3020), .CK(CLK), .Q(OUT2[26]), .QN(n2659) );
  DFF_X1 \OUT2_reg[25]  ( .D(n3021), .CK(CLK), .Q(OUT2[25]), .QN(n2660) );
  DFF_X1 \OUT2_reg[24]  ( .D(n3022), .CK(CLK), .Q(OUT2[24]), .QN(n2661) );
  DFF_X1 \OUT2_reg[23]  ( .D(n3023), .CK(CLK), .Q(OUT2[23]), .QN(n2662) );
  DFF_X1 \OUT2_reg[22]  ( .D(n3024), .CK(CLK), .Q(OUT2[22]), .QN(n2663) );
  DFF_X1 \OUT2_reg[21]  ( .D(n3025), .CK(CLK), .Q(OUT2[21]), .QN(n2664) );
  DFF_X1 \OUT2_reg[20]  ( .D(n3026), .CK(CLK), .Q(OUT2[20]), .QN(n2665) );
  DFF_X1 \OUT2_reg[19]  ( .D(n3027), .CK(CLK), .Q(OUT2[19]), .QN(n2666) );
  DFF_X1 \OUT2_reg[18]  ( .D(n3028), .CK(CLK), .Q(OUT2[18]), .QN(n2667) );
  DFF_X1 \OUT2_reg[17]  ( .D(n3029), .CK(CLK), .Q(OUT2[17]), .QN(n2668) );
  DFF_X1 \OUT2_reg[16]  ( .D(n3030), .CK(CLK), .Q(OUT2[16]), .QN(n2669) );
  DFF_X1 \OUT2_reg[15]  ( .D(n3031), .CK(CLK), .Q(OUT2[15]), .QN(n2670) );
  DFF_X1 \OUT2_reg[14]  ( .D(n3032), .CK(CLK), .Q(OUT2[14]), .QN(n2671) );
  DFF_X1 \OUT2_reg[13]  ( .D(n3033), .CK(CLK), .Q(OUT2[13]), .QN(n2672) );
  DFF_X1 \OUT2_reg[12]  ( .D(n3034), .CK(CLK), .Q(OUT2[12]), .QN(n2673) );
  DFF_X1 \OUT2_reg[11]  ( .D(n3035), .CK(CLK), .Q(OUT2[11]), .QN(n2674) );
  DFF_X1 \OUT2_reg[10]  ( .D(n3036), .CK(CLK), .Q(OUT2[10]), .QN(n2675) );
  DFF_X1 \OUT2_reg[9]  ( .D(n3037), .CK(CLK), .Q(OUT2[9]), .QN(n2676) );
  DFF_X1 \OUT2_reg[8]  ( .D(n3038), .CK(CLK), .Q(OUT2[8]), .QN(n2677) );
  DFF_X1 \OUT2_reg[7]  ( .D(n3039), .CK(CLK), .Q(OUT2[7]), .QN(n2678) );
  DFF_X1 \OUT2_reg[6]  ( .D(n3040), .CK(CLK), .Q(OUT2[6]), .QN(n2679) );
  DFF_X1 \OUT2_reg[5]  ( .D(n3041), .CK(CLK), .Q(OUT2[5]), .QN(n2680) );
  DFF_X1 \OUT2_reg[4]  ( .D(n3042), .CK(CLK), .Q(OUT2[4]), .QN(n2681) );
  DFF_X1 \OUT2_reg[3]  ( .D(n3043), .CK(CLK), .Q(OUT2[3]), .QN(n2682) );
  DFF_X1 \OUT2_reg[2]  ( .D(n3044), .CK(CLK), .Q(OUT2[2]), .QN(n2683) );
  DFF_X1 \OUT2_reg[1]  ( .D(n3045), .CK(CLK), .Q(OUT2[1]), .QN(n2684) );
  DFF_X1 \OUT2_reg[0]  ( .D(n3046), .CK(CLK), .Q(OUT2[0]), .QN(n2685) );
  DFF_X1 \OUT1_reg[31]  ( .D(n3014), .CK(CLK), .Q(OUT1[31]), .QN(n2653) );
  DFF_X1 \OUT1_reg[30]  ( .D(n3013), .CK(CLK), .Q(OUT1[30]), .QN(n2652) );
  DFF_X1 \OUT1_reg[29]  ( .D(n3012), .CK(CLK), .Q(OUT1[29]), .QN(n2651) );
  DFF_X1 \OUT1_reg[28]  ( .D(n3011), .CK(CLK), .Q(OUT1[28]), .QN(n2650) );
  DFF_X1 \OUT1_reg[27]  ( .D(n3010), .CK(CLK), .Q(OUT1[27]), .QN(n2649) );
  DFF_X1 \OUT1_reg[26]  ( .D(n3009), .CK(CLK), .Q(OUT1[26]), .QN(n2648) );
  DFF_X1 \OUT1_reg[25]  ( .D(n3008), .CK(CLK), .Q(OUT1[25]), .QN(n2647) );
  DFF_X1 \OUT1_reg[24]  ( .D(n3007), .CK(CLK), .Q(OUT1[24]), .QN(n2646) );
  DFF_X1 \OUT1_reg[23]  ( .D(n3006), .CK(CLK), .Q(OUT1[23]), .QN(n2645) );
  DFF_X1 \OUT1_reg[22]  ( .D(n3005), .CK(CLK), .Q(OUT1[22]), .QN(n2644) );
  DFF_X1 \OUT1_reg[21]  ( .D(n3004), .CK(CLK), .Q(OUT1[21]), .QN(n2643) );
  DFF_X1 \OUT1_reg[20]  ( .D(n3003), .CK(CLK), .Q(OUT1[20]), .QN(n2642) );
  DFF_X1 \OUT1_reg[19]  ( .D(n3002), .CK(CLK), .Q(OUT1[19]), .QN(n2641) );
  DFF_X1 \OUT1_reg[18]  ( .D(n3001), .CK(CLK), .Q(OUT1[18]), .QN(n2640) );
  DFF_X1 \OUT1_reg[17]  ( .D(n3000), .CK(CLK), .Q(OUT1[17]), .QN(n2639) );
  DFF_X1 \OUT1_reg[16]  ( .D(n2999), .CK(CLK), .Q(OUT1[16]), .QN(n2638) );
  DFF_X1 \OUT1_reg[15]  ( .D(n2998), .CK(CLK), .Q(OUT1[15]), .QN(n2637) );
  DFF_X1 \OUT1_reg[14]  ( .D(n2997), .CK(CLK), .Q(OUT1[14]), .QN(n2636) );
  DFF_X1 \OUT1_reg[13]  ( .D(n2996), .CK(CLK), .Q(OUT1[13]), .QN(n2635) );
  DFF_X1 \OUT1_reg[12]  ( .D(n2995), .CK(CLK), .Q(OUT1[12]), .QN(n2634) );
  DFF_X1 \OUT1_reg[11]  ( .D(n2994), .CK(CLK), .Q(OUT1[11]), .QN(n2633) );
  DFF_X1 \OUT1_reg[10]  ( .D(n2993), .CK(CLK), .Q(OUT1[10]), .QN(n2632) );
  DFF_X1 \OUT1_reg[9]  ( .D(n2992), .CK(CLK), .Q(OUT1[9]), .QN(n2631) );
  DFF_X1 \OUT1_reg[8]  ( .D(n2991), .CK(CLK), .Q(OUT1[8]), .QN(n2630) );
  DFF_X1 \OUT1_reg[7]  ( .D(n2990), .CK(CLK), .Q(OUT1[7]), .QN(n2629) );
  DFF_X1 \OUT1_reg[6]  ( .D(n2989), .CK(CLK), .Q(OUT1[6]), .QN(n2628) );
  DFF_X1 \OUT1_reg[5]  ( .D(n2988), .CK(CLK), .Q(OUT1[5]), .QN(n2627) );
  DFF_X1 \OUT1_reg[4]  ( .D(n2987), .CK(CLK), .Q(OUT1[4]), .QN(n2626) );
  DFF_X1 \OUT1_reg[3]  ( .D(n2986), .CK(CLK), .Q(OUT1[3]), .QN(n2625) );
  DFF_X1 \OUT1_reg[2]  ( .D(n2985), .CK(CLK), .Q(OUT1[2]), .QN(n2624) );
  DFF_X1 \OUT1_reg[1]  ( .D(n2984), .CK(CLK), .Q(OUT1[1]), .QN(n2623) );
  DFF_X1 \OUT1_reg[0]  ( .D(n2983), .CK(CLK), .Q(OUT1[0]), .QN(n2622) );
  DFFR_X1 \REGISTERS_reg[24][31]  ( .D(n3174), .CK(CLK), .RN(RST), .Q(n2877), 
        .QN(n1435) );
  DFFR_X1 \REGISTERS_reg[24][30]  ( .D(n3173), .CK(CLK), .RN(n471), .Q(n2876), 
        .QN(n1419) );
  DFFR_X1 \REGISTERS_reg[24][29]  ( .D(n3172), .CK(CLK), .RN(n471), .Q(n2875), 
        .QN(n1403) );
  DFFR_X1 \REGISTERS_reg[24][28]  ( .D(n3171), .CK(CLK), .RN(n471), .Q(n2874), 
        .QN(n1387) );
  DFFR_X1 \REGISTERS_reg[24][27]  ( .D(n3170), .CK(CLK), .RN(n471), .Q(n2873), 
        .QN(n1371) );
  DFFR_X1 \REGISTERS_reg[24][26]  ( .D(n3169), .CK(CLK), .RN(n471), .Q(n2872), 
        .QN(n1355) );
  DFFR_X1 \REGISTERS_reg[24][25]  ( .D(n3168), .CK(CLK), .RN(n471), .Q(n2871), 
        .QN(n1339) );
  DFFR_X1 \REGISTERS_reg[24][24]  ( .D(n3167), .CK(CLK), .RN(n471), .Q(n2870), 
        .QN(n1323) );
  DFFR_X1 \REGISTERS_reg[24][23]  ( .D(n3166), .CK(CLK), .RN(n472), .Q(n2869), 
        .QN(n1307) );
  DFFR_X1 \REGISTERS_reg[24][22]  ( .D(n3165), .CK(CLK), .RN(n472), .Q(n2868), 
        .QN(n1291) );
  DFFR_X1 \REGISTERS_reg[24][21]  ( .D(n3164), .CK(CLK), .RN(n472), .Q(n2867), 
        .QN(n1275) );
  DFFR_X1 \REGISTERS_reg[24][20]  ( .D(n3163), .CK(CLK), .RN(n472), .Q(n2866), 
        .QN(n1259) );
  DFFR_X1 \REGISTERS_reg[24][19]  ( .D(n3162), .CK(CLK), .RN(n472), .Q(n2865), 
        .QN(n1243) );
  DFFR_X1 \REGISTERS_reg[24][18]  ( .D(n3161), .CK(CLK), .RN(n472), .Q(n2864), 
        .QN(n1227) );
  DFFR_X1 \REGISTERS_reg[24][17]  ( .D(n3160), .CK(CLK), .RN(n472), .Q(n2863), 
        .QN(n1211) );
  DFFR_X1 \REGISTERS_reg[24][16]  ( .D(n3159), .CK(CLK), .RN(n472), .Q(n2862), 
        .QN(n1195) );
  DFFR_X1 \REGISTERS_reg[24][15]  ( .D(n3158), .CK(CLK), .RN(n472), .Q(n2861), 
        .QN(n1179) );
  DFFR_X1 \REGISTERS_reg[24][14]  ( .D(n3157), .CK(CLK), .RN(n472), .Q(n2860), 
        .QN(n1163) );
  DFFR_X1 \REGISTERS_reg[24][13]  ( .D(n3156), .CK(CLK), .RN(n472), .Q(n2859), 
        .QN(n1147) );
  DFFR_X1 \REGISTERS_reg[24][12]  ( .D(n3155), .CK(CLK), .RN(n472), .Q(n2858), 
        .QN(n1131) );
  DFFR_X1 \REGISTERS_reg[24][11]  ( .D(n3154), .CK(CLK), .RN(n473), .Q(n2857), 
        .QN(n1115) );
  DFFR_X1 \REGISTERS_reg[24][10]  ( .D(n3153), .CK(CLK), .RN(n473), .Q(n2856), 
        .QN(n1099) );
  DFFR_X1 \REGISTERS_reg[24][9]  ( .D(n3152), .CK(CLK), .RN(n473), .Q(n2855), 
        .QN(n1083) );
  DFFR_X1 \REGISTERS_reg[24][8]  ( .D(n3151), .CK(CLK), .RN(n473), .Q(n2854), 
        .QN(n1067) );
  DFFR_X1 \REGISTERS_reg[24][7]  ( .D(n3150), .CK(CLK), .RN(n473), .Q(n2853), 
        .QN(n1051) );
  DFFR_X1 \REGISTERS_reg[24][6]  ( .D(n3149), .CK(CLK), .RN(n473), .Q(n2852), 
        .QN(n1035) );
  DFFR_X1 \REGISTERS_reg[24][5]  ( .D(n3148), .CK(CLK), .RN(n473), .Q(n2851), 
        .QN(n1019) );
  DFFR_X1 \REGISTERS_reg[24][4]  ( .D(n3147), .CK(CLK), .RN(n473), .Q(n2850), 
        .QN(n1003) );
  DFFR_X1 \REGISTERS_reg[24][3]  ( .D(n3146), .CK(CLK), .RN(n473), .Q(n2849), 
        .QN(n987) );
  DFFR_X1 \REGISTERS_reg[24][2]  ( .D(n3145), .CK(CLK), .RN(n473), .Q(n2848), 
        .QN(n971) );
  DFFR_X1 \REGISTERS_reg[24][1]  ( .D(n3144), .CK(CLK), .RN(n473), .Q(n2847), 
        .QN(n955) );
  DFFR_X1 \REGISTERS_reg[24][0]  ( .D(n3143), .CK(CLK), .RN(n473), .Q(n2846), 
        .QN(n938) );
  DFFR_X1 \REGISTERS_reg[23][31]  ( .D(n3206), .CK(CLK), .RN(n468), .Q(n2909), 
        .QN(n1437) );
  DFFR_X1 \REGISTERS_reg[23][30]  ( .D(n3205), .CK(CLK), .RN(n468), .Q(n2908), 
        .QN(n1420) );
  DFFR_X1 \REGISTERS_reg[23][29]  ( .D(n3204), .CK(CLK), .RN(n468), .Q(n2907), 
        .QN(n1404) );
  DFFR_X1 \REGISTERS_reg[23][28]  ( .D(n3203), .CK(CLK), .RN(n468), .Q(n2906), 
        .QN(n1388) );
  DFFR_X1 \REGISTERS_reg[23][27]  ( .D(n3202), .CK(CLK), .RN(n469), .Q(n2905), 
        .QN(n1372) );
  DFFR_X1 \REGISTERS_reg[23][26]  ( .D(n3201), .CK(CLK), .RN(n469), .Q(n2904), 
        .QN(n1356) );
  DFFR_X1 \REGISTERS_reg[23][25]  ( .D(n3200), .CK(CLK), .RN(n469), .Q(n2903), 
        .QN(n1340) );
  DFFR_X1 \REGISTERS_reg[23][24]  ( .D(n3199), .CK(CLK), .RN(n469), .Q(n2902), 
        .QN(n1324) );
  DFFR_X1 \REGISTERS_reg[23][23]  ( .D(n3198), .CK(CLK), .RN(n469), .Q(n2901), 
        .QN(n1308) );
  DFFR_X1 \REGISTERS_reg[23][22]  ( .D(n3197), .CK(CLK), .RN(n469), .Q(n2900), 
        .QN(n1292) );
  DFFR_X1 \REGISTERS_reg[23][21]  ( .D(n3196), .CK(CLK), .RN(n469), .Q(n2899), 
        .QN(n1276) );
  DFFR_X1 \REGISTERS_reg[23][20]  ( .D(n3195), .CK(CLK), .RN(n469), .Q(n2898), 
        .QN(n1260) );
  DFFR_X1 \REGISTERS_reg[23][19]  ( .D(n3194), .CK(CLK), .RN(n469), .Q(n2897), 
        .QN(n1244) );
  DFFR_X1 \REGISTERS_reg[23][18]  ( .D(n3193), .CK(CLK), .RN(n469), .Q(n2896), 
        .QN(n1228) );
  DFFR_X1 \REGISTERS_reg[23][17]  ( .D(n3192), .CK(CLK), .RN(n469), .Q(n2895), 
        .QN(n1212) );
  DFFR_X1 \REGISTERS_reg[23][16]  ( .D(n3191), .CK(CLK), .RN(n469), .Q(n2894), 
        .QN(n1196) );
  DFFR_X1 \REGISTERS_reg[23][15]  ( .D(n3190), .CK(CLK), .RN(n470), .Q(n2893), 
        .QN(n1180) );
  DFFR_X1 \REGISTERS_reg[23][14]  ( .D(n3189), .CK(CLK), .RN(n470), .Q(n2892), 
        .QN(n1164) );
  DFFR_X1 \REGISTERS_reg[23][13]  ( .D(n3188), .CK(CLK), .RN(n470), .Q(n2891), 
        .QN(n1148) );
  DFFR_X1 \REGISTERS_reg[23][12]  ( .D(n3187), .CK(CLK), .RN(n470), .Q(n2890), 
        .QN(n1132) );
  DFFR_X1 \REGISTERS_reg[23][11]  ( .D(n3186), .CK(CLK), .RN(n470), .Q(n2889), 
        .QN(n1116) );
  DFFR_X1 \REGISTERS_reg[23][10]  ( .D(n3185), .CK(CLK), .RN(n470), .Q(n2888), 
        .QN(n1100) );
  DFFR_X1 \REGISTERS_reg[23][9]  ( .D(n3184), .CK(CLK), .RN(n470), .Q(n2887), 
        .QN(n1084) );
  DFFR_X1 \REGISTERS_reg[23][8]  ( .D(n3183), .CK(CLK), .RN(n470), .Q(n2886), 
        .QN(n1068) );
  DFFR_X1 \REGISTERS_reg[23][7]  ( .D(n3182), .CK(CLK), .RN(n470), .Q(n2885), 
        .QN(n1052) );
  DFFR_X1 \REGISTERS_reg[23][6]  ( .D(n3181), .CK(CLK), .RN(n470), .Q(n2884), 
        .QN(n1036) );
  DFFR_X1 \REGISTERS_reg[23][5]  ( .D(n3180), .CK(CLK), .RN(n470), .Q(n2883), 
        .QN(n1020) );
  DFFR_X1 \REGISTERS_reg[23][4]  ( .D(n3179), .CK(CLK), .RN(n470), .Q(n2882), 
        .QN(n1004) );
  DFFR_X1 \REGISTERS_reg[23][3]  ( .D(n3178), .CK(CLK), .RN(n471), .Q(n2881), 
        .QN(n988) );
  DFFR_X1 \REGISTERS_reg[23][2]  ( .D(n3177), .CK(CLK), .RN(n471), .Q(n2880), 
        .QN(n972) );
  DFFR_X1 \REGISTERS_reg[23][1]  ( .D(n3176), .CK(CLK), .RN(n471), .Q(n2879), 
        .QN(n956) );
  DFFR_X1 \REGISTERS_reg[23][0]  ( .D(n3175), .CK(CLK), .RN(n471), .Q(n2878), 
        .QN(n939) );
  DFFR_X1 \REGISTERS_reg[22][31]  ( .D(n3238), .CK(CLK), .RN(n466), .Q(n2941), 
        .QN(n2320) );
  DFFR_X1 \REGISTERS_reg[22][30]  ( .D(n3237), .CK(CLK), .RN(n466), .Q(n2940), 
        .QN(n2299) );
  DFFR_X1 \REGISTERS_reg[22][29]  ( .D(n3236), .CK(CLK), .RN(n466), .Q(n2939), 
        .QN(n2287) );
  DFFR_X1 \REGISTERS_reg[22][28]  ( .D(n3235), .CK(CLK), .RN(n466), .Q(n2938), 
        .QN(n2275) );
  DFFR_X1 \REGISTERS_reg[22][27]  ( .D(n3234), .CK(CLK), .RN(n466), .Q(n2937), 
        .QN(n2263) );
  DFFR_X1 \REGISTERS_reg[22][26]  ( .D(n3233), .CK(CLK), .RN(n466), .Q(n2936), 
        .QN(n2251) );
  DFFR_X1 \REGISTERS_reg[22][25]  ( .D(n3232), .CK(CLK), .RN(n466), .Q(n2935), 
        .QN(n2239) );
  DFFR_X1 \REGISTERS_reg[22][24]  ( .D(n3231), .CK(CLK), .RN(n466), .Q(n2934), 
        .QN(n2227) );
  DFFR_X1 \REGISTERS_reg[22][23]  ( .D(n3230), .CK(CLK), .RN(n466), .Q(n2933), 
        .QN(n2215) );
  DFFR_X1 \REGISTERS_reg[22][22]  ( .D(n3229), .CK(CLK), .RN(n466), .Q(n2932), 
        .QN(n2203) );
  DFFR_X1 \REGISTERS_reg[22][21]  ( .D(n3228), .CK(CLK), .RN(n466), .Q(n2931), 
        .QN(n2191) );
  DFFR_X1 \REGISTERS_reg[22][20]  ( .D(n3227), .CK(CLK), .RN(n466), .Q(n2930), 
        .QN(n2179) );
  DFFR_X1 \REGISTERS_reg[22][19]  ( .D(n3226), .CK(CLK), .RN(n467), .Q(n2929), 
        .QN(n2167) );
  DFFR_X1 \REGISTERS_reg[22][18]  ( .D(n3225), .CK(CLK), .RN(n467), .Q(n2928), 
        .QN(n2155) );
  DFFR_X1 \REGISTERS_reg[22][17]  ( .D(n3224), .CK(CLK), .RN(n467), .Q(n2927), 
        .QN(n2143) );
  DFFR_X1 \REGISTERS_reg[22][16]  ( .D(n3223), .CK(CLK), .RN(n467), .Q(n2926), 
        .QN(n2131) );
  DFFR_X1 \REGISTERS_reg[22][15]  ( .D(n3222), .CK(CLK), .RN(n467), .Q(n2925), 
        .QN(n2119) );
  DFFR_X1 \REGISTERS_reg[22][14]  ( .D(n3221), .CK(CLK), .RN(n467), .Q(n2924), 
        .QN(n2107) );
  DFFR_X1 \REGISTERS_reg[22][13]  ( .D(n3220), .CK(CLK), .RN(n467), .Q(n2923), 
        .QN(n2095) );
  DFFR_X1 \REGISTERS_reg[22][12]  ( .D(n3219), .CK(CLK), .RN(n467), .Q(n2922), 
        .QN(n2083) );
  DFFR_X1 \REGISTERS_reg[22][11]  ( .D(n3218), .CK(CLK), .RN(n467), .Q(n2921), 
        .QN(n2071) );
  DFFR_X1 \REGISTERS_reg[22][10]  ( .D(n3217), .CK(CLK), .RN(n467), .Q(n2920), 
        .QN(n2059) );
  DFFR_X1 \REGISTERS_reg[22][9]  ( .D(n3216), .CK(CLK), .RN(n467), .Q(n2919), 
        .QN(n2047) );
  DFFR_X1 \REGISTERS_reg[22][8]  ( .D(n3215), .CK(CLK), .RN(n467), .Q(n2918), 
        .QN(n2035) );
  DFFR_X1 \REGISTERS_reg[22][7]  ( .D(n3214), .CK(CLK), .RN(n468), .Q(n2917), 
        .QN(n2023) );
  DFFR_X1 \REGISTERS_reg[22][6]  ( .D(n3213), .CK(CLK), .RN(n468), .Q(n2916), 
        .QN(n2011) );
  DFFR_X1 \REGISTERS_reg[22][5]  ( .D(n3212), .CK(CLK), .RN(n468), .Q(n2915), 
        .QN(n1999) );
  DFFR_X1 \REGISTERS_reg[22][4]  ( .D(n3211), .CK(CLK), .RN(n468), .Q(n2914), 
        .QN(n1987) );
  DFFR_X1 \REGISTERS_reg[22][3]  ( .D(n3210), .CK(CLK), .RN(n468), .Q(n2913), 
        .QN(n1975) );
  DFFR_X1 \REGISTERS_reg[22][2]  ( .D(n3209), .CK(CLK), .RN(n468), .Q(n2912), 
        .QN(n1963) );
  DFFR_X1 \REGISTERS_reg[22][1]  ( .D(n3208), .CK(CLK), .RN(n468), .Q(n2911), 
        .QN(n1951) );
  DFFR_X1 \REGISTERS_reg[22][0]  ( .D(n3207), .CK(CLK), .RN(n468), .Q(n2910), 
        .QN(n1922) );
  DFFR_X1 \REGISTERS_reg[7][31]  ( .D(n3462), .CK(CLK), .RN(n426), .Q(n3965), 
        .QN(n2331) );
  DFFR_X1 \REGISTERS_reg[7][30]  ( .D(n3461), .CK(CLK), .RN(n426), .Q(n3964), 
        .QN(n2306) );
  DFFR_X1 \REGISTERS_reg[7][29]  ( .D(n3460), .CK(CLK), .RN(n426), .Q(n3963), 
        .QN(n2294) );
  DFFR_X1 \REGISTERS_reg[7][28]  ( .D(n3459), .CK(CLK), .RN(n426), .Q(n3962), 
        .QN(n2282) );
  DFFR_X1 \REGISTERS_reg[7][27]  ( .D(n3458), .CK(CLK), .RN(n426), .Q(n3961), 
        .QN(n2270) );
  DFFR_X1 \REGISTERS_reg[7][26]  ( .D(n3457), .CK(CLK), .RN(n426), .Q(n3960), 
        .QN(n2258) );
  DFFR_X1 \REGISTERS_reg[7][25]  ( .D(n3456), .CK(CLK), .RN(n426), .Q(n3959), 
        .QN(n2246) );
  DFFR_X1 \REGISTERS_reg[7][24]  ( .D(n3455), .CK(CLK), .RN(n426), .Q(n3958), 
        .QN(n2234) );
  DFFR_X1 \REGISTERS_reg[7][23]  ( .D(n3454), .CK(CLK), .RN(n426), .Q(n3957), 
        .QN(n2222) );
  DFFR_X1 \REGISTERS_reg[7][22]  ( .D(n3453), .CK(CLK), .RN(n426), .Q(n3956), 
        .QN(n2210) );
  DFFR_X1 \REGISTERS_reg[7][21]  ( .D(n3452), .CK(CLK), .RN(n426), .Q(n3955), 
        .QN(n2198) );
  DFFR_X1 \REGISTERS_reg[7][20]  ( .D(n3451), .CK(CLK), .RN(n426), .Q(n3954), 
        .QN(n2186) );
  DFFR_X1 \REGISTERS_reg[7][19]  ( .D(n3450), .CK(CLK), .RN(n427), .Q(n3953), 
        .QN(n2174) );
  DFFR_X1 \REGISTERS_reg[7][18]  ( .D(n3449), .CK(CLK), .RN(n427), .Q(n3952), 
        .QN(n2162) );
  DFFR_X1 \REGISTERS_reg[7][17]  ( .D(n3448), .CK(CLK), .RN(n427), .Q(n3951), 
        .QN(n2150) );
  DFFR_X1 \REGISTERS_reg[7][16]  ( .D(n3447), .CK(CLK), .RN(n427), .Q(n3950), 
        .QN(n2138) );
  DFFR_X1 \REGISTERS_reg[7][15]  ( .D(n3446), .CK(CLK), .RN(n427), .Q(n3949), 
        .QN(n2126) );
  DFFR_X1 \REGISTERS_reg[7][14]  ( .D(n3445), .CK(CLK), .RN(n427), .Q(n3948), 
        .QN(n2114) );
  DFFR_X1 \REGISTERS_reg[7][13]  ( .D(n3444), .CK(CLK), .RN(n427), .Q(n3947), 
        .QN(n2102) );
  DFFR_X1 \REGISTERS_reg[7][12]  ( .D(n3443), .CK(CLK), .RN(n427), .Q(n3946), 
        .QN(n2090) );
  DFFR_X1 \REGISTERS_reg[7][11]  ( .D(n3442), .CK(CLK), .RN(n427), .Q(n3945), 
        .QN(n2078) );
  DFFR_X1 \REGISTERS_reg[7][10]  ( .D(n3441), .CK(CLK), .RN(n427), .Q(n3944), 
        .QN(n2066) );
  DFFR_X1 \REGISTERS_reg[7][9]  ( .D(n3440), .CK(CLK), .RN(n427), .Q(n3943), 
        .QN(n2054) );
  DFFR_X1 \REGISTERS_reg[7][8]  ( .D(n3439), .CK(CLK), .RN(n427), .Q(n3942), 
        .QN(n2042) );
  DFFR_X1 \REGISTERS_reg[7][7]  ( .D(n3438), .CK(CLK), .RN(n428), .Q(n3941), 
        .QN(n2030) );
  DFFR_X1 \REGISTERS_reg[7][6]  ( .D(n3437), .CK(CLK), .RN(n428), .Q(n3940), 
        .QN(n2018) );
  DFFR_X1 \REGISTERS_reg[7][5]  ( .D(n3436), .CK(CLK), .RN(n428), .Q(n3939), 
        .QN(n2006) );
  DFFR_X1 \REGISTERS_reg[7][4]  ( .D(n3435), .CK(CLK), .RN(n428), .Q(n3938), 
        .QN(n1994) );
  DFFR_X1 \REGISTERS_reg[7][3]  ( .D(n3434), .CK(CLK), .RN(n428), .Q(n3937), 
        .QN(n1982) );
  DFFR_X1 \REGISTERS_reg[7][2]  ( .D(n3433), .CK(CLK), .RN(n428), .Q(n3936), 
        .QN(n1970) );
  DFFR_X1 \REGISTERS_reg[7][1]  ( .D(n3432), .CK(CLK), .RN(n428), .Q(n3935), 
        .QN(n1958) );
  DFFR_X1 \REGISTERS_reg[7][0]  ( .D(n3431), .CK(CLK), .RN(n428), .Q(n3934), 
        .QN(n1942) );
  DFFR_X1 \REGISTERS_reg[6][31]  ( .D(n3494), .CK(CLK), .RN(n423), .Q(n3997), 
        .QN(n2330) );
  DFFR_X1 \REGISTERS_reg[6][30]  ( .D(n3493), .CK(CLK), .RN(n423), .Q(n3996), 
        .QN(n2305) );
  DFFR_X1 \REGISTERS_reg[6][29]  ( .D(n3492), .CK(CLK), .RN(n423), .Q(n3995), 
        .QN(n2293) );
  DFFR_X1 \REGISTERS_reg[6][28]  ( .D(n3491), .CK(CLK), .RN(n423), .Q(n3994), 
        .QN(n2281) );
  DFFR_X1 \REGISTERS_reg[6][27]  ( .D(n3490), .CK(CLK), .RN(n423), .Q(n3993), 
        .QN(n2269) );
  DFFR_X1 \REGISTERS_reg[6][26]  ( .D(n3489), .CK(CLK), .RN(n423), .Q(n3992), 
        .QN(n2257) );
  DFFR_X1 \REGISTERS_reg[6][25]  ( .D(n3488), .CK(CLK), .RN(n423), .Q(n3991), 
        .QN(n2245) );
  DFFR_X1 \REGISTERS_reg[6][24]  ( .D(n3487), .CK(CLK), .RN(n423), .Q(n3990), 
        .QN(n2233) );
  DFFR_X1 \REGISTERS_reg[6][23]  ( .D(n3486), .CK(CLK), .RN(n424), .Q(n3989), 
        .QN(n2221) );
  DFFR_X1 \REGISTERS_reg[6][22]  ( .D(n3485), .CK(CLK), .RN(n424), .Q(n3988), 
        .QN(n2209) );
  DFFR_X1 \REGISTERS_reg[6][21]  ( .D(n3484), .CK(CLK), .RN(n424), .Q(n3987), 
        .QN(n2197) );
  DFFR_X1 \REGISTERS_reg[6][20]  ( .D(n3483), .CK(CLK), .RN(n424), .Q(n3986), 
        .QN(n2185) );
  DFFR_X1 \REGISTERS_reg[6][19]  ( .D(n3482), .CK(CLK), .RN(n424), .Q(n3985), 
        .QN(n2173) );
  DFFR_X1 \REGISTERS_reg[6][18]  ( .D(n3481), .CK(CLK), .RN(n424), .Q(n3984), 
        .QN(n2161) );
  DFFR_X1 \REGISTERS_reg[6][17]  ( .D(n3480), .CK(CLK), .RN(n424), .Q(n3983), 
        .QN(n2149) );
  DFFR_X1 \REGISTERS_reg[6][16]  ( .D(n3479), .CK(CLK), .RN(n424), .Q(n3982), 
        .QN(n2137) );
  DFFR_X1 \REGISTERS_reg[6][15]  ( .D(n3478), .CK(CLK), .RN(n424), .Q(n3981), 
        .QN(n2125) );
  DFFR_X1 \REGISTERS_reg[6][14]  ( .D(n3477), .CK(CLK), .RN(n424), .Q(n3980), 
        .QN(n2113) );
  DFFR_X1 \REGISTERS_reg[6][13]  ( .D(n3476), .CK(CLK), .RN(n424), .Q(n3979), 
        .QN(n2101) );
  DFFR_X1 \REGISTERS_reg[6][12]  ( .D(n3475), .CK(CLK), .RN(n424), .Q(n3978), 
        .QN(n2089) );
  DFFR_X1 \REGISTERS_reg[6][11]  ( .D(n3474), .CK(CLK), .RN(n425), .Q(n3977), 
        .QN(n2077) );
  DFFR_X1 \REGISTERS_reg[6][10]  ( .D(n3473), .CK(CLK), .RN(n425), .Q(n3976), 
        .QN(n2065) );
  DFFR_X1 \REGISTERS_reg[6][9]  ( .D(n3472), .CK(CLK), .RN(n425), .Q(n3975), 
        .QN(n2053) );
  DFFR_X1 \REGISTERS_reg[6][8]  ( .D(n3471), .CK(CLK), .RN(n425), .Q(n3974), 
        .QN(n2041) );
  DFFR_X1 \REGISTERS_reg[6][7]  ( .D(n3470), .CK(CLK), .RN(n425), .Q(n3973), 
        .QN(n2029) );
  DFFR_X1 \REGISTERS_reg[6][6]  ( .D(n3469), .CK(CLK), .RN(n425), .Q(n3972), 
        .QN(n2017) );
  DFFR_X1 \REGISTERS_reg[6][5]  ( .D(n3468), .CK(CLK), .RN(n425), .Q(n3971), 
        .QN(n2005) );
  DFFR_X1 \REGISTERS_reg[6][4]  ( .D(n3467), .CK(CLK), .RN(n425), .Q(n3970), 
        .QN(n1993) );
  DFFR_X1 \REGISTERS_reg[6][3]  ( .D(n3466), .CK(CLK), .RN(n425), .Q(n3969), 
        .QN(n1981) );
  DFFR_X1 \REGISTERS_reg[6][2]  ( .D(n3465), .CK(CLK), .RN(n425), .Q(n3968), 
        .QN(n1969) );
  DFFR_X1 \REGISTERS_reg[6][1]  ( .D(n3464), .CK(CLK), .RN(n425), .Q(n3967), 
        .QN(n1957) );
  DFFR_X1 \REGISTERS_reg[6][0]  ( .D(n3463), .CK(CLK), .RN(n425), .Q(n3966), 
        .QN(n1940) );
  DFFR_X1 \REGISTERS_reg[3][31]  ( .D(n3526), .CK(CLK), .RN(n415), .Q(n4061), 
        .QN(n2338) );
  DFFR_X1 \REGISTERS_reg[3][30]  ( .D(n3525), .CK(CLK), .RN(n415), .Q(n4060), 
        .QN(n2309) );
  DFFR_X1 \REGISTERS_reg[3][29]  ( .D(n3524), .CK(CLK), .RN(n415), .Q(n4059), 
        .QN(n2297) );
  DFFR_X1 \REGISTERS_reg[3][28]  ( .D(n3523), .CK(CLK), .RN(n415), .Q(n4058), 
        .QN(n2285) );
  DFFR_X1 \REGISTERS_reg[3][27]  ( .D(n3522), .CK(CLK), .RN(n415), .Q(n4057), 
        .QN(n2273) );
  DFFR_X1 \REGISTERS_reg[3][26]  ( .D(n3521), .CK(CLK), .RN(n415), .Q(n4056), 
        .QN(n2261) );
  DFFR_X1 \REGISTERS_reg[3][25]  ( .D(n3520), .CK(CLK), .RN(n415), .Q(n4055), 
        .QN(n2249) );
  DFFR_X1 \REGISTERS_reg[3][24]  ( .D(n3519), .CK(CLK), .RN(n415), .Q(n4054), 
        .QN(n2237) );
  DFFR_X1 \REGISTERS_reg[3][23]  ( .D(n3518), .CK(CLK), .RN(n416), .Q(n4053), 
        .QN(n2225) );
  DFFR_X1 \REGISTERS_reg[3][22]  ( .D(n3517), .CK(CLK), .RN(n416), .Q(n4052), 
        .QN(n2213) );
  DFFR_X1 \REGISTERS_reg[3][21]  ( .D(n3516), .CK(CLK), .RN(n416), .Q(n4051), 
        .QN(n2201) );
  DFFR_X1 \REGISTERS_reg[3][20]  ( .D(n3515), .CK(CLK), .RN(n416), .Q(n4050), 
        .QN(n2189) );
  DFFR_X1 \REGISTERS_reg[3][19]  ( .D(n3514), .CK(CLK), .RN(n416), .Q(n4049), 
        .QN(n2177) );
  DFFR_X1 \REGISTERS_reg[3][18]  ( .D(n3513), .CK(CLK), .RN(n416), .Q(n4048), 
        .QN(n2165) );
  DFFR_X1 \REGISTERS_reg[3][17]  ( .D(n3512), .CK(CLK), .RN(n416), .Q(n4047), 
        .QN(n2153) );
  DFFR_X1 \REGISTERS_reg[3][16]  ( .D(n3511), .CK(CLK), .RN(n416), .Q(n4046), 
        .QN(n2141) );
  DFFR_X1 \REGISTERS_reg[3][15]  ( .D(n3510), .CK(CLK), .RN(n416), .Q(n4045), 
        .QN(n2129) );
  DFFR_X1 \REGISTERS_reg[3][14]  ( .D(n3509), .CK(CLK), .RN(n416), .Q(n4044), 
        .QN(n2117) );
  DFFR_X1 \REGISTERS_reg[3][13]  ( .D(n3508), .CK(CLK), .RN(n416), .Q(n4043), 
        .QN(n2105) );
  DFFR_X1 \REGISTERS_reg[3][12]  ( .D(n3507), .CK(CLK), .RN(n416), .Q(n4042), 
        .QN(n2093) );
  DFFR_X1 \REGISTERS_reg[3][11]  ( .D(n3506), .CK(CLK), .RN(n417), .Q(n4041), 
        .QN(n2081) );
  DFFR_X1 \REGISTERS_reg[3][10]  ( .D(n3505), .CK(CLK), .RN(n417), .Q(n4040), 
        .QN(n2069) );
  DFFR_X1 \REGISTERS_reg[3][9]  ( .D(n3504), .CK(CLK), .RN(n417), .Q(n4039), 
        .QN(n2057) );
  DFFR_X1 \REGISTERS_reg[3][8]  ( .D(n3503), .CK(CLK), .RN(n417), .Q(n4038), 
        .QN(n2045) );
  DFFR_X1 \REGISTERS_reg[3][7]  ( .D(n3502), .CK(CLK), .RN(n417), .Q(n4037), 
        .QN(n2033) );
  DFFR_X1 \REGISTERS_reg[3][6]  ( .D(n3501), .CK(CLK), .RN(n417), .Q(n4036), 
        .QN(n2021) );
  DFFR_X1 \REGISTERS_reg[3][5]  ( .D(n3500), .CK(CLK), .RN(n417), .Q(n4035), 
        .QN(n2009) );
  DFFR_X1 \REGISTERS_reg[3][4]  ( .D(n3499), .CK(CLK), .RN(n417), .Q(n4034), 
        .QN(n1997) );
  DFFR_X1 \REGISTERS_reg[3][3]  ( .D(n3498), .CK(CLK), .RN(n417), .Q(n4033), 
        .QN(n1985) );
  DFFR_X1 \REGISTERS_reg[3][2]  ( .D(n3497), .CK(CLK), .RN(n417), .Q(n4032), 
        .QN(n1973) );
  DFFR_X1 \REGISTERS_reg[3][1]  ( .D(n3496), .CK(CLK), .RN(n417), .Q(n4031), 
        .QN(n1961) );
  DFFR_X1 \REGISTERS_reg[3][0]  ( .D(n3495), .CK(CLK), .RN(n417), .Q(n4030), 
        .QN(n1948) );
  DFFR_X1 \REGISTERS_reg[2][31]  ( .D(n3558), .CK(CLK), .RN(n412), .Q(n4093), 
        .QN(n2337) );
  DFFR_X1 \REGISTERS_reg[2][30]  ( .D(n3557), .CK(CLK), .RN(n412), .Q(n4092), 
        .QN(n2308) );
  DFFR_X1 \REGISTERS_reg[2][29]  ( .D(n3556), .CK(CLK), .RN(n412), .Q(n4091), 
        .QN(n2296) );
  DFFR_X1 \REGISTERS_reg[2][28]  ( .D(n3555), .CK(CLK), .RN(n412), .Q(n4090), 
        .QN(n2284) );
  DFFR_X1 \REGISTERS_reg[2][27]  ( .D(n3554), .CK(CLK), .RN(n413), .Q(n4089), 
        .QN(n2272) );
  DFFR_X1 \REGISTERS_reg[2][26]  ( .D(n3553), .CK(CLK), .RN(n413), .Q(n4088), 
        .QN(n2260) );
  DFFR_X1 \REGISTERS_reg[2][25]  ( .D(n3552), .CK(CLK), .RN(n413), .Q(n4087), 
        .QN(n2248) );
  DFFR_X1 \REGISTERS_reg[2][24]  ( .D(n3551), .CK(CLK), .RN(n413), .Q(n4086), 
        .QN(n2236) );
  DFFR_X1 \REGISTERS_reg[2][23]  ( .D(n3550), .CK(CLK), .RN(n413), .Q(n4085), 
        .QN(n2224) );
  DFFR_X1 \REGISTERS_reg[2][22]  ( .D(n3549), .CK(CLK), .RN(n413), .Q(n4084), 
        .QN(n2212) );
  DFFR_X1 \REGISTERS_reg[2][21]  ( .D(n3548), .CK(CLK), .RN(n413), .Q(n4083), 
        .QN(n2200) );
  DFFR_X1 \REGISTERS_reg[2][20]  ( .D(n3547), .CK(CLK), .RN(n413), .Q(n4082), 
        .QN(n2188) );
  DFFR_X1 \REGISTERS_reg[2][19]  ( .D(n3546), .CK(CLK), .RN(n413), .Q(n4081), 
        .QN(n2176) );
  DFFR_X1 \REGISTERS_reg[2][18]  ( .D(n3545), .CK(CLK), .RN(n413), .Q(n4080), 
        .QN(n2164) );
  DFFR_X1 \REGISTERS_reg[2][17]  ( .D(n3544), .CK(CLK), .RN(n413), .Q(n4079), 
        .QN(n2152) );
  DFFR_X1 \REGISTERS_reg[2][16]  ( .D(n3543), .CK(CLK), .RN(n413), .Q(n4078), 
        .QN(n2140) );
  DFFR_X1 \REGISTERS_reg[2][15]  ( .D(n3542), .CK(CLK), .RN(n414), .Q(n4077), 
        .QN(n2128) );
  DFFR_X1 \REGISTERS_reg[2][14]  ( .D(n3541), .CK(CLK), .RN(n414), .Q(n4076), 
        .QN(n2116) );
  DFFR_X1 \REGISTERS_reg[2][13]  ( .D(n3540), .CK(CLK), .RN(n414), .Q(n4075), 
        .QN(n2104) );
  DFFR_X1 \REGISTERS_reg[2][12]  ( .D(n3539), .CK(CLK), .RN(n414), .Q(n4074), 
        .QN(n2092) );
  DFFR_X1 \REGISTERS_reg[2][11]  ( .D(n3538), .CK(CLK), .RN(n414), .Q(n4073), 
        .QN(n2080) );
  DFFR_X1 \REGISTERS_reg[2][10]  ( .D(n3537), .CK(CLK), .RN(n414), .Q(n4072), 
        .QN(n2068) );
  DFFR_X1 \REGISTERS_reg[2][9]  ( .D(n3536), .CK(CLK), .RN(n414), .Q(n4071), 
        .QN(n2056) );
  DFFR_X1 \REGISTERS_reg[2][8]  ( .D(n3535), .CK(CLK), .RN(n414), .Q(n4070), 
        .QN(n2044) );
  DFFR_X1 \REGISTERS_reg[2][7]  ( .D(n3534), .CK(CLK), .RN(n414), .Q(n4069), 
        .QN(n2032) );
  DFFR_X1 \REGISTERS_reg[2][6]  ( .D(n3533), .CK(CLK), .RN(n414), .Q(n4068), 
        .QN(n2020) );
  DFFR_X1 \REGISTERS_reg[2][5]  ( .D(n3532), .CK(CLK), .RN(n414), .Q(n4067), 
        .QN(n2008) );
  DFFR_X1 \REGISTERS_reg[2][4]  ( .D(n3531), .CK(CLK), .RN(n414), .Q(n4066), 
        .QN(n1996) );
  DFFR_X1 \REGISTERS_reg[2][3]  ( .D(n3530), .CK(CLK), .RN(n415), .Q(n4065), 
        .QN(n1984) );
  DFFR_X1 \REGISTERS_reg[2][2]  ( .D(n3529), .CK(CLK), .RN(n415), .Q(n4064), 
        .QN(n1972) );
  DFFR_X1 \REGISTERS_reg[2][1]  ( .D(n3528), .CK(CLK), .RN(n415), .Q(n4063), 
        .QN(n1960) );
  DFFR_X1 \REGISTERS_reg[2][0]  ( .D(n3527), .CK(CLK), .RN(n415), .Q(n4062), 
        .QN(n1946) );
  DFFR_X1 \REGISTERS_reg[28][31]  ( .D(n3110), .CK(CLK), .RN(n482), .Q(n2813)
         );
  DFFR_X1 \REGISTERS_reg[28][30]  ( .D(n3109), .CK(CLK), .RN(n482), .Q(n2812)
         );
  DFFR_X1 \REGISTERS_reg[28][29]  ( .D(n3108), .CK(CLK), .RN(n482), .Q(n2811)
         );
  DFFR_X1 \REGISTERS_reg[28][28]  ( .D(n3107), .CK(CLK), .RN(n482), .Q(n2810)
         );
  DFFR_X1 \REGISTERS_reg[28][27]  ( .D(n3106), .CK(CLK), .RN(n482), .Q(n2809)
         );
  DFFR_X1 \REGISTERS_reg[28][26]  ( .D(n3105), .CK(CLK), .RN(n482), .Q(n2808)
         );
  DFFR_X1 \REGISTERS_reg[28][25]  ( .D(n3104), .CK(CLK), .RN(n482), .Q(n2807)
         );
  DFFR_X1 \REGISTERS_reg[28][24]  ( .D(n3103), .CK(CLK), .RN(n482), .Q(n2806)
         );
  DFFR_X1 \REGISTERS_reg[28][23]  ( .D(n3102), .CK(CLK), .RN(n482), .Q(n2805)
         );
  DFFR_X1 \REGISTERS_reg[28][22]  ( .D(n3101), .CK(CLK), .RN(n482), .Q(n2804)
         );
  DFFR_X1 \REGISTERS_reg[28][21]  ( .D(n3100), .CK(CLK), .RN(n482), .Q(n2803)
         );
  DFFR_X1 \REGISTERS_reg[28][20]  ( .D(n3099), .CK(CLK), .RN(n482), .Q(n2802)
         );
  DFFR_X1 \REGISTERS_reg[28][19]  ( .D(n3098), .CK(CLK), .RN(n483), .Q(n2801)
         );
  DFFR_X1 \REGISTERS_reg[28][18]  ( .D(n3097), .CK(CLK), .RN(n483), .Q(n2800)
         );
  DFFR_X1 \REGISTERS_reg[28][17]  ( .D(n3096), .CK(CLK), .RN(n483), .Q(n2799)
         );
  DFFR_X1 \REGISTERS_reg[28][16]  ( .D(n3095), .CK(CLK), .RN(n483), .Q(n2798)
         );
  DFFR_X1 \REGISTERS_reg[28][15]  ( .D(n3094), .CK(CLK), .RN(n483), .Q(n2797)
         );
  DFFR_X1 \REGISTERS_reg[28][14]  ( .D(n3093), .CK(CLK), .RN(n483), .Q(n2796)
         );
  DFFR_X1 \REGISTERS_reg[28][13]  ( .D(n3092), .CK(CLK), .RN(n483), .Q(n2795)
         );
  DFFR_X1 \REGISTERS_reg[28][12]  ( .D(n3091), .CK(CLK), .RN(n483), .Q(n2794)
         );
  DFFR_X1 \REGISTERS_reg[28][11]  ( .D(n3090), .CK(CLK), .RN(n483), .Q(n2793)
         );
  DFFR_X1 \REGISTERS_reg[28][10]  ( .D(n3089), .CK(CLK), .RN(n483), .Q(n2792)
         );
  DFFR_X1 \REGISTERS_reg[28][9]  ( .D(n3088), .CK(CLK), .RN(n483), .Q(n2791)
         );
  DFFR_X1 \REGISTERS_reg[28][8]  ( .D(n3087), .CK(CLK), .RN(n483), .Q(n2790)
         );
  DFFR_X1 \REGISTERS_reg[28][7]  ( .D(n3086), .CK(CLK), .RN(n484), .Q(n2789)
         );
  DFFR_X1 \REGISTERS_reg[28][6]  ( .D(n3085), .CK(CLK), .RN(n484), .Q(n2788)
         );
  DFFR_X1 \REGISTERS_reg[28][5]  ( .D(n3084), .CK(CLK), .RN(n484), .Q(n2787)
         );
  DFFR_X1 \REGISTERS_reg[28][4]  ( .D(n3083), .CK(CLK), .RN(n484), .Q(n2786)
         );
  DFFR_X1 \REGISTERS_reg[28][3]  ( .D(n3082), .CK(CLK), .RN(n484), .Q(n2785)
         );
  DFFR_X1 \REGISTERS_reg[28][2]  ( .D(n3081), .CK(CLK), .RN(n484), .Q(n2784)
         );
  DFFR_X1 \REGISTERS_reg[28][1]  ( .D(n3080), .CK(CLK), .RN(n484), .Q(n2783)
         );
  DFFR_X1 \REGISTERS_reg[28][0]  ( .D(n3079), .CK(CLK), .RN(n484), .Q(n2782)
         );
  DFFR_X1 \REGISTERS_reg[18][31]  ( .D(n3302), .CK(CLK), .RN(n455), .Q(n3645)
         );
  DFFR_X1 \REGISTERS_reg[27][31]  ( .D(n4541), .CK(CLK), .RN(RST), .Q(n1518)
         );
  DFFR_X1 \REGISTERS_reg[27][30]  ( .D(n4540), .CK(CLK), .RN(n479), .Q(n1517)
         );
  DFFR_X1 \REGISTERS_reg[27][29]  ( .D(n4539), .CK(CLK), .RN(n479), .Q(n1516)
         );
  DFFR_X1 \REGISTERS_reg[27][28]  ( .D(n4538), .CK(CLK), .RN(n479), .Q(n1515)
         );
  DFFR_X1 \REGISTERS_reg[27][27]  ( .D(n4537), .CK(CLK), .RN(n479), .Q(n1514)
         );
  DFFR_X1 \REGISTERS_reg[27][26]  ( .D(n4536), .CK(CLK), .RN(n479), .Q(n1513)
         );
  DFFR_X1 \REGISTERS_reg[27][25]  ( .D(n4535), .CK(CLK), .RN(n479), .Q(n1512)
         );
  DFFR_X1 \REGISTERS_reg[27][24]  ( .D(n4534), .CK(CLK), .RN(n479), .Q(n1511)
         );
  DFFR_X1 \REGISTERS_reg[27][23]  ( .D(n4533), .CK(CLK), .RN(n480), .Q(n1510)
         );
  DFFR_X1 \REGISTERS_reg[27][22]  ( .D(n4532), .CK(CLK), .RN(n480), .Q(n1509)
         );
  DFFR_X1 \REGISTERS_reg[27][21]  ( .D(n4531), .CK(CLK), .RN(n480), .Q(n1508)
         );
  DFFR_X1 \REGISTERS_reg[27][20]  ( .D(n4530), .CK(CLK), .RN(n480), .Q(n1507)
         );
  DFFR_X1 \REGISTERS_reg[27][19]  ( .D(n4529), .CK(CLK), .RN(n480), .Q(n1506)
         );
  DFFR_X1 \REGISTERS_reg[27][18]  ( .D(n4528), .CK(CLK), .RN(n480), .Q(n1505)
         );
  DFFR_X1 \REGISTERS_reg[27][17]  ( .D(n4527), .CK(CLK), .RN(n480), .Q(n1504)
         );
  DFFR_X1 \REGISTERS_reg[27][16]  ( .D(n4526), .CK(CLK), .RN(n480), .Q(n1503)
         );
  DFFR_X1 \REGISTERS_reg[27][15]  ( .D(n4525), .CK(CLK), .RN(n480), .Q(n1502)
         );
  DFFR_X1 \REGISTERS_reg[27][14]  ( .D(n4524), .CK(CLK), .RN(n480), .Q(n1501)
         );
  DFFR_X1 \REGISTERS_reg[27][13]  ( .D(n4523), .CK(CLK), .RN(n480), .Q(n1500)
         );
  DFFR_X1 \REGISTERS_reg[27][12]  ( .D(n4522), .CK(CLK), .RN(n480), .Q(n1499)
         );
  DFFR_X1 \REGISTERS_reg[27][11]  ( .D(n4521), .CK(CLK), .RN(n481), .Q(n1498)
         );
  DFFR_X1 \REGISTERS_reg[27][10]  ( .D(n4520), .CK(CLK), .RN(n481), .Q(n1497)
         );
  DFFR_X1 \REGISTERS_reg[27][9]  ( .D(n4519), .CK(CLK), .RN(n481), .Q(n1496)
         );
  DFFR_X1 \REGISTERS_reg[27][8]  ( .D(n4518), .CK(CLK), .RN(n481), .Q(n1495)
         );
  DFFR_X1 \REGISTERS_reg[27][7]  ( .D(n4517), .CK(CLK), .RN(n481), .Q(n1494)
         );
  DFFR_X1 \REGISTERS_reg[27][6]  ( .D(n4516), .CK(CLK), .RN(n481), .Q(n1493)
         );
  DFFR_X1 \REGISTERS_reg[27][5]  ( .D(n4515), .CK(CLK), .RN(n481), .Q(n1492)
         );
  DFFR_X1 \REGISTERS_reg[27][4]  ( .D(n4514), .CK(CLK), .RN(n481), .Q(n1491)
         );
  DFFR_X1 \REGISTERS_reg[27][3]  ( .D(n4513), .CK(CLK), .RN(n481), .Q(n1490)
         );
  DFFR_X1 \REGISTERS_reg[27][2]  ( .D(n4512), .CK(CLK), .RN(n481), .Q(n1489)
         );
  DFFR_X1 \REGISTERS_reg[27][1]  ( .D(n4511), .CK(CLK), .RN(n481), .Q(n1488)
         );
  DFFR_X1 \REGISTERS_reg[27][0]  ( .D(n4510), .CK(CLK), .RN(n481), .Q(n1487)
         );
  DFFR_X1 \REGISTERS_reg[4][31]  ( .D(n4317), .CK(CLK), .RN(n418), .Q(n1874)
         );
  DFFR_X1 \REGISTERS_reg[4][30]  ( .D(n4316), .CK(CLK), .RN(n418), .Q(n1873)
         );
  DFFR_X1 \REGISTERS_reg[4][29]  ( .D(n4315), .CK(CLK), .RN(n418), .Q(n1872)
         );
  DFFR_X1 \REGISTERS_reg[4][28]  ( .D(n4314), .CK(CLK), .RN(n418), .Q(n1871)
         );
  DFFR_X1 \REGISTERS_reg[4][27]  ( .D(n4313), .CK(CLK), .RN(n418), .Q(n1870)
         );
  DFFR_X1 \REGISTERS_reg[4][26]  ( .D(n4312), .CK(CLK), .RN(n418), .Q(n1869)
         );
  DFFR_X1 \REGISTERS_reg[4][25]  ( .D(n4311), .CK(CLK), .RN(n418), .Q(n1868)
         );
  DFFR_X1 \REGISTERS_reg[4][24]  ( .D(n4310), .CK(CLK), .RN(n418), .Q(n1867)
         );
  DFFR_X1 \REGISTERS_reg[4][23]  ( .D(n4309), .CK(CLK), .RN(n418), .Q(n1866)
         );
  DFFR_X1 \REGISTERS_reg[4][22]  ( .D(n4308), .CK(CLK), .RN(n418), .Q(n1865)
         );
  DFFR_X1 \REGISTERS_reg[4][21]  ( .D(n4307), .CK(CLK), .RN(n418), .Q(n1864)
         );
  DFFR_X1 \REGISTERS_reg[4][20]  ( .D(n4306), .CK(CLK), .RN(n418), .Q(n1863)
         );
  DFFR_X1 \REGISTERS_reg[4][19]  ( .D(n4305), .CK(CLK), .RN(n419), .Q(n1862)
         );
  DFFR_X1 \REGISTERS_reg[4][18]  ( .D(n4304), .CK(CLK), .RN(n419), .Q(n1861)
         );
  DFFR_X1 \REGISTERS_reg[4][17]  ( .D(n4303), .CK(CLK), .RN(n419), .Q(n1860)
         );
  DFFR_X1 \REGISTERS_reg[4][16]  ( .D(n4302), .CK(CLK), .RN(n419), .Q(n1859)
         );
  DFFR_X1 \REGISTERS_reg[4][15]  ( .D(n4301), .CK(CLK), .RN(n419), .Q(n1858)
         );
  DFFR_X1 \REGISTERS_reg[4][14]  ( .D(n4300), .CK(CLK), .RN(n419), .Q(n1857)
         );
  DFFR_X1 \REGISTERS_reg[4][13]  ( .D(n4299), .CK(CLK), .RN(n419), .Q(n1856)
         );
  DFFR_X1 \REGISTERS_reg[4][12]  ( .D(n4298), .CK(CLK), .RN(n419), .Q(n1855)
         );
  DFFR_X1 \REGISTERS_reg[4][11]  ( .D(n4297), .CK(CLK), .RN(n419), .Q(n1854)
         );
  DFFR_X1 \REGISTERS_reg[4][10]  ( .D(n4296), .CK(CLK), .RN(n419), .Q(n1853)
         );
  DFFR_X1 \REGISTERS_reg[4][9]  ( .D(n4295), .CK(CLK), .RN(n419), .Q(n1852) );
  DFFR_X1 \REGISTERS_reg[4][8]  ( .D(n4294), .CK(CLK), .RN(n419), .Q(n1851) );
  DFFR_X1 \REGISTERS_reg[4][7]  ( .D(n4293), .CK(CLK), .RN(n420), .Q(n1850) );
  DFFR_X1 \REGISTERS_reg[4][6]  ( .D(n4292), .CK(CLK), .RN(n420), .Q(n1849) );
  DFFR_X1 \REGISTERS_reg[4][5]  ( .D(n4291), .CK(CLK), .RN(n420), .Q(n1848) );
  DFFR_X1 \REGISTERS_reg[4][4]  ( .D(n4290), .CK(CLK), .RN(n420), .Q(n1847) );
  DFFR_X1 \REGISTERS_reg[4][3]  ( .D(n4289), .CK(CLK), .RN(n420), .Q(n1846) );
  DFFR_X1 \REGISTERS_reg[4][2]  ( .D(n4288), .CK(CLK), .RN(n420), .Q(n1845) );
  DFFR_X1 \REGISTERS_reg[4][1]  ( .D(n4287), .CK(CLK), .RN(n420), .Q(n1844) );
  DFFR_X1 \REGISTERS_reg[4][0]  ( .D(n4286), .CK(CLK), .RN(n420), .Q(n1843) );
  DFFR_X1 \REGISTERS_reg[26][31]  ( .D(n4509), .CK(CLK), .RN(n476), .Q(n1550)
         );
  DFFR_X1 \REGISTERS_reg[26][30]  ( .D(n4508), .CK(CLK), .RN(n476), .Q(n1549)
         );
  DFFR_X1 \REGISTERS_reg[26][29]  ( .D(n4507), .CK(CLK), .RN(n476), .Q(n1548)
         );
  DFFR_X1 \REGISTERS_reg[26][28]  ( .D(n4506), .CK(CLK), .RN(n476), .Q(n1547)
         );
  DFFR_X1 \REGISTERS_reg[26][27]  ( .D(n4505), .CK(CLK), .RN(n477), .Q(n1546)
         );
  DFFR_X1 \REGISTERS_reg[26][26]  ( .D(n4504), .CK(CLK), .RN(n477), .Q(n1545)
         );
  DFFR_X1 \REGISTERS_reg[26][25]  ( .D(n4503), .CK(CLK), .RN(n477), .Q(n1544)
         );
  DFFR_X1 \REGISTERS_reg[26][24]  ( .D(n4502), .CK(CLK), .RN(n477), .Q(n1543)
         );
  DFFR_X1 \REGISTERS_reg[26][23]  ( .D(n4501), .CK(CLK), .RN(n477), .Q(n1542)
         );
  DFFR_X1 \REGISTERS_reg[26][22]  ( .D(n4500), .CK(CLK), .RN(n477), .Q(n1541)
         );
  DFFR_X1 \REGISTERS_reg[26][21]  ( .D(n4499), .CK(CLK), .RN(n477), .Q(n1540)
         );
  DFFR_X1 \REGISTERS_reg[26][20]  ( .D(n4498), .CK(CLK), .RN(n477), .Q(n1539)
         );
  DFFR_X1 \REGISTERS_reg[26][19]  ( .D(n4497), .CK(CLK), .RN(n477), .Q(n1538)
         );
  DFFR_X1 \REGISTERS_reg[26][18]  ( .D(n4496), .CK(CLK), .RN(n477), .Q(n1537)
         );
  DFFR_X1 \REGISTERS_reg[26][17]  ( .D(n4495), .CK(CLK), .RN(n477), .Q(n1536)
         );
  DFFR_X1 \REGISTERS_reg[26][16]  ( .D(n4494), .CK(CLK), .RN(n477), .Q(n1535)
         );
  DFFR_X1 \REGISTERS_reg[26][15]  ( .D(n4493), .CK(CLK), .RN(n478), .Q(n1534)
         );
  DFFR_X1 \REGISTERS_reg[26][14]  ( .D(n4492), .CK(CLK), .RN(n478), .Q(n1533)
         );
  DFFR_X1 \REGISTERS_reg[26][13]  ( .D(n4491), .CK(CLK), .RN(n478), .Q(n1532)
         );
  DFFR_X1 \REGISTERS_reg[26][12]  ( .D(n4490), .CK(CLK), .RN(n478), .Q(n1531)
         );
  DFFR_X1 \REGISTERS_reg[26][11]  ( .D(n4489), .CK(CLK), .RN(n478), .Q(n1530)
         );
  DFFR_X1 \REGISTERS_reg[26][10]  ( .D(n4488), .CK(CLK), .RN(n478), .Q(n1529)
         );
  DFFR_X1 \REGISTERS_reg[26][9]  ( .D(n4487), .CK(CLK), .RN(n478), .Q(n1528)
         );
  DFFR_X1 \REGISTERS_reg[26][8]  ( .D(n4486), .CK(CLK), .RN(n478), .Q(n1527)
         );
  DFFR_X1 \REGISTERS_reg[26][7]  ( .D(n4485), .CK(CLK), .RN(n478), .Q(n1526)
         );
  DFFR_X1 \REGISTERS_reg[26][6]  ( .D(n4484), .CK(CLK), .RN(n478), .Q(n1525)
         );
  DFFR_X1 \REGISTERS_reg[26][5]  ( .D(n4483), .CK(CLK), .RN(n478), .Q(n1524)
         );
  DFFR_X1 \REGISTERS_reg[26][4]  ( .D(n4482), .CK(CLK), .RN(n478), .Q(n1523)
         );
  DFFR_X1 \REGISTERS_reg[26][3]  ( .D(n4481), .CK(CLK), .RN(n479), .Q(n1522)
         );
  DFFR_X1 \REGISTERS_reg[26][2]  ( .D(n4480), .CK(CLK), .RN(n479), .Q(n1521)
         );
  DFFR_X1 \REGISTERS_reg[26][1]  ( .D(n4479), .CK(CLK), .RN(n479), .Q(n1520)
         );
  DFFR_X1 \REGISTERS_reg[26][0]  ( .D(n4478), .CK(CLK), .RN(n479), .Q(n1519)
         );
  DFFR_X1 \REGISTERS_reg[17][31]  ( .D(n4413), .CK(CLK), .RN(n452), .Q(n1648)
         );
  DFFR_X1 \REGISTERS_reg[17][30]  ( .D(n4412), .CK(CLK), .RN(n452), .Q(n1647)
         );
  DFFR_X1 \REGISTERS_reg[17][29]  ( .D(n4411), .CK(CLK), .RN(n452), .Q(n1646)
         );
  DFFR_X1 \REGISTERS_reg[17][28]  ( .D(n4410), .CK(CLK), .RN(n452), .Q(n1645)
         );
  DFFR_X1 \REGISTERS_reg[17][27]  ( .D(n4409), .CK(CLK), .RN(n453), .Q(n1644)
         );
  DFFR_X1 \REGISTERS_reg[17][26]  ( .D(n4408), .CK(CLK), .RN(n453), .Q(n1643)
         );
  DFFR_X1 \REGISTERS_reg[17][25]  ( .D(n4407), .CK(CLK), .RN(n453), .Q(n1642)
         );
  DFFR_X1 \REGISTERS_reg[17][24]  ( .D(n4406), .CK(CLK), .RN(n453), .Q(n1641)
         );
  DFFR_X1 \REGISTERS_reg[17][23]  ( .D(n4405), .CK(CLK), .RN(n453), .Q(n1640)
         );
  DFFR_X1 \REGISTERS_reg[17][22]  ( .D(n4404), .CK(CLK), .RN(n453), .Q(n1639)
         );
  DFFR_X1 \REGISTERS_reg[17][21]  ( .D(n4403), .CK(CLK), .RN(n453), .Q(n1638)
         );
  DFFR_X1 \REGISTERS_reg[17][20]  ( .D(n4402), .CK(CLK), .RN(n453), .Q(n1637)
         );
  DFFR_X1 \REGISTERS_reg[17][19]  ( .D(n4401), .CK(CLK), .RN(n453), .Q(n1636)
         );
  DFFR_X1 \REGISTERS_reg[17][18]  ( .D(n4400), .CK(CLK), .RN(n453), .Q(n1635)
         );
  DFFR_X1 \REGISTERS_reg[17][17]  ( .D(n4399), .CK(CLK), .RN(n453), .Q(n1634)
         );
  DFFR_X1 \REGISTERS_reg[17][16]  ( .D(n4398), .CK(CLK), .RN(n453), .Q(n1633)
         );
  DFFR_X1 \REGISTERS_reg[17][15]  ( .D(n4397), .CK(CLK), .RN(n454), .Q(n1632)
         );
  DFFR_X1 \REGISTERS_reg[17][14]  ( .D(n4396), .CK(CLK), .RN(n454), .Q(n1631)
         );
  DFFR_X1 \REGISTERS_reg[17][13]  ( .D(n4395), .CK(CLK), .RN(n454), .Q(n1630)
         );
  DFFR_X1 \REGISTERS_reg[17][12]  ( .D(n4394), .CK(CLK), .RN(n454), .Q(n1629)
         );
  DFFR_X1 \REGISTERS_reg[17][11]  ( .D(n4393), .CK(CLK), .RN(n454), .Q(n1628)
         );
  DFFR_X1 \REGISTERS_reg[17][10]  ( .D(n4392), .CK(CLK), .RN(n454), .Q(n1627)
         );
  DFFR_X1 \REGISTERS_reg[17][9]  ( .D(n4391), .CK(CLK), .RN(n454), .Q(n1626)
         );
  DFFR_X1 \REGISTERS_reg[17][8]  ( .D(n4390), .CK(CLK), .RN(n454), .Q(n1625)
         );
  DFFR_X1 \REGISTERS_reg[17][7]  ( .D(n4389), .CK(CLK), .RN(n454), .Q(n1624)
         );
  DFFR_X1 \REGISTERS_reg[17][6]  ( .D(n4388), .CK(CLK), .RN(n454), .Q(n1623)
         );
  DFFR_X1 \REGISTERS_reg[17][5]  ( .D(n4387), .CK(CLK), .RN(n454), .Q(n1622)
         );
  DFFR_X1 \REGISTERS_reg[17][4]  ( .D(n4386), .CK(CLK), .RN(n454), .Q(n1621)
         );
  DFFR_X1 \REGISTERS_reg[17][3]  ( .D(n4385), .CK(CLK), .RN(n455), .Q(n1620)
         );
  DFFR_X1 \REGISTERS_reg[17][2]  ( .D(n4384), .CK(CLK), .RN(n455), .Q(n1619)
         );
  DFFR_X1 \REGISTERS_reg[17][1]  ( .D(n4383), .CK(CLK), .RN(n455), .Q(n1618)
         );
  DFFR_X1 \REGISTERS_reg[17][0]  ( .D(n4382), .CK(CLK), .RN(n455), .Q(n1617)
         );
  DFFR_X1 \REGISTERS_reg[5][31]  ( .D(n4349), .CK(CLK), .RN(n420), .Q(n1842), 
        .QN(n4029) );
  DFFR_X1 \REGISTERS_reg[5][30]  ( .D(n4348), .CK(CLK), .RN(n420), .Q(n1841), 
        .QN(n4028) );
  DFFR_X1 \REGISTERS_reg[5][29]  ( .D(n4347), .CK(CLK), .RN(n420), .Q(n1840), 
        .QN(n4027) );
  DFFR_X1 \REGISTERS_reg[5][28]  ( .D(n4346), .CK(CLK), .RN(n420), .Q(n1839), 
        .QN(n4026) );
  DFFR_X1 \REGISTERS_reg[5][27]  ( .D(n4345), .CK(CLK), .RN(n421), .Q(n1838), 
        .QN(n4025) );
  DFFR_X1 \REGISTERS_reg[5][26]  ( .D(n4344), .CK(CLK), .RN(n421), .Q(n1837), 
        .QN(n4024) );
  DFFR_X1 \REGISTERS_reg[5][25]  ( .D(n4343), .CK(CLK), .RN(n421), .Q(n1836), 
        .QN(n4023) );
  DFFR_X1 \REGISTERS_reg[5][24]  ( .D(n4342), .CK(CLK), .RN(n421), .Q(n1835), 
        .QN(n4022) );
  DFFR_X1 \REGISTERS_reg[5][23]  ( .D(n4341), .CK(CLK), .RN(n421), .Q(n1834), 
        .QN(n4021) );
  DFFR_X1 \REGISTERS_reg[5][22]  ( .D(n4340), .CK(CLK), .RN(n421), .Q(n1833), 
        .QN(n4020) );
  DFFR_X1 \REGISTERS_reg[5][21]  ( .D(n4339), .CK(CLK), .RN(n421), .Q(n1832), 
        .QN(n4019) );
  DFFR_X1 \REGISTERS_reg[5][20]  ( .D(n4338), .CK(CLK), .RN(n421), .Q(n1831), 
        .QN(n4018) );
  DFFR_X1 \REGISTERS_reg[5][19]  ( .D(n4337), .CK(CLK), .RN(n421), .Q(n1830), 
        .QN(n4017) );
  DFFR_X1 \REGISTERS_reg[5][18]  ( .D(n4336), .CK(CLK), .RN(n421), .Q(n1829), 
        .QN(n4016) );
  DFFR_X1 \REGISTERS_reg[5][17]  ( .D(n4335), .CK(CLK), .RN(n421), .Q(n1828), 
        .QN(n4015) );
  DFFR_X1 \REGISTERS_reg[5][16]  ( .D(n4334), .CK(CLK), .RN(n421), .Q(n1827), 
        .QN(n4014) );
  DFFR_X1 \REGISTERS_reg[5][15]  ( .D(n4333), .CK(CLK), .RN(n422), .Q(n1826), 
        .QN(n4013) );
  DFFR_X1 \REGISTERS_reg[5][14]  ( .D(n4332), .CK(CLK), .RN(n422), .Q(n1825), 
        .QN(n4012) );
  DFFR_X1 \REGISTERS_reg[5][13]  ( .D(n4331), .CK(CLK), .RN(n422), .Q(n1824), 
        .QN(n4011) );
  DFFR_X1 \REGISTERS_reg[5][12]  ( .D(n4330), .CK(CLK), .RN(n422), .Q(n1823), 
        .QN(n4010) );
  DFFR_X1 \REGISTERS_reg[5][11]  ( .D(n4329), .CK(CLK), .RN(n422), .Q(n1822), 
        .QN(n4009) );
  DFFR_X1 \REGISTERS_reg[5][10]  ( .D(n4328), .CK(CLK), .RN(n422), .Q(n1821), 
        .QN(n4008) );
  DFFR_X1 \REGISTERS_reg[5][9]  ( .D(n4327), .CK(CLK), .RN(n422), .Q(n1820), 
        .QN(n4007) );
  DFFR_X1 \REGISTERS_reg[5][8]  ( .D(n4326), .CK(CLK), .RN(n422), .Q(n1819), 
        .QN(n4006) );
  DFFR_X1 \REGISTERS_reg[5][7]  ( .D(n4325), .CK(CLK), .RN(n422), .Q(n1818), 
        .QN(n4005) );
  DFFR_X1 \REGISTERS_reg[5][6]  ( .D(n4324), .CK(CLK), .RN(n422), .Q(n1817), 
        .QN(n4004) );
  DFFR_X1 \REGISTERS_reg[5][5]  ( .D(n4323), .CK(CLK), .RN(n422), .Q(n1816), 
        .QN(n4003) );
  DFFR_X1 \REGISTERS_reg[5][4]  ( .D(n4322), .CK(CLK), .RN(n422), .Q(n1815), 
        .QN(n4002) );
  DFFR_X1 \REGISTERS_reg[5][3]  ( .D(n4321), .CK(CLK), .RN(n423), .Q(n1814), 
        .QN(n4001) );
  DFFR_X1 \REGISTERS_reg[5][2]  ( .D(n4320), .CK(CLK), .RN(n423), .Q(n1813), 
        .QN(n4000) );
  DFFR_X1 \REGISTERS_reg[5][1]  ( .D(n4319), .CK(CLK), .RN(n423), .Q(n1812), 
        .QN(n3999) );
  DFFR_X1 \REGISTERS_reg[5][0]  ( .D(n4318), .CK(CLK), .RN(n423), .Q(n1811), 
        .QN(n3998) );
  DFFR_X1 \REGISTERS_reg[31][31]  ( .D(n4605), .CK(CLK), .RN(n490), .Q(n1454), 
        .QN(n2717) );
  DFFR_X1 \REGISTERS_reg[31][30]  ( .D(n4604), .CK(CLK), .RN(n490), .Q(n1430), 
        .QN(n2716) );
  DFFR_X1 \REGISTERS_reg[31][29]  ( .D(n4603), .CK(CLK), .RN(n490), .Q(n1414), 
        .QN(n2715) );
  DFFR_X1 \REGISTERS_reg[31][28]  ( .D(n4602), .CK(CLK), .RN(n490), .Q(n1398), 
        .QN(n2714) );
  DFFR_X1 \REGISTERS_reg[31][27]  ( .D(n4601), .CK(CLK), .RN(n490), .Q(n1382), 
        .QN(n2713) );
  DFFR_X1 \REGISTERS_reg[31][26]  ( .D(n4600), .CK(CLK), .RN(n490), .Q(n1366), 
        .QN(n2712) );
  DFFR_X1 \REGISTERS_reg[31][25]  ( .D(n4599), .CK(CLK), .RN(n490), .Q(n1350), 
        .QN(n2711) );
  DFFR_X1 \REGISTERS_reg[31][24]  ( .D(n4598), .CK(CLK), .RN(n490), .Q(n1334), 
        .QN(n2710) );
  DFFR_X1 \REGISTERS_reg[31][23]  ( .D(n4597), .CK(CLK), .RN(n490), .Q(n1318), 
        .QN(n2709) );
  DFFR_X1 \REGISTERS_reg[31][22]  ( .D(n4596), .CK(CLK), .RN(n490), .Q(n1302), 
        .QN(n2708) );
  DFFR_X1 \REGISTERS_reg[31][21]  ( .D(n4595), .CK(CLK), .RN(n490), .Q(n1286), 
        .QN(n2707) );
  DFFR_X1 \REGISTERS_reg[31][20]  ( .D(n4594), .CK(CLK), .RN(n490), .Q(n1270), 
        .QN(n2706) );
  DFFR_X1 \REGISTERS_reg[31][19]  ( .D(n4593), .CK(CLK), .RN(n491), .Q(n1254), 
        .QN(n2705) );
  DFFR_X1 \REGISTERS_reg[31][18]  ( .D(n4592), .CK(CLK), .RN(n491), .Q(n1238), 
        .QN(n2704) );
  DFFR_X1 \REGISTERS_reg[31][17]  ( .D(n4591), .CK(CLK), .RN(n491), .Q(n1222), 
        .QN(n2703) );
  DFFR_X1 \REGISTERS_reg[31][16]  ( .D(n4590), .CK(CLK), .RN(n491), .Q(n1206), 
        .QN(n2702) );
  DFFR_X1 \REGISTERS_reg[31][15]  ( .D(n4589), .CK(CLK), .RN(n491), .Q(n1190), 
        .QN(n2701) );
  DFFR_X1 \REGISTERS_reg[31][14]  ( .D(n4588), .CK(CLK), .RN(n491), .Q(n1174), 
        .QN(n2700) );
  DFFR_X1 \REGISTERS_reg[31][13]  ( .D(n4587), .CK(CLK), .RN(n491), .Q(n1158), 
        .QN(n2699) );
  DFFR_X1 \REGISTERS_reg[31][12]  ( .D(n4586), .CK(CLK), .RN(n491), .Q(n1142), 
        .QN(n2698) );
  DFFR_X1 \REGISTERS_reg[31][11]  ( .D(n4585), .CK(CLK), .RN(n491), .Q(n1126), 
        .QN(n2697) );
  DFFR_X1 \REGISTERS_reg[31][10]  ( .D(n4584), .CK(CLK), .RN(n491), .Q(n1110), 
        .QN(n2696) );
  DFFR_X1 \REGISTERS_reg[31][9]  ( .D(n4583), .CK(CLK), .RN(n491), .Q(n1094), 
        .QN(n2695) );
  DFFR_X1 \REGISTERS_reg[31][8]  ( .D(n4582), .CK(CLK), .RN(n491), .Q(n1078), 
        .QN(n2694) );
  DFFR_X1 \REGISTERS_reg[31][7]  ( .D(n4581), .CK(CLK), .RN(n492), .Q(n1062), 
        .QN(n2693) );
  DFFR_X1 \REGISTERS_reg[31][6]  ( .D(n4580), .CK(CLK), .RN(n492), .Q(n1046), 
        .QN(n2692) );
  DFFR_X1 \REGISTERS_reg[31][5]  ( .D(n4579), .CK(CLK), .RN(n492), .Q(n1030), 
        .QN(n2691) );
  DFFR_X1 \REGISTERS_reg[31][4]  ( .D(n4578), .CK(CLK), .RN(n492), .Q(n1014), 
        .QN(n2690) );
  DFFR_X1 \REGISTERS_reg[31][3]  ( .D(n4577), .CK(CLK), .RN(n492), .Q(n998), 
        .QN(n2689) );
  DFFR_X1 \REGISTERS_reg[31][2]  ( .D(n4576), .CK(CLK), .RN(n492), .Q(n982), 
        .QN(n2688) );
  DFFR_X1 \REGISTERS_reg[31][1]  ( .D(n4575), .CK(CLK), .RN(n492), .Q(n966), 
        .QN(n2687) );
  DFFR_X1 \REGISTERS_reg[31][0]  ( .D(n4574), .CK(CLK), .RN(n492), .Q(n950), 
        .QN(n2686) );
  DFFR_X1 \REGISTERS_reg[21][31]  ( .D(n4477), .CK(CLK), .RN(n463), .Q(n1584), 
        .QN(n2973) );
  DFFR_X1 \REGISTERS_reg[21][30]  ( .D(n4476), .CK(CLK), .RN(n463), .Q(n1583), 
        .QN(n2972) );
  DFFR_X1 \REGISTERS_reg[21][29]  ( .D(n4475), .CK(CLK), .RN(n463), .Q(n1582), 
        .QN(n2971) );
  DFFR_X1 \REGISTERS_reg[21][28]  ( .D(n4474), .CK(CLK), .RN(n463), .Q(n1581), 
        .QN(n2970) );
  DFFR_X1 \REGISTERS_reg[21][27]  ( .D(n4473), .CK(CLK), .RN(n463), .Q(n1580), 
        .QN(n2969) );
  DFFR_X1 \REGISTERS_reg[21][26]  ( .D(n4472), .CK(CLK), .RN(n463), .Q(n1579), 
        .QN(n2968) );
  DFFR_X1 \REGISTERS_reg[21][25]  ( .D(n4471), .CK(CLK), .RN(n463), .Q(n1578), 
        .QN(n2967) );
  DFFR_X1 \REGISTERS_reg[21][24]  ( .D(n4470), .CK(CLK), .RN(n463), .Q(n1577), 
        .QN(n2966) );
  DFFR_X1 \REGISTERS_reg[21][23]  ( .D(n4469), .CK(CLK), .RN(n464), .Q(n1576), 
        .QN(n2965) );
  DFFR_X1 \REGISTERS_reg[21][22]  ( .D(n4468), .CK(CLK), .RN(n464), .Q(n1575), 
        .QN(n2964) );
  DFFR_X1 \REGISTERS_reg[21][21]  ( .D(n4467), .CK(CLK), .RN(n464), .Q(n1574), 
        .QN(n2963) );
  DFFR_X1 \REGISTERS_reg[21][20]  ( .D(n4466), .CK(CLK), .RN(n464), .Q(n1573), 
        .QN(n2962) );
  DFFR_X1 \REGISTERS_reg[21][19]  ( .D(n4465), .CK(CLK), .RN(n464), .Q(n1572), 
        .QN(n2961) );
  DFFR_X1 \REGISTERS_reg[21][18]  ( .D(n4464), .CK(CLK), .RN(n464), .Q(n1571), 
        .QN(n2960) );
  DFFR_X1 \REGISTERS_reg[21][17]  ( .D(n4463), .CK(CLK), .RN(n464), .Q(n1570), 
        .QN(n2959) );
  DFFR_X1 \REGISTERS_reg[21][16]  ( .D(n4462), .CK(CLK), .RN(n464), .Q(n1569), 
        .QN(n2958) );
  DFFR_X1 \REGISTERS_reg[21][15]  ( .D(n4461), .CK(CLK), .RN(n464), .Q(n1568), 
        .QN(n2957) );
  DFFR_X1 \REGISTERS_reg[21][14]  ( .D(n4460), .CK(CLK), .RN(n464), .Q(n1567), 
        .QN(n2956) );
  DFFR_X1 \REGISTERS_reg[21][13]  ( .D(n4459), .CK(CLK), .RN(n464), .Q(n1566), 
        .QN(n2955) );
  DFFR_X1 \REGISTERS_reg[21][12]  ( .D(n4458), .CK(CLK), .RN(n464), .Q(n1565), 
        .QN(n2954) );
  DFFR_X1 \REGISTERS_reg[21][11]  ( .D(n4457), .CK(CLK), .RN(n465), .Q(n1564), 
        .QN(n2953) );
  DFFR_X1 \REGISTERS_reg[21][10]  ( .D(n4456), .CK(CLK), .RN(n465), .Q(n1563), 
        .QN(n2952) );
  DFFR_X1 \REGISTERS_reg[21][9]  ( .D(n4455), .CK(CLK), .RN(n465), .Q(n1562), 
        .QN(n2951) );
  DFFR_X1 \REGISTERS_reg[21][8]  ( .D(n4454), .CK(CLK), .RN(n465), .Q(n1561), 
        .QN(n2950) );
  DFFR_X1 \REGISTERS_reg[21][7]  ( .D(n4453), .CK(CLK), .RN(n465), .Q(n1560), 
        .QN(n2949) );
  DFFR_X1 \REGISTERS_reg[21][6]  ( .D(n4452), .CK(CLK), .RN(n465), .Q(n1559), 
        .QN(n2948) );
  DFFR_X1 \REGISTERS_reg[21][5]  ( .D(n4451), .CK(CLK), .RN(n465), .Q(n1558), 
        .QN(n2947) );
  DFFR_X1 \REGISTERS_reg[21][4]  ( .D(n4450), .CK(CLK), .RN(n465), .Q(n1557), 
        .QN(n2946) );
  DFFR_X1 \REGISTERS_reg[21][3]  ( .D(n4449), .CK(CLK), .RN(n465), .Q(n1556), 
        .QN(n2945) );
  DFFR_X1 \REGISTERS_reg[21][2]  ( .D(n4448), .CK(CLK), .RN(n465), .Q(n1555), 
        .QN(n2944) );
  DFFR_X1 \REGISTERS_reg[21][1]  ( .D(n4447), .CK(CLK), .RN(n465), .Q(n1554), 
        .QN(n2943) );
  DFFR_X1 \REGISTERS_reg[21][0]  ( .D(n4446), .CK(CLK), .RN(n465), .Q(n1553), 
        .QN(n2942) );
  DFFR_X1 \REGISTERS_reg[12][31]  ( .D(n4221), .CK(CLK), .RN(n439), .Q(n1744), 
        .QN(n3805) );
  DFFR_X1 \REGISTERS_reg[12][30]  ( .D(n4220), .CK(CLK), .RN(n439), .Q(n1743), 
        .QN(n3804) );
  DFFR_X1 \REGISTERS_reg[12][29]  ( .D(n4219), .CK(CLK), .RN(n439), .Q(n1742), 
        .QN(n3803) );
  DFFR_X1 \REGISTERS_reg[12][28]  ( .D(n4218), .CK(CLK), .RN(n439), .Q(n1741), 
        .QN(n3802) );
  DFFR_X1 \REGISTERS_reg[12][27]  ( .D(n4217), .CK(CLK), .RN(n439), .Q(n1740), 
        .QN(n3801) );
  DFFR_X1 \REGISTERS_reg[12][26]  ( .D(n4216), .CK(CLK), .RN(n439), .Q(n1739), 
        .QN(n3800) );
  DFFR_X1 \REGISTERS_reg[12][25]  ( .D(n4215), .CK(CLK), .RN(n439), .Q(n1738), 
        .QN(n3799) );
  DFFR_X1 \REGISTERS_reg[12][24]  ( .D(n4214), .CK(CLK), .RN(n439), .Q(n1737), 
        .QN(n3798) );
  DFFR_X1 \REGISTERS_reg[12][23]  ( .D(n4213), .CK(CLK), .RN(n440), .Q(n1736), 
        .QN(n3797) );
  DFFR_X1 \REGISTERS_reg[12][22]  ( .D(n4212), .CK(CLK), .RN(n440), .Q(n1735), 
        .QN(n3796) );
  DFFR_X1 \REGISTERS_reg[12][21]  ( .D(n4211), .CK(CLK), .RN(n440), .Q(n1734), 
        .QN(n3795) );
  DFFR_X1 \REGISTERS_reg[12][20]  ( .D(n4210), .CK(CLK), .RN(n440), .Q(n1733), 
        .QN(n3794) );
  DFFR_X1 \REGISTERS_reg[12][19]  ( .D(n4209), .CK(CLK), .RN(n440), .Q(n1732), 
        .QN(n3793) );
  DFFR_X1 \REGISTERS_reg[12][18]  ( .D(n4208), .CK(CLK), .RN(n440), .Q(n1731), 
        .QN(n3792) );
  DFFR_X1 \REGISTERS_reg[12][17]  ( .D(n4207), .CK(CLK), .RN(n440), .Q(n1730), 
        .QN(n3791) );
  DFFR_X1 \REGISTERS_reg[12][16]  ( .D(n4206), .CK(CLK), .RN(n440), .Q(n1729), 
        .QN(n3790) );
  DFFR_X1 \REGISTERS_reg[12][15]  ( .D(n4205), .CK(CLK), .RN(n440), .Q(n1728), 
        .QN(n3789) );
  DFFR_X1 \REGISTERS_reg[12][14]  ( .D(n4204), .CK(CLK), .RN(n440), .Q(n1727), 
        .QN(n3788) );
  DFFR_X1 \REGISTERS_reg[12][13]  ( .D(n4203), .CK(CLK), .RN(n440), .Q(n1726), 
        .QN(n3787) );
  DFFR_X1 \REGISTERS_reg[12][12]  ( .D(n4202), .CK(CLK), .RN(n440), .Q(n1725), 
        .QN(n3786) );
  DFFR_X1 \REGISTERS_reg[12][11]  ( .D(n4201), .CK(CLK), .RN(n441), .Q(n1724), 
        .QN(n3785) );
  DFFR_X1 \REGISTERS_reg[12][10]  ( .D(n4200), .CK(CLK), .RN(n441), .Q(n1723), 
        .QN(n3784) );
  DFFR_X1 \REGISTERS_reg[12][9]  ( .D(n4199), .CK(CLK), .RN(n441), .Q(n1722), 
        .QN(n3783) );
  DFFR_X1 \REGISTERS_reg[12][8]  ( .D(n4198), .CK(CLK), .RN(n441), .Q(n1721), 
        .QN(n3782) );
  DFFR_X1 \REGISTERS_reg[12][7]  ( .D(n4197), .CK(CLK), .RN(n441), .Q(n1720), 
        .QN(n3781) );
  DFFR_X1 \REGISTERS_reg[12][6]  ( .D(n4196), .CK(CLK), .RN(n441), .Q(n1719), 
        .QN(n3780) );
  DFFR_X1 \REGISTERS_reg[12][5]  ( .D(n4195), .CK(CLK), .RN(n441), .Q(n1718), 
        .QN(n3779) );
  DFFR_X1 \REGISTERS_reg[12][4]  ( .D(n4194), .CK(CLK), .RN(n441), .Q(n1717), 
        .QN(n3778) );
  DFFR_X1 \REGISTERS_reg[12][3]  ( .D(n4193), .CK(CLK), .RN(n441), .Q(n1716), 
        .QN(n3777) );
  DFFR_X1 \REGISTERS_reg[12][2]  ( .D(n4192), .CK(CLK), .RN(n441), .Q(n1715), 
        .QN(n3776) );
  DFFR_X1 \REGISTERS_reg[12][1]  ( .D(n4191), .CK(CLK), .RN(n441), .Q(n1714), 
        .QN(n3775) );
  DFFR_X1 \REGISTERS_reg[12][0]  ( .D(n4190), .CK(CLK), .RN(n441), .Q(n1713), 
        .QN(n3774) );
  DFFR_X1 \REGISTERS_reg[8][31]  ( .D(n4157), .CK(CLK), .RN(n428), .Q(n1808), 
        .QN(n3933) );
  DFFR_X1 \REGISTERS_reg[8][30]  ( .D(n4156), .CK(CLK), .RN(n428), .Q(n1807), 
        .QN(n3932) );
  DFFR_X1 \REGISTERS_reg[8][29]  ( .D(n4155), .CK(CLK), .RN(n428), .Q(n1806), 
        .QN(n3931) );
  DFFR_X1 \REGISTERS_reg[8][28]  ( .D(n4154), .CK(CLK), .RN(n428), .Q(n1805), 
        .QN(n3930) );
  DFFR_X1 \REGISTERS_reg[8][27]  ( .D(n4153), .CK(CLK), .RN(n429), .Q(n1804), 
        .QN(n3929) );
  DFFR_X1 \REGISTERS_reg[8][26]  ( .D(n4152), .CK(CLK), .RN(n429), .Q(n1803), 
        .QN(n3928) );
  DFFR_X1 \REGISTERS_reg[8][25]  ( .D(n4151), .CK(CLK), .RN(n429), .Q(n1802), 
        .QN(n3927) );
  DFFR_X1 \REGISTERS_reg[8][24]  ( .D(n4150), .CK(CLK), .RN(n429), .Q(n1801), 
        .QN(n3926) );
  DFFR_X1 \REGISTERS_reg[8][23]  ( .D(n4149), .CK(CLK), .RN(n429), .Q(n1800), 
        .QN(n3925) );
  DFFR_X1 \REGISTERS_reg[8][22]  ( .D(n4148), .CK(CLK), .RN(n429), .Q(n1799), 
        .QN(n3924) );
  DFFR_X1 \REGISTERS_reg[8][21]  ( .D(n4147), .CK(CLK), .RN(n429), .Q(n1798), 
        .QN(n3923) );
  DFFR_X1 \REGISTERS_reg[8][20]  ( .D(n4146), .CK(CLK), .RN(n429), .Q(n1797), 
        .QN(n3922) );
  DFFR_X1 \REGISTERS_reg[8][19]  ( .D(n4145), .CK(CLK), .RN(n429), .Q(n1796), 
        .QN(n3921) );
  DFFR_X1 \REGISTERS_reg[8][18]  ( .D(n4144), .CK(CLK), .RN(n429), .Q(n1795), 
        .QN(n3920) );
  DFFR_X1 \REGISTERS_reg[8][17]  ( .D(n4143), .CK(CLK), .RN(n429), .Q(n1794), 
        .QN(n3919) );
  DFFR_X1 \REGISTERS_reg[8][16]  ( .D(n4142), .CK(CLK), .RN(n429), .Q(n1793), 
        .QN(n3918) );
  DFFR_X1 \REGISTERS_reg[8][15]  ( .D(n4141), .CK(CLK), .RN(n430), .Q(n1792), 
        .QN(n3917) );
  DFFR_X1 \REGISTERS_reg[8][14]  ( .D(n4140), .CK(CLK), .RN(n430), .Q(n1791), 
        .QN(n3916) );
  DFFR_X1 \REGISTERS_reg[8][13]  ( .D(n4139), .CK(CLK), .RN(n430), .Q(n1790), 
        .QN(n3915) );
  DFFR_X1 \REGISTERS_reg[8][12]  ( .D(n4138), .CK(CLK), .RN(n430), .Q(n1789), 
        .QN(n3914) );
  DFFR_X1 \REGISTERS_reg[8][11]  ( .D(n4137), .CK(CLK), .RN(n430), .Q(n1788), 
        .QN(n3913) );
  DFFR_X1 \REGISTERS_reg[8][10]  ( .D(n4136), .CK(CLK), .RN(n430), .Q(n1787), 
        .QN(n3912) );
  DFFR_X1 \REGISTERS_reg[8][9]  ( .D(n4135), .CK(CLK), .RN(n430), .Q(n1786), 
        .QN(n3911) );
  DFFR_X1 \REGISTERS_reg[8][8]  ( .D(n4134), .CK(CLK), .RN(n430), .Q(n1785), 
        .QN(n3910) );
  DFFR_X1 \REGISTERS_reg[8][7]  ( .D(n4133), .CK(CLK), .RN(n430), .Q(n1784), 
        .QN(n3909) );
  DFFR_X1 \REGISTERS_reg[8][6]  ( .D(n4132), .CK(CLK), .RN(n430), .Q(n1783), 
        .QN(n3908) );
  DFFR_X1 \REGISTERS_reg[8][5]  ( .D(n4131), .CK(CLK), .RN(n430), .Q(n1782), 
        .QN(n3907) );
  DFFR_X1 \REGISTERS_reg[8][4]  ( .D(n4130), .CK(CLK), .RN(n430), .Q(n1781), 
        .QN(n3906) );
  DFFR_X1 \REGISTERS_reg[8][3]  ( .D(n4129), .CK(CLK), .RN(n431), .Q(n1780), 
        .QN(n3905) );
  DFFR_X1 \REGISTERS_reg[8][2]  ( .D(n4128), .CK(CLK), .RN(n431), .Q(n1779), 
        .QN(n3904) );
  DFFR_X1 \REGISTERS_reg[8][1]  ( .D(n4127), .CK(CLK), .RN(n431), .Q(n1778), 
        .QN(n3903) );
  DFFR_X1 \REGISTERS_reg[8][0]  ( .D(n4126), .CK(CLK), .RN(n431), .Q(n1777), 
        .QN(n3902) );
  DFFR_X1 \REGISTERS_reg[30][31]  ( .D(n4573), .CK(CLK), .RN(n487), .Q(n1486), 
        .QN(n2749) );
  DFFR_X1 \REGISTERS_reg[30][30]  ( .D(n4572), .CK(CLK), .RN(n487), .Q(n1485), 
        .QN(n2748) );
  DFFR_X1 \REGISTERS_reg[30][29]  ( .D(n4571), .CK(CLK), .RN(n487), .Q(n1484), 
        .QN(n2747) );
  DFFR_X1 \REGISTERS_reg[30][28]  ( .D(n4570), .CK(CLK), .RN(n487), .Q(n1483), 
        .QN(n2746) );
  DFFR_X1 \REGISTERS_reg[30][27]  ( .D(n4569), .CK(CLK), .RN(n487), .Q(n1482), 
        .QN(n2745) );
  DFFR_X1 \REGISTERS_reg[30][26]  ( .D(n4568), .CK(CLK), .RN(n487), .Q(n1481), 
        .QN(n2744) );
  DFFR_X1 \REGISTERS_reg[30][25]  ( .D(n4567), .CK(CLK), .RN(n487), .Q(n1480), 
        .QN(n2743) );
  DFFR_X1 \REGISTERS_reg[30][24]  ( .D(n4566), .CK(CLK), .RN(n487), .Q(n1479), 
        .QN(n2742) );
  DFFR_X1 \REGISTERS_reg[30][23]  ( .D(n4565), .CK(CLK), .RN(n488), .Q(n1478), 
        .QN(n2741) );
  DFFR_X1 \REGISTERS_reg[30][22]  ( .D(n4564), .CK(CLK), .RN(n488), .Q(n1477), 
        .QN(n2740) );
  DFFR_X1 \REGISTERS_reg[30][21]  ( .D(n4563), .CK(CLK), .RN(n488), .Q(n1476), 
        .QN(n2739) );
  DFFR_X1 \REGISTERS_reg[30][20]  ( .D(n4562), .CK(CLK), .RN(n488), .Q(n1475), 
        .QN(n2738) );
  DFFR_X1 \REGISTERS_reg[30][19]  ( .D(n4561), .CK(CLK), .RN(n488), .Q(n1474), 
        .QN(n2737) );
  DFFR_X1 \REGISTERS_reg[30][18]  ( .D(n4560), .CK(CLK), .RN(n488), .Q(n1473), 
        .QN(n2736) );
  DFFR_X1 \REGISTERS_reg[30][17]  ( .D(n4559), .CK(CLK), .RN(n488), .Q(n1472), 
        .QN(n2735) );
  DFFR_X1 \REGISTERS_reg[30][16]  ( .D(n4558), .CK(CLK), .RN(n488), .Q(n1471), 
        .QN(n2734) );
  DFFR_X1 \REGISTERS_reg[30][15]  ( .D(n4557), .CK(CLK), .RN(n488), .Q(n1470), 
        .QN(n2733) );
  DFFR_X1 \REGISTERS_reg[30][14]  ( .D(n4556), .CK(CLK), .RN(n488), .Q(n1469), 
        .QN(n2732) );
  DFFR_X1 \REGISTERS_reg[30][13]  ( .D(n4555), .CK(CLK), .RN(n488), .Q(n1468), 
        .QN(n2731) );
  DFFR_X1 \REGISTERS_reg[30][12]  ( .D(n4554), .CK(CLK), .RN(n488), .Q(n1467), 
        .QN(n2730) );
  DFFR_X1 \REGISTERS_reg[30][11]  ( .D(n4553), .CK(CLK), .RN(n489), .Q(n1466), 
        .QN(n2729) );
  DFFR_X1 \REGISTERS_reg[30][10]  ( .D(n4552), .CK(CLK), .RN(n489), .Q(n1465), 
        .QN(n2728) );
  DFFR_X1 \REGISTERS_reg[30][9]  ( .D(n4551), .CK(CLK), .RN(n489), .Q(n1464), 
        .QN(n2727) );
  DFFR_X1 \REGISTERS_reg[30][8]  ( .D(n4550), .CK(CLK), .RN(n489), .Q(n1463), 
        .QN(n2726) );
  DFFR_X1 \REGISTERS_reg[30][7]  ( .D(n4549), .CK(CLK), .RN(n489), .Q(n1462), 
        .QN(n2725) );
  DFFR_X1 \REGISTERS_reg[30][6]  ( .D(n4548), .CK(CLK), .RN(n489), .Q(n1461), 
        .QN(n2724) );
  DFFR_X1 \REGISTERS_reg[30][5]  ( .D(n4547), .CK(CLK), .RN(n489), .Q(n1460), 
        .QN(n2723) );
  DFFR_X1 \REGISTERS_reg[30][4]  ( .D(n4546), .CK(CLK), .RN(n489), .Q(n1459), 
        .QN(n2722) );
  DFFR_X1 \REGISTERS_reg[30][3]  ( .D(n4545), .CK(CLK), .RN(n489), .Q(n1458), 
        .QN(n2721) );
  DFFR_X1 \REGISTERS_reg[30][2]  ( .D(n4544), .CK(CLK), .RN(n489), .Q(n1457), 
        .QN(n2720) );
  DFFR_X1 \REGISTERS_reg[30][1]  ( .D(n4543), .CK(CLK), .RN(n489), .Q(n1456), 
        .QN(n2719) );
  DFFR_X1 \REGISTERS_reg[30][0]  ( .D(n4542), .CK(CLK), .RN(n489), .Q(n1455), 
        .QN(n2718) );
  DFFR_X1 \REGISTERS_reg[20][31]  ( .D(n4445), .CK(CLK), .RN(n460), .Q(n1616), 
        .QN(n3581) );
  DFFR_X1 \REGISTERS_reg[20][30]  ( .D(n4444), .CK(CLK), .RN(n460), .Q(n1615), 
        .QN(n3580) );
  DFFR_X1 \REGISTERS_reg[20][29]  ( .D(n4443), .CK(CLK), .RN(n460), .Q(n1614), 
        .QN(n3579) );
  DFFR_X1 \REGISTERS_reg[20][28]  ( .D(n4442), .CK(CLK), .RN(n460), .Q(n1613), 
        .QN(n3578) );
  DFFR_X1 \REGISTERS_reg[20][27]  ( .D(n4441), .CK(CLK), .RN(n461), .Q(n1612), 
        .QN(n3577) );
  DFFR_X1 \REGISTERS_reg[20][26]  ( .D(n4440), .CK(CLK), .RN(n461), .Q(n1611), 
        .QN(n3576) );
  DFFR_X1 \REGISTERS_reg[20][25]  ( .D(n4439), .CK(CLK), .RN(n461), .Q(n1610), 
        .QN(n3575) );
  DFFR_X1 \REGISTERS_reg[20][24]  ( .D(n4438), .CK(CLK), .RN(n461), .Q(n1609), 
        .QN(n3574) );
  DFFR_X1 \REGISTERS_reg[20][23]  ( .D(n4437), .CK(CLK), .RN(n461), .Q(n1608), 
        .QN(n3573) );
  DFFR_X1 \REGISTERS_reg[20][22]  ( .D(n4436), .CK(CLK), .RN(n461), .Q(n1607), 
        .QN(n3572) );
  DFFR_X1 \REGISTERS_reg[20][21]  ( .D(n4435), .CK(CLK), .RN(n461), .Q(n1606), 
        .QN(n3571) );
  DFFR_X1 \REGISTERS_reg[20][20]  ( .D(n4434), .CK(CLK), .RN(n461), .Q(n1605), 
        .QN(n3570) );
  DFFR_X1 \REGISTERS_reg[20][19]  ( .D(n4433), .CK(CLK), .RN(n461), .Q(n1604), 
        .QN(n3569) );
  DFFR_X1 \REGISTERS_reg[20][18]  ( .D(n4432), .CK(CLK), .RN(n461), .Q(n1603), 
        .QN(n3568) );
  DFFR_X1 \REGISTERS_reg[20][17]  ( .D(n4431), .CK(CLK), .RN(n461), .Q(n1602), 
        .QN(n3567) );
  DFFR_X1 \REGISTERS_reg[20][16]  ( .D(n4430), .CK(CLK), .RN(n461), .Q(n1601), 
        .QN(n3566) );
  DFFR_X1 \REGISTERS_reg[20][15]  ( .D(n4429), .CK(CLK), .RN(n462), .Q(n1600), 
        .QN(n3565) );
  DFFR_X1 \REGISTERS_reg[20][14]  ( .D(n4428), .CK(CLK), .RN(n462), .Q(n1599), 
        .QN(n3564) );
  DFFR_X1 \REGISTERS_reg[20][13]  ( .D(n4427), .CK(CLK), .RN(n462), .Q(n1598), 
        .QN(n3563) );
  DFFR_X1 \REGISTERS_reg[20][12]  ( .D(n4426), .CK(CLK), .RN(n462), .Q(n1597), 
        .QN(n3562) );
  DFFR_X1 \REGISTERS_reg[20][11]  ( .D(n4425), .CK(CLK), .RN(n462), .Q(n1596), 
        .QN(n3561) );
  DFFR_X1 \REGISTERS_reg[20][10]  ( .D(n4424), .CK(CLK), .RN(n462), .Q(n1595), 
        .QN(n3560) );
  DFFR_X1 \REGISTERS_reg[20][9]  ( .D(n4423), .CK(CLK), .RN(n462), .Q(n1594), 
        .QN(n3559) );
  DFFR_X1 \REGISTERS_reg[20][8]  ( .D(n4422), .CK(CLK), .RN(n462), .Q(n1593), 
        .QN(n2982) );
  DFFR_X1 \REGISTERS_reg[20][7]  ( .D(n4421), .CK(CLK), .RN(n462), .Q(n1592), 
        .QN(n2981) );
  DFFR_X1 \REGISTERS_reg[20][6]  ( .D(n4420), .CK(CLK), .RN(n462), .Q(n1591), 
        .QN(n2980) );
  DFFR_X1 \REGISTERS_reg[20][5]  ( .D(n4419), .CK(CLK), .RN(n462), .Q(n1590), 
        .QN(n2979) );
  DFFR_X1 \REGISTERS_reg[20][4]  ( .D(n4418), .CK(CLK), .RN(n462), .Q(n1589), 
        .QN(n2978) );
  DFFR_X1 \REGISTERS_reg[20][3]  ( .D(n4417), .CK(CLK), .RN(n463), .Q(n1588), 
        .QN(n2977) );
  DFFR_X1 \REGISTERS_reg[20][2]  ( .D(n4416), .CK(CLK), .RN(n463), .Q(n1587), 
        .QN(n2976) );
  DFFR_X1 \REGISTERS_reg[20][1]  ( .D(n4415), .CK(CLK), .RN(n463), .Q(n1586), 
        .QN(n2975) );
  DFFR_X1 \REGISTERS_reg[20][0]  ( .D(n4414), .CK(CLK), .RN(n463), .Q(n1585), 
        .QN(n2974) );
  DFFR_X1 \REGISTERS_reg[16][31]  ( .D(n4381), .CK(CLK), .RN(n450), .Q(n1680), 
        .QN(n3677) );
  DFFR_X1 \REGISTERS_reg[16][30]  ( .D(n4380), .CK(CLK), .RN(n450), .Q(n1679), 
        .QN(n3676) );
  DFFR_X1 \REGISTERS_reg[16][29]  ( .D(n4379), .CK(CLK), .RN(n450), .Q(n1678), 
        .QN(n3675) );
  DFFR_X1 \REGISTERS_reg[16][28]  ( .D(n4378), .CK(CLK), .RN(n450), .Q(n1677), 
        .QN(n3674) );
  DFFR_X1 \REGISTERS_reg[16][27]  ( .D(n4377), .CK(CLK), .RN(n450), .Q(n1676), 
        .QN(n3673) );
  DFFR_X1 \REGISTERS_reg[16][26]  ( .D(n4376), .CK(CLK), .RN(n450), .Q(n1675), 
        .QN(n3672) );
  DFFR_X1 \REGISTERS_reg[16][25]  ( .D(n4375), .CK(CLK), .RN(n450), .Q(n1674), 
        .QN(n3671) );
  DFFR_X1 \REGISTERS_reg[16][24]  ( .D(n4374), .CK(CLK), .RN(n450), .Q(n1673), 
        .QN(n3670) );
  DFFR_X1 \REGISTERS_reg[16][23]  ( .D(n4373), .CK(CLK), .RN(n450), .Q(n1672), 
        .QN(n3669) );
  DFFR_X1 \REGISTERS_reg[16][22]  ( .D(n4372), .CK(CLK), .RN(n450), .Q(n1671), 
        .QN(n3668) );
  DFFR_X1 \REGISTERS_reg[16][21]  ( .D(n4371), .CK(CLK), .RN(n450), .Q(n1670), 
        .QN(n3667) );
  DFFR_X1 \REGISTERS_reg[16][20]  ( .D(n4370), .CK(CLK), .RN(n450), .Q(n1669), 
        .QN(n3666) );
  DFFR_X1 \REGISTERS_reg[16][19]  ( .D(n4369), .CK(CLK), .RN(n451), .Q(n1668), 
        .QN(n3665) );
  DFFR_X1 \REGISTERS_reg[16][18]  ( .D(n4368), .CK(CLK), .RN(n451), .Q(n1667), 
        .QN(n3664) );
  DFFR_X1 \REGISTERS_reg[16][17]  ( .D(n4367), .CK(CLK), .RN(n451), .Q(n1666), 
        .QN(n3663) );
  DFFR_X1 \REGISTERS_reg[16][16]  ( .D(n4366), .CK(CLK), .RN(n451), .Q(n1665), 
        .QN(n3662) );
  DFFR_X1 \REGISTERS_reg[16][15]  ( .D(n4365), .CK(CLK), .RN(n451), .Q(n1664), 
        .QN(n3661) );
  DFFR_X1 \REGISTERS_reg[16][14]  ( .D(n4364), .CK(CLK), .RN(n451), .Q(n1663), 
        .QN(n3660) );
  DFFR_X1 \REGISTERS_reg[16][13]  ( .D(n4363), .CK(CLK), .RN(n451), .Q(n1662), 
        .QN(n3659) );
  DFFR_X1 \REGISTERS_reg[16][12]  ( .D(n4362), .CK(CLK), .RN(n451), .Q(n1661), 
        .QN(n3658) );
  DFFR_X1 \REGISTERS_reg[16][11]  ( .D(n4361), .CK(CLK), .RN(n451), .Q(n1660), 
        .QN(n3657) );
  DFFR_X1 \REGISTERS_reg[16][10]  ( .D(n4360), .CK(CLK), .RN(n451), .Q(n1659), 
        .QN(n3656) );
  DFFR_X1 \REGISTERS_reg[16][9]  ( .D(n4359), .CK(CLK), .RN(n451), .Q(n1658), 
        .QN(n3655) );
  DFFR_X1 \REGISTERS_reg[16][8]  ( .D(n4358), .CK(CLK), .RN(n451), .Q(n1657), 
        .QN(n3654) );
  DFFR_X1 \REGISTERS_reg[16][7]  ( .D(n4357), .CK(CLK), .RN(n452), .Q(n1656), 
        .QN(n3653) );
  DFFR_X1 \REGISTERS_reg[16][6]  ( .D(n4356), .CK(CLK), .RN(n452), .Q(n1655), 
        .QN(n3652) );
  DFFR_X1 \REGISTERS_reg[16][5]  ( .D(n4355), .CK(CLK), .RN(n452), .Q(n1654), 
        .QN(n3651) );
  DFFR_X1 \REGISTERS_reg[16][4]  ( .D(n4354), .CK(CLK), .RN(n452), .Q(n1653), 
        .QN(n3650) );
  DFFR_X1 \REGISTERS_reg[16][3]  ( .D(n4353), .CK(CLK), .RN(n452), .Q(n1652), 
        .QN(n3649) );
  DFFR_X1 \REGISTERS_reg[16][2]  ( .D(n4352), .CK(CLK), .RN(n452), .Q(n1651), 
        .QN(n3648) );
  DFFR_X1 \REGISTERS_reg[16][1]  ( .D(n4351), .CK(CLK), .RN(n452), .Q(n1650), 
        .QN(n3647) );
  DFFR_X1 \REGISTERS_reg[16][0]  ( .D(n4350), .CK(CLK), .RN(n452), .Q(n1649), 
        .QN(n3646) );
  DFFR_X1 \REGISTERS_reg[13][31]  ( .D(n4253), .CK(CLK), .RN(n442), .Q(n1712), 
        .QN(n3773) );
  DFFR_X1 \REGISTERS_reg[13][30]  ( .D(n4252), .CK(CLK), .RN(n442), .Q(n1711), 
        .QN(n3772) );
  DFFR_X1 \REGISTERS_reg[13][29]  ( .D(n4251), .CK(CLK), .RN(n442), .Q(n1710), 
        .QN(n3771) );
  DFFR_X1 \REGISTERS_reg[13][28]  ( .D(n4250), .CK(CLK), .RN(n442), .Q(n1709), 
        .QN(n3770) );
  DFFR_X1 \REGISTERS_reg[13][27]  ( .D(n4249), .CK(CLK), .RN(n442), .Q(n1708), 
        .QN(n3769) );
  DFFR_X1 \REGISTERS_reg[13][26]  ( .D(n4248), .CK(CLK), .RN(n442), .Q(n1707), 
        .QN(n3768) );
  DFFR_X1 \REGISTERS_reg[13][25]  ( .D(n4247), .CK(CLK), .RN(n442), .Q(n1706), 
        .QN(n3767) );
  DFFR_X1 \REGISTERS_reg[13][24]  ( .D(n4246), .CK(CLK), .RN(n442), .Q(n1705), 
        .QN(n3766) );
  DFFR_X1 \REGISTERS_reg[13][23]  ( .D(n4245), .CK(CLK), .RN(n442), .Q(n1704), 
        .QN(n3765) );
  DFFR_X1 \REGISTERS_reg[13][22]  ( .D(n4244), .CK(CLK), .RN(n442), .Q(n1703), 
        .QN(n3764) );
  DFFR_X1 \REGISTERS_reg[13][21]  ( .D(n4243), .CK(CLK), .RN(n442), .Q(n1702), 
        .QN(n3763) );
  DFFR_X1 \REGISTERS_reg[13][20]  ( .D(n4242), .CK(CLK), .RN(n442), .Q(n1701), 
        .QN(n3762) );
  DFFR_X1 \REGISTERS_reg[13][19]  ( .D(n4241), .CK(CLK), .RN(n443), .Q(n1700), 
        .QN(n3761) );
  DFFR_X1 \REGISTERS_reg[13][18]  ( .D(n4240), .CK(CLK), .RN(n443), .Q(n1699), 
        .QN(n3760) );
  DFFR_X1 \REGISTERS_reg[13][17]  ( .D(n4239), .CK(CLK), .RN(n443), .Q(n1698), 
        .QN(n3759) );
  DFFR_X1 \REGISTERS_reg[13][16]  ( .D(n4238), .CK(CLK), .RN(n443), .Q(n1697), 
        .QN(n3758) );
  DFFR_X1 \REGISTERS_reg[13][15]  ( .D(n4237), .CK(CLK), .RN(n443), .Q(n1696), 
        .QN(n3757) );
  DFFR_X1 \REGISTERS_reg[13][14]  ( .D(n4236), .CK(CLK), .RN(n443), .Q(n1695), 
        .QN(n3756) );
  DFFR_X1 \REGISTERS_reg[13][13]  ( .D(n4235), .CK(CLK), .RN(n443), .Q(n1694), 
        .QN(n3755) );
  DFFR_X1 \REGISTERS_reg[13][12]  ( .D(n4234), .CK(CLK), .RN(n443), .Q(n1693), 
        .QN(n3754) );
  DFFR_X1 \REGISTERS_reg[13][11]  ( .D(n4233), .CK(CLK), .RN(n443), .Q(n1692), 
        .QN(n3753) );
  DFFR_X1 \REGISTERS_reg[13][10]  ( .D(n4232), .CK(CLK), .RN(n443), .Q(n1691), 
        .QN(n3752) );
  DFFR_X1 \REGISTERS_reg[13][9]  ( .D(n4231), .CK(CLK), .RN(n443), .Q(n1690), 
        .QN(n3751) );
  DFFR_X1 \REGISTERS_reg[13][8]  ( .D(n4230), .CK(CLK), .RN(n443), .Q(n1689), 
        .QN(n3750) );
  DFFR_X1 \REGISTERS_reg[13][7]  ( .D(n4229), .CK(CLK), .RN(n444), .Q(n1688), 
        .QN(n3749) );
  DFFR_X1 \REGISTERS_reg[13][6]  ( .D(n4228), .CK(CLK), .RN(n444), .Q(n1687), 
        .QN(n3748) );
  DFFR_X1 \REGISTERS_reg[13][5]  ( .D(n4227), .CK(CLK), .RN(n444), .Q(n1686), 
        .QN(n3747) );
  DFFR_X1 \REGISTERS_reg[13][4]  ( .D(n4226), .CK(CLK), .RN(n444), .Q(n1685), 
        .QN(n3746) );
  DFFR_X1 \REGISTERS_reg[13][3]  ( .D(n4225), .CK(CLK), .RN(n444), .Q(n1684), 
        .QN(n3745) );
  DFFR_X1 \REGISTERS_reg[13][2]  ( .D(n4224), .CK(CLK), .RN(n444), .Q(n1683), 
        .QN(n3744) );
  DFFR_X1 \REGISTERS_reg[13][1]  ( .D(n4223), .CK(CLK), .RN(n444), .Q(n1682), 
        .QN(n3743) );
  DFFR_X1 \REGISTERS_reg[13][0]  ( .D(n4222), .CK(CLK), .RN(n444), .Q(n1681), 
        .QN(n3742) );
  DFFR_X1 \REGISTERS_reg[9][31]  ( .D(n4189), .CK(CLK), .RN(n431), .Q(n1776), 
        .QN(n3901) );
  DFFR_X1 \REGISTERS_reg[9][30]  ( .D(n4188), .CK(CLK), .RN(n431), .Q(n1775), 
        .QN(n3900) );
  DFFR_X1 \REGISTERS_reg[9][29]  ( .D(n4187), .CK(CLK), .RN(n431), .Q(n1774), 
        .QN(n3899) );
  DFFR_X1 \REGISTERS_reg[9][28]  ( .D(n4186), .CK(CLK), .RN(n431), .Q(n1773), 
        .QN(n3898) );
  DFFR_X1 \REGISTERS_reg[9][27]  ( .D(n4185), .CK(CLK), .RN(n431), .Q(n1772), 
        .QN(n3897) );
  DFFR_X1 \REGISTERS_reg[9][26]  ( .D(n4184), .CK(CLK), .RN(n431), .Q(n1771), 
        .QN(n3896) );
  DFFR_X1 \REGISTERS_reg[9][25]  ( .D(n4183), .CK(CLK), .RN(n431), .Q(n1770), 
        .QN(n3895) );
  DFFR_X1 \REGISTERS_reg[9][24]  ( .D(n4182), .CK(CLK), .RN(n431), .Q(n1769), 
        .QN(n3894) );
  DFFR_X1 \REGISTERS_reg[9][23]  ( .D(n4181), .CK(CLK), .RN(n432), .Q(n1768), 
        .QN(n3893) );
  DFFR_X1 \REGISTERS_reg[9][22]  ( .D(n4180), .CK(CLK), .RN(n432), .Q(n1767), 
        .QN(n3892) );
  DFFR_X1 \REGISTERS_reg[9][21]  ( .D(n4179), .CK(CLK), .RN(n432), .Q(n1766), 
        .QN(n3891) );
  DFFR_X1 \REGISTERS_reg[9][20]  ( .D(n4178), .CK(CLK), .RN(n432), .Q(n1765), 
        .QN(n3890) );
  DFFR_X1 \REGISTERS_reg[9][19]  ( .D(n4177), .CK(CLK), .RN(n432), .Q(n1764), 
        .QN(n3889) );
  DFFR_X1 \REGISTERS_reg[9][18]  ( .D(n4176), .CK(CLK), .RN(n432), .Q(n1763), 
        .QN(n3888) );
  DFFR_X1 \REGISTERS_reg[9][17]  ( .D(n4175), .CK(CLK), .RN(n432), .Q(n1762), 
        .QN(n3887) );
  DFFR_X1 \REGISTERS_reg[9][16]  ( .D(n4174), .CK(CLK), .RN(n432), .Q(n1761), 
        .QN(n3886) );
  DFFR_X1 \REGISTERS_reg[9][15]  ( .D(n4173), .CK(CLK), .RN(n432), .Q(n1760), 
        .QN(n3885) );
  DFFR_X1 \REGISTERS_reg[9][14]  ( .D(n4172), .CK(CLK), .RN(n432), .Q(n1759), 
        .QN(n3884) );
  DFFR_X1 \REGISTERS_reg[9][13]  ( .D(n4171), .CK(CLK), .RN(n432), .Q(n1758), 
        .QN(n3883) );
  DFFR_X1 \REGISTERS_reg[9][12]  ( .D(n4170), .CK(CLK), .RN(n432), .Q(n1757), 
        .QN(n3882) );
  DFFR_X1 \REGISTERS_reg[9][11]  ( .D(n4169), .CK(CLK), .RN(n433), .Q(n1756), 
        .QN(n3881) );
  DFFR_X1 \REGISTERS_reg[9][10]  ( .D(n4168), .CK(CLK), .RN(n433), .Q(n1755), 
        .QN(n3880) );
  DFFR_X1 \REGISTERS_reg[9][9]  ( .D(n4167), .CK(CLK), .RN(n433), .Q(n1754), 
        .QN(n3879) );
  DFFR_X1 \REGISTERS_reg[9][8]  ( .D(n4166), .CK(CLK), .RN(n433), .Q(n1753), 
        .QN(n3878) );
  DFFR_X1 \REGISTERS_reg[9][7]  ( .D(n4165), .CK(CLK), .RN(n433), .Q(n1752), 
        .QN(n3877) );
  DFFR_X1 \REGISTERS_reg[9][6]  ( .D(n4164), .CK(CLK), .RN(n433), .Q(n1751), 
        .QN(n3876) );
  DFFR_X1 \REGISTERS_reg[9][5]  ( .D(n4163), .CK(CLK), .RN(n433), .Q(n1750), 
        .QN(n3875) );
  DFFR_X1 \REGISTERS_reg[9][4]  ( .D(n4162), .CK(CLK), .RN(n433), .Q(n1749), 
        .QN(n3874) );
  DFFR_X1 \REGISTERS_reg[9][3]  ( .D(n4161), .CK(CLK), .RN(n433), .Q(n1748), 
        .QN(n3873) );
  DFFR_X1 \REGISTERS_reg[9][2]  ( .D(n4160), .CK(CLK), .RN(n433), .Q(n1747), 
        .QN(n3872) );
  DFFR_X1 \REGISTERS_reg[9][1]  ( .D(n4159), .CK(CLK), .RN(n433), .Q(n1746), 
        .QN(n3871) );
  DFFR_X1 \REGISTERS_reg[9][0]  ( .D(n4158), .CK(CLK), .RN(n433), .Q(n1745), 
        .QN(n3870) );
  DFFR_X1 \REGISTERS_reg[1][31]  ( .D(n4285), .CK(CLK), .RN(n410), .Q(n1906), 
        .QN(n4094) );
  DFFR_X1 \REGISTERS_reg[1][30]  ( .D(n4284), .CK(CLK), .RN(n410), .Q(n1905), 
        .QN(n4095) );
  DFFR_X1 \REGISTERS_reg[1][29]  ( .D(n4283), .CK(CLK), .RN(n410), .Q(n1904), 
        .QN(n4096) );
  DFFR_X1 \REGISTERS_reg[1][28]  ( .D(n4282), .CK(CLK), .RN(n410), .Q(n1903), 
        .QN(n4097) );
  DFFR_X1 \REGISTERS_reg[1][27]  ( .D(n4281), .CK(CLK), .RN(n410), .Q(n1902), 
        .QN(n4098) );
  DFFR_X1 \REGISTERS_reg[1][26]  ( .D(n4280), .CK(CLK), .RN(n410), .Q(n1901), 
        .QN(n4099) );
  DFFR_X1 \REGISTERS_reg[1][25]  ( .D(n4279), .CK(CLK), .RN(n410), .Q(n1900), 
        .QN(n4100) );
  DFFR_X1 \REGISTERS_reg[1][24]  ( .D(n4278), .CK(CLK), .RN(n410), .Q(n1899), 
        .QN(n4101) );
  DFFR_X1 \REGISTERS_reg[1][23]  ( .D(n4277), .CK(CLK), .RN(n410), .Q(n1898), 
        .QN(n4102) );
  DFFR_X1 \REGISTERS_reg[1][22]  ( .D(n4276), .CK(CLK), .RN(n410), .Q(n1897), 
        .QN(n4103) );
  DFFR_X1 \REGISTERS_reg[1][21]  ( .D(n4275), .CK(CLK), .RN(n410), .Q(n1896), 
        .QN(n4104) );
  DFFR_X1 \REGISTERS_reg[1][20]  ( .D(n4274), .CK(CLK), .RN(n410), .Q(n1895), 
        .QN(n4105) );
  DFFR_X1 \REGISTERS_reg[1][19]  ( .D(n4273), .CK(CLK), .RN(n411), .Q(n1894), 
        .QN(n4106) );
  DFFR_X1 \REGISTERS_reg[1][18]  ( .D(n4272), .CK(CLK), .RN(n411), .Q(n1893), 
        .QN(n4107) );
  DFFR_X1 \REGISTERS_reg[1][17]  ( .D(n4271), .CK(CLK), .RN(n411), .Q(n1892), 
        .QN(n4108) );
  DFFR_X1 \REGISTERS_reg[1][16]  ( .D(n4270), .CK(CLK), .RN(n411), .Q(n1891), 
        .QN(n4109) );
  DFFR_X1 \REGISTERS_reg[1][15]  ( .D(n4269), .CK(CLK), .RN(n411), .Q(n1890), 
        .QN(n4110) );
  DFFR_X1 \REGISTERS_reg[1][14]  ( .D(n4268), .CK(CLK), .RN(n411), .Q(n1889), 
        .QN(n4111) );
  DFFR_X1 \REGISTERS_reg[1][13]  ( .D(n4267), .CK(CLK), .RN(n411), .Q(n1888), 
        .QN(n4112) );
  DFFR_X1 \REGISTERS_reg[1][12]  ( .D(n4266), .CK(CLK), .RN(n411), .Q(n1887), 
        .QN(n4113) );
  DFFR_X1 \REGISTERS_reg[1][11]  ( .D(n4265), .CK(CLK), .RN(n411), .Q(n1886), 
        .QN(n4114) );
  DFFR_X1 \REGISTERS_reg[1][10]  ( .D(n4264), .CK(CLK), .RN(n411), .Q(n1885), 
        .QN(n4115) );
  DFFR_X1 \REGISTERS_reg[1][9]  ( .D(n4263), .CK(CLK), .RN(n411), .Q(n1884), 
        .QN(n4116) );
  DFFR_X1 \REGISTERS_reg[1][8]  ( .D(n4262), .CK(CLK), .RN(n411), .Q(n1883), 
        .QN(n4117) );
  DFFR_X1 \REGISTERS_reg[1][7]  ( .D(n4261), .CK(CLK), .RN(n412), .Q(n1882), 
        .QN(n4118) );
  DFFR_X1 \REGISTERS_reg[1][6]  ( .D(n4260), .CK(CLK), .RN(n412), .Q(n1881), 
        .QN(n4119) );
  DFFR_X1 \REGISTERS_reg[1][5]  ( .D(n4259), .CK(CLK), .RN(n412), .Q(n1880), 
        .QN(n4120) );
  DFFR_X1 \REGISTERS_reg[1][4]  ( .D(n4258), .CK(CLK), .RN(n412), .Q(n1879), 
        .QN(n4121) );
  DFFR_X1 \REGISTERS_reg[1][3]  ( .D(n4257), .CK(CLK), .RN(n412), .Q(n1878), 
        .QN(n4122) );
  DFFR_X1 \REGISTERS_reg[1][2]  ( .D(n4256), .CK(CLK), .RN(n412), .Q(n1877), 
        .QN(n4123) );
  DFFR_X1 \REGISTERS_reg[1][1]  ( .D(n4255), .CK(CLK), .RN(n412), .Q(n1876), 
        .QN(n4124) );
  DFFR_X1 \REGISTERS_reg[1][0]  ( .D(n4254), .CK(CLK), .RN(n412), .Q(n1875), 
        .QN(n4125) );
  AND3_X1 U2 ( .A1(ADD_WR[4]), .A2(ADD_WR[3]), .A3(n1908), .ZN(n1) );
  AND3_X1 U3 ( .A1(ADD_WR[4]), .A2(n1908), .A3(n1810), .ZN(n2) );
  AND3_X1 U4 ( .A1(ADD_WR[3]), .A2(n1908), .A3(n1809), .ZN(n3) );
  AND3_X1 U5 ( .A1(n1908), .A2(n1810), .A3(n1809), .ZN(n4) );
  AND2_X1 U6 ( .A1(n45), .A2(ADD_WR[0]), .ZN(n5) );
  AND2_X1 U7 ( .A1(n45), .A2(n1907), .ZN(n6) );
  AND3_X1 U8 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(n1551), .ZN(n7) );
  AND3_X1 U9 ( .A1(ADD_WR[1]), .A2(n1907), .A3(n1551), .ZN(n8) );
  AND3_X1 U10 ( .A1(ADD_WR[2]), .A2(ADD_WR[0]), .A3(n1552), .ZN(n9) );
  AND3_X1 U11 ( .A1(ADD_WR[2]), .A2(n1907), .A3(n1552), .ZN(n10) );
  AND3_X1 U12 ( .A1(ADD_WR[0]), .A2(n1552), .A3(n1551), .ZN(n11) );
  AND3_X1 U13 ( .A1(n1907), .A2(n1552), .A3(n1551), .ZN(n12) );
  AND2_X1 U14 ( .A1(n1), .A2(n5), .ZN(n13) );
  AND2_X1 U15 ( .A1(n1), .A2(n6), .ZN(n14) );
  AND2_X1 U16 ( .A1(n1), .A2(n9), .ZN(n15) );
  AND2_X1 U17 ( .A1(n1), .A2(n10), .ZN(n16) );
  AND2_X1 U18 ( .A1(n1), .A2(n7), .ZN(n17) );
  AND2_X1 U19 ( .A1(n1), .A2(n8), .ZN(n18) );
  AND2_X1 U20 ( .A1(n1), .A2(n11), .ZN(n19) );
  AND2_X1 U21 ( .A1(n1), .A2(n12), .ZN(n20) );
  AND2_X1 U22 ( .A1(n2), .A2(n5), .ZN(n21) );
  AND2_X1 U23 ( .A1(n2), .A2(n6), .ZN(n22) );
  AND2_X1 U24 ( .A1(n2), .A2(n9), .ZN(n23) );
  AND2_X1 U25 ( .A1(n2), .A2(n10), .ZN(n24) );
  AND2_X1 U26 ( .A1(n2), .A2(n7), .ZN(n25) );
  AND2_X1 U27 ( .A1(n2), .A2(n8), .ZN(n26) );
  AND2_X1 U28 ( .A1(n2), .A2(n11), .ZN(n27) );
  AND2_X1 U29 ( .A1(n2), .A2(n12), .ZN(n28) );
  AND2_X1 U30 ( .A1(n3), .A2(n5), .ZN(n29) );
  AND2_X1 U31 ( .A1(n3), .A2(n6), .ZN(n30) );
  AND2_X1 U32 ( .A1(n3), .A2(n9), .ZN(n31) );
  AND2_X1 U33 ( .A1(n3), .A2(n10), .ZN(n32) );
  AND2_X1 U34 ( .A1(n3), .A2(n7), .ZN(n33) );
  AND2_X1 U35 ( .A1(n3), .A2(n8), .ZN(n34) );
  AND2_X1 U36 ( .A1(n3), .A2(n11), .ZN(n35) );
  AND2_X1 U37 ( .A1(n3), .A2(n12), .ZN(n36) );
  AND2_X1 U38 ( .A1(n2349), .A2(n85), .ZN(n37) );
  AND2_X1 U39 ( .A1(n2353), .A2(n85), .ZN(n38) );
  AND2_X1 U40 ( .A1(n2356), .A2(n85), .ZN(n39) );
  AND2_X1 U41 ( .A1(n2360), .A2(n85), .ZN(n40) );
  AND2_X1 U42 ( .A1(n1912), .A2(n142), .ZN(n41) );
  AND2_X1 U43 ( .A1(n1916), .A2(n142), .ZN(n42) );
  AND2_X1 U44 ( .A1(n1919), .A2(n142), .ZN(n43) );
  AND2_X1 U45 ( .A1(n1924), .A2(n142), .ZN(n44) );
  AND2_X1 U46 ( .A1(ADD_WR[2]), .A2(ADD_WR[1]), .ZN(n45) );
  AND2_X1 U47 ( .A1(ENABLE), .A2(n492), .ZN(n46) );
  AND2_X1 U48 ( .A1(n5), .A2(n4), .ZN(n47) );
  AND2_X1 U49 ( .A1(n6), .A2(n4), .ZN(n48) );
  AND2_X1 U50 ( .A1(n9), .A2(n4), .ZN(n49) );
  AND2_X1 U51 ( .A1(n10), .A2(n4), .ZN(n50) );
  AND2_X1 U52 ( .A1(n7), .A2(n4), .ZN(n51) );
  AND2_X1 U53 ( .A1(n8), .A2(n4), .ZN(n52) );
  AND2_X1 U54 ( .A1(n11), .A2(n4), .ZN(n53) );
  NOR2_X1 U55 ( .A1(n2346), .A2(n516), .ZN(n54) );
  NOR2_X1 U56 ( .A1(n2350), .A2(n516), .ZN(n55) );
  NOR2_X1 U57 ( .A1(n2354), .A2(n516), .ZN(n56) );
  NOR2_X1 U58 ( .A1(n1909), .A2(n944), .ZN(n57) );
  NOR2_X1 U59 ( .A1(n1913), .A2(n944), .ZN(n58) );
  NOR2_X1 U60 ( .A1(n1917), .A2(n944), .ZN(n59) );
  AND2_X1 U61 ( .A1(RD1), .A2(n46), .ZN(n60) );
  AND2_X1 U62 ( .A1(RD2), .A2(n46), .ZN(n61) );
  NAND2_X1 U63 ( .A1(n2611), .A2(n2594), .ZN(n62) );
  NAND2_X1 U64 ( .A1(n2332), .A2(n2312), .ZN(n63) );
  NAND2_X1 U65 ( .A1(n2611), .A2(n2598), .ZN(n64) );
  NAND2_X1 U66 ( .A1(n2332), .A2(n2316), .ZN(n65) );
  AND2_X1 U67 ( .A1(n2617), .A2(n2616), .ZN(n66) );
  AND2_X1 U68 ( .A1(n2340), .A2(n2339), .ZN(n67) );
  BUF_X1 U69 ( .A(n493), .Z(n492) );
  BUF_X1 U70 ( .A(n1442), .Z(n146) );
  BUF_X1 U71 ( .A(n1442), .Z(n147) );
  BUF_X1 U72 ( .A(n1442), .Z(n148) );
  BUF_X1 U73 ( .A(n1944), .Z(n314) );
  BUF_X1 U74 ( .A(n1944), .Z(n315) );
  BUF_X1 U75 ( .A(n43), .Z(n164) );
  BUF_X1 U76 ( .A(n42), .Z(n152) );
  BUF_X1 U77 ( .A(n43), .Z(n165) );
  BUF_X1 U78 ( .A(n42), .Z(n153) );
  BUF_X1 U79 ( .A(n1436), .Z(n131) );
  BUF_X1 U80 ( .A(n1436), .Z(n132) );
  BUF_X1 U81 ( .A(n63), .Z(n128) );
  BUF_X1 U82 ( .A(n63), .Z(n129) );
  BUF_X1 U83 ( .A(n1934), .Z(n297) );
  BUF_X1 U84 ( .A(n1934), .Z(n296) );
  BUF_X1 U85 ( .A(n1929), .Z(n285) );
  BUF_X1 U86 ( .A(n1929), .Z(n284) );
  BUF_X1 U87 ( .A(n2378), .Z(n362) );
  BUF_X1 U88 ( .A(n2378), .Z(n363) );
  BUF_X1 U89 ( .A(n39), .Z(n107) );
  BUF_X1 U90 ( .A(n38), .Z(n95) );
  BUF_X1 U91 ( .A(n37), .Z(n80) );
  BUF_X1 U92 ( .A(n39), .Z(n108) );
  BUF_X1 U93 ( .A(n38), .Z(n96) );
  BUF_X1 U94 ( .A(n37), .Z(n81) );
  BUF_X1 U95 ( .A(n41), .Z(n137) );
  BUF_X1 U96 ( .A(n41), .Z(n138) );
  BUF_X1 U97 ( .A(n44), .Z(n179) );
  BUF_X1 U98 ( .A(n44), .Z(n180) );
  BUF_X1 U99 ( .A(n1949), .Z(n321) );
  BUF_X1 U100 ( .A(n1949), .Z(n320) );
  BUF_X1 U101 ( .A(n1937), .Z(n303) );
  BUF_X1 U102 ( .A(n1932), .Z(n291) );
  BUF_X1 U103 ( .A(n1937), .Z(n302) );
  BUF_X1 U104 ( .A(n1932), .Z(n290) );
  BUF_X1 U105 ( .A(n2359), .Z(n326) );
  BUF_X1 U106 ( .A(n2359), .Z(n327) );
  BUF_X1 U107 ( .A(n1943), .Z(n312) );
  BUF_X1 U108 ( .A(n1923), .Z(n279) );
  BUF_X1 U109 ( .A(n1943), .Z(n311) );
  BUF_X1 U110 ( .A(n1923), .Z(n278) );
  BUF_X1 U111 ( .A(n924), .Z(n101) );
  BUF_X1 U112 ( .A(n921), .Z(n89) );
  BUF_X1 U113 ( .A(n916), .Z(n74) );
  BUF_X1 U114 ( .A(n924), .Z(n102) );
  BUF_X1 U115 ( .A(n921), .Z(n90) );
  BUF_X1 U116 ( .A(n916), .Z(n75) );
  BUF_X1 U117 ( .A(n1445), .Z(n158) );
  BUF_X1 U118 ( .A(n1445), .Z(n159) );
  BUF_X1 U119 ( .A(n1947), .Z(n318) );
  BUF_X1 U120 ( .A(n1947), .Z(n317) );
  BUF_X1 U121 ( .A(n2358), .Z(n323) );
  BUF_X1 U122 ( .A(n2358), .Z(n324) );
  BUF_X1 U123 ( .A(n1921), .Z(n276) );
  BUF_X1 U124 ( .A(n1921), .Z(n275) );
  BUF_X1 U125 ( .A(n1936), .Z(n300) );
  BUF_X1 U126 ( .A(n1931), .Z(n288) );
  BUF_X1 U127 ( .A(n1936), .Z(n299) );
  BUF_X1 U128 ( .A(n1931), .Z(n287) );
  BUF_X1 U129 ( .A(n1941), .Z(n309) );
  BUF_X1 U130 ( .A(n1941), .Z(n308) );
  BUF_X1 U131 ( .A(n925), .Z(n104) );
  BUF_X1 U132 ( .A(n925), .Z(n105) );
  BUF_X1 U133 ( .A(n1446), .Z(n161) );
  BUF_X1 U134 ( .A(n1446), .Z(n162) );
  BUF_X1 U135 ( .A(n1928), .Z(n282) );
  BUF_X1 U136 ( .A(n1928), .Z(n281) );
  BUF_X1 U137 ( .A(n1933), .Z(n294) );
  BUF_X1 U138 ( .A(n1933), .Z(n293) );
  BUF_X1 U139 ( .A(n1938), .Z(n305) );
  BUF_X1 U140 ( .A(n1938), .Z(n306) );
  BUF_X1 U141 ( .A(n40), .Z(n122) );
  BUF_X1 U142 ( .A(n40), .Z(n123) );
  BUF_X1 U143 ( .A(n65), .Z(n125) );
  BUF_X1 U144 ( .A(n65), .Z(n126) );
  BUF_X1 U145 ( .A(n83), .Z(n85) );
  BUF_X1 U146 ( .A(n140), .Z(n142) );
  BUF_X1 U147 ( .A(n43), .Z(n166) );
  BUF_X1 U148 ( .A(n42), .Z(n154) );
  BUF_X1 U149 ( .A(n1944), .Z(n316) );
  BUF_X1 U150 ( .A(n83), .Z(n86) );
  BUF_X1 U151 ( .A(n140), .Z(n143) );
  BUF_X1 U152 ( .A(n84), .Z(n87) );
  BUF_X1 U153 ( .A(n141), .Z(n144) );
  BUF_X1 U154 ( .A(n1436), .Z(n133) );
  BUF_X1 U155 ( .A(n63), .Z(n130) );
  BUF_X1 U156 ( .A(n1934), .Z(n298) );
  BUF_X1 U157 ( .A(n1929), .Z(n286) );
  BUF_X1 U158 ( .A(n2378), .Z(n364) );
  BUF_X1 U159 ( .A(n39), .Z(n109) );
  BUF_X1 U160 ( .A(n38), .Z(n97) );
  BUF_X1 U161 ( .A(n37), .Z(n82) );
  BUF_X1 U162 ( .A(n41), .Z(n139) );
  BUF_X1 U163 ( .A(n44), .Z(n181) );
  BUF_X1 U164 ( .A(n1949), .Z(n322) );
  BUF_X1 U165 ( .A(n2359), .Z(n328) );
  BUF_X1 U166 ( .A(n1943), .Z(n313) );
  BUF_X1 U167 ( .A(n1923), .Z(n280) );
  BUF_X1 U168 ( .A(n1937), .Z(n304) );
  BUF_X1 U169 ( .A(n1932), .Z(n292) );
  BUF_X1 U170 ( .A(n924), .Z(n103) );
  BUF_X1 U171 ( .A(n921), .Z(n91) );
  BUF_X1 U172 ( .A(n916), .Z(n76) );
  BUF_X1 U173 ( .A(n1445), .Z(n160) );
  BUF_X1 U174 ( .A(n1947), .Z(n319) );
  BUF_X1 U175 ( .A(n2358), .Z(n325) );
  BUF_X1 U176 ( .A(n1921), .Z(n277) );
  BUF_X1 U177 ( .A(n1941), .Z(n310) );
  BUF_X1 U178 ( .A(n1936), .Z(n301) );
  BUF_X1 U179 ( .A(n1931), .Z(n289) );
  BUF_X1 U180 ( .A(n925), .Z(n106) );
  BUF_X1 U181 ( .A(n1446), .Z(n163) );
  BUF_X1 U182 ( .A(n1928), .Z(n283) );
  BUF_X1 U183 ( .A(n1933), .Z(n295) );
  BUF_X1 U184 ( .A(n1938), .Z(n307) );
  BUF_X1 U185 ( .A(n40), .Z(n124) );
  BUF_X1 U186 ( .A(n65), .Z(n127) );
  BUF_X1 U187 ( .A(n403), .Z(n493) );
  BUF_X1 U188 ( .A(n84), .Z(n88) );
  BUF_X1 U189 ( .A(n141), .Z(n145) );
  BUF_X1 U190 ( .A(n403), .Z(n494) );
  BUF_X1 U191 ( .A(n403), .Z(n495) );
  BUF_X1 U192 ( .A(n404), .Z(n496) );
  BUF_X1 U193 ( .A(n404), .Z(n497) );
  BUF_X1 U194 ( .A(n404), .Z(n498) );
  BUF_X1 U195 ( .A(n405), .Z(n499) );
  BUF_X1 U196 ( .A(n405), .Z(n500) );
  BUF_X1 U197 ( .A(n405), .Z(n501) );
  BUF_X1 U198 ( .A(n406), .Z(n502) );
  BUF_X1 U199 ( .A(n406), .Z(n503) );
  BUF_X1 U200 ( .A(n406), .Z(n504) );
  BUF_X1 U201 ( .A(n407), .Z(n505) );
  BUF_X1 U202 ( .A(n407), .Z(n506) );
  BUF_X1 U203 ( .A(n48), .Z(n257) );
  BUF_X1 U204 ( .A(n48), .Z(n258) );
  BUF_X1 U205 ( .A(n1438), .Z(n134) );
  BUF_X1 U206 ( .A(n1438), .Z(n135) );
  BUF_X1 U207 ( .A(n62), .Z(n71) );
  BUF_X1 U208 ( .A(n62), .Z(n72) );
  BUF_X1 U209 ( .A(n2370), .Z(n344) );
  BUF_X1 U210 ( .A(n2370), .Z(n345) );
  BUF_X1 U211 ( .A(n2365), .Z(n332) );
  BUF_X1 U212 ( .A(n2365), .Z(n333) );
  BUF_X1 U213 ( .A(n56), .Z(n119) );
  BUF_X1 U214 ( .A(n56), .Z(n120) );
  BUF_X1 U215 ( .A(n59), .Z(n176) );
  BUF_X1 U216 ( .A(n59), .Z(n177) );
  BUF_X1 U217 ( .A(n58), .Z(n167) );
  BUF_X1 U218 ( .A(n58), .Z(n168) );
  BUF_X1 U219 ( .A(n2381), .Z(n368) );
  BUF_X1 U220 ( .A(n2381), .Z(n369) );
  BUF_X1 U221 ( .A(n2373), .Z(n350) );
  BUF_X1 U222 ( .A(n2368), .Z(n338) );
  BUF_X1 U223 ( .A(n2373), .Z(n351) );
  BUF_X1 U224 ( .A(n2368), .Z(n339) );
  BUF_X1 U225 ( .A(n2377), .Z(n359) );
  BUF_X1 U226 ( .A(n2377), .Z(n360) );
  BUF_X1 U227 ( .A(n2380), .Z(n365) );
  BUF_X1 U228 ( .A(n2380), .Z(n366) );
  BUF_X1 U229 ( .A(n2372), .Z(n347) );
  BUF_X1 U230 ( .A(n2367), .Z(n335) );
  BUF_X1 U231 ( .A(n2372), .Z(n348) );
  BUF_X1 U232 ( .A(n2367), .Z(n336) );
  BUF_X1 U233 ( .A(n2376), .Z(n356) );
  BUF_X1 U234 ( .A(n2376), .Z(n357) );
  BUF_X1 U235 ( .A(n922), .Z(n92) );
  BUF_X1 U236 ( .A(n917), .Z(n77) );
  BUF_X1 U237 ( .A(n922), .Z(n93) );
  BUF_X1 U238 ( .A(n917), .Z(n78) );
  BUF_X1 U239 ( .A(n1443), .Z(n149) );
  BUF_X1 U240 ( .A(n1443), .Z(n150) );
  BUF_X1 U241 ( .A(n2364), .Z(n329) );
  BUF_X1 U242 ( .A(n2364), .Z(n330) );
  BUF_X1 U243 ( .A(n2369), .Z(n341) );
  BUF_X1 U244 ( .A(n2369), .Z(n342) );
  BUF_X1 U245 ( .A(n2374), .Z(n353) );
  BUF_X1 U246 ( .A(n2374), .Z(n354) );
  BUF_X1 U247 ( .A(n55), .Z(n110) );
  BUF_X1 U248 ( .A(n54), .Z(n98) );
  BUF_X1 U249 ( .A(n55), .Z(n111) );
  BUF_X1 U250 ( .A(n54), .Z(n99) );
  BUF_X1 U251 ( .A(n57), .Z(n155) );
  BUF_X1 U252 ( .A(n57), .Z(n156) );
  BUF_X1 U253 ( .A(n64), .Z(n68) );
  BUF_X1 U254 ( .A(n64), .Z(n69) );
  BUF_X1 U255 ( .A(n48), .Z(n259) );
  BUF_X1 U256 ( .A(n1438), .Z(n136) );
  BUF_X1 U257 ( .A(n62), .Z(n73) );
  BUF_X1 U258 ( .A(n2370), .Z(n346) );
  BUF_X1 U259 ( .A(n2365), .Z(n334) );
  BUF_X1 U260 ( .A(n56), .Z(n121) );
  BUF_X1 U261 ( .A(n59), .Z(n178) );
  BUF_X1 U262 ( .A(n58), .Z(n169) );
  BUF_X1 U263 ( .A(n2381), .Z(n370) );
  BUF_X1 U264 ( .A(n2377), .Z(n361) );
  BUF_X1 U265 ( .A(n2373), .Z(n352) );
  BUF_X1 U266 ( .A(n2368), .Z(n340) );
  BUF_X1 U267 ( .A(n2380), .Z(n367) );
  BUF_X1 U268 ( .A(n2376), .Z(n358) );
  BUF_X1 U269 ( .A(n2372), .Z(n349) );
  BUF_X1 U270 ( .A(n2367), .Z(n337) );
  BUF_X1 U271 ( .A(n922), .Z(n94) );
  BUF_X1 U272 ( .A(n917), .Z(n79) );
  BUF_X1 U273 ( .A(n1443), .Z(n151) );
  BUF_X1 U274 ( .A(n2364), .Z(n331) );
  BUF_X1 U275 ( .A(n2369), .Z(n343) );
  BUF_X1 U276 ( .A(n2374), .Z(n355) );
  BUF_X1 U277 ( .A(n55), .Z(n112) );
  BUF_X1 U278 ( .A(n54), .Z(n100) );
  BUF_X1 U279 ( .A(n57), .Z(n157) );
  BUF_X1 U280 ( .A(n64), .Z(n70) );
  BUF_X1 U281 ( .A(n920), .Z(n83) );
  BUF_X1 U282 ( .A(n1441), .Z(n140) );
  BUF_X1 U283 ( .A(n920), .Z(n84) );
  BUF_X1 U284 ( .A(n1441), .Z(n141) );
  BUF_X1 U285 ( .A(n408), .Z(n405) );
  BUF_X1 U286 ( .A(n408), .Z(n406) );
  BUF_X1 U287 ( .A(n409), .Z(n403) );
  BUF_X1 U288 ( .A(n409), .Z(n404) );
  BUF_X1 U289 ( .A(n408), .Z(n407) );
  BUF_X1 U290 ( .A(n13), .Z(n182) );
  BUF_X1 U291 ( .A(n13), .Z(n183) );
  BUF_X1 U292 ( .A(n14), .Z(n185) );
  BUF_X1 U293 ( .A(n14), .Z(n186) );
  BUF_X1 U294 ( .A(n15), .Z(n188) );
  BUF_X1 U295 ( .A(n15), .Z(n189) );
  BUF_X1 U296 ( .A(n16), .Z(n191) );
  BUF_X1 U297 ( .A(n16), .Z(n192) );
  BUF_X1 U298 ( .A(n17), .Z(n194) );
  BUF_X1 U299 ( .A(n17), .Z(n195) );
  BUF_X1 U300 ( .A(n18), .Z(n197) );
  BUF_X1 U301 ( .A(n18), .Z(n198) );
  BUF_X1 U302 ( .A(n19), .Z(n200) );
  BUF_X1 U303 ( .A(n19), .Z(n201) );
  BUF_X1 U304 ( .A(n20), .Z(n203) );
  BUF_X1 U305 ( .A(n20), .Z(n204) );
  BUF_X1 U306 ( .A(n21), .Z(n206) );
  BUF_X1 U307 ( .A(n21), .Z(n207) );
  BUF_X1 U308 ( .A(n22), .Z(n209) );
  BUF_X1 U309 ( .A(n22), .Z(n210) );
  BUF_X1 U310 ( .A(n23), .Z(n212) );
  BUF_X1 U311 ( .A(n23), .Z(n213) );
  BUF_X1 U312 ( .A(n24), .Z(n215) );
  BUF_X1 U313 ( .A(n24), .Z(n216) );
  BUF_X1 U314 ( .A(n25), .Z(n218) );
  BUF_X1 U315 ( .A(n25), .Z(n219) );
  BUF_X1 U316 ( .A(n26), .Z(n221) );
  BUF_X1 U317 ( .A(n26), .Z(n222) );
  BUF_X1 U318 ( .A(n27), .Z(n224) );
  BUF_X1 U319 ( .A(n27), .Z(n225) );
  BUF_X1 U320 ( .A(n28), .Z(n227) );
  BUF_X1 U321 ( .A(n28), .Z(n228) );
  BUF_X1 U322 ( .A(n29), .Z(n230) );
  BUF_X1 U323 ( .A(n29), .Z(n231) );
  BUF_X1 U324 ( .A(n30), .Z(n233) );
  BUF_X1 U325 ( .A(n30), .Z(n234) );
  BUF_X1 U326 ( .A(n31), .Z(n236) );
  BUF_X1 U327 ( .A(n31), .Z(n237) );
  BUF_X1 U328 ( .A(n32), .Z(n239) );
  BUF_X1 U329 ( .A(n32), .Z(n240) );
  BUF_X1 U330 ( .A(n33), .Z(n242) );
  BUF_X1 U331 ( .A(n33), .Z(n243) );
  BUF_X1 U332 ( .A(n34), .Z(n245) );
  BUF_X1 U333 ( .A(n34), .Z(n246) );
  BUF_X1 U334 ( .A(n35), .Z(n248) );
  BUF_X1 U335 ( .A(n35), .Z(n249) );
  BUF_X1 U336 ( .A(n36), .Z(n251) );
  BUF_X1 U337 ( .A(n36), .Z(n252) );
  BUF_X1 U338 ( .A(n47), .Z(n254) );
  BUF_X1 U339 ( .A(n47), .Z(n255) );
  BUF_X1 U340 ( .A(n49), .Z(n260) );
  BUF_X1 U341 ( .A(n49), .Z(n261) );
  BUF_X1 U342 ( .A(n50), .Z(n263) );
  BUF_X1 U343 ( .A(n50), .Z(n264) );
  BUF_X1 U344 ( .A(n51), .Z(n266) );
  BUF_X1 U345 ( .A(n51), .Z(n267) );
  BUF_X1 U346 ( .A(n52), .Z(n269) );
  BUF_X1 U347 ( .A(n52), .Z(n270) );
  BUF_X1 U348 ( .A(n53), .Z(n272) );
  BUF_X1 U349 ( .A(n53), .Z(n273) );
  BUF_X1 U350 ( .A(n1448), .Z(n170) );
  BUF_X1 U351 ( .A(n1448), .Z(n171) );
  BUF_X1 U352 ( .A(n927), .Z(n113) );
  BUF_X1 U353 ( .A(n927), .Z(n114) );
  BUF_X1 U354 ( .A(n13), .Z(n184) );
  BUF_X1 U355 ( .A(n14), .Z(n187) );
  BUF_X1 U356 ( .A(n15), .Z(n190) );
  BUF_X1 U357 ( .A(n16), .Z(n193) );
  BUF_X1 U358 ( .A(n17), .Z(n196) );
  BUF_X1 U359 ( .A(n18), .Z(n199) );
  BUF_X1 U360 ( .A(n19), .Z(n202) );
  BUF_X1 U361 ( .A(n20), .Z(n205) );
  BUF_X1 U362 ( .A(n21), .Z(n208) );
  BUF_X1 U363 ( .A(n22), .Z(n211) );
  BUF_X1 U364 ( .A(n23), .Z(n214) );
  BUF_X1 U365 ( .A(n24), .Z(n217) );
  BUF_X1 U366 ( .A(n25), .Z(n220) );
  BUF_X1 U367 ( .A(n26), .Z(n223) );
  BUF_X1 U368 ( .A(n27), .Z(n226) );
  BUF_X1 U369 ( .A(n28), .Z(n229) );
  BUF_X1 U370 ( .A(n29), .Z(n232) );
  BUF_X1 U371 ( .A(n30), .Z(n235) );
  BUF_X1 U372 ( .A(n31), .Z(n238) );
  BUF_X1 U373 ( .A(n32), .Z(n241) );
  BUF_X1 U374 ( .A(n33), .Z(n244) );
  BUF_X1 U375 ( .A(n34), .Z(n247) );
  BUF_X1 U376 ( .A(n35), .Z(n250) );
  BUF_X1 U377 ( .A(n36), .Z(n253) );
  BUF_X1 U378 ( .A(n47), .Z(n256) );
  BUF_X1 U379 ( .A(n49), .Z(n262) );
  BUF_X1 U380 ( .A(n50), .Z(n265) );
  BUF_X1 U381 ( .A(n51), .Z(n268) );
  BUF_X1 U382 ( .A(n52), .Z(n271) );
  BUF_X1 U383 ( .A(n53), .Z(n274) );
  BUF_X1 U384 ( .A(n1448), .Z(n172) );
  BUF_X1 U385 ( .A(n927), .Z(n115) );
  BUF_X1 U386 ( .A(RST), .Z(n408) );
  BUF_X1 U387 ( .A(RST), .Z(n409) );
  BUF_X1 U388 ( .A(n60), .Z(n116) );
  BUF_X1 U389 ( .A(n61), .Z(n173) );
  BUF_X1 U390 ( .A(n60), .Z(n117) );
  BUF_X1 U391 ( .A(n61), .Z(n174) );
  BUF_X1 U392 ( .A(n60), .Z(n118) );
  BUF_X1 U393 ( .A(n61), .Z(n175) );
  INV_X1 U394 ( .A(DATAIN[0]), .ZN(n371) );
  INV_X1 U395 ( .A(DATAIN[1]), .ZN(n372) );
  INV_X1 U396 ( .A(DATAIN[2]), .ZN(n373) );
  INV_X1 U397 ( .A(DATAIN[3]), .ZN(n374) );
  INV_X1 U398 ( .A(DATAIN[4]), .ZN(n375) );
  INV_X1 U399 ( .A(DATAIN[5]), .ZN(n376) );
  INV_X1 U400 ( .A(DATAIN[6]), .ZN(n377) );
  INV_X1 U401 ( .A(DATAIN[7]), .ZN(n378) );
  INV_X1 U402 ( .A(DATAIN[8]), .ZN(n379) );
  INV_X1 U403 ( .A(DATAIN[10]), .ZN(n381) );
  INV_X1 U404 ( .A(DATAIN[11]), .ZN(n382) );
  INV_X1 U405 ( .A(DATAIN[12]), .ZN(n383) );
  INV_X1 U406 ( .A(DATAIN[13]), .ZN(n384) );
  INV_X1 U407 ( .A(DATAIN[14]), .ZN(n385) );
  INV_X1 U408 ( .A(DATAIN[15]), .ZN(n386) );
  INV_X1 U409 ( .A(DATAIN[16]), .ZN(n387) );
  INV_X1 U410 ( .A(DATAIN[17]), .ZN(n388) );
  INV_X1 U411 ( .A(DATAIN[18]), .ZN(n389) );
  INV_X1 U412 ( .A(DATAIN[19]), .ZN(n390) );
  INV_X1 U413 ( .A(DATAIN[20]), .ZN(n391) );
  INV_X1 U414 ( .A(DATAIN[21]), .ZN(n392) );
  INV_X1 U415 ( .A(DATAIN[22]), .ZN(n393) );
  INV_X1 U416 ( .A(DATAIN[23]), .ZN(n394) );
  INV_X1 U417 ( .A(DATAIN[24]), .ZN(n395) );
  INV_X1 U418 ( .A(DATAIN[25]), .ZN(n396) );
  INV_X1 U419 ( .A(DATAIN[26]), .ZN(n397) );
  INV_X1 U420 ( .A(DATAIN[27]), .ZN(n398) );
  INV_X1 U421 ( .A(DATAIN[28]), .ZN(n399) );
  INV_X1 U422 ( .A(DATAIN[29]), .ZN(n400) );
  INV_X1 U423 ( .A(DATAIN[30]), .ZN(n401) );
  INV_X1 U424 ( .A(DATAIN[31]), .ZN(n402) );
  INV_X1 U425 ( .A(DATAIN[9]), .ZN(n380) );
  CLKBUF_X1 U426 ( .A(n506), .Z(n410) );
  CLKBUF_X1 U427 ( .A(n506), .Z(n411) );
  CLKBUF_X1 U428 ( .A(n506), .Z(n412) );
  CLKBUF_X1 U429 ( .A(n506), .Z(n413) );
  CLKBUF_X1 U430 ( .A(n506), .Z(n414) );
  CLKBUF_X1 U431 ( .A(n505), .Z(n415) );
  CLKBUF_X1 U432 ( .A(n505), .Z(n416) );
  CLKBUF_X1 U433 ( .A(n505), .Z(n417) );
  CLKBUF_X1 U434 ( .A(n505), .Z(n418) );
  CLKBUF_X1 U435 ( .A(n505), .Z(n419) );
  CLKBUF_X1 U436 ( .A(n505), .Z(n420) );
  CLKBUF_X1 U437 ( .A(n504), .Z(n421) );
  CLKBUF_X1 U438 ( .A(n504), .Z(n422) );
  CLKBUF_X1 U439 ( .A(n504), .Z(n423) );
  CLKBUF_X1 U440 ( .A(n504), .Z(n424) );
  CLKBUF_X1 U441 ( .A(n504), .Z(n425) );
  CLKBUF_X1 U442 ( .A(n504), .Z(n426) );
  CLKBUF_X1 U443 ( .A(n503), .Z(n427) );
  CLKBUF_X1 U444 ( .A(n503), .Z(n428) );
  CLKBUF_X1 U445 ( .A(n503), .Z(n429) );
  CLKBUF_X1 U446 ( .A(n503), .Z(n430) );
  CLKBUF_X1 U447 ( .A(n503), .Z(n431) );
  CLKBUF_X1 U448 ( .A(n503), .Z(n432) );
  CLKBUF_X1 U449 ( .A(n502), .Z(n433) );
  CLKBUF_X1 U450 ( .A(n502), .Z(n434) );
  CLKBUF_X1 U451 ( .A(n502), .Z(n435) );
  CLKBUF_X1 U452 ( .A(n502), .Z(n436) );
  CLKBUF_X1 U453 ( .A(n502), .Z(n437) );
  CLKBUF_X1 U454 ( .A(n502), .Z(n438) );
  CLKBUF_X1 U455 ( .A(n501), .Z(n439) );
  CLKBUF_X1 U456 ( .A(n501), .Z(n440) );
  CLKBUF_X1 U457 ( .A(n501), .Z(n441) );
  CLKBUF_X1 U458 ( .A(n501), .Z(n442) );
  CLKBUF_X1 U459 ( .A(n501), .Z(n443) );
  CLKBUF_X1 U460 ( .A(n501), .Z(n444) );
  CLKBUF_X1 U461 ( .A(n500), .Z(n445) );
  CLKBUF_X1 U462 ( .A(n500), .Z(n446) );
  CLKBUF_X1 U463 ( .A(n500), .Z(n447) );
  CLKBUF_X1 U464 ( .A(n500), .Z(n448) );
  CLKBUF_X1 U465 ( .A(n500), .Z(n449) );
  CLKBUF_X1 U466 ( .A(n500), .Z(n450) );
  CLKBUF_X1 U467 ( .A(n499), .Z(n451) );
  CLKBUF_X1 U468 ( .A(n499), .Z(n452) );
  CLKBUF_X1 U469 ( .A(n499), .Z(n453) );
  CLKBUF_X1 U470 ( .A(n499), .Z(n454) );
  CLKBUF_X1 U471 ( .A(n499), .Z(n455) );
  CLKBUF_X1 U472 ( .A(n499), .Z(n456) );
  CLKBUF_X1 U473 ( .A(n498), .Z(n457) );
  CLKBUF_X1 U474 ( .A(n498), .Z(n458) );
  CLKBUF_X1 U475 ( .A(n498), .Z(n459) );
  CLKBUF_X1 U476 ( .A(n498), .Z(n460) );
  CLKBUF_X1 U477 ( .A(n498), .Z(n461) );
  CLKBUF_X1 U478 ( .A(n498), .Z(n462) );
  CLKBUF_X1 U479 ( .A(n497), .Z(n463) );
  CLKBUF_X1 U480 ( .A(n497), .Z(n464) );
  CLKBUF_X1 U481 ( .A(n497), .Z(n465) );
  CLKBUF_X1 U482 ( .A(n497), .Z(n466) );
  CLKBUF_X1 U483 ( .A(n497), .Z(n467) );
  CLKBUF_X1 U484 ( .A(n497), .Z(n468) );
  CLKBUF_X1 U485 ( .A(n496), .Z(n469) );
  CLKBUF_X1 U486 ( .A(n496), .Z(n470) );
  CLKBUF_X1 U487 ( .A(n496), .Z(n471) );
  CLKBUF_X1 U488 ( .A(n496), .Z(n472) );
  CLKBUF_X1 U489 ( .A(n496), .Z(n473) );
  CLKBUF_X1 U490 ( .A(n496), .Z(n474) );
  CLKBUF_X1 U491 ( .A(n495), .Z(n475) );
  CLKBUF_X1 U492 ( .A(n495), .Z(n476) );
  CLKBUF_X1 U493 ( .A(n495), .Z(n477) );
  CLKBUF_X1 U494 ( .A(n495), .Z(n478) );
  CLKBUF_X1 U495 ( .A(n495), .Z(n479) );
  CLKBUF_X1 U496 ( .A(n495), .Z(n480) );
  CLKBUF_X1 U497 ( .A(n494), .Z(n481) );
  CLKBUF_X1 U498 ( .A(n494), .Z(n482) );
  CLKBUF_X1 U499 ( .A(n494), .Z(n483) );
  CLKBUF_X1 U500 ( .A(n494), .Z(n484) );
  CLKBUF_X1 U501 ( .A(n494), .Z(n485) );
  CLKBUF_X1 U502 ( .A(n494), .Z(n486) );
  CLKBUF_X1 U503 ( .A(n493), .Z(n487) );
  CLKBUF_X1 U504 ( .A(n493), .Z(n488) );
  CLKBUF_X1 U505 ( .A(n493), .Z(n489) );
  CLKBUF_X1 U506 ( .A(n493), .Z(n490) );
  CLKBUF_X1 U507 ( .A(n493), .Z(n491) );
  INV_X1 U508 ( .A(ADD_WR[0]), .ZN(n1907) );
  NAND3_X1 U509 ( .A1(n2619), .A2(n2618), .A3(n66), .ZN(n507) );
  NAND2_X1 U510 ( .A1(n116), .A2(n507), .ZN(n516) );
  INV_X1 U511 ( .A(n516), .ZN(n920) );
  OAI211_X1 U512 ( .C1(n3998), .C2(n68), .A(n2605), .B(n2604), .ZN(n508) );
  AOI221_X1 U513 ( .B1(n353), .B2(n1843), .C1(n362), .C2(n2750), .A(n508), 
        .ZN(n511) );
  NOR2_X1 U514 ( .A1(n4125), .A2(n71), .ZN(n509) );
  NOR4_X1 U515 ( .A1(n2615), .A2(n2610), .A3(n2601), .A4(n509), .ZN(n510) );
  NAND2_X1 U516 ( .A1(n511), .A2(n510), .ZN(n513) );
  OR2_X1 U517 ( .A1(n2347), .A2(n516), .ZN(n917) );
  NAND2_X1 U518 ( .A1(n2348), .A2(n85), .ZN(n916) );
  OAI22_X1 U519 ( .A1(n939), .A2(n77), .B1(n938), .B2(n74), .ZN(n512) );
  AOI221_X1 U520 ( .B1(n85), .B2(n513), .C1(n80), .C2(n1519), .A(n512), .ZN(
        n521) );
  OR2_X1 U521 ( .A1(n2351), .A2(n516), .ZN(n922) );
  NAND2_X1 U522 ( .A1(n2352), .A2(n85), .ZN(n921) );
  OAI22_X1 U523 ( .A1(n2718), .A2(n92), .B1(n2686), .B2(n89), .ZN(n514) );
  AOI221_X1 U524 ( .B1(n98), .B2(n1487), .C1(n95), .C2(n2814), .A(n514), .ZN(
        n520) );
  NAND2_X1 U525 ( .A1(n2361), .A2(n85), .ZN(n925) );
  NAND2_X1 U526 ( .A1(n2355), .A2(n85), .ZN(n924) );
  OAI22_X1 U527 ( .A1(n3646), .A2(n104), .B1(n2942), .B2(n101), .ZN(n515) );
  AOI221_X1 U528 ( .B1(n110), .B2(n2782), .C1(n107), .C2(n3582), .A(n515), 
        .ZN(n519) );
  NAND4_X1 U529 ( .A1(n66), .A2(n2618), .A3(n116), .A4(n2619), .ZN(n927) );
  OAI22_X1 U530 ( .A1(n2622), .A2(n116), .B1(n371), .B2(n113), .ZN(n517) );
  AOI221_X1 U531 ( .B1(n122), .B2(n3614), .C1(n119), .C2(n1617), .A(n517), 
        .ZN(n518) );
  NAND4_X1 U532 ( .A1(n521), .A2(n520), .A3(n519), .A4(n518), .ZN(n2983) );
  OAI211_X1 U533 ( .C1(n3999), .C2(n68), .A(n2587), .B(n2586), .ZN(n522) );
  AOI221_X1 U534 ( .B1(n353), .B2(n1844), .C1(n362), .C2(n2751), .A(n522), 
        .ZN(n525) );
  NOR2_X1 U535 ( .A1(n4124), .A2(n71), .ZN(n523) );
  NOR4_X1 U536 ( .A1(n2591), .A2(n2590), .A3(n2585), .A4(n523), .ZN(n524) );
  NAND2_X1 U537 ( .A1(n525), .A2(n524), .ZN(n527) );
  OAI22_X1 U538 ( .A1(n956), .A2(n77), .B1(n955), .B2(n74), .ZN(n526) );
  AOI221_X1 U539 ( .B1(n88), .B2(n527), .C1(n80), .C2(n1520), .A(n526), .ZN(
        n534) );
  OAI22_X1 U540 ( .A1(n2719), .A2(n92), .B1(n2687), .B2(n89), .ZN(n528) );
  AOI221_X1 U541 ( .B1(n98), .B2(n1488), .C1(n95), .C2(n2815), .A(n528), .ZN(
        n533) );
  OAI22_X1 U542 ( .A1(n3647), .A2(n104), .B1(n2943), .B2(n101), .ZN(n529) );
  AOI221_X1 U543 ( .B1(n110), .B2(n2783), .C1(n107), .C2(n3583), .A(n529), 
        .ZN(n532) );
  OAI22_X1 U544 ( .A1(n2623), .A2(n118), .B1(n372), .B2(n113), .ZN(n530) );
  AOI221_X1 U545 ( .B1(n122), .B2(n3615), .C1(n119), .C2(n1618), .A(n530), 
        .ZN(n531) );
  NAND4_X1 U546 ( .A1(n534), .A2(n533), .A3(n532), .A4(n531), .ZN(n2984) );
  OAI211_X1 U547 ( .C1(n4000), .C2(n68), .A(n2580), .B(n2579), .ZN(n535) );
  AOI221_X1 U548 ( .B1(n353), .B2(n1845), .C1(n362), .C2(n2752), .A(n535), 
        .ZN(n538) );
  NOR2_X1 U549 ( .A1(n4123), .A2(n71), .ZN(n536) );
  NOR4_X1 U550 ( .A1(n2584), .A2(n2583), .A3(n2578), .A4(n536), .ZN(n537) );
  NAND2_X1 U551 ( .A1(n538), .A2(n537), .ZN(n540) );
  OAI22_X1 U552 ( .A1(n972), .A2(n77), .B1(n971), .B2(n74), .ZN(n539) );
  AOI221_X1 U553 ( .B1(n88), .B2(n540), .C1(n80), .C2(n1521), .A(n539), .ZN(
        n547) );
  OAI22_X1 U554 ( .A1(n2720), .A2(n92), .B1(n2688), .B2(n89), .ZN(n541) );
  AOI221_X1 U555 ( .B1(n98), .B2(n1489), .C1(n95), .C2(n2816), .A(n541), .ZN(
        n546) );
  OAI22_X1 U556 ( .A1(n3648), .A2(n104), .B1(n2944), .B2(n101), .ZN(n542) );
  AOI221_X1 U557 ( .B1(n110), .B2(n2784), .C1(n107), .C2(n3584), .A(n542), 
        .ZN(n545) );
  OAI22_X1 U558 ( .A1(n2624), .A2(n118), .B1(n373), .B2(n113), .ZN(n543) );
  AOI221_X1 U559 ( .B1(n122), .B2(n3616), .C1(n119), .C2(n1619), .A(n543), 
        .ZN(n544) );
  NAND4_X1 U560 ( .A1(n547), .A2(n546), .A3(n545), .A4(n544), .ZN(n2985) );
  OAI211_X1 U561 ( .C1(n4001), .C2(n68), .A(n2573), .B(n2572), .ZN(n548) );
  AOI221_X1 U562 ( .B1(n353), .B2(n1846), .C1(n362), .C2(n2753), .A(n548), 
        .ZN(n551) );
  NOR2_X1 U563 ( .A1(n4122), .A2(n71), .ZN(n549) );
  NOR4_X1 U564 ( .A1(n2577), .A2(n2576), .A3(n2571), .A4(n549), .ZN(n550) );
  NAND2_X1 U565 ( .A1(n551), .A2(n550), .ZN(n553) );
  OAI22_X1 U566 ( .A1(n988), .A2(n77), .B1(n987), .B2(n74), .ZN(n552) );
  AOI221_X1 U567 ( .B1(n88), .B2(n553), .C1(n80), .C2(n1522), .A(n552), .ZN(
        n560) );
  OAI22_X1 U568 ( .A1(n2721), .A2(n92), .B1(n2689), .B2(n89), .ZN(n554) );
  AOI221_X1 U569 ( .B1(n98), .B2(n1490), .C1(n95), .C2(n2817), .A(n554), .ZN(
        n559) );
  OAI22_X1 U570 ( .A1(n3649), .A2(n104), .B1(n2945), .B2(n101), .ZN(n555) );
  AOI221_X1 U571 ( .B1(n110), .B2(n2785), .C1(n107), .C2(n3585), .A(n555), 
        .ZN(n558) );
  OAI22_X1 U572 ( .A1(n2625), .A2(n118), .B1(n374), .B2(n113), .ZN(n556) );
  AOI221_X1 U573 ( .B1(n122), .B2(n3617), .C1(n119), .C2(n1620), .A(n556), 
        .ZN(n557) );
  NAND4_X1 U574 ( .A1(n560), .A2(n559), .A3(n558), .A4(n557), .ZN(n2986) );
  OAI211_X1 U575 ( .C1(n4002), .C2(n68), .A(n2566), .B(n2565), .ZN(n561) );
  AOI221_X1 U576 ( .B1(n353), .B2(n1847), .C1(n362), .C2(n2754), .A(n561), 
        .ZN(n564) );
  NOR2_X1 U577 ( .A1(n4121), .A2(n71), .ZN(n562) );
  NOR4_X1 U578 ( .A1(n2570), .A2(n2569), .A3(n2564), .A4(n562), .ZN(n563) );
  NAND2_X1 U579 ( .A1(n564), .A2(n563), .ZN(n566) );
  OAI22_X1 U580 ( .A1(n1004), .A2(n77), .B1(n1003), .B2(n74), .ZN(n565) );
  AOI221_X1 U581 ( .B1(n88), .B2(n566), .C1(n80), .C2(n1523), .A(n565), .ZN(
        n573) );
  OAI22_X1 U582 ( .A1(n2722), .A2(n92), .B1(n2690), .B2(n89), .ZN(n567) );
  AOI221_X1 U583 ( .B1(n98), .B2(n1491), .C1(n95), .C2(n2818), .A(n567), .ZN(
        n572) );
  OAI22_X1 U584 ( .A1(n3650), .A2(n104), .B1(n2946), .B2(n101), .ZN(n568) );
  AOI221_X1 U585 ( .B1(n110), .B2(n2786), .C1(n107), .C2(n3586), .A(n568), 
        .ZN(n571) );
  OAI22_X1 U586 ( .A1(n2626), .A2(n118), .B1(n375), .B2(n113), .ZN(n569) );
  AOI221_X1 U587 ( .B1(n122), .B2(n3618), .C1(n119), .C2(n1621), .A(n569), 
        .ZN(n570) );
  NAND4_X1 U588 ( .A1(n573), .A2(n572), .A3(n571), .A4(n570), .ZN(n2987) );
  OAI211_X1 U589 ( .C1(n4003), .C2(n68), .A(n2559), .B(n2558), .ZN(n574) );
  AOI221_X1 U590 ( .B1(n353), .B2(n1848), .C1(n362), .C2(n2755), .A(n574), 
        .ZN(n577) );
  NOR2_X1 U591 ( .A1(n4120), .A2(n71), .ZN(n575) );
  NOR4_X1 U592 ( .A1(n2563), .A2(n2562), .A3(n2557), .A4(n575), .ZN(n576) );
  NAND2_X1 U593 ( .A1(n577), .A2(n576), .ZN(n579) );
  OAI22_X1 U594 ( .A1(n1020), .A2(n77), .B1(n1019), .B2(n74), .ZN(n578) );
  AOI221_X1 U595 ( .B1(n87), .B2(n579), .C1(n80), .C2(n1524), .A(n578), .ZN(
        n586) );
  OAI22_X1 U596 ( .A1(n2723), .A2(n92), .B1(n2691), .B2(n89), .ZN(n580) );
  AOI221_X1 U597 ( .B1(n98), .B2(n1492), .C1(n95), .C2(n2819), .A(n580), .ZN(
        n585) );
  OAI22_X1 U598 ( .A1(n3651), .A2(n104), .B1(n2947), .B2(n101), .ZN(n581) );
  AOI221_X1 U599 ( .B1(n110), .B2(n2787), .C1(n107), .C2(n3587), .A(n581), 
        .ZN(n584) );
  OAI22_X1 U600 ( .A1(n2627), .A2(n118), .B1(n376), .B2(n113), .ZN(n582) );
  AOI221_X1 U601 ( .B1(n122), .B2(n3619), .C1(n119), .C2(n1622), .A(n582), 
        .ZN(n583) );
  NAND4_X1 U602 ( .A1(n586), .A2(n585), .A3(n584), .A4(n583), .ZN(n2988) );
  OAI211_X1 U603 ( .C1(n4004), .C2(n68), .A(n2552), .B(n2551), .ZN(n587) );
  AOI221_X1 U604 ( .B1(n353), .B2(n1849), .C1(n362), .C2(n2756), .A(n587), 
        .ZN(n590) );
  NOR2_X1 U605 ( .A1(n4119), .A2(n71), .ZN(n588) );
  NOR4_X1 U606 ( .A1(n2556), .A2(n2555), .A3(n2550), .A4(n588), .ZN(n589) );
  NAND2_X1 U607 ( .A1(n590), .A2(n589), .ZN(n592) );
  OAI22_X1 U608 ( .A1(n1036), .A2(n77), .B1(n1035), .B2(n74), .ZN(n591) );
  AOI221_X1 U609 ( .B1(n87), .B2(n592), .C1(n80), .C2(n1525), .A(n591), .ZN(
        n599) );
  OAI22_X1 U610 ( .A1(n2724), .A2(n92), .B1(n2692), .B2(n89), .ZN(n593) );
  AOI221_X1 U611 ( .B1(n98), .B2(n1493), .C1(n95), .C2(n2820), .A(n593), .ZN(
        n598) );
  OAI22_X1 U612 ( .A1(n3652), .A2(n104), .B1(n2948), .B2(n101), .ZN(n594) );
  AOI221_X1 U613 ( .B1(n110), .B2(n2788), .C1(n107), .C2(n3588), .A(n594), 
        .ZN(n597) );
  OAI22_X1 U614 ( .A1(n2628), .A2(n118), .B1(n377), .B2(n113), .ZN(n595) );
  AOI221_X1 U615 ( .B1(n122), .B2(n3620), .C1(n119), .C2(n1623), .A(n595), 
        .ZN(n596) );
  NAND4_X1 U616 ( .A1(n599), .A2(n598), .A3(n597), .A4(n596), .ZN(n2989) );
  OAI211_X1 U617 ( .C1(n4005), .C2(n68), .A(n2545), .B(n2544), .ZN(n600) );
  AOI221_X1 U618 ( .B1(n353), .B2(n1850), .C1(n362), .C2(n2757), .A(n600), 
        .ZN(n603) );
  NOR2_X1 U619 ( .A1(n4118), .A2(n71), .ZN(n601) );
  NOR4_X1 U620 ( .A1(n2549), .A2(n2548), .A3(n2543), .A4(n601), .ZN(n602) );
  NAND2_X1 U621 ( .A1(n603), .A2(n602), .ZN(n605) );
  OAI22_X1 U622 ( .A1(n1052), .A2(n77), .B1(n1051), .B2(n74), .ZN(n604) );
  AOI221_X1 U623 ( .B1(n87), .B2(n605), .C1(n80), .C2(n1526), .A(n604), .ZN(
        n612) );
  OAI22_X1 U624 ( .A1(n2725), .A2(n92), .B1(n2693), .B2(n89), .ZN(n606) );
  AOI221_X1 U625 ( .B1(n98), .B2(n1494), .C1(n95), .C2(n2821), .A(n606), .ZN(
        n611) );
  OAI22_X1 U626 ( .A1(n3653), .A2(n104), .B1(n2949), .B2(n101), .ZN(n607) );
  AOI221_X1 U627 ( .B1(n110), .B2(n2789), .C1(n107), .C2(n3589), .A(n607), 
        .ZN(n610) );
  OAI22_X1 U628 ( .A1(n2629), .A2(n118), .B1(n378), .B2(n113), .ZN(n608) );
  AOI221_X1 U629 ( .B1(n122), .B2(n3621), .C1(n119), .C2(n1624), .A(n608), 
        .ZN(n609) );
  NAND4_X1 U630 ( .A1(n612), .A2(n611), .A3(n610), .A4(n609), .ZN(n2990) );
  OAI211_X1 U631 ( .C1(n4006), .C2(n68), .A(n2538), .B(n2537), .ZN(n613) );
  AOI221_X1 U632 ( .B1(n353), .B2(n1851), .C1(n362), .C2(n2758), .A(n613), 
        .ZN(n616) );
  NOR2_X1 U633 ( .A1(n4117), .A2(n71), .ZN(n614) );
  NOR4_X1 U634 ( .A1(n2542), .A2(n2541), .A3(n2536), .A4(n614), .ZN(n615) );
  NAND2_X1 U635 ( .A1(n616), .A2(n615), .ZN(n618) );
  OAI22_X1 U636 ( .A1(n1068), .A2(n77), .B1(n1067), .B2(n74), .ZN(n617) );
  AOI221_X1 U637 ( .B1(n87), .B2(n618), .C1(n80), .C2(n1527), .A(n617), .ZN(
        n625) );
  OAI22_X1 U638 ( .A1(n2726), .A2(n92), .B1(n2694), .B2(n89), .ZN(n619) );
  AOI221_X1 U639 ( .B1(n98), .B2(n1495), .C1(n95), .C2(n2822), .A(n619), .ZN(
        n624) );
  OAI22_X1 U640 ( .A1(n3654), .A2(n104), .B1(n2950), .B2(n101), .ZN(n620) );
  AOI221_X1 U641 ( .B1(n110), .B2(n2790), .C1(n107), .C2(n3590), .A(n620), 
        .ZN(n623) );
  OAI22_X1 U642 ( .A1(n2630), .A2(n118), .B1(n379), .B2(n113), .ZN(n621) );
  AOI221_X1 U643 ( .B1(n122), .B2(n3622), .C1(n119), .C2(n1625), .A(n621), 
        .ZN(n622) );
  NAND4_X1 U644 ( .A1(n625), .A2(n624), .A3(n623), .A4(n622), .ZN(n2991) );
  OAI211_X1 U645 ( .C1(n4007), .C2(n68), .A(n2531), .B(n2530), .ZN(n626) );
  AOI221_X1 U646 ( .B1(n353), .B2(n1852), .C1(n362), .C2(n2759), .A(n626), 
        .ZN(n629) );
  NOR2_X1 U647 ( .A1(n4116), .A2(n71), .ZN(n627) );
  NOR4_X1 U648 ( .A1(n2535), .A2(n2534), .A3(n2529), .A4(n627), .ZN(n628) );
  NAND2_X1 U649 ( .A1(n629), .A2(n628), .ZN(n631) );
  OAI22_X1 U650 ( .A1(n1084), .A2(n77), .B1(n1083), .B2(n74), .ZN(n630) );
  AOI221_X1 U651 ( .B1(n87), .B2(n631), .C1(n80), .C2(n1528), .A(n630), .ZN(
        n638) );
  OAI22_X1 U652 ( .A1(n2727), .A2(n92), .B1(n2695), .B2(n89), .ZN(n632) );
  AOI221_X1 U653 ( .B1(n98), .B2(n1496), .C1(n95), .C2(n2823), .A(n632), .ZN(
        n637) );
  OAI22_X1 U654 ( .A1(n3655), .A2(n104), .B1(n2951), .B2(n101), .ZN(n633) );
  AOI221_X1 U655 ( .B1(n110), .B2(n2791), .C1(n107), .C2(n3591), .A(n633), 
        .ZN(n636) );
  OAI22_X1 U656 ( .A1(n2631), .A2(n118), .B1(n380), .B2(n113), .ZN(n634) );
  AOI221_X1 U657 ( .B1(n122), .B2(n3623), .C1(n119), .C2(n1626), .A(n634), 
        .ZN(n635) );
  NAND4_X1 U658 ( .A1(n638), .A2(n637), .A3(n636), .A4(n635), .ZN(n2992) );
  OAI211_X1 U659 ( .C1(n4008), .C2(n68), .A(n2524), .B(n2523), .ZN(n639) );
  AOI221_X1 U660 ( .B1(n353), .B2(n1853), .C1(n362), .C2(n2760), .A(n639), 
        .ZN(n642) );
  NOR2_X1 U661 ( .A1(n4115), .A2(n71), .ZN(n640) );
  NOR4_X1 U662 ( .A1(n2528), .A2(n2527), .A3(n2522), .A4(n640), .ZN(n641) );
  NAND2_X1 U663 ( .A1(n642), .A2(n641), .ZN(n644) );
  OAI22_X1 U664 ( .A1(n1100), .A2(n77), .B1(n1099), .B2(n74), .ZN(n643) );
  AOI221_X1 U665 ( .B1(n87), .B2(n644), .C1(n80), .C2(n1529), .A(n643), .ZN(
        n651) );
  OAI22_X1 U666 ( .A1(n2728), .A2(n92), .B1(n2696), .B2(n89), .ZN(n645) );
  AOI221_X1 U667 ( .B1(n98), .B2(n1497), .C1(n95), .C2(n2824), .A(n645), .ZN(
        n650) );
  OAI22_X1 U668 ( .A1(n3656), .A2(n104), .B1(n2952), .B2(n101), .ZN(n646) );
  AOI221_X1 U669 ( .B1(n110), .B2(n2792), .C1(n107), .C2(n3592), .A(n646), 
        .ZN(n649) );
  OAI22_X1 U670 ( .A1(n2632), .A2(n118), .B1(n381), .B2(n113), .ZN(n647) );
  AOI221_X1 U671 ( .B1(n122), .B2(n3624), .C1(n119), .C2(n1627), .A(n647), 
        .ZN(n648) );
  NAND4_X1 U672 ( .A1(n651), .A2(n650), .A3(n649), .A4(n648), .ZN(n2993) );
  OAI211_X1 U673 ( .C1(n4009), .C2(n68), .A(n2517), .B(n2516), .ZN(n652) );
  AOI221_X1 U674 ( .B1(n353), .B2(n1854), .C1(n362), .C2(n2761), .A(n652), 
        .ZN(n655) );
  NOR2_X1 U675 ( .A1(n4114), .A2(n71), .ZN(n653) );
  NOR4_X1 U676 ( .A1(n2521), .A2(n2520), .A3(n2515), .A4(n653), .ZN(n654) );
  NAND2_X1 U677 ( .A1(n655), .A2(n654), .ZN(n657) );
  OAI22_X1 U678 ( .A1(n1116), .A2(n77), .B1(n1115), .B2(n74), .ZN(n656) );
  AOI221_X1 U679 ( .B1(n87), .B2(n657), .C1(n80), .C2(n1530), .A(n656), .ZN(
        n664) );
  OAI22_X1 U680 ( .A1(n2729), .A2(n92), .B1(n2697), .B2(n89), .ZN(n658) );
  AOI221_X1 U681 ( .B1(n98), .B2(n1498), .C1(n95), .C2(n2825), .A(n658), .ZN(
        n663) );
  OAI22_X1 U682 ( .A1(n3657), .A2(n104), .B1(n2953), .B2(n101), .ZN(n659) );
  AOI221_X1 U683 ( .B1(n110), .B2(n2793), .C1(n107), .C2(n3593), .A(n659), 
        .ZN(n662) );
  OAI22_X1 U684 ( .A1(n2633), .A2(n117), .B1(n382), .B2(n113), .ZN(n660) );
  AOI221_X1 U685 ( .B1(n122), .B2(n3625), .C1(n119), .C2(n1628), .A(n660), 
        .ZN(n661) );
  NAND4_X1 U686 ( .A1(n664), .A2(n663), .A3(n662), .A4(n661), .ZN(n2994) );
  OAI211_X1 U687 ( .C1(n4010), .C2(n69), .A(n2510), .B(n2509), .ZN(n665) );
  AOI221_X1 U688 ( .B1(n354), .B2(n1855), .C1(n363), .C2(n2762), .A(n665), 
        .ZN(n668) );
  NOR2_X1 U689 ( .A1(n4113), .A2(n72), .ZN(n666) );
  NOR4_X1 U690 ( .A1(n2514), .A2(n2513), .A3(n2508), .A4(n666), .ZN(n667) );
  NAND2_X1 U691 ( .A1(n668), .A2(n667), .ZN(n670) );
  OAI22_X1 U692 ( .A1(n1132), .A2(n78), .B1(n1131), .B2(n75), .ZN(n669) );
  AOI221_X1 U693 ( .B1(n87), .B2(n670), .C1(n81), .C2(n1531), .A(n669), .ZN(
        n677) );
  OAI22_X1 U694 ( .A1(n2730), .A2(n93), .B1(n2698), .B2(n90), .ZN(n671) );
  AOI221_X1 U695 ( .B1(n99), .B2(n1499), .C1(n96), .C2(n2826), .A(n671), .ZN(
        n676) );
  OAI22_X1 U696 ( .A1(n3658), .A2(n105), .B1(n2954), .B2(n102), .ZN(n672) );
  AOI221_X1 U697 ( .B1(n111), .B2(n2794), .C1(n108), .C2(n3594), .A(n672), 
        .ZN(n675) );
  OAI22_X1 U698 ( .A1(n2634), .A2(n117), .B1(n383), .B2(n114), .ZN(n673) );
  AOI221_X1 U699 ( .B1(n123), .B2(n3626), .C1(n120), .C2(n1629), .A(n673), 
        .ZN(n674) );
  NAND4_X1 U700 ( .A1(n677), .A2(n676), .A3(n675), .A4(n674), .ZN(n2995) );
  OAI211_X1 U701 ( .C1(n4011), .C2(n69), .A(n2503), .B(n2502), .ZN(n678) );
  AOI221_X1 U702 ( .B1(n354), .B2(n1856), .C1(n363), .C2(n2763), .A(n678), 
        .ZN(n681) );
  NOR2_X1 U703 ( .A1(n4112), .A2(n72), .ZN(n679) );
  NOR4_X1 U704 ( .A1(n2507), .A2(n2506), .A3(n2501), .A4(n679), .ZN(n680) );
  NAND2_X1 U705 ( .A1(n681), .A2(n680), .ZN(n683) );
  OAI22_X1 U706 ( .A1(n1148), .A2(n78), .B1(n1147), .B2(n75), .ZN(n682) );
  AOI221_X1 U707 ( .B1(n87), .B2(n683), .C1(n81), .C2(n1532), .A(n682), .ZN(
        n690) );
  OAI22_X1 U708 ( .A1(n2731), .A2(n93), .B1(n2699), .B2(n90), .ZN(n684) );
  AOI221_X1 U709 ( .B1(n99), .B2(n1500), .C1(n96), .C2(n2827), .A(n684), .ZN(
        n689) );
  OAI22_X1 U710 ( .A1(n3659), .A2(n105), .B1(n2955), .B2(n102), .ZN(n685) );
  AOI221_X1 U711 ( .B1(n111), .B2(n2795), .C1(n108), .C2(n3595), .A(n685), 
        .ZN(n688) );
  OAI22_X1 U712 ( .A1(n2635), .A2(n117), .B1(n384), .B2(n114), .ZN(n686) );
  AOI221_X1 U713 ( .B1(n123), .B2(n3627), .C1(n120), .C2(n1630), .A(n686), 
        .ZN(n687) );
  NAND4_X1 U714 ( .A1(n690), .A2(n689), .A3(n688), .A4(n687), .ZN(n2996) );
  OAI211_X1 U715 ( .C1(n4012), .C2(n69), .A(n2496), .B(n2495), .ZN(n691) );
  AOI221_X1 U716 ( .B1(n354), .B2(n1857), .C1(n363), .C2(n2764), .A(n691), 
        .ZN(n694) );
  NOR2_X1 U717 ( .A1(n4111), .A2(n72), .ZN(n692) );
  NOR4_X1 U718 ( .A1(n2500), .A2(n2499), .A3(n2494), .A4(n692), .ZN(n693) );
  NAND2_X1 U719 ( .A1(n694), .A2(n693), .ZN(n696) );
  OAI22_X1 U720 ( .A1(n1164), .A2(n78), .B1(n1163), .B2(n75), .ZN(n695) );
  AOI221_X1 U721 ( .B1(n87), .B2(n696), .C1(n81), .C2(n1533), .A(n695), .ZN(
        n703) );
  OAI22_X1 U722 ( .A1(n2732), .A2(n93), .B1(n2700), .B2(n90), .ZN(n697) );
  AOI221_X1 U723 ( .B1(n99), .B2(n1501), .C1(n96), .C2(n2828), .A(n697), .ZN(
        n702) );
  OAI22_X1 U724 ( .A1(n3660), .A2(n105), .B1(n2956), .B2(n102), .ZN(n698) );
  AOI221_X1 U725 ( .B1(n111), .B2(n2796), .C1(n108), .C2(n3596), .A(n698), 
        .ZN(n701) );
  OAI22_X1 U726 ( .A1(n2636), .A2(n117), .B1(n385), .B2(n114), .ZN(n699) );
  AOI221_X1 U727 ( .B1(n123), .B2(n3628), .C1(n120), .C2(n1631), .A(n699), 
        .ZN(n700) );
  NAND4_X1 U728 ( .A1(n703), .A2(n702), .A3(n701), .A4(n700), .ZN(n2997) );
  OAI211_X1 U729 ( .C1(n4013), .C2(n69), .A(n2489), .B(n2488), .ZN(n704) );
  AOI221_X1 U730 ( .B1(n354), .B2(n1858), .C1(n363), .C2(n2765), .A(n704), 
        .ZN(n707) );
  NOR2_X1 U731 ( .A1(n4110), .A2(n72), .ZN(n705) );
  NOR4_X1 U732 ( .A1(n2493), .A2(n2492), .A3(n2487), .A4(n705), .ZN(n706) );
  NAND2_X1 U733 ( .A1(n707), .A2(n706), .ZN(n709) );
  OAI22_X1 U734 ( .A1(n1180), .A2(n78), .B1(n1179), .B2(n75), .ZN(n708) );
  AOI221_X1 U735 ( .B1(n87), .B2(n709), .C1(n81), .C2(n1534), .A(n708), .ZN(
        n716) );
  OAI22_X1 U736 ( .A1(n2733), .A2(n93), .B1(n2701), .B2(n90), .ZN(n710) );
  AOI221_X1 U737 ( .B1(n99), .B2(n1502), .C1(n96), .C2(n2829), .A(n710), .ZN(
        n715) );
  OAI22_X1 U738 ( .A1(n3661), .A2(n105), .B1(n2957), .B2(n102), .ZN(n711) );
  AOI221_X1 U739 ( .B1(n111), .B2(n2797), .C1(n108), .C2(n3597), .A(n711), 
        .ZN(n714) );
  OAI22_X1 U740 ( .A1(n2637), .A2(n117), .B1(n386), .B2(n114), .ZN(n712) );
  AOI221_X1 U741 ( .B1(n123), .B2(n3629), .C1(n120), .C2(n1632), .A(n712), 
        .ZN(n713) );
  NAND4_X1 U742 ( .A1(n716), .A2(n715), .A3(n714), .A4(n713), .ZN(n2998) );
  OAI211_X1 U743 ( .C1(n4014), .C2(n69), .A(n2482), .B(n2481), .ZN(n717) );
  AOI221_X1 U744 ( .B1(n354), .B2(n1859), .C1(n363), .C2(n2766), .A(n717), 
        .ZN(n720) );
  NOR2_X1 U745 ( .A1(n4109), .A2(n72), .ZN(n718) );
  NOR4_X1 U746 ( .A1(n2486), .A2(n2485), .A3(n2480), .A4(n718), .ZN(n719) );
  NAND2_X1 U747 ( .A1(n720), .A2(n719), .ZN(n722) );
  OAI22_X1 U748 ( .A1(n1196), .A2(n78), .B1(n1195), .B2(n75), .ZN(n721) );
  AOI221_X1 U749 ( .B1(n86), .B2(n722), .C1(n81), .C2(n1535), .A(n721), .ZN(
        n729) );
  OAI22_X1 U750 ( .A1(n2734), .A2(n93), .B1(n2702), .B2(n90), .ZN(n723) );
  AOI221_X1 U751 ( .B1(n99), .B2(n1503), .C1(n96), .C2(n2830), .A(n723), .ZN(
        n728) );
  OAI22_X1 U752 ( .A1(n3662), .A2(n105), .B1(n2958), .B2(n102), .ZN(n724) );
  AOI221_X1 U753 ( .B1(n111), .B2(n2798), .C1(n108), .C2(n3598), .A(n724), 
        .ZN(n727) );
  OAI22_X1 U754 ( .A1(n2638), .A2(n117), .B1(n387), .B2(n114), .ZN(n725) );
  AOI221_X1 U755 ( .B1(n123), .B2(n3630), .C1(n120), .C2(n1633), .A(n725), 
        .ZN(n726) );
  NAND4_X1 U756 ( .A1(n729), .A2(n728), .A3(n727), .A4(n726), .ZN(n2999) );
  OAI211_X1 U757 ( .C1(n4015), .C2(n69), .A(n2475), .B(n2474), .ZN(n730) );
  AOI221_X1 U758 ( .B1(n354), .B2(n1860), .C1(n363), .C2(n2767), .A(n730), 
        .ZN(n733) );
  NOR2_X1 U759 ( .A1(n4108), .A2(n72), .ZN(n731) );
  NOR4_X1 U760 ( .A1(n2479), .A2(n2478), .A3(n2473), .A4(n731), .ZN(n732) );
  NAND2_X1 U761 ( .A1(n733), .A2(n732), .ZN(n735) );
  OAI22_X1 U762 ( .A1(n1212), .A2(n78), .B1(n1211), .B2(n75), .ZN(n734) );
  AOI221_X1 U763 ( .B1(n86), .B2(n735), .C1(n81), .C2(n1536), .A(n734), .ZN(
        n742) );
  OAI22_X1 U764 ( .A1(n2735), .A2(n93), .B1(n2703), .B2(n90), .ZN(n736) );
  AOI221_X1 U765 ( .B1(n99), .B2(n1504), .C1(n96), .C2(n2831), .A(n736), .ZN(
        n741) );
  OAI22_X1 U766 ( .A1(n3663), .A2(n105), .B1(n2959), .B2(n102), .ZN(n737) );
  AOI221_X1 U767 ( .B1(n111), .B2(n2799), .C1(n108), .C2(n3599), .A(n737), 
        .ZN(n740) );
  OAI22_X1 U768 ( .A1(n2639), .A2(n117), .B1(n388), .B2(n114), .ZN(n738) );
  AOI221_X1 U769 ( .B1(n123), .B2(n3631), .C1(n120), .C2(n1634), .A(n738), 
        .ZN(n739) );
  NAND4_X1 U770 ( .A1(n742), .A2(n741), .A3(n740), .A4(n739), .ZN(n3000) );
  OAI211_X1 U771 ( .C1(n4016), .C2(n69), .A(n2468), .B(n2467), .ZN(n743) );
  AOI221_X1 U772 ( .B1(n354), .B2(n1861), .C1(n363), .C2(n2768), .A(n743), 
        .ZN(n746) );
  NOR2_X1 U773 ( .A1(n4107), .A2(n72), .ZN(n744) );
  NOR4_X1 U774 ( .A1(n2472), .A2(n2471), .A3(n2466), .A4(n744), .ZN(n745) );
  NAND2_X1 U775 ( .A1(n746), .A2(n745), .ZN(n748) );
  OAI22_X1 U776 ( .A1(n1228), .A2(n78), .B1(n1227), .B2(n75), .ZN(n747) );
  AOI221_X1 U777 ( .B1(n86), .B2(n748), .C1(n81), .C2(n1537), .A(n747), .ZN(
        n755) );
  OAI22_X1 U778 ( .A1(n2736), .A2(n93), .B1(n2704), .B2(n90), .ZN(n749) );
  AOI221_X1 U779 ( .B1(n99), .B2(n1505), .C1(n96), .C2(n2832), .A(n749), .ZN(
        n754) );
  OAI22_X1 U780 ( .A1(n3664), .A2(n105), .B1(n2960), .B2(n102), .ZN(n750) );
  AOI221_X1 U781 ( .B1(n111), .B2(n2800), .C1(n108), .C2(n3600), .A(n750), 
        .ZN(n753) );
  OAI22_X1 U782 ( .A1(n2640), .A2(n117), .B1(n389), .B2(n114), .ZN(n751) );
  AOI221_X1 U783 ( .B1(n123), .B2(n3632), .C1(n120), .C2(n1635), .A(n751), 
        .ZN(n752) );
  NAND4_X1 U784 ( .A1(n755), .A2(n754), .A3(n753), .A4(n752), .ZN(n3001) );
  OAI211_X1 U785 ( .C1(n4017), .C2(n69), .A(n2461), .B(n2460), .ZN(n756) );
  AOI221_X1 U786 ( .B1(n354), .B2(n1862), .C1(n363), .C2(n2769), .A(n756), 
        .ZN(n759) );
  NOR2_X1 U787 ( .A1(n4106), .A2(n72), .ZN(n757) );
  NOR4_X1 U788 ( .A1(n2465), .A2(n2464), .A3(n2459), .A4(n757), .ZN(n758) );
  NAND2_X1 U789 ( .A1(n759), .A2(n758), .ZN(n761) );
  OAI22_X1 U790 ( .A1(n1244), .A2(n78), .B1(n1243), .B2(n75), .ZN(n760) );
  AOI221_X1 U791 ( .B1(n86), .B2(n761), .C1(n81), .C2(n1538), .A(n760), .ZN(
        n768) );
  OAI22_X1 U792 ( .A1(n2737), .A2(n93), .B1(n2705), .B2(n90), .ZN(n762) );
  AOI221_X1 U793 ( .B1(n99), .B2(n1506), .C1(n96), .C2(n2833), .A(n762), .ZN(
        n767) );
  OAI22_X1 U794 ( .A1(n3665), .A2(n105), .B1(n2961), .B2(n102), .ZN(n763) );
  AOI221_X1 U795 ( .B1(n111), .B2(n2801), .C1(n108), .C2(n3601), .A(n763), 
        .ZN(n766) );
  OAI22_X1 U796 ( .A1(n2641), .A2(n117), .B1(n390), .B2(n114), .ZN(n764) );
  AOI221_X1 U797 ( .B1(n123), .B2(n3633), .C1(n120), .C2(n1636), .A(n764), 
        .ZN(n765) );
  NAND4_X1 U798 ( .A1(n768), .A2(n767), .A3(n766), .A4(n765), .ZN(n3002) );
  OAI211_X1 U799 ( .C1(n4018), .C2(n69), .A(n2454), .B(n2453), .ZN(n769) );
  AOI221_X1 U800 ( .B1(n354), .B2(n1863), .C1(n363), .C2(n2770), .A(n769), 
        .ZN(n772) );
  NOR2_X1 U801 ( .A1(n4105), .A2(n72), .ZN(n770) );
  NOR4_X1 U802 ( .A1(n2458), .A2(n2457), .A3(n2452), .A4(n770), .ZN(n771) );
  NAND2_X1 U803 ( .A1(n772), .A2(n771), .ZN(n774) );
  OAI22_X1 U804 ( .A1(n1260), .A2(n78), .B1(n1259), .B2(n75), .ZN(n773) );
  AOI221_X1 U805 ( .B1(n86), .B2(n774), .C1(n81), .C2(n1539), .A(n773), .ZN(
        n781) );
  OAI22_X1 U806 ( .A1(n2738), .A2(n93), .B1(n2706), .B2(n90), .ZN(n775) );
  AOI221_X1 U807 ( .B1(n99), .B2(n1507), .C1(n96), .C2(n2834), .A(n775), .ZN(
        n780) );
  OAI22_X1 U808 ( .A1(n3666), .A2(n105), .B1(n2962), .B2(n102), .ZN(n776) );
  AOI221_X1 U809 ( .B1(n111), .B2(n2802), .C1(n108), .C2(n3602), .A(n776), 
        .ZN(n779) );
  OAI22_X1 U810 ( .A1(n2642), .A2(n117), .B1(n391), .B2(n114), .ZN(n777) );
  AOI221_X1 U811 ( .B1(n123), .B2(n3634), .C1(n120), .C2(n1637), .A(n777), 
        .ZN(n778) );
  NAND4_X1 U812 ( .A1(n781), .A2(n780), .A3(n779), .A4(n778), .ZN(n3003) );
  OAI211_X1 U813 ( .C1(n4019), .C2(n69), .A(n2447), .B(n2446), .ZN(n782) );
  AOI221_X1 U814 ( .B1(n354), .B2(n1864), .C1(n363), .C2(n2771), .A(n782), 
        .ZN(n785) );
  NOR2_X1 U815 ( .A1(n4104), .A2(n72), .ZN(n783) );
  NOR4_X1 U816 ( .A1(n2451), .A2(n2450), .A3(n2445), .A4(n783), .ZN(n784) );
  NAND2_X1 U817 ( .A1(n785), .A2(n784), .ZN(n787) );
  OAI22_X1 U818 ( .A1(n1276), .A2(n78), .B1(n1275), .B2(n75), .ZN(n786) );
  AOI221_X1 U819 ( .B1(n86), .B2(n787), .C1(n81), .C2(n1540), .A(n786), .ZN(
        n794) );
  OAI22_X1 U820 ( .A1(n2739), .A2(n93), .B1(n2707), .B2(n90), .ZN(n788) );
  AOI221_X1 U821 ( .B1(n99), .B2(n1508), .C1(n96), .C2(n2835), .A(n788), .ZN(
        n793) );
  OAI22_X1 U822 ( .A1(n3667), .A2(n105), .B1(n2963), .B2(n102), .ZN(n789) );
  AOI221_X1 U823 ( .B1(n111), .B2(n2803), .C1(n108), .C2(n3603), .A(n789), 
        .ZN(n792) );
  OAI22_X1 U824 ( .A1(n2643), .A2(n117), .B1(n392), .B2(n114), .ZN(n790) );
  AOI221_X1 U825 ( .B1(n123), .B2(n3635), .C1(n120), .C2(n1638), .A(n790), 
        .ZN(n791) );
  NAND4_X1 U826 ( .A1(n794), .A2(n793), .A3(n792), .A4(n791), .ZN(n3004) );
  OAI211_X1 U827 ( .C1(n4020), .C2(n69), .A(n2440), .B(n2439), .ZN(n795) );
  AOI221_X1 U828 ( .B1(n354), .B2(n1865), .C1(n363), .C2(n2772), .A(n795), 
        .ZN(n798) );
  NOR2_X1 U829 ( .A1(n4103), .A2(n72), .ZN(n796) );
  NOR4_X1 U830 ( .A1(n2444), .A2(n2443), .A3(n2438), .A4(n796), .ZN(n797) );
  NAND2_X1 U831 ( .A1(n798), .A2(n797), .ZN(n800) );
  OAI22_X1 U832 ( .A1(n1292), .A2(n78), .B1(n1291), .B2(n75), .ZN(n799) );
  AOI221_X1 U833 ( .B1(n86), .B2(n800), .C1(n81), .C2(n1541), .A(n799), .ZN(
        n807) );
  OAI22_X1 U834 ( .A1(n2740), .A2(n93), .B1(n2708), .B2(n90), .ZN(n801) );
  AOI221_X1 U835 ( .B1(n99), .B2(n1509), .C1(n96), .C2(n2836), .A(n801), .ZN(
        n806) );
  OAI22_X1 U836 ( .A1(n3668), .A2(n105), .B1(n2964), .B2(n102), .ZN(n802) );
  AOI221_X1 U837 ( .B1(n111), .B2(n2804), .C1(n108), .C2(n3604), .A(n802), 
        .ZN(n805) );
  OAI22_X1 U838 ( .A1(n2644), .A2(n116), .B1(n393), .B2(n114), .ZN(n803) );
  AOI221_X1 U839 ( .B1(n123), .B2(n3636), .C1(n120), .C2(n1639), .A(n803), 
        .ZN(n804) );
  NAND4_X1 U840 ( .A1(n807), .A2(n806), .A3(n805), .A4(n804), .ZN(n3005) );
  OAI211_X1 U841 ( .C1(n4021), .C2(n69), .A(n2433), .B(n2432), .ZN(n808) );
  AOI221_X1 U842 ( .B1(n354), .B2(n1866), .C1(n363), .C2(n2773), .A(n808), 
        .ZN(n811) );
  NOR2_X1 U843 ( .A1(n4102), .A2(n72), .ZN(n809) );
  NOR4_X1 U844 ( .A1(n2437), .A2(n2436), .A3(n2431), .A4(n809), .ZN(n810) );
  NAND2_X1 U845 ( .A1(n811), .A2(n810), .ZN(n813) );
  OAI22_X1 U846 ( .A1(n1308), .A2(n78), .B1(n1307), .B2(n75), .ZN(n812) );
  AOI221_X1 U847 ( .B1(n86), .B2(n813), .C1(n81), .C2(n1542), .A(n812), .ZN(
        n820) );
  OAI22_X1 U848 ( .A1(n2741), .A2(n93), .B1(n2709), .B2(n90), .ZN(n814) );
  AOI221_X1 U849 ( .B1(n99), .B2(n1510), .C1(n96), .C2(n2837), .A(n814), .ZN(
        n819) );
  OAI22_X1 U850 ( .A1(n3669), .A2(n105), .B1(n2965), .B2(n102), .ZN(n815) );
  AOI221_X1 U851 ( .B1(n111), .B2(n2805), .C1(n108), .C2(n3605), .A(n815), 
        .ZN(n818) );
  OAI22_X1 U852 ( .A1(n2645), .A2(n116), .B1(n394), .B2(n114), .ZN(n816) );
  AOI221_X1 U853 ( .B1(n123), .B2(n3637), .C1(n120), .C2(n1640), .A(n816), 
        .ZN(n817) );
  NAND4_X1 U854 ( .A1(n820), .A2(n819), .A3(n818), .A4(n817), .ZN(n3006) );
  OAI211_X1 U855 ( .C1(n4022), .C2(n70), .A(n2426), .B(n2425), .ZN(n821) );
  AOI221_X1 U856 ( .B1(n355), .B2(n1867), .C1(n364), .C2(n2774), .A(n821), 
        .ZN(n824) );
  NOR2_X1 U857 ( .A1(n4101), .A2(n73), .ZN(n822) );
  NOR4_X1 U858 ( .A1(n2430), .A2(n2429), .A3(n2424), .A4(n822), .ZN(n823) );
  NAND2_X1 U859 ( .A1(n824), .A2(n823), .ZN(n826) );
  OAI22_X1 U860 ( .A1(n1324), .A2(n79), .B1(n1323), .B2(n76), .ZN(n825) );
  AOI221_X1 U861 ( .B1(n86), .B2(n826), .C1(n82), .C2(n1543), .A(n825), .ZN(
        n833) );
  OAI22_X1 U862 ( .A1(n2742), .A2(n94), .B1(n2710), .B2(n91), .ZN(n827) );
  AOI221_X1 U863 ( .B1(n100), .B2(n1511), .C1(n97), .C2(n2838), .A(n827), .ZN(
        n832) );
  OAI22_X1 U864 ( .A1(n3670), .A2(n106), .B1(n2966), .B2(n103), .ZN(n828) );
  AOI221_X1 U865 ( .B1(n112), .B2(n2806), .C1(n109), .C2(n3606), .A(n828), 
        .ZN(n831) );
  OAI22_X1 U866 ( .A1(n2646), .A2(n116), .B1(n395), .B2(n115), .ZN(n829) );
  AOI221_X1 U867 ( .B1(n124), .B2(n3638), .C1(n121), .C2(n1641), .A(n829), 
        .ZN(n830) );
  NAND4_X1 U868 ( .A1(n833), .A2(n832), .A3(n831), .A4(n830), .ZN(n3007) );
  OAI211_X1 U869 ( .C1(n4023), .C2(n70), .A(n2419), .B(n2418), .ZN(n834) );
  AOI221_X1 U870 ( .B1(n355), .B2(n1868), .C1(n364), .C2(n2775), .A(n834), 
        .ZN(n837) );
  NOR2_X1 U871 ( .A1(n4100), .A2(n73), .ZN(n835) );
  NOR4_X1 U872 ( .A1(n2423), .A2(n2422), .A3(n2417), .A4(n835), .ZN(n836) );
  NAND2_X1 U873 ( .A1(n837), .A2(n836), .ZN(n839) );
  OAI22_X1 U874 ( .A1(n1340), .A2(n79), .B1(n1339), .B2(n76), .ZN(n838) );
  AOI221_X1 U875 ( .B1(n86), .B2(n839), .C1(n82), .C2(n1544), .A(n838), .ZN(
        n846) );
  OAI22_X1 U876 ( .A1(n2743), .A2(n94), .B1(n2711), .B2(n91), .ZN(n840) );
  AOI221_X1 U877 ( .B1(n100), .B2(n1512), .C1(n97), .C2(n2839), .A(n840), .ZN(
        n845) );
  OAI22_X1 U878 ( .A1(n3671), .A2(n106), .B1(n2967), .B2(n103), .ZN(n841) );
  AOI221_X1 U879 ( .B1(n112), .B2(n2807), .C1(n109), .C2(n3607), .A(n841), 
        .ZN(n844) );
  OAI22_X1 U880 ( .A1(n2647), .A2(n116), .B1(n396), .B2(n115), .ZN(n842) );
  AOI221_X1 U881 ( .B1(n124), .B2(n3639), .C1(n121), .C2(n1642), .A(n842), 
        .ZN(n843) );
  NAND4_X1 U882 ( .A1(n846), .A2(n845), .A3(n844), .A4(n843), .ZN(n3008) );
  OAI211_X1 U883 ( .C1(n4024), .C2(n70), .A(n2412), .B(n2411), .ZN(n847) );
  AOI221_X1 U884 ( .B1(n355), .B2(n1869), .C1(n364), .C2(n2776), .A(n847), 
        .ZN(n850) );
  NOR2_X1 U885 ( .A1(n4099), .A2(n73), .ZN(n848) );
  NOR4_X1 U886 ( .A1(n2416), .A2(n2415), .A3(n2410), .A4(n848), .ZN(n849) );
  NAND2_X1 U887 ( .A1(n850), .A2(n849), .ZN(n852) );
  OAI22_X1 U888 ( .A1(n1356), .A2(n79), .B1(n1355), .B2(n76), .ZN(n851) );
  AOI221_X1 U889 ( .B1(n86), .B2(n852), .C1(n82), .C2(n1545), .A(n851), .ZN(
        n859) );
  OAI22_X1 U890 ( .A1(n2744), .A2(n94), .B1(n2712), .B2(n91), .ZN(n853) );
  AOI221_X1 U891 ( .B1(n100), .B2(n1513), .C1(n97), .C2(n2840), .A(n853), .ZN(
        n858) );
  OAI22_X1 U892 ( .A1(n3672), .A2(n106), .B1(n2968), .B2(n103), .ZN(n854) );
  AOI221_X1 U893 ( .B1(n112), .B2(n2808), .C1(n109), .C2(n3608), .A(n854), 
        .ZN(n857) );
  OAI22_X1 U894 ( .A1(n2648), .A2(n116), .B1(n397), .B2(n115), .ZN(n855) );
  AOI221_X1 U895 ( .B1(n124), .B2(n3640), .C1(n121), .C2(n1643), .A(n855), 
        .ZN(n856) );
  NAND4_X1 U896 ( .A1(n859), .A2(n858), .A3(n857), .A4(n856), .ZN(n3009) );
  OAI211_X1 U897 ( .C1(n4025), .C2(n70), .A(n2405), .B(n2404), .ZN(n860) );
  AOI221_X1 U898 ( .B1(n355), .B2(n1870), .C1(n364), .C2(n2777), .A(n860), 
        .ZN(n863) );
  NOR2_X1 U899 ( .A1(n4098), .A2(n73), .ZN(n861) );
  NOR4_X1 U900 ( .A1(n2409), .A2(n2408), .A3(n2403), .A4(n861), .ZN(n862) );
  NAND2_X1 U901 ( .A1(n863), .A2(n862), .ZN(n865) );
  OAI22_X1 U902 ( .A1(n1372), .A2(n79), .B1(n1371), .B2(n76), .ZN(n864) );
  AOI221_X1 U903 ( .B1(n86), .B2(n865), .C1(n82), .C2(n1546), .A(n864), .ZN(
        n872) );
  OAI22_X1 U904 ( .A1(n2745), .A2(n94), .B1(n2713), .B2(n91), .ZN(n866) );
  AOI221_X1 U905 ( .B1(n100), .B2(n1514), .C1(n97), .C2(n2841), .A(n866), .ZN(
        n871) );
  OAI22_X1 U906 ( .A1(n3673), .A2(n106), .B1(n2969), .B2(n103), .ZN(n867) );
  AOI221_X1 U907 ( .B1(n112), .B2(n2809), .C1(n109), .C2(n3609), .A(n867), 
        .ZN(n870) );
  OAI22_X1 U908 ( .A1(n2649), .A2(n116), .B1(n398), .B2(n115), .ZN(n868) );
  AOI221_X1 U909 ( .B1(n124), .B2(n3641), .C1(n121), .C2(n1644), .A(n868), 
        .ZN(n869) );
  NAND4_X1 U910 ( .A1(n872), .A2(n871), .A3(n870), .A4(n869), .ZN(n3010) );
  OAI211_X1 U911 ( .C1(n4026), .C2(n70), .A(n2398), .B(n2397), .ZN(n873) );
  AOI221_X1 U912 ( .B1(n355), .B2(n1871), .C1(n364), .C2(n2778), .A(n873), 
        .ZN(n876) );
  NOR2_X1 U913 ( .A1(n4097), .A2(n73), .ZN(n874) );
  NOR4_X1 U914 ( .A1(n2402), .A2(n2401), .A3(n2396), .A4(n874), .ZN(n875) );
  NAND2_X1 U915 ( .A1(n876), .A2(n875), .ZN(n878) );
  OAI22_X1 U916 ( .A1(n1388), .A2(n79), .B1(n1387), .B2(n76), .ZN(n877) );
  AOI221_X1 U917 ( .B1(n85), .B2(n878), .C1(n82), .C2(n1547), .A(n877), .ZN(
        n885) );
  OAI22_X1 U918 ( .A1(n2746), .A2(n94), .B1(n2714), .B2(n91), .ZN(n879) );
  AOI221_X1 U919 ( .B1(n100), .B2(n1515), .C1(n97), .C2(n2842), .A(n879), .ZN(
        n884) );
  OAI22_X1 U920 ( .A1(n3674), .A2(n106), .B1(n2970), .B2(n103), .ZN(n880) );
  AOI221_X1 U921 ( .B1(n112), .B2(n2810), .C1(n109), .C2(n3610), .A(n880), 
        .ZN(n883) );
  OAI22_X1 U922 ( .A1(n2650), .A2(n116), .B1(n399), .B2(n115), .ZN(n881) );
  AOI221_X1 U923 ( .B1(n124), .B2(n3642), .C1(n121), .C2(n1645), .A(n881), 
        .ZN(n882) );
  NAND4_X1 U924 ( .A1(n885), .A2(n884), .A3(n883), .A4(n882), .ZN(n3011) );
  OAI211_X1 U925 ( .C1(n4027), .C2(n70), .A(n2391), .B(n2390), .ZN(n886) );
  AOI221_X1 U926 ( .B1(n355), .B2(n1872), .C1(n364), .C2(n2779), .A(n886), 
        .ZN(n889) );
  NOR2_X1 U927 ( .A1(n4096), .A2(n73), .ZN(n887) );
  NOR4_X1 U928 ( .A1(n2395), .A2(n2394), .A3(n2389), .A4(n887), .ZN(n888) );
  NAND2_X1 U929 ( .A1(n889), .A2(n888), .ZN(n891) );
  OAI22_X1 U930 ( .A1(n1404), .A2(n79), .B1(n1403), .B2(n76), .ZN(n890) );
  AOI221_X1 U931 ( .B1(n85), .B2(n891), .C1(n82), .C2(n1548), .A(n890), .ZN(
        n898) );
  OAI22_X1 U932 ( .A1(n2747), .A2(n94), .B1(n2715), .B2(n91), .ZN(n892) );
  AOI221_X1 U933 ( .B1(n100), .B2(n1516), .C1(n97), .C2(n2843), .A(n892), .ZN(
        n897) );
  OAI22_X1 U934 ( .A1(n3675), .A2(n106), .B1(n2971), .B2(n103), .ZN(n893) );
  AOI221_X1 U935 ( .B1(n112), .B2(n2811), .C1(n109), .C2(n3611), .A(n893), 
        .ZN(n896) );
  OAI22_X1 U936 ( .A1(n2651), .A2(n116), .B1(n400), .B2(n115), .ZN(n894) );
  AOI221_X1 U937 ( .B1(n124), .B2(n3643), .C1(n121), .C2(n1646), .A(n894), 
        .ZN(n895) );
  NAND4_X1 U938 ( .A1(n898), .A2(n897), .A3(n896), .A4(n895), .ZN(n3012) );
  OAI211_X1 U939 ( .C1(n4028), .C2(n70), .A(n2384), .B(n2383), .ZN(n899) );
  AOI221_X1 U940 ( .B1(n355), .B2(n1873), .C1(n364), .C2(n2780), .A(n899), 
        .ZN(n902) );
  NOR2_X1 U941 ( .A1(n4095), .A2(n73), .ZN(n900) );
  NOR4_X1 U942 ( .A1(n2388), .A2(n2387), .A3(n2382), .A4(n900), .ZN(n901) );
  NAND2_X1 U943 ( .A1(n902), .A2(n901), .ZN(n904) );
  OAI22_X1 U944 ( .A1(n1420), .A2(n79), .B1(n1419), .B2(n76), .ZN(n903) );
  AOI221_X1 U945 ( .B1(n85), .B2(n904), .C1(n82), .C2(n1549), .A(n903), .ZN(
        n911) );
  OAI22_X1 U946 ( .A1(n2748), .A2(n94), .B1(n2716), .B2(n91), .ZN(n905) );
  AOI221_X1 U947 ( .B1(n100), .B2(n1517), .C1(n97), .C2(n2844), .A(n905), .ZN(
        n910) );
  OAI22_X1 U948 ( .A1(n3676), .A2(n106), .B1(n2972), .B2(n103), .ZN(n906) );
  AOI221_X1 U949 ( .B1(n112), .B2(n2812), .C1(n109), .C2(n3612), .A(n906), 
        .ZN(n909) );
  OAI22_X1 U950 ( .A1(n2652), .A2(n116), .B1(n401), .B2(n115), .ZN(n907) );
  AOI221_X1 U951 ( .B1(n124), .B2(n3644), .C1(n121), .C2(n1647), .A(n907), 
        .ZN(n908) );
  NAND4_X1 U952 ( .A1(n911), .A2(n910), .A3(n909), .A4(n908), .ZN(n3013) );
  OAI211_X1 U953 ( .C1(n4029), .C2(n70), .A(n2363), .B(n2362), .ZN(n912) );
  AOI221_X1 U954 ( .B1(n355), .B2(n1874), .C1(n364), .C2(n2781), .A(n912), 
        .ZN(n915) );
  NOR2_X1 U955 ( .A1(n4094), .A2(n73), .ZN(n913) );
  NOR4_X1 U956 ( .A1(n2379), .A2(n2375), .A3(n2357), .A4(n913), .ZN(n914) );
  NAND2_X1 U957 ( .A1(n915), .A2(n914), .ZN(n919) );
  OAI22_X1 U958 ( .A1(n1437), .A2(n79), .B1(n1435), .B2(n76), .ZN(n918) );
  AOI221_X1 U959 ( .B1(n87), .B2(n919), .C1(n82), .C2(n1550), .A(n918), .ZN(
        n932) );
  OAI22_X1 U960 ( .A1(n2749), .A2(n94), .B1(n2717), .B2(n91), .ZN(n923) );
  AOI221_X1 U961 ( .B1(n100), .B2(n1518), .C1(n97), .C2(n2845), .A(n923), .ZN(
        n931) );
  OAI22_X1 U962 ( .A1(n3677), .A2(n106), .B1(n2973), .B2(n103), .ZN(n926) );
  AOI221_X1 U963 ( .B1(n112), .B2(n2813), .C1(n109), .C2(n3613), .A(n926), 
        .ZN(n930) );
  OAI22_X1 U964 ( .A1(n2653), .A2(n117), .B1(n402), .B2(n115), .ZN(n928) );
  AOI221_X1 U965 ( .B1(n124), .B2(n3645), .C1(n121), .C2(n1648), .A(n928), 
        .ZN(n929) );
  NAND4_X1 U966 ( .A1(n932), .A2(n931), .A3(n930), .A4(n929), .ZN(n3014) );
  NAND3_X1 U967 ( .A1(n2342), .A2(n2341), .A3(n67), .ZN(n933) );
  NAND2_X1 U968 ( .A1(n173), .A2(n933), .ZN(n944) );
  INV_X1 U969 ( .A(n944), .ZN(n1441) );
  OAI211_X1 U970 ( .C1(n3998), .C2(n125), .A(n1927), .B(n1926), .ZN(n934) );
  AOI221_X1 U971 ( .B1(n305), .B2(n1843), .C1(n2750), .C2(n314), .A(n934), 
        .ZN(n937) );
  NOR2_X1 U972 ( .A1(n4125), .A2(n128), .ZN(n935) );
  NOR4_X1 U973 ( .A1(n1945), .A2(n1939), .A3(n1920), .A4(n935), .ZN(n936) );
  NAND2_X1 U974 ( .A1(n937), .A2(n936), .ZN(n941) );
  OR2_X1 U975 ( .A1(n1910), .A2(n944), .ZN(n1438) );
  NAND2_X1 U976 ( .A1(n1911), .A2(n142), .ZN(n1436) );
  OAI22_X1 U977 ( .A1(n134), .A2(n939), .B1(n131), .B2(n938), .ZN(n940) );
  AOI221_X1 U978 ( .B1(n142), .B2(n941), .C1(n137), .C2(n1519), .A(n940), .ZN(
        n949) );
  OR2_X1 U979 ( .A1(n1914), .A2(n944), .ZN(n1443) );
  NAND2_X1 U980 ( .A1(n1915), .A2(n142), .ZN(n1442) );
  OAI22_X1 U981 ( .A1(n2718), .A2(n149), .B1(n2686), .B2(n146), .ZN(n942) );
  AOI221_X1 U982 ( .B1(n155), .B2(n1487), .C1(n2814), .C2(n152), .A(n942), 
        .ZN(n948) );
  NAND2_X1 U983 ( .A1(n1925), .A2(n142), .ZN(n1446) );
  NAND2_X1 U984 ( .A1(n1918), .A2(n142), .ZN(n1445) );
  OAI22_X1 U985 ( .A1(n3646), .A2(n161), .B1(n2942), .B2(n158), .ZN(n943) );
  AOI221_X1 U986 ( .B1(n2782), .B2(n167), .C1(n3582), .C2(n164), .A(n943), 
        .ZN(n947) );
  NAND4_X1 U987 ( .A1(n67), .A2(n2341), .A3(n173), .A4(n2342), .ZN(n1448) );
  OAI22_X1 U988 ( .A1(n2685), .A2(n173), .B1(n170), .B2(n371), .ZN(n945) );
  AOI221_X1 U989 ( .B1(n3614), .B2(n179), .C1(n176), .C2(n1617), .A(n945), 
        .ZN(n946) );
  NAND4_X1 U990 ( .A1(n949), .A2(n948), .A3(n947), .A4(n946), .ZN(n3046) );
  MUX2_X1 U991 ( .A(n950), .B(DATAIN[0]), .S(n182), .Z(n4574) );
  OAI211_X1 U992 ( .C1(n3999), .C2(n125), .A(n1953), .B(n1952), .ZN(n951) );
  AOI221_X1 U993 ( .B1(n305), .B2(n1844), .C1(n2751), .C2(n314), .A(n951), 
        .ZN(n954) );
  NOR2_X1 U994 ( .A1(n4124), .A2(n128), .ZN(n952) );
  NOR4_X1 U995 ( .A1(n1959), .A2(n1956), .A3(n1950), .A4(n952), .ZN(n953) );
  NAND2_X1 U996 ( .A1(n954), .A2(n953), .ZN(n958) );
  OAI22_X1 U997 ( .A1(n134), .A2(n956), .B1(n131), .B2(n955), .ZN(n957) );
  AOI221_X1 U998 ( .B1(n145), .B2(n958), .C1(n137), .C2(n1520), .A(n957), .ZN(
        n965) );
  OAI22_X1 U999 ( .A1(n2719), .A2(n149), .B1(n2687), .B2(n146), .ZN(n959) );
  AOI221_X1 U1000 ( .B1(n155), .B2(n1488), .C1(n2815), .C2(n152), .A(n959), 
        .ZN(n964) );
  OAI22_X1 U1001 ( .A1(n3647), .A2(n161), .B1(n2943), .B2(n158), .ZN(n960) );
  AOI221_X1 U1002 ( .B1(n2783), .B2(n167), .C1(n3583), .C2(n164), .A(n960), 
        .ZN(n963) );
  OAI22_X1 U1003 ( .A1(n2684), .A2(n175), .B1(n170), .B2(n372), .ZN(n961) );
  AOI221_X1 U1004 ( .B1(n3615), .B2(n179), .C1(n176), .C2(n1618), .A(n961), 
        .ZN(n962) );
  NAND4_X1 U1005 ( .A1(n965), .A2(n964), .A3(n963), .A4(n962), .ZN(n3045) );
  MUX2_X1 U1006 ( .A(n966), .B(DATAIN[1]), .S(n182), .Z(n4575) );
  OAI211_X1 U1007 ( .C1(n4000), .C2(n125), .A(n1965), .B(n1964), .ZN(n967) );
  AOI221_X1 U1008 ( .B1(n305), .B2(n1845), .C1(n2752), .C2(n314), .A(n967), 
        .ZN(n970) );
  NOR2_X1 U1009 ( .A1(n4123), .A2(n128), .ZN(n968) );
  NOR4_X1 U1010 ( .A1(n1971), .A2(n1968), .A3(n1962), .A4(n968), .ZN(n969) );
  NAND2_X1 U1011 ( .A1(n970), .A2(n969), .ZN(n974) );
  OAI22_X1 U1012 ( .A1(n134), .A2(n972), .B1(n131), .B2(n971), .ZN(n973) );
  AOI221_X1 U1013 ( .B1(n145), .B2(n974), .C1(n137), .C2(n1521), .A(n973), 
        .ZN(n981) );
  OAI22_X1 U1014 ( .A1(n2720), .A2(n149), .B1(n2688), .B2(n146), .ZN(n975) );
  AOI221_X1 U1015 ( .B1(n155), .B2(n1489), .C1(n2816), .C2(n152), .A(n975), 
        .ZN(n980) );
  OAI22_X1 U1016 ( .A1(n3648), .A2(n161), .B1(n2944), .B2(n158), .ZN(n976) );
  AOI221_X1 U1017 ( .B1(n2784), .B2(n167), .C1(n3584), .C2(n164), .A(n976), 
        .ZN(n979) );
  OAI22_X1 U1018 ( .A1(n2683), .A2(n175), .B1(n170), .B2(n373), .ZN(n977) );
  AOI221_X1 U1019 ( .B1(n3616), .B2(n179), .C1(n176), .C2(n1619), .A(n977), 
        .ZN(n978) );
  NAND4_X1 U1020 ( .A1(n981), .A2(n980), .A3(n979), .A4(n978), .ZN(n3044) );
  MUX2_X1 U1021 ( .A(n982), .B(DATAIN[2]), .S(n182), .Z(n4576) );
  OAI211_X1 U1022 ( .C1(n4001), .C2(n125), .A(n1977), .B(n1976), .ZN(n983) );
  AOI221_X1 U1023 ( .B1(n305), .B2(n1846), .C1(n2753), .C2(n314), .A(n983), 
        .ZN(n986) );
  NOR2_X1 U1024 ( .A1(n4122), .A2(n128), .ZN(n984) );
  NOR4_X1 U1025 ( .A1(n1983), .A2(n1980), .A3(n1974), .A4(n984), .ZN(n985) );
  NAND2_X1 U1026 ( .A1(n986), .A2(n985), .ZN(n990) );
  OAI22_X1 U1027 ( .A1(n134), .A2(n988), .B1(n131), .B2(n987), .ZN(n989) );
  AOI221_X1 U1028 ( .B1(n145), .B2(n990), .C1(n137), .C2(n1522), .A(n989), 
        .ZN(n997) );
  OAI22_X1 U1029 ( .A1(n2721), .A2(n149), .B1(n2689), .B2(n146), .ZN(n991) );
  AOI221_X1 U1030 ( .B1(n155), .B2(n1490), .C1(n2817), .C2(n152), .A(n991), 
        .ZN(n996) );
  OAI22_X1 U1031 ( .A1(n3649), .A2(n161), .B1(n2945), .B2(n158), .ZN(n992) );
  AOI221_X1 U1032 ( .B1(n2785), .B2(n167), .C1(n3585), .C2(n164), .A(n992), 
        .ZN(n995) );
  OAI22_X1 U1033 ( .A1(n2682), .A2(n175), .B1(n170), .B2(n374), .ZN(n993) );
  AOI221_X1 U1034 ( .B1(n3617), .B2(n179), .C1(n176), .C2(n1620), .A(n993), 
        .ZN(n994) );
  NAND4_X1 U1035 ( .A1(n997), .A2(n996), .A3(n995), .A4(n994), .ZN(n3043) );
  MUX2_X1 U1036 ( .A(n998), .B(DATAIN[3]), .S(n182), .Z(n4577) );
  OAI211_X1 U1037 ( .C1(n4002), .C2(n125), .A(n1989), .B(n1988), .ZN(n999) );
  AOI221_X1 U1038 ( .B1(n305), .B2(n1847), .C1(n2754), .C2(n314), .A(n999), 
        .ZN(n1002) );
  NOR2_X1 U1039 ( .A1(n4121), .A2(n128), .ZN(n1000) );
  NOR4_X1 U1040 ( .A1(n1995), .A2(n1992), .A3(n1986), .A4(n1000), .ZN(n1001)
         );
  NAND2_X1 U1041 ( .A1(n1002), .A2(n1001), .ZN(n1006) );
  OAI22_X1 U1042 ( .A1(n134), .A2(n1004), .B1(n131), .B2(n1003), .ZN(n1005) );
  AOI221_X1 U1043 ( .B1(n145), .B2(n1006), .C1(n137), .C2(n1523), .A(n1005), 
        .ZN(n1013) );
  OAI22_X1 U1044 ( .A1(n2722), .A2(n149), .B1(n2690), .B2(n146), .ZN(n1007) );
  AOI221_X1 U1045 ( .B1(n155), .B2(n1491), .C1(n2818), .C2(n152), .A(n1007), 
        .ZN(n1012) );
  OAI22_X1 U1046 ( .A1(n3650), .A2(n161), .B1(n2946), .B2(n158), .ZN(n1008) );
  AOI221_X1 U1047 ( .B1(n2786), .B2(n167), .C1(n3586), .C2(n164), .A(n1008), 
        .ZN(n1011) );
  OAI22_X1 U1048 ( .A1(n2681), .A2(n175), .B1(n170), .B2(n375), .ZN(n1009) );
  AOI221_X1 U1049 ( .B1(n3618), .B2(n179), .C1(n176), .C2(n1621), .A(n1009), 
        .ZN(n1010) );
  NAND4_X1 U1050 ( .A1(n1013), .A2(n1012), .A3(n1011), .A4(n1010), .ZN(n3042)
         );
  MUX2_X1 U1051 ( .A(n1014), .B(DATAIN[4]), .S(n182), .Z(n4578) );
  OAI211_X1 U1052 ( .C1(n4003), .C2(n125), .A(n2001), .B(n2000), .ZN(n1015) );
  AOI221_X1 U1053 ( .B1(n305), .B2(n1848), .C1(n2755), .C2(n314), .A(n1015), 
        .ZN(n1018) );
  NOR2_X1 U1054 ( .A1(n4120), .A2(n128), .ZN(n1016) );
  NOR4_X1 U1055 ( .A1(n2007), .A2(n2004), .A3(n1998), .A4(n1016), .ZN(n1017)
         );
  NAND2_X1 U1056 ( .A1(n1018), .A2(n1017), .ZN(n1022) );
  OAI22_X1 U1057 ( .A1(n134), .A2(n1020), .B1(n131), .B2(n1019), .ZN(n1021) );
  AOI221_X1 U1058 ( .B1(n144), .B2(n1022), .C1(n137), .C2(n1524), .A(n1021), 
        .ZN(n1029) );
  OAI22_X1 U1059 ( .A1(n2723), .A2(n149), .B1(n2691), .B2(n146), .ZN(n1023) );
  AOI221_X1 U1060 ( .B1(n155), .B2(n1492), .C1(n2819), .C2(n152), .A(n1023), 
        .ZN(n1028) );
  OAI22_X1 U1061 ( .A1(n3651), .A2(n161), .B1(n2947), .B2(n158), .ZN(n1024) );
  AOI221_X1 U1062 ( .B1(n2787), .B2(n167), .C1(n3587), .C2(n164), .A(n1024), 
        .ZN(n1027) );
  OAI22_X1 U1063 ( .A1(n2680), .A2(n175), .B1(n170), .B2(n376), .ZN(n1025) );
  AOI221_X1 U1064 ( .B1(n3619), .B2(n179), .C1(n176), .C2(n1622), .A(n1025), 
        .ZN(n1026) );
  NAND4_X1 U1065 ( .A1(n1029), .A2(n1028), .A3(n1027), .A4(n1026), .ZN(n3041)
         );
  MUX2_X1 U1066 ( .A(n1030), .B(DATAIN[5]), .S(n182), .Z(n4579) );
  OAI211_X1 U1067 ( .C1(n4004), .C2(n125), .A(n2013), .B(n2012), .ZN(n1031) );
  AOI221_X1 U1068 ( .B1(n305), .B2(n1849), .C1(n2756), .C2(n314), .A(n1031), 
        .ZN(n1034) );
  NOR2_X1 U1069 ( .A1(n4119), .A2(n128), .ZN(n1032) );
  NOR4_X1 U1070 ( .A1(n2019), .A2(n2016), .A3(n2010), .A4(n1032), .ZN(n1033)
         );
  NAND2_X1 U1071 ( .A1(n1034), .A2(n1033), .ZN(n1038) );
  OAI22_X1 U1072 ( .A1(n134), .A2(n1036), .B1(n131), .B2(n1035), .ZN(n1037) );
  AOI221_X1 U1073 ( .B1(n144), .B2(n1038), .C1(n137), .C2(n1525), .A(n1037), 
        .ZN(n1045) );
  OAI22_X1 U1074 ( .A1(n2724), .A2(n149), .B1(n2692), .B2(n146), .ZN(n1039) );
  AOI221_X1 U1075 ( .B1(n155), .B2(n1493), .C1(n2820), .C2(n152), .A(n1039), 
        .ZN(n1044) );
  OAI22_X1 U1076 ( .A1(n3652), .A2(n161), .B1(n2948), .B2(n158), .ZN(n1040) );
  AOI221_X1 U1077 ( .B1(n2788), .B2(n167), .C1(n3588), .C2(n164), .A(n1040), 
        .ZN(n1043) );
  OAI22_X1 U1078 ( .A1(n2679), .A2(n175), .B1(n170), .B2(n377), .ZN(n1041) );
  AOI221_X1 U1079 ( .B1(n3620), .B2(n179), .C1(n176), .C2(n1623), .A(n1041), 
        .ZN(n1042) );
  NAND4_X1 U1080 ( .A1(n1045), .A2(n1044), .A3(n1043), .A4(n1042), .ZN(n3040)
         );
  MUX2_X1 U1081 ( .A(n1046), .B(DATAIN[6]), .S(n182), .Z(n4580) );
  OAI211_X1 U1082 ( .C1(n4005), .C2(n125), .A(n2025), .B(n2024), .ZN(n1047) );
  AOI221_X1 U1083 ( .B1(n305), .B2(n1850), .C1(n2757), .C2(n314), .A(n1047), 
        .ZN(n1050) );
  NOR2_X1 U1084 ( .A1(n4118), .A2(n128), .ZN(n1048) );
  NOR4_X1 U1085 ( .A1(n2031), .A2(n2028), .A3(n2022), .A4(n1048), .ZN(n1049)
         );
  NAND2_X1 U1086 ( .A1(n1050), .A2(n1049), .ZN(n1054) );
  OAI22_X1 U1087 ( .A1(n134), .A2(n1052), .B1(n131), .B2(n1051), .ZN(n1053) );
  AOI221_X1 U1088 ( .B1(n144), .B2(n1054), .C1(n137), .C2(n1526), .A(n1053), 
        .ZN(n1061) );
  OAI22_X1 U1089 ( .A1(n2725), .A2(n149), .B1(n2693), .B2(n146), .ZN(n1055) );
  AOI221_X1 U1090 ( .B1(n155), .B2(n1494), .C1(n2821), .C2(n152), .A(n1055), 
        .ZN(n1060) );
  OAI22_X1 U1091 ( .A1(n3653), .A2(n161), .B1(n2949), .B2(n158), .ZN(n1056) );
  AOI221_X1 U1092 ( .B1(n2789), .B2(n167), .C1(n3589), .C2(n164), .A(n1056), 
        .ZN(n1059) );
  OAI22_X1 U1093 ( .A1(n2678), .A2(n175), .B1(n170), .B2(n378), .ZN(n1057) );
  AOI221_X1 U1094 ( .B1(n3621), .B2(n179), .C1(n176), .C2(n1624), .A(n1057), 
        .ZN(n1058) );
  NAND4_X1 U1095 ( .A1(n1061), .A2(n1060), .A3(n1059), .A4(n1058), .ZN(n3039)
         );
  MUX2_X1 U1096 ( .A(n1062), .B(DATAIN[7]), .S(n182), .Z(n4581) );
  OAI211_X1 U1097 ( .C1(n4006), .C2(n125), .A(n2037), .B(n2036), .ZN(n1063) );
  AOI221_X1 U1098 ( .B1(n305), .B2(n1851), .C1(n2758), .C2(n314), .A(n1063), 
        .ZN(n1066) );
  NOR2_X1 U1099 ( .A1(n4117), .A2(n128), .ZN(n1064) );
  NOR4_X1 U1100 ( .A1(n2043), .A2(n2040), .A3(n2034), .A4(n1064), .ZN(n1065)
         );
  NAND2_X1 U1101 ( .A1(n1066), .A2(n1065), .ZN(n1070) );
  OAI22_X1 U1102 ( .A1(n134), .A2(n1068), .B1(n131), .B2(n1067), .ZN(n1069) );
  AOI221_X1 U1103 ( .B1(n144), .B2(n1070), .C1(n137), .C2(n1527), .A(n1069), 
        .ZN(n1077) );
  OAI22_X1 U1104 ( .A1(n2726), .A2(n149), .B1(n2694), .B2(n146), .ZN(n1071) );
  AOI221_X1 U1105 ( .B1(n155), .B2(n1495), .C1(n2822), .C2(n152), .A(n1071), 
        .ZN(n1076) );
  OAI22_X1 U1106 ( .A1(n3654), .A2(n161), .B1(n2950), .B2(n158), .ZN(n1072) );
  AOI221_X1 U1107 ( .B1(n2790), .B2(n167), .C1(n3590), .C2(n164), .A(n1072), 
        .ZN(n1075) );
  OAI22_X1 U1108 ( .A1(n2677), .A2(n175), .B1(n170), .B2(n379), .ZN(n1073) );
  AOI221_X1 U1109 ( .B1(n3622), .B2(n179), .C1(n176), .C2(n1625), .A(n1073), 
        .ZN(n1074) );
  NAND4_X1 U1110 ( .A1(n1077), .A2(n1076), .A3(n1075), .A4(n1074), .ZN(n3038)
         );
  MUX2_X1 U1111 ( .A(n1078), .B(DATAIN[8]), .S(n182), .Z(n4582) );
  OAI211_X1 U1112 ( .C1(n4007), .C2(n125), .A(n2049), .B(n2048), .ZN(n1079) );
  AOI221_X1 U1113 ( .B1(n305), .B2(n1852), .C1(n2759), .C2(n314), .A(n1079), 
        .ZN(n1082) );
  NOR2_X1 U1114 ( .A1(n4116), .A2(n128), .ZN(n1080) );
  NOR4_X1 U1115 ( .A1(n2055), .A2(n2052), .A3(n2046), .A4(n1080), .ZN(n1081)
         );
  NAND2_X1 U1116 ( .A1(n1082), .A2(n1081), .ZN(n1086) );
  OAI22_X1 U1117 ( .A1(n134), .A2(n1084), .B1(n131), .B2(n1083), .ZN(n1085) );
  AOI221_X1 U1118 ( .B1(n144), .B2(n1086), .C1(n137), .C2(n1528), .A(n1085), 
        .ZN(n1093) );
  OAI22_X1 U1119 ( .A1(n2727), .A2(n149), .B1(n2695), .B2(n146), .ZN(n1087) );
  AOI221_X1 U1120 ( .B1(n155), .B2(n1496), .C1(n2823), .C2(n152), .A(n1087), 
        .ZN(n1092) );
  OAI22_X1 U1121 ( .A1(n3655), .A2(n161), .B1(n2951), .B2(n158), .ZN(n1088) );
  AOI221_X1 U1122 ( .B1(n2791), .B2(n167), .C1(n3591), .C2(n164), .A(n1088), 
        .ZN(n1091) );
  OAI22_X1 U1123 ( .A1(n2676), .A2(n175), .B1(n170), .B2(n380), .ZN(n1089) );
  AOI221_X1 U1124 ( .B1(n3623), .B2(n179), .C1(n176), .C2(n1626), .A(n1089), 
        .ZN(n1090) );
  NAND4_X1 U1125 ( .A1(n1093), .A2(n1092), .A3(n1091), .A4(n1090), .ZN(n3037)
         );
  MUX2_X1 U1126 ( .A(n1094), .B(DATAIN[9]), .S(n182), .Z(n4583) );
  OAI211_X1 U1127 ( .C1(n4008), .C2(n125), .A(n2061), .B(n2060), .ZN(n1095) );
  AOI221_X1 U1128 ( .B1(n305), .B2(n1853), .C1(n2760), .C2(n314), .A(n1095), 
        .ZN(n1098) );
  NOR2_X1 U1129 ( .A1(n4115), .A2(n128), .ZN(n1096) );
  NOR4_X1 U1130 ( .A1(n2067), .A2(n2064), .A3(n2058), .A4(n1096), .ZN(n1097)
         );
  NAND2_X1 U1131 ( .A1(n1098), .A2(n1097), .ZN(n1102) );
  OAI22_X1 U1132 ( .A1(n134), .A2(n1100), .B1(n131), .B2(n1099), .ZN(n1101) );
  AOI221_X1 U1133 ( .B1(n144), .B2(n1102), .C1(n137), .C2(n1529), .A(n1101), 
        .ZN(n1109) );
  OAI22_X1 U1134 ( .A1(n2728), .A2(n149), .B1(n2696), .B2(n146), .ZN(n1103) );
  AOI221_X1 U1135 ( .B1(n155), .B2(n1497), .C1(n2824), .C2(n152), .A(n1103), 
        .ZN(n1108) );
  OAI22_X1 U1136 ( .A1(n3656), .A2(n161), .B1(n2952), .B2(n158), .ZN(n1104) );
  AOI221_X1 U1137 ( .B1(n2792), .B2(n167), .C1(n3592), .C2(n164), .A(n1104), 
        .ZN(n1107) );
  OAI22_X1 U1138 ( .A1(n2675), .A2(n175), .B1(n170), .B2(n381), .ZN(n1105) );
  AOI221_X1 U1139 ( .B1(n3624), .B2(n179), .C1(n176), .C2(n1627), .A(n1105), 
        .ZN(n1106) );
  NAND4_X1 U1140 ( .A1(n1109), .A2(n1108), .A3(n1107), .A4(n1106), .ZN(n3036)
         );
  MUX2_X1 U1141 ( .A(n1110), .B(DATAIN[10]), .S(n182), .Z(n4584) );
  OAI211_X1 U1142 ( .C1(n4009), .C2(n125), .A(n2073), .B(n2072), .ZN(n1111) );
  AOI221_X1 U1143 ( .B1(n305), .B2(n1854), .C1(n2761), .C2(n314), .A(n1111), 
        .ZN(n1114) );
  NOR2_X1 U1144 ( .A1(n4114), .A2(n128), .ZN(n1112) );
  NOR4_X1 U1145 ( .A1(n2079), .A2(n2076), .A3(n2070), .A4(n1112), .ZN(n1113)
         );
  NAND2_X1 U1146 ( .A1(n1114), .A2(n1113), .ZN(n1118) );
  OAI22_X1 U1147 ( .A1(n134), .A2(n1116), .B1(n131), .B2(n1115), .ZN(n1117) );
  AOI221_X1 U1148 ( .B1(n144), .B2(n1118), .C1(n137), .C2(n1530), .A(n1117), 
        .ZN(n1125) );
  OAI22_X1 U1149 ( .A1(n2729), .A2(n149), .B1(n2697), .B2(n146), .ZN(n1119) );
  AOI221_X1 U1150 ( .B1(n155), .B2(n1498), .C1(n2825), .C2(n152), .A(n1119), 
        .ZN(n1124) );
  OAI22_X1 U1151 ( .A1(n3657), .A2(n161), .B1(n2953), .B2(n158), .ZN(n1120) );
  AOI221_X1 U1152 ( .B1(n2793), .B2(n167), .C1(n3593), .C2(n164), .A(n1120), 
        .ZN(n1123) );
  OAI22_X1 U1153 ( .A1(n2674), .A2(n174), .B1(n170), .B2(n382), .ZN(n1121) );
  AOI221_X1 U1154 ( .B1(n3625), .B2(n179), .C1(n176), .C2(n1628), .A(n1121), 
        .ZN(n1122) );
  NAND4_X1 U1155 ( .A1(n1125), .A2(n1124), .A3(n1123), .A4(n1122), .ZN(n3035)
         );
  MUX2_X1 U1156 ( .A(n1126), .B(DATAIN[11]), .S(n182), .Z(n4585) );
  OAI211_X1 U1157 ( .C1(n4010), .C2(n126), .A(n2085), .B(n2084), .ZN(n1127) );
  AOI221_X1 U1158 ( .B1(n306), .B2(n1855), .C1(n2762), .C2(n315), .A(n1127), 
        .ZN(n1130) );
  NOR2_X1 U1159 ( .A1(n4113), .A2(n129), .ZN(n1128) );
  NOR4_X1 U1160 ( .A1(n2091), .A2(n2088), .A3(n2082), .A4(n1128), .ZN(n1129)
         );
  NAND2_X1 U1161 ( .A1(n1130), .A2(n1129), .ZN(n1134) );
  OAI22_X1 U1162 ( .A1(n135), .A2(n1132), .B1(n132), .B2(n1131), .ZN(n1133) );
  AOI221_X1 U1163 ( .B1(n144), .B2(n1134), .C1(n138), .C2(n1531), .A(n1133), 
        .ZN(n1141) );
  OAI22_X1 U1164 ( .A1(n2730), .A2(n150), .B1(n2698), .B2(n147), .ZN(n1135) );
  AOI221_X1 U1165 ( .B1(n156), .B2(n1499), .C1(n2826), .C2(n153), .A(n1135), 
        .ZN(n1140) );
  OAI22_X1 U1166 ( .A1(n3658), .A2(n162), .B1(n2954), .B2(n159), .ZN(n1136) );
  AOI221_X1 U1167 ( .B1(n2794), .B2(n168), .C1(n3594), .C2(n165), .A(n1136), 
        .ZN(n1139) );
  OAI22_X1 U1168 ( .A1(n2673), .A2(n174), .B1(n171), .B2(n383), .ZN(n1137) );
  AOI221_X1 U1169 ( .B1(n3626), .B2(n180), .C1(n177), .C2(n1629), .A(n1137), 
        .ZN(n1138) );
  NAND4_X1 U1170 ( .A1(n1141), .A2(n1140), .A3(n1139), .A4(n1138), .ZN(n3034)
         );
  MUX2_X1 U1171 ( .A(n1142), .B(DATAIN[12]), .S(n183), .Z(n4586) );
  OAI211_X1 U1172 ( .C1(n4011), .C2(n126), .A(n2097), .B(n2096), .ZN(n1143) );
  AOI221_X1 U1173 ( .B1(n306), .B2(n1856), .C1(n2763), .C2(n315), .A(n1143), 
        .ZN(n1146) );
  NOR2_X1 U1174 ( .A1(n4112), .A2(n129), .ZN(n1144) );
  NOR4_X1 U1175 ( .A1(n2103), .A2(n2100), .A3(n2094), .A4(n1144), .ZN(n1145)
         );
  NAND2_X1 U1176 ( .A1(n1146), .A2(n1145), .ZN(n1150) );
  OAI22_X1 U1177 ( .A1(n135), .A2(n1148), .B1(n132), .B2(n1147), .ZN(n1149) );
  AOI221_X1 U1178 ( .B1(n144), .B2(n1150), .C1(n138), .C2(n1532), .A(n1149), 
        .ZN(n1157) );
  OAI22_X1 U1179 ( .A1(n2731), .A2(n150), .B1(n2699), .B2(n147), .ZN(n1151) );
  AOI221_X1 U1180 ( .B1(n156), .B2(n1500), .C1(n2827), .C2(n153), .A(n1151), 
        .ZN(n1156) );
  OAI22_X1 U1181 ( .A1(n3659), .A2(n162), .B1(n2955), .B2(n159), .ZN(n1152) );
  AOI221_X1 U1182 ( .B1(n2795), .B2(n168), .C1(n3595), .C2(n165), .A(n1152), 
        .ZN(n1155) );
  OAI22_X1 U1183 ( .A1(n2672), .A2(n174), .B1(n171), .B2(n384), .ZN(n1153) );
  AOI221_X1 U1184 ( .B1(n3627), .B2(n180), .C1(n177), .C2(n1630), .A(n1153), 
        .ZN(n1154) );
  NAND4_X1 U1185 ( .A1(n1157), .A2(n1156), .A3(n1155), .A4(n1154), .ZN(n3033)
         );
  MUX2_X1 U1186 ( .A(n1158), .B(DATAIN[13]), .S(n183), .Z(n4587) );
  OAI211_X1 U1187 ( .C1(n4012), .C2(n126), .A(n2109), .B(n2108), .ZN(n1159) );
  AOI221_X1 U1188 ( .B1(n306), .B2(n1857), .C1(n2764), .C2(n315), .A(n1159), 
        .ZN(n1162) );
  NOR2_X1 U1189 ( .A1(n4111), .A2(n129), .ZN(n1160) );
  NOR4_X1 U1190 ( .A1(n2115), .A2(n2112), .A3(n2106), .A4(n1160), .ZN(n1161)
         );
  NAND2_X1 U1191 ( .A1(n1162), .A2(n1161), .ZN(n1166) );
  OAI22_X1 U1192 ( .A1(n135), .A2(n1164), .B1(n132), .B2(n1163), .ZN(n1165) );
  AOI221_X1 U1193 ( .B1(n144), .B2(n1166), .C1(n138), .C2(n1533), .A(n1165), 
        .ZN(n1173) );
  OAI22_X1 U1194 ( .A1(n2732), .A2(n150), .B1(n2700), .B2(n147), .ZN(n1167) );
  AOI221_X1 U1195 ( .B1(n156), .B2(n1501), .C1(n2828), .C2(n153), .A(n1167), 
        .ZN(n1172) );
  OAI22_X1 U1196 ( .A1(n3660), .A2(n162), .B1(n2956), .B2(n159), .ZN(n1168) );
  AOI221_X1 U1197 ( .B1(n2796), .B2(n168), .C1(n3596), .C2(n165), .A(n1168), 
        .ZN(n1171) );
  OAI22_X1 U1198 ( .A1(n2671), .A2(n174), .B1(n171), .B2(n385), .ZN(n1169) );
  AOI221_X1 U1199 ( .B1(n3628), .B2(n180), .C1(n177), .C2(n1631), .A(n1169), 
        .ZN(n1170) );
  NAND4_X1 U1200 ( .A1(n1173), .A2(n1172), .A3(n1171), .A4(n1170), .ZN(n3032)
         );
  MUX2_X1 U1201 ( .A(n1174), .B(DATAIN[14]), .S(n183), .Z(n4588) );
  OAI211_X1 U1202 ( .C1(n4013), .C2(n126), .A(n2121), .B(n2120), .ZN(n1175) );
  AOI221_X1 U1203 ( .B1(n306), .B2(n1858), .C1(n2765), .C2(n315), .A(n1175), 
        .ZN(n1178) );
  NOR2_X1 U1204 ( .A1(n4110), .A2(n129), .ZN(n1176) );
  NOR4_X1 U1205 ( .A1(n2127), .A2(n2124), .A3(n2118), .A4(n1176), .ZN(n1177)
         );
  NAND2_X1 U1206 ( .A1(n1178), .A2(n1177), .ZN(n1182) );
  OAI22_X1 U1207 ( .A1(n135), .A2(n1180), .B1(n132), .B2(n1179), .ZN(n1181) );
  AOI221_X1 U1208 ( .B1(n144), .B2(n1182), .C1(n138), .C2(n1534), .A(n1181), 
        .ZN(n1189) );
  OAI22_X1 U1209 ( .A1(n2733), .A2(n150), .B1(n2701), .B2(n147), .ZN(n1183) );
  AOI221_X1 U1210 ( .B1(n156), .B2(n1502), .C1(n2829), .C2(n153), .A(n1183), 
        .ZN(n1188) );
  OAI22_X1 U1211 ( .A1(n3661), .A2(n162), .B1(n2957), .B2(n159), .ZN(n1184) );
  AOI221_X1 U1212 ( .B1(n2797), .B2(n168), .C1(n3597), .C2(n165), .A(n1184), 
        .ZN(n1187) );
  OAI22_X1 U1213 ( .A1(n2670), .A2(n174), .B1(n171), .B2(n386), .ZN(n1185) );
  AOI221_X1 U1214 ( .B1(n3629), .B2(n180), .C1(n177), .C2(n1632), .A(n1185), 
        .ZN(n1186) );
  NAND4_X1 U1215 ( .A1(n1189), .A2(n1188), .A3(n1187), .A4(n1186), .ZN(n3031)
         );
  MUX2_X1 U1216 ( .A(n1190), .B(DATAIN[15]), .S(n183), .Z(n4589) );
  OAI211_X1 U1217 ( .C1(n4014), .C2(n126), .A(n2133), .B(n2132), .ZN(n1191) );
  AOI221_X1 U1218 ( .B1(n306), .B2(n1859), .C1(n2766), .C2(n315), .A(n1191), 
        .ZN(n1194) );
  NOR2_X1 U1219 ( .A1(n4109), .A2(n129), .ZN(n1192) );
  NOR4_X1 U1220 ( .A1(n2139), .A2(n2136), .A3(n2130), .A4(n1192), .ZN(n1193)
         );
  NAND2_X1 U1221 ( .A1(n1194), .A2(n1193), .ZN(n1198) );
  OAI22_X1 U1222 ( .A1(n135), .A2(n1196), .B1(n132), .B2(n1195), .ZN(n1197) );
  AOI221_X1 U1223 ( .B1(n143), .B2(n1198), .C1(n138), .C2(n1535), .A(n1197), 
        .ZN(n1205) );
  OAI22_X1 U1224 ( .A1(n2734), .A2(n150), .B1(n2702), .B2(n147), .ZN(n1199) );
  AOI221_X1 U1225 ( .B1(n156), .B2(n1503), .C1(n2830), .C2(n153), .A(n1199), 
        .ZN(n1204) );
  OAI22_X1 U1226 ( .A1(n3662), .A2(n162), .B1(n2958), .B2(n159), .ZN(n1200) );
  AOI221_X1 U1227 ( .B1(n2798), .B2(n168), .C1(n3598), .C2(n165), .A(n1200), 
        .ZN(n1203) );
  OAI22_X1 U1228 ( .A1(n2669), .A2(n174), .B1(n171), .B2(n387), .ZN(n1201) );
  AOI221_X1 U1229 ( .B1(n3630), .B2(n180), .C1(n177), .C2(n1633), .A(n1201), 
        .ZN(n1202) );
  NAND4_X1 U1230 ( .A1(n1205), .A2(n1204), .A3(n1203), .A4(n1202), .ZN(n3030)
         );
  MUX2_X1 U1231 ( .A(n1206), .B(DATAIN[16]), .S(n183), .Z(n4590) );
  OAI211_X1 U1232 ( .C1(n4015), .C2(n126), .A(n2145), .B(n2144), .ZN(n1207) );
  AOI221_X1 U1233 ( .B1(n306), .B2(n1860), .C1(n2767), .C2(n315), .A(n1207), 
        .ZN(n1210) );
  NOR2_X1 U1234 ( .A1(n4108), .A2(n129), .ZN(n1208) );
  NOR4_X1 U1235 ( .A1(n2151), .A2(n2148), .A3(n2142), .A4(n1208), .ZN(n1209)
         );
  NAND2_X1 U1236 ( .A1(n1210), .A2(n1209), .ZN(n1214) );
  OAI22_X1 U1237 ( .A1(n135), .A2(n1212), .B1(n132), .B2(n1211), .ZN(n1213) );
  AOI221_X1 U1238 ( .B1(n143), .B2(n1214), .C1(n138), .C2(n1536), .A(n1213), 
        .ZN(n1221) );
  OAI22_X1 U1239 ( .A1(n2735), .A2(n150), .B1(n2703), .B2(n147), .ZN(n1215) );
  AOI221_X1 U1240 ( .B1(n156), .B2(n1504), .C1(n2831), .C2(n153), .A(n1215), 
        .ZN(n1220) );
  OAI22_X1 U1241 ( .A1(n3663), .A2(n162), .B1(n2959), .B2(n159), .ZN(n1216) );
  AOI221_X1 U1242 ( .B1(n2799), .B2(n168), .C1(n3599), .C2(n165), .A(n1216), 
        .ZN(n1219) );
  OAI22_X1 U1243 ( .A1(n2668), .A2(n174), .B1(n171), .B2(n388), .ZN(n1217) );
  AOI221_X1 U1244 ( .B1(n3631), .B2(n180), .C1(n177), .C2(n1634), .A(n1217), 
        .ZN(n1218) );
  NAND4_X1 U1245 ( .A1(n1221), .A2(n1220), .A3(n1219), .A4(n1218), .ZN(n3029)
         );
  MUX2_X1 U1246 ( .A(n1222), .B(DATAIN[17]), .S(n183), .Z(n4591) );
  OAI211_X1 U1247 ( .C1(n4016), .C2(n126), .A(n2157), .B(n2156), .ZN(n1223) );
  AOI221_X1 U1248 ( .B1(n306), .B2(n1861), .C1(n2768), .C2(n315), .A(n1223), 
        .ZN(n1226) );
  NOR2_X1 U1249 ( .A1(n4107), .A2(n129), .ZN(n1224) );
  NOR4_X1 U1250 ( .A1(n2163), .A2(n2160), .A3(n2154), .A4(n1224), .ZN(n1225)
         );
  NAND2_X1 U1251 ( .A1(n1226), .A2(n1225), .ZN(n1230) );
  OAI22_X1 U1252 ( .A1(n135), .A2(n1228), .B1(n132), .B2(n1227), .ZN(n1229) );
  AOI221_X1 U1253 ( .B1(n143), .B2(n1230), .C1(n138), .C2(n1537), .A(n1229), 
        .ZN(n1237) );
  OAI22_X1 U1254 ( .A1(n2736), .A2(n150), .B1(n2704), .B2(n147), .ZN(n1231) );
  AOI221_X1 U1255 ( .B1(n156), .B2(n1505), .C1(n2832), .C2(n153), .A(n1231), 
        .ZN(n1236) );
  OAI22_X1 U1256 ( .A1(n3664), .A2(n162), .B1(n2960), .B2(n159), .ZN(n1232) );
  AOI221_X1 U1257 ( .B1(n2800), .B2(n168), .C1(n3600), .C2(n165), .A(n1232), 
        .ZN(n1235) );
  OAI22_X1 U1258 ( .A1(n2667), .A2(n174), .B1(n171), .B2(n389), .ZN(n1233) );
  AOI221_X1 U1259 ( .B1(n3632), .B2(n180), .C1(n177), .C2(n1635), .A(n1233), 
        .ZN(n1234) );
  NAND4_X1 U1260 ( .A1(n1237), .A2(n1236), .A3(n1235), .A4(n1234), .ZN(n3028)
         );
  MUX2_X1 U1261 ( .A(n1238), .B(DATAIN[18]), .S(n183), .Z(n4592) );
  OAI211_X1 U1262 ( .C1(n4017), .C2(n126), .A(n2169), .B(n2168), .ZN(n1239) );
  AOI221_X1 U1263 ( .B1(n306), .B2(n1862), .C1(n2769), .C2(n315), .A(n1239), 
        .ZN(n1242) );
  NOR2_X1 U1264 ( .A1(n4106), .A2(n129), .ZN(n1240) );
  NOR4_X1 U1265 ( .A1(n2175), .A2(n2172), .A3(n2166), .A4(n1240), .ZN(n1241)
         );
  NAND2_X1 U1266 ( .A1(n1242), .A2(n1241), .ZN(n1246) );
  OAI22_X1 U1267 ( .A1(n135), .A2(n1244), .B1(n132), .B2(n1243), .ZN(n1245) );
  AOI221_X1 U1268 ( .B1(n143), .B2(n1246), .C1(n138), .C2(n1538), .A(n1245), 
        .ZN(n1253) );
  OAI22_X1 U1269 ( .A1(n2737), .A2(n150), .B1(n2705), .B2(n147), .ZN(n1247) );
  AOI221_X1 U1270 ( .B1(n156), .B2(n1506), .C1(n2833), .C2(n153), .A(n1247), 
        .ZN(n1252) );
  OAI22_X1 U1271 ( .A1(n3665), .A2(n162), .B1(n2961), .B2(n159), .ZN(n1248) );
  AOI221_X1 U1272 ( .B1(n2801), .B2(n168), .C1(n3601), .C2(n165), .A(n1248), 
        .ZN(n1251) );
  OAI22_X1 U1273 ( .A1(n2666), .A2(n174), .B1(n171), .B2(n390), .ZN(n1249) );
  AOI221_X1 U1274 ( .B1(n3633), .B2(n180), .C1(n177), .C2(n1636), .A(n1249), 
        .ZN(n1250) );
  NAND4_X1 U1275 ( .A1(n1253), .A2(n1252), .A3(n1251), .A4(n1250), .ZN(n3027)
         );
  MUX2_X1 U1276 ( .A(n1254), .B(DATAIN[19]), .S(n183), .Z(n4593) );
  OAI211_X1 U1277 ( .C1(n4018), .C2(n126), .A(n2181), .B(n2180), .ZN(n1255) );
  AOI221_X1 U1278 ( .B1(n306), .B2(n1863), .C1(n2770), .C2(n315), .A(n1255), 
        .ZN(n1258) );
  NOR2_X1 U1279 ( .A1(n4105), .A2(n129), .ZN(n1256) );
  NOR4_X1 U1280 ( .A1(n2187), .A2(n2184), .A3(n2178), .A4(n1256), .ZN(n1257)
         );
  NAND2_X1 U1281 ( .A1(n1258), .A2(n1257), .ZN(n1262) );
  OAI22_X1 U1282 ( .A1(n135), .A2(n1260), .B1(n132), .B2(n1259), .ZN(n1261) );
  AOI221_X1 U1283 ( .B1(n143), .B2(n1262), .C1(n138), .C2(n1539), .A(n1261), 
        .ZN(n1269) );
  OAI22_X1 U1284 ( .A1(n2738), .A2(n150), .B1(n2706), .B2(n147), .ZN(n1263) );
  AOI221_X1 U1285 ( .B1(n156), .B2(n1507), .C1(n2834), .C2(n153), .A(n1263), 
        .ZN(n1268) );
  OAI22_X1 U1286 ( .A1(n3666), .A2(n162), .B1(n2962), .B2(n159), .ZN(n1264) );
  AOI221_X1 U1287 ( .B1(n2802), .B2(n168), .C1(n3602), .C2(n165), .A(n1264), 
        .ZN(n1267) );
  OAI22_X1 U1288 ( .A1(n2665), .A2(n174), .B1(n171), .B2(n391), .ZN(n1265) );
  AOI221_X1 U1289 ( .B1(n3634), .B2(n180), .C1(n177), .C2(n1637), .A(n1265), 
        .ZN(n1266) );
  NAND4_X1 U1290 ( .A1(n1269), .A2(n1268), .A3(n1267), .A4(n1266), .ZN(n3026)
         );
  MUX2_X1 U1291 ( .A(n1270), .B(DATAIN[20]), .S(n183), .Z(n4594) );
  OAI211_X1 U1292 ( .C1(n4019), .C2(n126), .A(n2193), .B(n2192), .ZN(n1271) );
  AOI221_X1 U1293 ( .B1(n306), .B2(n1864), .C1(n2771), .C2(n315), .A(n1271), 
        .ZN(n1274) );
  NOR2_X1 U1294 ( .A1(n4104), .A2(n129), .ZN(n1272) );
  NOR4_X1 U1295 ( .A1(n2199), .A2(n2196), .A3(n2190), .A4(n1272), .ZN(n1273)
         );
  NAND2_X1 U1296 ( .A1(n1274), .A2(n1273), .ZN(n1278) );
  OAI22_X1 U1297 ( .A1(n135), .A2(n1276), .B1(n132), .B2(n1275), .ZN(n1277) );
  AOI221_X1 U1298 ( .B1(n143), .B2(n1278), .C1(n138), .C2(n1540), .A(n1277), 
        .ZN(n1285) );
  OAI22_X1 U1299 ( .A1(n2739), .A2(n150), .B1(n2707), .B2(n147), .ZN(n1279) );
  AOI221_X1 U1300 ( .B1(n156), .B2(n1508), .C1(n2835), .C2(n153), .A(n1279), 
        .ZN(n1284) );
  OAI22_X1 U1301 ( .A1(n3667), .A2(n162), .B1(n2963), .B2(n159), .ZN(n1280) );
  AOI221_X1 U1302 ( .B1(n2803), .B2(n168), .C1(n3603), .C2(n165), .A(n1280), 
        .ZN(n1283) );
  OAI22_X1 U1303 ( .A1(n2664), .A2(n174), .B1(n171), .B2(n392), .ZN(n1281) );
  AOI221_X1 U1304 ( .B1(n3635), .B2(n180), .C1(n177), .C2(n1638), .A(n1281), 
        .ZN(n1282) );
  NAND4_X1 U1305 ( .A1(n1285), .A2(n1284), .A3(n1283), .A4(n1282), .ZN(n3025)
         );
  MUX2_X1 U1306 ( .A(n1286), .B(DATAIN[21]), .S(n183), .Z(n4595) );
  OAI211_X1 U1307 ( .C1(n4020), .C2(n126), .A(n2205), .B(n2204), .ZN(n1287) );
  AOI221_X1 U1308 ( .B1(n306), .B2(n1865), .C1(n2772), .C2(n315), .A(n1287), 
        .ZN(n1290) );
  NOR2_X1 U1309 ( .A1(n4103), .A2(n129), .ZN(n1288) );
  NOR4_X1 U1310 ( .A1(n2211), .A2(n2208), .A3(n2202), .A4(n1288), .ZN(n1289)
         );
  NAND2_X1 U1311 ( .A1(n1290), .A2(n1289), .ZN(n1294) );
  OAI22_X1 U1312 ( .A1(n135), .A2(n1292), .B1(n132), .B2(n1291), .ZN(n1293) );
  AOI221_X1 U1313 ( .B1(n143), .B2(n1294), .C1(n138), .C2(n1541), .A(n1293), 
        .ZN(n1301) );
  OAI22_X1 U1314 ( .A1(n2740), .A2(n150), .B1(n2708), .B2(n147), .ZN(n1295) );
  AOI221_X1 U1315 ( .B1(n156), .B2(n1509), .C1(n2836), .C2(n153), .A(n1295), 
        .ZN(n1300) );
  OAI22_X1 U1316 ( .A1(n3668), .A2(n162), .B1(n2964), .B2(n159), .ZN(n1296) );
  AOI221_X1 U1317 ( .B1(n2804), .B2(n168), .C1(n3604), .C2(n165), .A(n1296), 
        .ZN(n1299) );
  OAI22_X1 U1318 ( .A1(n2663), .A2(n173), .B1(n171), .B2(n393), .ZN(n1297) );
  AOI221_X1 U1319 ( .B1(n3636), .B2(n180), .C1(n177), .C2(n1639), .A(n1297), 
        .ZN(n1298) );
  NAND4_X1 U1320 ( .A1(n1301), .A2(n1300), .A3(n1299), .A4(n1298), .ZN(n3024)
         );
  MUX2_X1 U1321 ( .A(n1302), .B(DATAIN[22]), .S(n183), .Z(n4596) );
  OAI211_X1 U1322 ( .C1(n4021), .C2(n126), .A(n2217), .B(n2216), .ZN(n1303) );
  AOI221_X1 U1323 ( .B1(n306), .B2(n1866), .C1(n2773), .C2(n315), .A(n1303), 
        .ZN(n1306) );
  NOR2_X1 U1324 ( .A1(n4102), .A2(n129), .ZN(n1304) );
  NOR4_X1 U1325 ( .A1(n2223), .A2(n2220), .A3(n2214), .A4(n1304), .ZN(n1305)
         );
  NAND2_X1 U1326 ( .A1(n1306), .A2(n1305), .ZN(n1310) );
  OAI22_X1 U1327 ( .A1(n135), .A2(n1308), .B1(n132), .B2(n1307), .ZN(n1309) );
  AOI221_X1 U1328 ( .B1(n143), .B2(n1310), .C1(n138), .C2(n1542), .A(n1309), 
        .ZN(n1317) );
  OAI22_X1 U1329 ( .A1(n2741), .A2(n150), .B1(n2709), .B2(n147), .ZN(n1311) );
  AOI221_X1 U1330 ( .B1(n156), .B2(n1510), .C1(n2837), .C2(n153), .A(n1311), 
        .ZN(n1316) );
  OAI22_X1 U1331 ( .A1(n3669), .A2(n162), .B1(n2965), .B2(n159), .ZN(n1312) );
  AOI221_X1 U1332 ( .B1(n2805), .B2(n168), .C1(n3605), .C2(n165), .A(n1312), 
        .ZN(n1315) );
  OAI22_X1 U1333 ( .A1(n2662), .A2(n173), .B1(n171), .B2(n394), .ZN(n1313) );
  AOI221_X1 U1334 ( .B1(n3637), .B2(n180), .C1(n177), .C2(n1640), .A(n1313), 
        .ZN(n1314) );
  NAND4_X1 U1335 ( .A1(n1317), .A2(n1316), .A3(n1315), .A4(n1314), .ZN(n3023)
         );
  MUX2_X1 U1336 ( .A(n1318), .B(DATAIN[23]), .S(n183), .Z(n4597) );
  OAI211_X1 U1337 ( .C1(n4022), .C2(n127), .A(n2229), .B(n2228), .ZN(n1319) );
  AOI221_X1 U1338 ( .B1(n307), .B2(n1867), .C1(n2774), .C2(n316), .A(n1319), 
        .ZN(n1322) );
  NOR2_X1 U1339 ( .A1(n4101), .A2(n130), .ZN(n1320) );
  NOR4_X1 U1340 ( .A1(n2235), .A2(n2232), .A3(n2226), .A4(n1320), .ZN(n1321)
         );
  NAND2_X1 U1341 ( .A1(n1322), .A2(n1321), .ZN(n1326) );
  OAI22_X1 U1342 ( .A1(n136), .A2(n1324), .B1(n133), .B2(n1323), .ZN(n1325) );
  AOI221_X1 U1343 ( .B1(n143), .B2(n1326), .C1(n139), .C2(n1543), .A(n1325), 
        .ZN(n1333) );
  OAI22_X1 U1344 ( .A1(n2742), .A2(n151), .B1(n2710), .B2(n148), .ZN(n1327) );
  AOI221_X1 U1345 ( .B1(n157), .B2(n1511), .C1(n2838), .C2(n154), .A(n1327), 
        .ZN(n1332) );
  OAI22_X1 U1346 ( .A1(n3670), .A2(n163), .B1(n2966), .B2(n160), .ZN(n1328) );
  AOI221_X1 U1347 ( .B1(n2806), .B2(n169), .C1(n3606), .C2(n166), .A(n1328), 
        .ZN(n1331) );
  OAI22_X1 U1348 ( .A1(n2661), .A2(n173), .B1(n172), .B2(n395), .ZN(n1329) );
  AOI221_X1 U1349 ( .B1(n3638), .B2(n181), .C1(n178), .C2(n1641), .A(n1329), 
        .ZN(n1330) );
  NAND4_X1 U1350 ( .A1(n1333), .A2(n1332), .A3(n1331), .A4(n1330), .ZN(n3022)
         );
  MUX2_X1 U1351 ( .A(n1334), .B(DATAIN[24]), .S(n184), .Z(n4598) );
  OAI211_X1 U1352 ( .C1(n4023), .C2(n127), .A(n2241), .B(n2240), .ZN(n1335) );
  AOI221_X1 U1353 ( .B1(n307), .B2(n1868), .C1(n2775), .C2(n316), .A(n1335), 
        .ZN(n1338) );
  NOR2_X1 U1354 ( .A1(n4100), .A2(n130), .ZN(n1336) );
  NOR4_X1 U1355 ( .A1(n2247), .A2(n2244), .A3(n2238), .A4(n1336), .ZN(n1337)
         );
  NAND2_X1 U1356 ( .A1(n1338), .A2(n1337), .ZN(n1342) );
  OAI22_X1 U1357 ( .A1(n136), .A2(n1340), .B1(n133), .B2(n1339), .ZN(n1341) );
  AOI221_X1 U1358 ( .B1(n143), .B2(n1342), .C1(n139), .C2(n1544), .A(n1341), 
        .ZN(n1349) );
  OAI22_X1 U1359 ( .A1(n2743), .A2(n151), .B1(n2711), .B2(n148), .ZN(n1343) );
  AOI221_X1 U1360 ( .B1(n157), .B2(n1512), .C1(n2839), .C2(n154), .A(n1343), 
        .ZN(n1348) );
  OAI22_X1 U1361 ( .A1(n3671), .A2(n163), .B1(n2967), .B2(n160), .ZN(n1344) );
  AOI221_X1 U1362 ( .B1(n2807), .B2(n169), .C1(n3607), .C2(n166), .A(n1344), 
        .ZN(n1347) );
  OAI22_X1 U1363 ( .A1(n2660), .A2(n173), .B1(n172), .B2(n396), .ZN(n1345) );
  AOI221_X1 U1364 ( .B1(n3639), .B2(n181), .C1(n178), .C2(n1642), .A(n1345), 
        .ZN(n1346) );
  NAND4_X1 U1365 ( .A1(n1349), .A2(n1348), .A3(n1347), .A4(n1346), .ZN(n3021)
         );
  MUX2_X1 U1366 ( .A(n1350), .B(DATAIN[25]), .S(n184), .Z(n4599) );
  OAI211_X1 U1367 ( .C1(n4024), .C2(n127), .A(n2253), .B(n2252), .ZN(n1351) );
  AOI221_X1 U1368 ( .B1(n307), .B2(n1869), .C1(n2776), .C2(n316), .A(n1351), 
        .ZN(n1354) );
  NOR2_X1 U1369 ( .A1(n4099), .A2(n130), .ZN(n1352) );
  NOR4_X1 U1370 ( .A1(n2259), .A2(n2256), .A3(n2250), .A4(n1352), .ZN(n1353)
         );
  NAND2_X1 U1371 ( .A1(n1354), .A2(n1353), .ZN(n1358) );
  OAI22_X1 U1372 ( .A1(n136), .A2(n1356), .B1(n133), .B2(n1355), .ZN(n1357) );
  AOI221_X1 U1373 ( .B1(n143), .B2(n1358), .C1(n139), .C2(n1545), .A(n1357), 
        .ZN(n1365) );
  OAI22_X1 U1374 ( .A1(n2744), .A2(n151), .B1(n2712), .B2(n148), .ZN(n1359) );
  AOI221_X1 U1375 ( .B1(n157), .B2(n1513), .C1(n2840), .C2(n154), .A(n1359), 
        .ZN(n1364) );
  OAI22_X1 U1376 ( .A1(n3672), .A2(n163), .B1(n2968), .B2(n160), .ZN(n1360) );
  AOI221_X1 U1377 ( .B1(n2808), .B2(n169), .C1(n3608), .C2(n166), .A(n1360), 
        .ZN(n1363) );
  OAI22_X1 U1378 ( .A1(n2659), .A2(n173), .B1(n172), .B2(n397), .ZN(n1361) );
  AOI221_X1 U1379 ( .B1(n3640), .B2(n181), .C1(n178), .C2(n1643), .A(n1361), 
        .ZN(n1362) );
  NAND4_X1 U1380 ( .A1(n1365), .A2(n1364), .A3(n1363), .A4(n1362), .ZN(n3020)
         );
  MUX2_X1 U1381 ( .A(n1366), .B(DATAIN[26]), .S(n184), .Z(n4600) );
  OAI211_X1 U1382 ( .C1(n4025), .C2(n127), .A(n2265), .B(n2264), .ZN(n1367) );
  AOI221_X1 U1383 ( .B1(n307), .B2(n1870), .C1(n2777), .C2(n316), .A(n1367), 
        .ZN(n1370) );
  NOR2_X1 U1384 ( .A1(n4098), .A2(n130), .ZN(n1368) );
  NOR4_X1 U1385 ( .A1(n2271), .A2(n2268), .A3(n2262), .A4(n1368), .ZN(n1369)
         );
  NAND2_X1 U1386 ( .A1(n1370), .A2(n1369), .ZN(n1374) );
  OAI22_X1 U1387 ( .A1(n136), .A2(n1372), .B1(n133), .B2(n1371), .ZN(n1373) );
  AOI221_X1 U1388 ( .B1(n143), .B2(n1374), .C1(n139), .C2(n1546), .A(n1373), 
        .ZN(n1381) );
  OAI22_X1 U1389 ( .A1(n2745), .A2(n151), .B1(n2713), .B2(n148), .ZN(n1375) );
  AOI221_X1 U1390 ( .B1(n157), .B2(n1514), .C1(n2841), .C2(n154), .A(n1375), 
        .ZN(n1380) );
  OAI22_X1 U1391 ( .A1(n3673), .A2(n163), .B1(n2969), .B2(n160), .ZN(n1376) );
  AOI221_X1 U1392 ( .B1(n2809), .B2(n169), .C1(n3609), .C2(n166), .A(n1376), 
        .ZN(n1379) );
  OAI22_X1 U1393 ( .A1(n2658), .A2(n173), .B1(n172), .B2(n398), .ZN(n1377) );
  AOI221_X1 U1394 ( .B1(n3641), .B2(n181), .C1(n178), .C2(n1644), .A(n1377), 
        .ZN(n1378) );
  NAND4_X1 U1395 ( .A1(n1381), .A2(n1380), .A3(n1379), .A4(n1378), .ZN(n3019)
         );
  MUX2_X1 U1396 ( .A(n1382), .B(DATAIN[27]), .S(n184), .Z(n4601) );
  OAI211_X1 U1397 ( .C1(n4026), .C2(n127), .A(n2277), .B(n2276), .ZN(n1383) );
  AOI221_X1 U1398 ( .B1(n307), .B2(n1871), .C1(n2778), .C2(n316), .A(n1383), 
        .ZN(n1386) );
  NOR2_X1 U1399 ( .A1(n4097), .A2(n130), .ZN(n1384) );
  NOR4_X1 U1400 ( .A1(n2283), .A2(n2280), .A3(n2274), .A4(n1384), .ZN(n1385)
         );
  NAND2_X1 U1401 ( .A1(n1386), .A2(n1385), .ZN(n1390) );
  OAI22_X1 U1402 ( .A1(n136), .A2(n1388), .B1(n133), .B2(n1387), .ZN(n1389) );
  AOI221_X1 U1403 ( .B1(n142), .B2(n1390), .C1(n139), .C2(n1547), .A(n1389), 
        .ZN(n1397) );
  OAI22_X1 U1404 ( .A1(n2746), .A2(n151), .B1(n2714), .B2(n148), .ZN(n1391) );
  AOI221_X1 U1405 ( .B1(n157), .B2(n1515), .C1(n2842), .C2(n154), .A(n1391), 
        .ZN(n1396) );
  OAI22_X1 U1406 ( .A1(n3674), .A2(n163), .B1(n2970), .B2(n160), .ZN(n1392) );
  AOI221_X1 U1407 ( .B1(n2810), .B2(n169), .C1(n3610), .C2(n166), .A(n1392), 
        .ZN(n1395) );
  OAI22_X1 U1408 ( .A1(n2657), .A2(n173), .B1(n172), .B2(n399), .ZN(n1393) );
  AOI221_X1 U1409 ( .B1(n3642), .B2(n181), .C1(n178), .C2(n1645), .A(n1393), 
        .ZN(n1394) );
  NAND4_X1 U1410 ( .A1(n1397), .A2(n1396), .A3(n1395), .A4(n1394), .ZN(n3018)
         );
  MUX2_X1 U1411 ( .A(n1398), .B(DATAIN[28]), .S(n184), .Z(n4602) );
  OAI211_X1 U1412 ( .C1(n4027), .C2(n127), .A(n2289), .B(n2288), .ZN(n1399) );
  AOI221_X1 U1413 ( .B1(n307), .B2(n1872), .C1(n2779), .C2(n316), .A(n1399), 
        .ZN(n1402) );
  NOR2_X1 U1414 ( .A1(n4096), .A2(n130), .ZN(n1400) );
  NOR4_X1 U1415 ( .A1(n2295), .A2(n2292), .A3(n2286), .A4(n1400), .ZN(n1401)
         );
  NAND2_X1 U1416 ( .A1(n1402), .A2(n1401), .ZN(n1406) );
  OAI22_X1 U1417 ( .A1(n136), .A2(n1404), .B1(n133), .B2(n1403), .ZN(n1405) );
  AOI221_X1 U1418 ( .B1(n142), .B2(n1406), .C1(n139), .C2(n1548), .A(n1405), 
        .ZN(n1413) );
  OAI22_X1 U1419 ( .A1(n2747), .A2(n151), .B1(n2715), .B2(n148), .ZN(n1407) );
  AOI221_X1 U1420 ( .B1(n157), .B2(n1516), .C1(n2843), .C2(n154), .A(n1407), 
        .ZN(n1412) );
  OAI22_X1 U1421 ( .A1(n3675), .A2(n163), .B1(n2971), .B2(n160), .ZN(n1408) );
  AOI221_X1 U1422 ( .B1(n2811), .B2(n169), .C1(n3611), .C2(n166), .A(n1408), 
        .ZN(n1411) );
  OAI22_X1 U1423 ( .A1(n2656), .A2(n173), .B1(n172), .B2(n400), .ZN(n1409) );
  AOI221_X1 U1424 ( .B1(n3643), .B2(n181), .C1(n178), .C2(n1646), .A(n1409), 
        .ZN(n1410) );
  NAND4_X1 U1425 ( .A1(n1413), .A2(n1412), .A3(n1411), .A4(n1410), .ZN(n3017)
         );
  MUX2_X1 U1426 ( .A(n1414), .B(DATAIN[29]), .S(n184), .Z(n4603) );
  OAI211_X1 U1427 ( .C1(n4028), .C2(n127), .A(n2301), .B(n2300), .ZN(n1415) );
  AOI221_X1 U1428 ( .B1(n307), .B2(n1873), .C1(n2780), .C2(n316), .A(n1415), 
        .ZN(n1418) );
  NOR2_X1 U1429 ( .A1(n4095), .A2(n130), .ZN(n1416) );
  NOR4_X1 U1430 ( .A1(n2307), .A2(n2304), .A3(n2298), .A4(n1416), .ZN(n1417)
         );
  NAND2_X1 U1431 ( .A1(n1418), .A2(n1417), .ZN(n1422) );
  OAI22_X1 U1432 ( .A1(n136), .A2(n1420), .B1(n133), .B2(n1419), .ZN(n1421) );
  AOI221_X1 U1433 ( .B1(n142), .B2(n1422), .C1(n139), .C2(n1549), .A(n1421), 
        .ZN(n1429) );
  OAI22_X1 U1434 ( .A1(n2748), .A2(n151), .B1(n2716), .B2(n148), .ZN(n1423) );
  AOI221_X1 U1435 ( .B1(n157), .B2(n1517), .C1(n2844), .C2(n154), .A(n1423), 
        .ZN(n1428) );
  OAI22_X1 U1436 ( .A1(n3676), .A2(n163), .B1(n2972), .B2(n160), .ZN(n1424) );
  AOI221_X1 U1437 ( .B1(n2812), .B2(n169), .C1(n3612), .C2(n166), .A(n1424), 
        .ZN(n1427) );
  OAI22_X1 U1438 ( .A1(n2655), .A2(n173), .B1(n172), .B2(n401), .ZN(n1425) );
  AOI221_X1 U1439 ( .B1(n3644), .B2(n181), .C1(n178), .C2(n1647), .A(n1425), 
        .ZN(n1426) );
  NAND4_X1 U1440 ( .A1(n1429), .A2(n1428), .A3(n1427), .A4(n1426), .ZN(n3016)
         );
  MUX2_X1 U1441 ( .A(n1430), .B(DATAIN[30]), .S(n184), .Z(n4604) );
  OAI211_X1 U1442 ( .C1(n4029), .C2(n127), .A(n2324), .B(n2323), .ZN(n1431) );
  AOI221_X1 U1443 ( .B1(n307), .B2(n1874), .C1(n316), .C2(n2781), .A(n1431), 
        .ZN(n1434) );
  NOR2_X1 U1444 ( .A1(n4094), .A2(n130), .ZN(n1432) );
  NOR4_X1 U1445 ( .A1(n2336), .A2(n2329), .A3(n2319), .A4(n1432), .ZN(n1433)
         );
  NAND2_X1 U1446 ( .A1(n1434), .A2(n1433), .ZN(n1440) );
  OAI22_X1 U1447 ( .A1(n136), .A2(n1437), .B1(n133), .B2(n1435), .ZN(n1439) );
  AOI221_X1 U1448 ( .B1(n144), .B2(n1440), .C1(n139), .C2(n1550), .A(n1439), 
        .ZN(n1453) );
  OAI22_X1 U1449 ( .A1(n2749), .A2(n151), .B1(n2717), .B2(n148), .ZN(n1444) );
  AOI221_X1 U1450 ( .B1(n157), .B2(n1518), .C1(n2845), .C2(n154), .A(n1444), 
        .ZN(n1452) );
  OAI22_X1 U1451 ( .A1(n3677), .A2(n163), .B1(n2973), .B2(n160), .ZN(n1447) );
  AOI221_X1 U1452 ( .B1(n2813), .B2(n169), .C1(n3613), .C2(n166), .A(n1447), 
        .ZN(n1451) );
  OAI22_X1 U1453 ( .A1(n2654), .A2(n174), .B1(n172), .B2(n402), .ZN(n1449) );
  AOI221_X1 U1454 ( .B1(n3645), .B2(n181), .C1(n178), .C2(n1648), .A(n1449), 
        .ZN(n1450) );
  NAND4_X1 U1455 ( .A1(n1453), .A2(n1452), .A3(n1451), .A4(n1450), .ZN(n3015)
         );
  MUX2_X1 U1456 ( .A(n1454), .B(DATAIN[31]), .S(n184), .Z(n4605) );
  MUX2_X1 U1457 ( .A(n1455), .B(DATAIN[0]), .S(n185), .Z(n4542) );
  MUX2_X1 U1458 ( .A(n1456), .B(DATAIN[1]), .S(n185), .Z(n4543) );
  MUX2_X1 U1459 ( .A(n1457), .B(DATAIN[2]), .S(n185), .Z(n4544) );
  MUX2_X1 U1460 ( .A(n1458), .B(DATAIN[3]), .S(n185), .Z(n4545) );
  MUX2_X1 U1461 ( .A(n1459), .B(DATAIN[4]), .S(n185), .Z(n4546) );
  MUX2_X1 U1462 ( .A(n1460), .B(DATAIN[5]), .S(n185), .Z(n4547) );
  MUX2_X1 U1463 ( .A(n1461), .B(DATAIN[6]), .S(n185), .Z(n4548) );
  MUX2_X1 U1464 ( .A(n1462), .B(DATAIN[7]), .S(n185), .Z(n4549) );
  MUX2_X1 U1465 ( .A(n1463), .B(DATAIN[8]), .S(n185), .Z(n4550) );
  MUX2_X1 U1466 ( .A(n1464), .B(DATAIN[9]), .S(n185), .Z(n4551) );
  MUX2_X1 U1467 ( .A(n1465), .B(DATAIN[10]), .S(n185), .Z(n4552) );
  MUX2_X1 U1468 ( .A(n1466), .B(DATAIN[11]), .S(n185), .Z(n4553) );
  MUX2_X1 U1469 ( .A(n1467), .B(DATAIN[12]), .S(n186), .Z(n4554) );
  MUX2_X1 U1470 ( .A(n1468), .B(DATAIN[13]), .S(n186), .Z(n4555) );
  MUX2_X1 U1471 ( .A(n1469), .B(DATAIN[14]), .S(n186), .Z(n4556) );
  MUX2_X1 U1472 ( .A(n1470), .B(DATAIN[15]), .S(n186), .Z(n4557) );
  MUX2_X1 U1473 ( .A(n1471), .B(DATAIN[16]), .S(n186), .Z(n4558) );
  MUX2_X1 U1474 ( .A(n1472), .B(DATAIN[17]), .S(n186), .Z(n4559) );
  MUX2_X1 U1475 ( .A(n1473), .B(DATAIN[18]), .S(n186), .Z(n4560) );
  MUX2_X1 U1476 ( .A(n1474), .B(DATAIN[19]), .S(n186), .Z(n4561) );
  MUX2_X1 U1477 ( .A(n1475), .B(DATAIN[20]), .S(n186), .Z(n4562) );
  MUX2_X1 U1478 ( .A(n1476), .B(DATAIN[21]), .S(n186), .Z(n4563) );
  MUX2_X1 U1479 ( .A(n1477), .B(DATAIN[22]), .S(n186), .Z(n4564) );
  MUX2_X1 U1480 ( .A(n1478), .B(DATAIN[23]), .S(n186), .Z(n4565) );
  MUX2_X1 U1481 ( .A(n1479), .B(DATAIN[24]), .S(n187), .Z(n4566) );
  MUX2_X1 U1482 ( .A(n1480), .B(DATAIN[25]), .S(n187), .Z(n4567) );
  MUX2_X1 U1483 ( .A(n1481), .B(DATAIN[26]), .S(n187), .Z(n4568) );
  MUX2_X1 U1484 ( .A(n1482), .B(DATAIN[27]), .S(n187), .Z(n4569) );
  MUX2_X1 U1485 ( .A(n1483), .B(DATAIN[28]), .S(n187), .Z(n4570) );
  MUX2_X1 U1486 ( .A(n1484), .B(DATAIN[29]), .S(n187), .Z(n4571) );
  MUX2_X1 U1487 ( .A(n1485), .B(DATAIN[30]), .S(n187), .Z(n4572) );
  MUX2_X1 U1488 ( .A(n1486), .B(DATAIN[31]), .S(n187), .Z(n4573) );
  INV_X1 U1489 ( .A(ADD_WR[1]), .ZN(n1552) );
  MUX2_X1 U1490 ( .A(n2750), .B(DATAIN[0]), .S(n188), .Z(n3047) );
  MUX2_X1 U1491 ( .A(n2751), .B(DATAIN[1]), .S(n188), .Z(n3048) );
  MUX2_X1 U1492 ( .A(n2752), .B(DATAIN[2]), .S(n188), .Z(n3049) );
  MUX2_X1 U1493 ( .A(n2753), .B(DATAIN[3]), .S(n188), .Z(n3050) );
  MUX2_X1 U1494 ( .A(n2754), .B(DATAIN[4]), .S(n188), .Z(n3051) );
  MUX2_X1 U1495 ( .A(n2755), .B(DATAIN[5]), .S(n188), .Z(n3052) );
  MUX2_X1 U1496 ( .A(n2756), .B(DATAIN[6]), .S(n188), .Z(n3053) );
  MUX2_X1 U1497 ( .A(n2757), .B(DATAIN[7]), .S(n188), .Z(n3054) );
  MUX2_X1 U1498 ( .A(n2758), .B(DATAIN[8]), .S(n188), .Z(n3055) );
  MUX2_X1 U1499 ( .A(n2759), .B(DATAIN[9]), .S(n188), .Z(n3056) );
  MUX2_X1 U1500 ( .A(n2760), .B(DATAIN[10]), .S(n188), .Z(n3057) );
  MUX2_X1 U1501 ( .A(n2761), .B(DATAIN[11]), .S(n188), .Z(n3058) );
  MUX2_X1 U1502 ( .A(n2762), .B(DATAIN[12]), .S(n189), .Z(n3059) );
  MUX2_X1 U1503 ( .A(n2763), .B(DATAIN[13]), .S(n189), .Z(n3060) );
  MUX2_X1 U1504 ( .A(n2764), .B(DATAIN[14]), .S(n189), .Z(n3061) );
  MUX2_X1 U1505 ( .A(n2765), .B(DATAIN[15]), .S(n189), .Z(n3062) );
  MUX2_X1 U1506 ( .A(n2766), .B(DATAIN[16]), .S(n189), .Z(n3063) );
  MUX2_X1 U1507 ( .A(n2767), .B(DATAIN[17]), .S(n189), .Z(n3064) );
  MUX2_X1 U1508 ( .A(n2768), .B(DATAIN[18]), .S(n189), .Z(n3065) );
  MUX2_X1 U1509 ( .A(n2769), .B(DATAIN[19]), .S(n189), .Z(n3066) );
  MUX2_X1 U1510 ( .A(n2770), .B(DATAIN[20]), .S(n189), .Z(n3067) );
  MUX2_X1 U1511 ( .A(n2771), .B(DATAIN[21]), .S(n189), .Z(n3068) );
  MUX2_X1 U1512 ( .A(n2772), .B(DATAIN[22]), .S(n189), .Z(n3069) );
  MUX2_X1 U1513 ( .A(n2773), .B(DATAIN[23]), .S(n189), .Z(n3070) );
  MUX2_X1 U1514 ( .A(n2774), .B(DATAIN[24]), .S(n190), .Z(n3071) );
  MUX2_X1 U1515 ( .A(n2775), .B(DATAIN[25]), .S(n190), .Z(n3072) );
  MUX2_X1 U1516 ( .A(n2776), .B(DATAIN[26]), .S(n190), .Z(n3073) );
  MUX2_X1 U1517 ( .A(n2777), .B(DATAIN[27]), .S(n190), .Z(n3074) );
  MUX2_X1 U1518 ( .A(n2778), .B(DATAIN[28]), .S(n190), .Z(n3075) );
  MUX2_X1 U1519 ( .A(n2779), .B(DATAIN[29]), .S(n190), .Z(n3076) );
  MUX2_X1 U1520 ( .A(n2780), .B(DATAIN[30]), .S(n190), .Z(n3077) );
  MUX2_X1 U1521 ( .A(n2781), .B(DATAIN[31]), .S(n190), .Z(n3078) );
  MUX2_X1 U1522 ( .A(n2782), .B(DATAIN[0]), .S(n191), .Z(n3079) );
  MUX2_X1 U1523 ( .A(n2783), .B(DATAIN[1]), .S(n191), .Z(n3080) );
  MUX2_X1 U1524 ( .A(n2784), .B(DATAIN[2]), .S(n191), .Z(n3081) );
  MUX2_X1 U1525 ( .A(n2785), .B(DATAIN[3]), .S(n191), .Z(n3082) );
  MUX2_X1 U1526 ( .A(n2786), .B(DATAIN[4]), .S(n191), .Z(n3083) );
  MUX2_X1 U1527 ( .A(n2787), .B(DATAIN[5]), .S(n191), .Z(n3084) );
  MUX2_X1 U1528 ( .A(n2788), .B(DATAIN[6]), .S(n191), .Z(n3085) );
  MUX2_X1 U1529 ( .A(n2789), .B(DATAIN[7]), .S(n191), .Z(n3086) );
  MUX2_X1 U1530 ( .A(n2790), .B(DATAIN[8]), .S(n191), .Z(n3087) );
  MUX2_X1 U1531 ( .A(n2791), .B(DATAIN[9]), .S(n191), .Z(n3088) );
  MUX2_X1 U1532 ( .A(n2792), .B(DATAIN[10]), .S(n191), .Z(n3089) );
  MUX2_X1 U1533 ( .A(n2793), .B(DATAIN[11]), .S(n191), .Z(n3090) );
  MUX2_X1 U1534 ( .A(n2794), .B(DATAIN[12]), .S(n192), .Z(n3091) );
  MUX2_X1 U1535 ( .A(n2795), .B(DATAIN[13]), .S(n192), .Z(n3092) );
  MUX2_X1 U1536 ( .A(n2796), .B(DATAIN[14]), .S(n192), .Z(n3093) );
  MUX2_X1 U1537 ( .A(n2797), .B(DATAIN[15]), .S(n192), .Z(n3094) );
  MUX2_X1 U1538 ( .A(n2798), .B(DATAIN[16]), .S(n192), .Z(n3095) );
  MUX2_X1 U1539 ( .A(n2799), .B(DATAIN[17]), .S(n192), .Z(n3096) );
  MUX2_X1 U1540 ( .A(n2800), .B(DATAIN[18]), .S(n192), .Z(n3097) );
  MUX2_X1 U1541 ( .A(n2801), .B(DATAIN[19]), .S(n192), .Z(n3098) );
  MUX2_X1 U1542 ( .A(n2802), .B(DATAIN[20]), .S(n192), .Z(n3099) );
  MUX2_X1 U1543 ( .A(n2803), .B(DATAIN[21]), .S(n192), .Z(n3100) );
  MUX2_X1 U1544 ( .A(n2804), .B(DATAIN[22]), .S(n192), .Z(n3101) );
  MUX2_X1 U1545 ( .A(n2805), .B(DATAIN[23]), .S(n192), .Z(n3102) );
  MUX2_X1 U1546 ( .A(n2806), .B(DATAIN[24]), .S(n193), .Z(n3103) );
  MUX2_X1 U1547 ( .A(n2807), .B(DATAIN[25]), .S(n193), .Z(n3104) );
  MUX2_X1 U1548 ( .A(n2808), .B(DATAIN[26]), .S(n193), .Z(n3105) );
  MUX2_X1 U1549 ( .A(n2809), .B(DATAIN[27]), .S(n193), .Z(n3106) );
  MUX2_X1 U1550 ( .A(n2810), .B(DATAIN[28]), .S(n193), .Z(n3107) );
  MUX2_X1 U1551 ( .A(n2811), .B(DATAIN[29]), .S(n193), .Z(n3108) );
  MUX2_X1 U1552 ( .A(n2812), .B(DATAIN[30]), .S(n193), .Z(n3109) );
  MUX2_X1 U1553 ( .A(n2813), .B(DATAIN[31]), .S(n193), .Z(n3110) );
  INV_X1 U1554 ( .A(ADD_WR[2]), .ZN(n1551) );
  MUX2_X1 U1555 ( .A(n1487), .B(DATAIN[0]), .S(n194), .Z(n4510) );
  MUX2_X1 U1556 ( .A(n1488), .B(DATAIN[1]), .S(n194), .Z(n4511) );
  MUX2_X1 U1557 ( .A(n1489), .B(DATAIN[2]), .S(n194), .Z(n4512) );
  MUX2_X1 U1558 ( .A(n1490), .B(DATAIN[3]), .S(n194), .Z(n4513) );
  MUX2_X1 U1559 ( .A(n1491), .B(DATAIN[4]), .S(n194), .Z(n4514) );
  MUX2_X1 U1560 ( .A(n1492), .B(DATAIN[5]), .S(n194), .Z(n4515) );
  MUX2_X1 U1561 ( .A(n1493), .B(DATAIN[6]), .S(n194), .Z(n4516) );
  MUX2_X1 U1562 ( .A(n1494), .B(DATAIN[7]), .S(n194), .Z(n4517) );
  MUX2_X1 U1563 ( .A(n1495), .B(DATAIN[8]), .S(n194), .Z(n4518) );
  MUX2_X1 U1564 ( .A(n1496), .B(DATAIN[9]), .S(n194), .Z(n4519) );
  MUX2_X1 U1565 ( .A(n1497), .B(DATAIN[10]), .S(n194), .Z(n4520) );
  MUX2_X1 U1566 ( .A(n1498), .B(DATAIN[11]), .S(n194), .Z(n4521) );
  MUX2_X1 U1567 ( .A(n1499), .B(DATAIN[12]), .S(n195), .Z(n4522) );
  MUX2_X1 U1568 ( .A(n1500), .B(DATAIN[13]), .S(n195), .Z(n4523) );
  MUX2_X1 U1569 ( .A(n1501), .B(DATAIN[14]), .S(n195), .Z(n4524) );
  MUX2_X1 U1570 ( .A(n1502), .B(DATAIN[15]), .S(n195), .Z(n4525) );
  MUX2_X1 U1571 ( .A(n1503), .B(DATAIN[16]), .S(n195), .Z(n4526) );
  MUX2_X1 U1572 ( .A(n1504), .B(DATAIN[17]), .S(n195), .Z(n4527) );
  MUX2_X1 U1573 ( .A(n1505), .B(DATAIN[18]), .S(n195), .Z(n4528) );
  MUX2_X1 U1574 ( .A(n1506), .B(DATAIN[19]), .S(n195), .Z(n4529) );
  MUX2_X1 U1575 ( .A(n1507), .B(DATAIN[20]), .S(n195), .Z(n4530) );
  MUX2_X1 U1576 ( .A(n1508), .B(DATAIN[21]), .S(n195), .Z(n4531) );
  MUX2_X1 U1577 ( .A(n1509), .B(DATAIN[22]), .S(n195), .Z(n4532) );
  MUX2_X1 U1578 ( .A(n1510), .B(DATAIN[23]), .S(n195), .Z(n4533) );
  MUX2_X1 U1579 ( .A(n1511), .B(DATAIN[24]), .S(n196), .Z(n4534) );
  MUX2_X1 U1580 ( .A(n1512), .B(DATAIN[25]), .S(n196), .Z(n4535) );
  MUX2_X1 U1581 ( .A(n1513), .B(DATAIN[26]), .S(n196), .Z(n4536) );
  MUX2_X1 U1582 ( .A(n1514), .B(DATAIN[27]), .S(n196), .Z(n4537) );
  MUX2_X1 U1583 ( .A(n1515), .B(DATAIN[28]), .S(n196), .Z(n4538) );
  MUX2_X1 U1584 ( .A(n1516), .B(DATAIN[29]), .S(n196), .Z(n4539) );
  MUX2_X1 U1585 ( .A(n1517), .B(DATAIN[30]), .S(n196), .Z(n4540) );
  MUX2_X1 U1586 ( .A(n1518), .B(DATAIN[31]), .S(n196), .Z(n4541) );
  MUX2_X1 U1587 ( .A(n1519), .B(DATAIN[0]), .S(n197), .Z(n4478) );
  MUX2_X1 U1588 ( .A(n1520), .B(DATAIN[1]), .S(n197), .Z(n4479) );
  MUX2_X1 U1589 ( .A(n1521), .B(DATAIN[2]), .S(n197), .Z(n4480) );
  MUX2_X1 U1590 ( .A(n1522), .B(DATAIN[3]), .S(n197), .Z(n4481) );
  MUX2_X1 U1591 ( .A(n1523), .B(DATAIN[4]), .S(n197), .Z(n4482) );
  MUX2_X1 U1592 ( .A(n1524), .B(DATAIN[5]), .S(n197), .Z(n4483) );
  MUX2_X1 U1593 ( .A(n1525), .B(DATAIN[6]), .S(n197), .Z(n4484) );
  MUX2_X1 U1594 ( .A(n1526), .B(DATAIN[7]), .S(n197), .Z(n4485) );
  MUX2_X1 U1595 ( .A(n1527), .B(DATAIN[8]), .S(n197), .Z(n4486) );
  MUX2_X1 U1596 ( .A(n1528), .B(DATAIN[9]), .S(n197), .Z(n4487) );
  MUX2_X1 U1597 ( .A(n1529), .B(DATAIN[10]), .S(n197), .Z(n4488) );
  MUX2_X1 U1598 ( .A(n1530), .B(DATAIN[11]), .S(n197), .Z(n4489) );
  MUX2_X1 U1599 ( .A(n1531), .B(DATAIN[12]), .S(n198), .Z(n4490) );
  MUX2_X1 U1600 ( .A(n1532), .B(DATAIN[13]), .S(n198), .Z(n4491) );
  MUX2_X1 U1601 ( .A(n1533), .B(DATAIN[14]), .S(n198), .Z(n4492) );
  MUX2_X1 U1602 ( .A(n1534), .B(DATAIN[15]), .S(n198), .Z(n4493) );
  MUX2_X1 U1603 ( .A(n1535), .B(DATAIN[16]), .S(n198), .Z(n4494) );
  MUX2_X1 U1604 ( .A(n1536), .B(DATAIN[17]), .S(n198), .Z(n4495) );
  MUX2_X1 U1605 ( .A(n1537), .B(DATAIN[18]), .S(n198), .Z(n4496) );
  MUX2_X1 U1606 ( .A(n1538), .B(DATAIN[19]), .S(n198), .Z(n4497) );
  MUX2_X1 U1607 ( .A(n1539), .B(DATAIN[20]), .S(n198), .Z(n4498) );
  MUX2_X1 U1608 ( .A(n1540), .B(DATAIN[21]), .S(n198), .Z(n4499) );
  MUX2_X1 U1609 ( .A(n1541), .B(DATAIN[22]), .S(n198), .Z(n4500) );
  MUX2_X1 U1610 ( .A(n1542), .B(DATAIN[23]), .S(n198), .Z(n4501) );
  MUX2_X1 U1611 ( .A(n1543), .B(DATAIN[24]), .S(n199), .Z(n4502) );
  MUX2_X1 U1612 ( .A(n1544), .B(DATAIN[25]), .S(n199), .Z(n4503) );
  MUX2_X1 U1613 ( .A(n1545), .B(DATAIN[26]), .S(n199), .Z(n4504) );
  MUX2_X1 U1614 ( .A(n1546), .B(DATAIN[27]), .S(n199), .Z(n4505) );
  MUX2_X1 U1615 ( .A(n1547), .B(DATAIN[28]), .S(n199), .Z(n4506) );
  MUX2_X1 U1616 ( .A(n1548), .B(DATAIN[29]), .S(n199), .Z(n4507) );
  MUX2_X1 U1617 ( .A(n1549), .B(DATAIN[30]), .S(n199), .Z(n4508) );
  MUX2_X1 U1618 ( .A(n1550), .B(DATAIN[31]), .S(n199), .Z(n4509) );
  MUX2_X1 U1619 ( .A(n2814), .B(DATAIN[0]), .S(n200), .Z(n3111) );
  MUX2_X1 U1620 ( .A(n2815), .B(DATAIN[1]), .S(n200), .Z(n3112) );
  MUX2_X1 U1621 ( .A(n2816), .B(DATAIN[2]), .S(n200), .Z(n3113) );
  MUX2_X1 U1622 ( .A(n2817), .B(DATAIN[3]), .S(n200), .Z(n3114) );
  MUX2_X1 U1623 ( .A(n2818), .B(DATAIN[4]), .S(n200), .Z(n3115) );
  MUX2_X1 U1624 ( .A(n2819), .B(DATAIN[5]), .S(n200), .Z(n3116) );
  MUX2_X1 U1625 ( .A(n2820), .B(DATAIN[6]), .S(n200), .Z(n3117) );
  MUX2_X1 U1626 ( .A(n2821), .B(DATAIN[7]), .S(n200), .Z(n3118) );
  MUX2_X1 U1627 ( .A(n2822), .B(DATAIN[8]), .S(n200), .Z(n3119) );
  MUX2_X1 U1628 ( .A(n2823), .B(DATAIN[9]), .S(n200), .Z(n3120) );
  MUX2_X1 U1629 ( .A(n2824), .B(DATAIN[10]), .S(n200), .Z(n3121) );
  MUX2_X1 U1630 ( .A(n2825), .B(DATAIN[11]), .S(n200), .Z(n3122) );
  MUX2_X1 U1631 ( .A(n2826), .B(DATAIN[12]), .S(n201), .Z(n3123) );
  MUX2_X1 U1632 ( .A(n2827), .B(DATAIN[13]), .S(n201), .Z(n3124) );
  MUX2_X1 U1633 ( .A(n2828), .B(DATAIN[14]), .S(n201), .Z(n3125) );
  MUX2_X1 U1634 ( .A(n2829), .B(DATAIN[15]), .S(n201), .Z(n3126) );
  MUX2_X1 U1635 ( .A(n2830), .B(DATAIN[16]), .S(n201), .Z(n3127) );
  MUX2_X1 U1636 ( .A(n2831), .B(DATAIN[17]), .S(n201), .Z(n3128) );
  MUX2_X1 U1637 ( .A(n2832), .B(DATAIN[18]), .S(n201), .Z(n3129) );
  MUX2_X1 U1638 ( .A(n2833), .B(DATAIN[19]), .S(n201), .Z(n3130) );
  MUX2_X1 U1639 ( .A(n2834), .B(DATAIN[20]), .S(n201), .Z(n3131) );
  MUX2_X1 U1640 ( .A(n2835), .B(DATAIN[21]), .S(n201), .Z(n3132) );
  MUX2_X1 U1641 ( .A(n2836), .B(DATAIN[22]), .S(n201), .Z(n3133) );
  MUX2_X1 U1642 ( .A(n2837), .B(DATAIN[23]), .S(n201), .Z(n3134) );
  MUX2_X1 U1643 ( .A(n2838), .B(DATAIN[24]), .S(n202), .Z(n3135) );
  MUX2_X1 U1644 ( .A(n2839), .B(DATAIN[25]), .S(n202), .Z(n3136) );
  MUX2_X1 U1645 ( .A(n2840), .B(DATAIN[26]), .S(n202), .Z(n3137) );
  MUX2_X1 U1646 ( .A(n2841), .B(DATAIN[27]), .S(n202), .Z(n3138) );
  MUX2_X1 U1647 ( .A(n2842), .B(DATAIN[28]), .S(n202), .Z(n3139) );
  MUX2_X1 U1648 ( .A(n2843), .B(DATAIN[29]), .S(n202), .Z(n3140) );
  MUX2_X1 U1649 ( .A(n2844), .B(DATAIN[30]), .S(n202), .Z(n3141) );
  MUX2_X1 U1650 ( .A(n2845), .B(DATAIN[31]), .S(n202), .Z(n3142) );
  MUX2_X1 U1651 ( .A(n2846), .B(DATAIN[0]), .S(n203), .Z(n3143) );
  MUX2_X1 U1652 ( .A(n2847), .B(DATAIN[1]), .S(n203), .Z(n3144) );
  MUX2_X1 U1653 ( .A(n2848), .B(DATAIN[2]), .S(n203), .Z(n3145) );
  MUX2_X1 U1654 ( .A(n2849), .B(DATAIN[3]), .S(n203), .Z(n3146) );
  MUX2_X1 U1655 ( .A(n2850), .B(DATAIN[4]), .S(n203), .Z(n3147) );
  MUX2_X1 U1656 ( .A(n2851), .B(DATAIN[5]), .S(n203), .Z(n3148) );
  MUX2_X1 U1657 ( .A(n2852), .B(DATAIN[6]), .S(n203), .Z(n3149) );
  MUX2_X1 U1658 ( .A(n2853), .B(DATAIN[7]), .S(n203), .Z(n3150) );
  MUX2_X1 U1659 ( .A(n2854), .B(DATAIN[8]), .S(n203), .Z(n3151) );
  MUX2_X1 U1660 ( .A(n2855), .B(DATAIN[9]), .S(n203), .Z(n3152) );
  MUX2_X1 U1661 ( .A(n2856), .B(DATAIN[10]), .S(n203), .Z(n3153) );
  MUX2_X1 U1662 ( .A(n2857), .B(DATAIN[11]), .S(n203), .Z(n3154) );
  MUX2_X1 U1663 ( .A(n2858), .B(DATAIN[12]), .S(n204), .Z(n3155) );
  MUX2_X1 U1664 ( .A(n2859), .B(DATAIN[13]), .S(n204), .Z(n3156) );
  MUX2_X1 U1665 ( .A(n2860), .B(DATAIN[14]), .S(n204), .Z(n3157) );
  MUX2_X1 U1666 ( .A(n2861), .B(DATAIN[15]), .S(n204), .Z(n3158) );
  MUX2_X1 U1667 ( .A(n2862), .B(DATAIN[16]), .S(n204), .Z(n3159) );
  MUX2_X1 U1668 ( .A(n2863), .B(DATAIN[17]), .S(n204), .Z(n3160) );
  MUX2_X1 U1669 ( .A(n2864), .B(DATAIN[18]), .S(n204), .Z(n3161) );
  MUX2_X1 U1670 ( .A(n2865), .B(DATAIN[19]), .S(n204), .Z(n3162) );
  MUX2_X1 U1671 ( .A(n2866), .B(DATAIN[20]), .S(n204), .Z(n3163) );
  MUX2_X1 U1672 ( .A(n2867), .B(DATAIN[21]), .S(n204), .Z(n3164) );
  MUX2_X1 U1673 ( .A(n2868), .B(DATAIN[22]), .S(n204), .Z(n3165) );
  MUX2_X1 U1674 ( .A(n2869), .B(DATAIN[23]), .S(n204), .Z(n3166) );
  MUX2_X1 U1675 ( .A(n2870), .B(DATAIN[24]), .S(n205), .Z(n3167) );
  MUX2_X1 U1676 ( .A(n2871), .B(DATAIN[25]), .S(n205), .Z(n3168) );
  MUX2_X1 U1677 ( .A(n2872), .B(DATAIN[26]), .S(n205), .Z(n3169) );
  MUX2_X1 U1678 ( .A(n2873), .B(DATAIN[27]), .S(n205), .Z(n3170) );
  MUX2_X1 U1679 ( .A(n2874), .B(DATAIN[28]), .S(n205), .Z(n3171) );
  MUX2_X1 U1680 ( .A(n2875), .B(DATAIN[29]), .S(n205), .Z(n3172) );
  MUX2_X1 U1681 ( .A(n2876), .B(DATAIN[30]), .S(n205), .Z(n3173) );
  MUX2_X1 U1682 ( .A(n2877), .B(DATAIN[31]), .S(n205), .Z(n3174) );
  INV_X1 U1683 ( .A(ADD_WR[3]), .ZN(n1810) );
  MUX2_X1 U1684 ( .A(n2878), .B(DATAIN[0]), .S(n206), .Z(n3175) );
  MUX2_X1 U1685 ( .A(n2879), .B(DATAIN[1]), .S(n206), .Z(n3176) );
  MUX2_X1 U1686 ( .A(n2880), .B(DATAIN[2]), .S(n206), .Z(n3177) );
  MUX2_X1 U1687 ( .A(n2881), .B(DATAIN[3]), .S(n206), .Z(n3178) );
  MUX2_X1 U1688 ( .A(n2882), .B(DATAIN[4]), .S(n206), .Z(n3179) );
  MUX2_X1 U1689 ( .A(n2883), .B(DATAIN[5]), .S(n206), .Z(n3180) );
  MUX2_X1 U1690 ( .A(n2884), .B(DATAIN[6]), .S(n206), .Z(n3181) );
  MUX2_X1 U1691 ( .A(n2885), .B(DATAIN[7]), .S(n206), .Z(n3182) );
  MUX2_X1 U1692 ( .A(n2886), .B(DATAIN[8]), .S(n206), .Z(n3183) );
  MUX2_X1 U1693 ( .A(n2887), .B(DATAIN[9]), .S(n206), .Z(n3184) );
  MUX2_X1 U1694 ( .A(n2888), .B(DATAIN[10]), .S(n206), .Z(n3185) );
  MUX2_X1 U1695 ( .A(n2889), .B(DATAIN[11]), .S(n206), .Z(n3186) );
  MUX2_X1 U1696 ( .A(n2890), .B(DATAIN[12]), .S(n207), .Z(n3187) );
  MUX2_X1 U1697 ( .A(n2891), .B(DATAIN[13]), .S(n207), .Z(n3188) );
  MUX2_X1 U1698 ( .A(n2892), .B(DATAIN[14]), .S(n207), .Z(n3189) );
  MUX2_X1 U1699 ( .A(n2893), .B(DATAIN[15]), .S(n207), .Z(n3190) );
  MUX2_X1 U1700 ( .A(n2894), .B(DATAIN[16]), .S(n207), .Z(n3191) );
  MUX2_X1 U1701 ( .A(n2895), .B(DATAIN[17]), .S(n207), .Z(n3192) );
  MUX2_X1 U1702 ( .A(n2896), .B(DATAIN[18]), .S(n207), .Z(n3193) );
  MUX2_X1 U1703 ( .A(n2897), .B(DATAIN[19]), .S(n207), .Z(n3194) );
  MUX2_X1 U1704 ( .A(n2898), .B(DATAIN[20]), .S(n207), .Z(n3195) );
  MUX2_X1 U1705 ( .A(n2899), .B(DATAIN[21]), .S(n207), .Z(n3196) );
  MUX2_X1 U1706 ( .A(n2900), .B(DATAIN[22]), .S(n207), .Z(n3197) );
  MUX2_X1 U1707 ( .A(n2901), .B(DATAIN[23]), .S(n207), .Z(n3198) );
  MUX2_X1 U1708 ( .A(n2902), .B(DATAIN[24]), .S(n208), .Z(n3199) );
  MUX2_X1 U1709 ( .A(n2903), .B(DATAIN[25]), .S(n208), .Z(n3200) );
  MUX2_X1 U1710 ( .A(n2904), .B(DATAIN[26]), .S(n208), .Z(n3201) );
  MUX2_X1 U1711 ( .A(n2905), .B(DATAIN[27]), .S(n208), .Z(n3202) );
  MUX2_X1 U1712 ( .A(n2906), .B(DATAIN[28]), .S(n208), .Z(n3203) );
  MUX2_X1 U1713 ( .A(n2907), .B(DATAIN[29]), .S(n208), .Z(n3204) );
  MUX2_X1 U1714 ( .A(n2908), .B(DATAIN[30]), .S(n208), .Z(n3205) );
  MUX2_X1 U1715 ( .A(n2909), .B(DATAIN[31]), .S(n208), .Z(n3206) );
  MUX2_X1 U1716 ( .A(n2910), .B(DATAIN[0]), .S(n209), .Z(n3207) );
  MUX2_X1 U1717 ( .A(n2911), .B(DATAIN[1]), .S(n209), .Z(n3208) );
  MUX2_X1 U1718 ( .A(n2912), .B(DATAIN[2]), .S(n209), .Z(n3209) );
  MUX2_X1 U1719 ( .A(n2913), .B(DATAIN[3]), .S(n209), .Z(n3210) );
  MUX2_X1 U1720 ( .A(n2914), .B(DATAIN[4]), .S(n209), .Z(n3211) );
  MUX2_X1 U1721 ( .A(n2915), .B(DATAIN[5]), .S(n209), .Z(n3212) );
  MUX2_X1 U1722 ( .A(n2916), .B(DATAIN[6]), .S(n209), .Z(n3213) );
  MUX2_X1 U1723 ( .A(n2917), .B(DATAIN[7]), .S(n209), .Z(n3214) );
  MUX2_X1 U1724 ( .A(n2918), .B(DATAIN[8]), .S(n209), .Z(n3215) );
  MUX2_X1 U1725 ( .A(n2919), .B(DATAIN[9]), .S(n209), .Z(n3216) );
  MUX2_X1 U1726 ( .A(n2920), .B(DATAIN[10]), .S(n209), .Z(n3217) );
  MUX2_X1 U1727 ( .A(n2921), .B(DATAIN[11]), .S(n209), .Z(n3218) );
  MUX2_X1 U1728 ( .A(n2922), .B(DATAIN[12]), .S(n210), .Z(n3219) );
  MUX2_X1 U1729 ( .A(n2923), .B(DATAIN[13]), .S(n210), .Z(n3220) );
  MUX2_X1 U1730 ( .A(n2924), .B(DATAIN[14]), .S(n210), .Z(n3221) );
  MUX2_X1 U1731 ( .A(n2925), .B(DATAIN[15]), .S(n210), .Z(n3222) );
  MUX2_X1 U1732 ( .A(n2926), .B(DATAIN[16]), .S(n210), .Z(n3223) );
  MUX2_X1 U1733 ( .A(n2927), .B(DATAIN[17]), .S(n210), .Z(n3224) );
  MUX2_X1 U1734 ( .A(n2928), .B(DATAIN[18]), .S(n210), .Z(n3225) );
  MUX2_X1 U1735 ( .A(n2929), .B(DATAIN[19]), .S(n210), .Z(n3226) );
  MUX2_X1 U1736 ( .A(n2930), .B(DATAIN[20]), .S(n210), .Z(n3227) );
  MUX2_X1 U1737 ( .A(n2931), .B(DATAIN[21]), .S(n210), .Z(n3228) );
  MUX2_X1 U1738 ( .A(n2932), .B(DATAIN[22]), .S(n210), .Z(n3229) );
  MUX2_X1 U1739 ( .A(n2933), .B(DATAIN[23]), .S(n210), .Z(n3230) );
  MUX2_X1 U1740 ( .A(n2934), .B(DATAIN[24]), .S(n211), .Z(n3231) );
  MUX2_X1 U1741 ( .A(n2935), .B(DATAIN[25]), .S(n211), .Z(n3232) );
  MUX2_X1 U1742 ( .A(n2936), .B(DATAIN[26]), .S(n211), .Z(n3233) );
  MUX2_X1 U1743 ( .A(n2937), .B(DATAIN[27]), .S(n211), .Z(n3234) );
  MUX2_X1 U1744 ( .A(n2938), .B(DATAIN[28]), .S(n211), .Z(n3235) );
  MUX2_X1 U1745 ( .A(n2939), .B(DATAIN[29]), .S(n211), .Z(n3236) );
  MUX2_X1 U1746 ( .A(n2940), .B(DATAIN[30]), .S(n211), .Z(n3237) );
  MUX2_X1 U1747 ( .A(n2941), .B(DATAIN[31]), .S(n211), .Z(n3238) );
  MUX2_X1 U1748 ( .A(n1553), .B(DATAIN[0]), .S(n212), .Z(n4446) );
  MUX2_X1 U1749 ( .A(n1554), .B(DATAIN[1]), .S(n212), .Z(n4447) );
  MUX2_X1 U1750 ( .A(n1555), .B(DATAIN[2]), .S(n212), .Z(n4448) );
  MUX2_X1 U1751 ( .A(n1556), .B(DATAIN[3]), .S(n212), .Z(n4449) );
  MUX2_X1 U1752 ( .A(n1557), .B(DATAIN[4]), .S(n212), .Z(n4450) );
  MUX2_X1 U1753 ( .A(n1558), .B(DATAIN[5]), .S(n212), .Z(n4451) );
  MUX2_X1 U1754 ( .A(n1559), .B(DATAIN[6]), .S(n212), .Z(n4452) );
  MUX2_X1 U1755 ( .A(n1560), .B(DATAIN[7]), .S(n212), .Z(n4453) );
  MUX2_X1 U1756 ( .A(n1561), .B(DATAIN[8]), .S(n212), .Z(n4454) );
  MUX2_X1 U1757 ( .A(n1562), .B(DATAIN[9]), .S(n212), .Z(n4455) );
  MUX2_X1 U1758 ( .A(n1563), .B(DATAIN[10]), .S(n212), .Z(n4456) );
  MUX2_X1 U1759 ( .A(n1564), .B(DATAIN[11]), .S(n212), .Z(n4457) );
  MUX2_X1 U1760 ( .A(n1565), .B(DATAIN[12]), .S(n213), .Z(n4458) );
  MUX2_X1 U1761 ( .A(n1566), .B(DATAIN[13]), .S(n213), .Z(n4459) );
  MUX2_X1 U1762 ( .A(n1567), .B(DATAIN[14]), .S(n213), .Z(n4460) );
  MUX2_X1 U1763 ( .A(n1568), .B(DATAIN[15]), .S(n213), .Z(n4461) );
  MUX2_X1 U1764 ( .A(n1569), .B(DATAIN[16]), .S(n213), .Z(n4462) );
  MUX2_X1 U1765 ( .A(n1570), .B(DATAIN[17]), .S(n213), .Z(n4463) );
  MUX2_X1 U1766 ( .A(n1571), .B(DATAIN[18]), .S(n213), .Z(n4464) );
  MUX2_X1 U1767 ( .A(n1572), .B(DATAIN[19]), .S(n213), .Z(n4465) );
  MUX2_X1 U1768 ( .A(n1573), .B(DATAIN[20]), .S(n213), .Z(n4466) );
  MUX2_X1 U1769 ( .A(n1574), .B(DATAIN[21]), .S(n213), .Z(n4467) );
  MUX2_X1 U1770 ( .A(n1575), .B(DATAIN[22]), .S(n213), .Z(n4468) );
  MUX2_X1 U1771 ( .A(n1576), .B(DATAIN[23]), .S(n213), .Z(n4469) );
  MUX2_X1 U1772 ( .A(n1577), .B(DATAIN[24]), .S(n214), .Z(n4470) );
  MUX2_X1 U1773 ( .A(n1578), .B(DATAIN[25]), .S(n214), .Z(n4471) );
  MUX2_X1 U1774 ( .A(n1579), .B(DATAIN[26]), .S(n214), .Z(n4472) );
  MUX2_X1 U1775 ( .A(n1580), .B(DATAIN[27]), .S(n214), .Z(n4473) );
  MUX2_X1 U1776 ( .A(n1581), .B(DATAIN[28]), .S(n214), .Z(n4474) );
  MUX2_X1 U1777 ( .A(n1582), .B(DATAIN[29]), .S(n214), .Z(n4475) );
  MUX2_X1 U1778 ( .A(n1583), .B(DATAIN[30]), .S(n214), .Z(n4476) );
  MUX2_X1 U1779 ( .A(n1584), .B(DATAIN[31]), .S(n214), .Z(n4477) );
  MUX2_X1 U1780 ( .A(n1585), .B(DATAIN[0]), .S(n215), .Z(n4414) );
  MUX2_X1 U1781 ( .A(n1586), .B(DATAIN[1]), .S(n215), .Z(n4415) );
  MUX2_X1 U1782 ( .A(n1587), .B(DATAIN[2]), .S(n215), .Z(n4416) );
  MUX2_X1 U1783 ( .A(n1588), .B(DATAIN[3]), .S(n215), .Z(n4417) );
  MUX2_X1 U1784 ( .A(n1589), .B(DATAIN[4]), .S(n215), .Z(n4418) );
  MUX2_X1 U1785 ( .A(n1590), .B(DATAIN[5]), .S(n215), .Z(n4419) );
  MUX2_X1 U1786 ( .A(n1591), .B(DATAIN[6]), .S(n215), .Z(n4420) );
  MUX2_X1 U1787 ( .A(n1592), .B(DATAIN[7]), .S(n215), .Z(n4421) );
  MUX2_X1 U1788 ( .A(n1593), .B(DATAIN[8]), .S(n215), .Z(n4422) );
  MUX2_X1 U1789 ( .A(n1594), .B(DATAIN[9]), .S(n215), .Z(n4423) );
  MUX2_X1 U1790 ( .A(n1595), .B(DATAIN[10]), .S(n215), .Z(n4424) );
  MUX2_X1 U1791 ( .A(n1596), .B(DATAIN[11]), .S(n215), .Z(n4425) );
  MUX2_X1 U1792 ( .A(n1597), .B(DATAIN[12]), .S(n216), .Z(n4426) );
  MUX2_X1 U1793 ( .A(n1598), .B(DATAIN[13]), .S(n216), .Z(n4427) );
  MUX2_X1 U1794 ( .A(n1599), .B(DATAIN[14]), .S(n216), .Z(n4428) );
  MUX2_X1 U1795 ( .A(n1600), .B(DATAIN[15]), .S(n216), .Z(n4429) );
  MUX2_X1 U1796 ( .A(n1601), .B(DATAIN[16]), .S(n216), .Z(n4430) );
  MUX2_X1 U1797 ( .A(n1602), .B(DATAIN[17]), .S(n216), .Z(n4431) );
  MUX2_X1 U1798 ( .A(n1603), .B(DATAIN[18]), .S(n216), .Z(n4432) );
  MUX2_X1 U1799 ( .A(n1604), .B(DATAIN[19]), .S(n216), .Z(n4433) );
  MUX2_X1 U1800 ( .A(n1605), .B(DATAIN[20]), .S(n216), .Z(n4434) );
  MUX2_X1 U1801 ( .A(n1606), .B(DATAIN[21]), .S(n216), .Z(n4435) );
  MUX2_X1 U1802 ( .A(n1607), .B(DATAIN[22]), .S(n216), .Z(n4436) );
  MUX2_X1 U1803 ( .A(n1608), .B(DATAIN[23]), .S(n216), .Z(n4437) );
  MUX2_X1 U1804 ( .A(n1609), .B(DATAIN[24]), .S(n217), .Z(n4438) );
  MUX2_X1 U1805 ( .A(n1610), .B(DATAIN[25]), .S(n217), .Z(n4439) );
  MUX2_X1 U1806 ( .A(n1611), .B(DATAIN[26]), .S(n217), .Z(n4440) );
  MUX2_X1 U1807 ( .A(n1612), .B(DATAIN[27]), .S(n217), .Z(n4441) );
  MUX2_X1 U1808 ( .A(n1613), .B(DATAIN[28]), .S(n217), .Z(n4442) );
  MUX2_X1 U1809 ( .A(n1614), .B(DATAIN[29]), .S(n217), .Z(n4443) );
  MUX2_X1 U1810 ( .A(n1615), .B(DATAIN[30]), .S(n217), .Z(n4444) );
  MUX2_X1 U1811 ( .A(n1616), .B(DATAIN[31]), .S(n217), .Z(n4445) );
  MUX2_X1 U1812 ( .A(n3582), .B(DATAIN[0]), .S(n218), .Z(n3239) );
  MUX2_X1 U1813 ( .A(n3583), .B(DATAIN[1]), .S(n218), .Z(n3240) );
  MUX2_X1 U1814 ( .A(n3584), .B(DATAIN[2]), .S(n218), .Z(n3241) );
  MUX2_X1 U1815 ( .A(n3585), .B(DATAIN[3]), .S(n218), .Z(n3242) );
  MUX2_X1 U1816 ( .A(n3586), .B(DATAIN[4]), .S(n218), .Z(n3243) );
  MUX2_X1 U1817 ( .A(n3587), .B(DATAIN[5]), .S(n218), .Z(n3244) );
  MUX2_X1 U1818 ( .A(n3588), .B(DATAIN[6]), .S(n218), .Z(n3245) );
  MUX2_X1 U1819 ( .A(n3589), .B(DATAIN[7]), .S(n218), .Z(n3246) );
  MUX2_X1 U1820 ( .A(n3590), .B(DATAIN[8]), .S(n218), .Z(n3247) );
  MUX2_X1 U1821 ( .A(n3591), .B(DATAIN[9]), .S(n218), .Z(n3248) );
  MUX2_X1 U1822 ( .A(n3592), .B(DATAIN[10]), .S(n218), .Z(n3249) );
  MUX2_X1 U1823 ( .A(n3593), .B(DATAIN[11]), .S(n218), .Z(n3250) );
  MUX2_X1 U1824 ( .A(n3594), .B(DATAIN[12]), .S(n219), .Z(n3251) );
  MUX2_X1 U1825 ( .A(n3595), .B(DATAIN[13]), .S(n219), .Z(n3252) );
  MUX2_X1 U1826 ( .A(n3596), .B(DATAIN[14]), .S(n219), .Z(n3253) );
  MUX2_X1 U1827 ( .A(n3597), .B(DATAIN[15]), .S(n219), .Z(n3254) );
  MUX2_X1 U1828 ( .A(n3598), .B(DATAIN[16]), .S(n219), .Z(n3255) );
  MUX2_X1 U1829 ( .A(n3599), .B(DATAIN[17]), .S(n219), .Z(n3256) );
  MUX2_X1 U1830 ( .A(n3600), .B(DATAIN[18]), .S(n219), .Z(n3257) );
  MUX2_X1 U1831 ( .A(n3601), .B(DATAIN[19]), .S(n219), .Z(n3258) );
  MUX2_X1 U1832 ( .A(n3602), .B(DATAIN[20]), .S(n219), .Z(n3259) );
  MUX2_X1 U1833 ( .A(n3603), .B(DATAIN[21]), .S(n219), .Z(n3260) );
  MUX2_X1 U1834 ( .A(n3604), .B(DATAIN[22]), .S(n219), .Z(n3261) );
  MUX2_X1 U1835 ( .A(n3605), .B(DATAIN[23]), .S(n219), .Z(n3262) );
  MUX2_X1 U1836 ( .A(n3606), .B(DATAIN[24]), .S(n220), .Z(n3263) );
  MUX2_X1 U1837 ( .A(n3607), .B(DATAIN[25]), .S(n220), .Z(n3264) );
  MUX2_X1 U1838 ( .A(n3608), .B(DATAIN[26]), .S(n220), .Z(n3265) );
  MUX2_X1 U1839 ( .A(n3609), .B(DATAIN[27]), .S(n220), .Z(n3266) );
  MUX2_X1 U1840 ( .A(n3610), .B(DATAIN[28]), .S(n220), .Z(n3267) );
  MUX2_X1 U1841 ( .A(n3611), .B(DATAIN[29]), .S(n220), .Z(n3268) );
  MUX2_X1 U1842 ( .A(n3612), .B(DATAIN[30]), .S(n220), .Z(n3269) );
  MUX2_X1 U1843 ( .A(n3613), .B(DATAIN[31]), .S(n220), .Z(n3270) );
  MUX2_X1 U1844 ( .A(n3614), .B(DATAIN[0]), .S(n221), .Z(n3271) );
  MUX2_X1 U1845 ( .A(n3615), .B(DATAIN[1]), .S(n221), .Z(n3272) );
  MUX2_X1 U1846 ( .A(n3616), .B(DATAIN[2]), .S(n221), .Z(n3273) );
  MUX2_X1 U1847 ( .A(n3617), .B(DATAIN[3]), .S(n221), .Z(n3274) );
  MUX2_X1 U1848 ( .A(n3618), .B(DATAIN[4]), .S(n221), .Z(n3275) );
  MUX2_X1 U1849 ( .A(n3619), .B(DATAIN[5]), .S(n221), .Z(n3276) );
  MUX2_X1 U1850 ( .A(n3620), .B(DATAIN[6]), .S(n221), .Z(n3277) );
  MUX2_X1 U1851 ( .A(n3621), .B(DATAIN[7]), .S(n221), .Z(n3278) );
  MUX2_X1 U1852 ( .A(n3622), .B(DATAIN[8]), .S(n221), .Z(n3279) );
  MUX2_X1 U1853 ( .A(n3623), .B(DATAIN[9]), .S(n221), .Z(n3280) );
  MUX2_X1 U1854 ( .A(n3624), .B(DATAIN[10]), .S(n221), .Z(n3281) );
  MUX2_X1 U1855 ( .A(n3625), .B(DATAIN[11]), .S(n221), .Z(n3282) );
  MUX2_X1 U1856 ( .A(n3626), .B(DATAIN[12]), .S(n222), .Z(n3283) );
  MUX2_X1 U1857 ( .A(n3627), .B(DATAIN[13]), .S(n222), .Z(n3284) );
  MUX2_X1 U1858 ( .A(n3628), .B(DATAIN[14]), .S(n222), .Z(n3285) );
  MUX2_X1 U1859 ( .A(n3629), .B(DATAIN[15]), .S(n222), .Z(n3286) );
  MUX2_X1 U1860 ( .A(n3630), .B(DATAIN[16]), .S(n222), .Z(n3287) );
  MUX2_X1 U1861 ( .A(n3631), .B(DATAIN[17]), .S(n222), .Z(n3288) );
  MUX2_X1 U1862 ( .A(n3632), .B(DATAIN[18]), .S(n222), .Z(n3289) );
  MUX2_X1 U1863 ( .A(n3633), .B(DATAIN[19]), .S(n222), .Z(n3290) );
  MUX2_X1 U1864 ( .A(n3634), .B(DATAIN[20]), .S(n222), .Z(n3291) );
  MUX2_X1 U1865 ( .A(n3635), .B(DATAIN[21]), .S(n222), .Z(n3292) );
  MUX2_X1 U1866 ( .A(n3636), .B(DATAIN[22]), .S(n222), .Z(n3293) );
  MUX2_X1 U1867 ( .A(n3637), .B(DATAIN[23]), .S(n222), .Z(n3294) );
  MUX2_X1 U1868 ( .A(n3638), .B(DATAIN[24]), .S(n223), .Z(n3295) );
  MUX2_X1 U1869 ( .A(n3639), .B(DATAIN[25]), .S(n223), .Z(n3296) );
  MUX2_X1 U1870 ( .A(n3640), .B(DATAIN[26]), .S(n223), .Z(n3297) );
  MUX2_X1 U1871 ( .A(n3641), .B(DATAIN[27]), .S(n223), .Z(n3298) );
  MUX2_X1 U1872 ( .A(n3642), .B(DATAIN[28]), .S(n223), .Z(n3299) );
  MUX2_X1 U1873 ( .A(n3643), .B(DATAIN[29]), .S(n223), .Z(n3300) );
  MUX2_X1 U1874 ( .A(n3644), .B(DATAIN[30]), .S(n223), .Z(n3301) );
  MUX2_X1 U1875 ( .A(n3645), .B(DATAIN[31]), .S(n223), .Z(n3302) );
  MUX2_X1 U1876 ( .A(n1617), .B(DATAIN[0]), .S(n224), .Z(n4382) );
  MUX2_X1 U1877 ( .A(n1618), .B(DATAIN[1]), .S(n224), .Z(n4383) );
  MUX2_X1 U1878 ( .A(n1619), .B(DATAIN[2]), .S(n224), .Z(n4384) );
  MUX2_X1 U1879 ( .A(n1620), .B(DATAIN[3]), .S(n224), .Z(n4385) );
  MUX2_X1 U1880 ( .A(n1621), .B(DATAIN[4]), .S(n224), .Z(n4386) );
  MUX2_X1 U1881 ( .A(n1622), .B(DATAIN[5]), .S(n224), .Z(n4387) );
  MUX2_X1 U1882 ( .A(n1623), .B(DATAIN[6]), .S(n224), .Z(n4388) );
  MUX2_X1 U1883 ( .A(n1624), .B(DATAIN[7]), .S(n224), .Z(n4389) );
  MUX2_X1 U1884 ( .A(n1625), .B(DATAIN[8]), .S(n224), .Z(n4390) );
  MUX2_X1 U1885 ( .A(n1626), .B(DATAIN[9]), .S(n224), .Z(n4391) );
  MUX2_X1 U1886 ( .A(n1627), .B(DATAIN[10]), .S(n224), .Z(n4392) );
  MUX2_X1 U1887 ( .A(n1628), .B(DATAIN[11]), .S(n224), .Z(n4393) );
  MUX2_X1 U1888 ( .A(n1629), .B(DATAIN[12]), .S(n225), .Z(n4394) );
  MUX2_X1 U1889 ( .A(n1630), .B(DATAIN[13]), .S(n225), .Z(n4395) );
  MUX2_X1 U1890 ( .A(n1631), .B(DATAIN[14]), .S(n225), .Z(n4396) );
  MUX2_X1 U1891 ( .A(n1632), .B(DATAIN[15]), .S(n225), .Z(n4397) );
  MUX2_X1 U1892 ( .A(n1633), .B(DATAIN[16]), .S(n225), .Z(n4398) );
  MUX2_X1 U1893 ( .A(n1634), .B(DATAIN[17]), .S(n225), .Z(n4399) );
  MUX2_X1 U1894 ( .A(n1635), .B(DATAIN[18]), .S(n225), .Z(n4400) );
  MUX2_X1 U1895 ( .A(n1636), .B(DATAIN[19]), .S(n225), .Z(n4401) );
  MUX2_X1 U1896 ( .A(n1637), .B(DATAIN[20]), .S(n225), .Z(n4402) );
  MUX2_X1 U1897 ( .A(n1638), .B(DATAIN[21]), .S(n225), .Z(n4403) );
  MUX2_X1 U1898 ( .A(n1639), .B(DATAIN[22]), .S(n225), .Z(n4404) );
  MUX2_X1 U1899 ( .A(n1640), .B(DATAIN[23]), .S(n225), .Z(n4405) );
  MUX2_X1 U1900 ( .A(n1641), .B(DATAIN[24]), .S(n226), .Z(n4406) );
  MUX2_X1 U1901 ( .A(n1642), .B(DATAIN[25]), .S(n226), .Z(n4407) );
  MUX2_X1 U1902 ( .A(n1643), .B(DATAIN[26]), .S(n226), .Z(n4408) );
  MUX2_X1 U1903 ( .A(n1644), .B(DATAIN[27]), .S(n226), .Z(n4409) );
  MUX2_X1 U1904 ( .A(n1645), .B(DATAIN[28]), .S(n226), .Z(n4410) );
  MUX2_X1 U1905 ( .A(n1646), .B(DATAIN[29]), .S(n226), .Z(n4411) );
  MUX2_X1 U1906 ( .A(n1647), .B(DATAIN[30]), .S(n226), .Z(n4412) );
  MUX2_X1 U1907 ( .A(n1648), .B(DATAIN[31]), .S(n226), .Z(n4413) );
  MUX2_X1 U1908 ( .A(n1649), .B(DATAIN[0]), .S(n227), .Z(n4350) );
  MUX2_X1 U1909 ( .A(n1650), .B(DATAIN[1]), .S(n227), .Z(n4351) );
  MUX2_X1 U1910 ( .A(n1651), .B(DATAIN[2]), .S(n227), .Z(n4352) );
  MUX2_X1 U1911 ( .A(n1652), .B(DATAIN[3]), .S(n227), .Z(n4353) );
  MUX2_X1 U1912 ( .A(n1653), .B(DATAIN[4]), .S(n227), .Z(n4354) );
  MUX2_X1 U1913 ( .A(n1654), .B(DATAIN[5]), .S(n227), .Z(n4355) );
  MUX2_X1 U1914 ( .A(n1655), .B(DATAIN[6]), .S(n227), .Z(n4356) );
  MUX2_X1 U1915 ( .A(n1656), .B(DATAIN[7]), .S(n227), .Z(n4357) );
  MUX2_X1 U1916 ( .A(n1657), .B(DATAIN[8]), .S(n227), .Z(n4358) );
  MUX2_X1 U1917 ( .A(n1658), .B(DATAIN[9]), .S(n227), .Z(n4359) );
  MUX2_X1 U1918 ( .A(n1659), .B(DATAIN[10]), .S(n227), .Z(n4360) );
  MUX2_X1 U1919 ( .A(n1660), .B(DATAIN[11]), .S(n227), .Z(n4361) );
  MUX2_X1 U1920 ( .A(n1661), .B(DATAIN[12]), .S(n228), .Z(n4362) );
  MUX2_X1 U1921 ( .A(n1662), .B(DATAIN[13]), .S(n228), .Z(n4363) );
  MUX2_X1 U1922 ( .A(n1663), .B(DATAIN[14]), .S(n228), .Z(n4364) );
  MUX2_X1 U1923 ( .A(n1664), .B(DATAIN[15]), .S(n228), .Z(n4365) );
  MUX2_X1 U1924 ( .A(n1665), .B(DATAIN[16]), .S(n228), .Z(n4366) );
  MUX2_X1 U1925 ( .A(n1666), .B(DATAIN[17]), .S(n228), .Z(n4367) );
  MUX2_X1 U1926 ( .A(n1667), .B(DATAIN[18]), .S(n228), .Z(n4368) );
  MUX2_X1 U1927 ( .A(n1668), .B(DATAIN[19]), .S(n228), .Z(n4369) );
  MUX2_X1 U1928 ( .A(n1669), .B(DATAIN[20]), .S(n228), .Z(n4370) );
  MUX2_X1 U1929 ( .A(n1670), .B(DATAIN[21]), .S(n228), .Z(n4371) );
  MUX2_X1 U1930 ( .A(n1671), .B(DATAIN[22]), .S(n228), .Z(n4372) );
  MUX2_X1 U1931 ( .A(n1672), .B(DATAIN[23]), .S(n228), .Z(n4373) );
  MUX2_X1 U1932 ( .A(n1673), .B(DATAIN[24]), .S(n229), .Z(n4374) );
  MUX2_X1 U1933 ( .A(n1674), .B(DATAIN[25]), .S(n229), .Z(n4375) );
  MUX2_X1 U1934 ( .A(n1675), .B(DATAIN[26]), .S(n229), .Z(n4376) );
  MUX2_X1 U1935 ( .A(n1676), .B(DATAIN[27]), .S(n229), .Z(n4377) );
  MUX2_X1 U1936 ( .A(n1677), .B(DATAIN[28]), .S(n229), .Z(n4378) );
  MUX2_X1 U1937 ( .A(n1678), .B(DATAIN[29]), .S(n229), .Z(n4379) );
  MUX2_X1 U1938 ( .A(n1679), .B(DATAIN[30]), .S(n229), .Z(n4380) );
  MUX2_X1 U1939 ( .A(n1680), .B(DATAIN[31]), .S(n229), .Z(n4381) );
  INV_X1 U1940 ( .A(ADD_WR[4]), .ZN(n1809) );
  MUX2_X1 U1941 ( .A(n3678), .B(DATAIN[0]), .S(n230), .Z(n3303) );
  MUX2_X1 U1942 ( .A(n3679), .B(DATAIN[1]), .S(n230), .Z(n3304) );
  MUX2_X1 U1943 ( .A(n3680), .B(DATAIN[2]), .S(n230), .Z(n3305) );
  MUX2_X1 U1944 ( .A(n3681), .B(DATAIN[3]), .S(n230), .Z(n3306) );
  MUX2_X1 U1945 ( .A(n3682), .B(DATAIN[4]), .S(n230), .Z(n3307) );
  MUX2_X1 U1946 ( .A(n3683), .B(DATAIN[5]), .S(n230), .Z(n3308) );
  MUX2_X1 U1947 ( .A(n3684), .B(DATAIN[6]), .S(n230), .Z(n3309) );
  MUX2_X1 U1948 ( .A(n3685), .B(DATAIN[7]), .S(n230), .Z(n3310) );
  MUX2_X1 U1949 ( .A(n3686), .B(DATAIN[8]), .S(n230), .Z(n3311) );
  MUX2_X1 U1950 ( .A(n3687), .B(DATAIN[9]), .S(n230), .Z(n3312) );
  MUX2_X1 U1951 ( .A(n3688), .B(DATAIN[10]), .S(n230), .Z(n3313) );
  MUX2_X1 U1952 ( .A(n3689), .B(DATAIN[11]), .S(n230), .Z(n3314) );
  MUX2_X1 U1953 ( .A(n3690), .B(DATAIN[12]), .S(n231), .Z(n3315) );
  MUX2_X1 U1954 ( .A(n3691), .B(DATAIN[13]), .S(n231), .Z(n3316) );
  MUX2_X1 U1955 ( .A(n3692), .B(DATAIN[14]), .S(n231), .Z(n3317) );
  MUX2_X1 U1956 ( .A(n3693), .B(DATAIN[15]), .S(n231), .Z(n3318) );
  MUX2_X1 U1957 ( .A(n3694), .B(DATAIN[16]), .S(n231), .Z(n3319) );
  MUX2_X1 U1958 ( .A(n3695), .B(DATAIN[17]), .S(n231), .Z(n3320) );
  MUX2_X1 U1959 ( .A(n3696), .B(DATAIN[18]), .S(n231), .Z(n3321) );
  MUX2_X1 U1960 ( .A(n3697), .B(DATAIN[19]), .S(n231), .Z(n3322) );
  MUX2_X1 U1961 ( .A(n3698), .B(DATAIN[20]), .S(n231), .Z(n3323) );
  MUX2_X1 U1962 ( .A(n3699), .B(DATAIN[21]), .S(n231), .Z(n3324) );
  MUX2_X1 U1963 ( .A(n3700), .B(DATAIN[22]), .S(n231), .Z(n3325) );
  MUX2_X1 U1964 ( .A(n3701), .B(DATAIN[23]), .S(n231), .Z(n3326) );
  MUX2_X1 U1965 ( .A(n3702), .B(DATAIN[24]), .S(n232), .Z(n3327) );
  MUX2_X1 U1966 ( .A(n3703), .B(DATAIN[25]), .S(n232), .Z(n3328) );
  MUX2_X1 U1967 ( .A(n3704), .B(DATAIN[26]), .S(n232), .Z(n3329) );
  MUX2_X1 U1968 ( .A(n3705), .B(DATAIN[27]), .S(n232), .Z(n3330) );
  MUX2_X1 U1969 ( .A(n3706), .B(DATAIN[28]), .S(n232), .Z(n3331) );
  MUX2_X1 U1970 ( .A(n3707), .B(DATAIN[29]), .S(n232), .Z(n3332) );
  MUX2_X1 U1971 ( .A(n3708), .B(DATAIN[30]), .S(n232), .Z(n3333) );
  MUX2_X1 U1972 ( .A(n3709), .B(DATAIN[31]), .S(n232), .Z(n3334) );
  MUX2_X1 U1973 ( .A(n3710), .B(DATAIN[0]), .S(n233), .Z(n3335) );
  MUX2_X1 U1974 ( .A(n3711), .B(DATAIN[1]), .S(n233), .Z(n3336) );
  MUX2_X1 U1975 ( .A(n3712), .B(DATAIN[2]), .S(n233), .Z(n3337) );
  MUX2_X1 U1976 ( .A(n3713), .B(DATAIN[3]), .S(n233), .Z(n3338) );
  MUX2_X1 U1977 ( .A(n3714), .B(DATAIN[4]), .S(n233), .Z(n3339) );
  MUX2_X1 U1978 ( .A(n3715), .B(DATAIN[5]), .S(n233), .Z(n3340) );
  MUX2_X1 U1979 ( .A(n3716), .B(DATAIN[6]), .S(n233), .Z(n3341) );
  MUX2_X1 U1980 ( .A(n3717), .B(DATAIN[7]), .S(n233), .Z(n3342) );
  MUX2_X1 U1981 ( .A(n3718), .B(DATAIN[8]), .S(n233), .Z(n3343) );
  MUX2_X1 U1982 ( .A(n3719), .B(DATAIN[9]), .S(n233), .Z(n3344) );
  MUX2_X1 U1983 ( .A(n3720), .B(DATAIN[10]), .S(n233), .Z(n3345) );
  MUX2_X1 U1984 ( .A(n3721), .B(DATAIN[11]), .S(n233), .Z(n3346) );
  MUX2_X1 U1985 ( .A(n3722), .B(DATAIN[12]), .S(n234), .Z(n3347) );
  MUX2_X1 U1986 ( .A(n3723), .B(DATAIN[13]), .S(n234), .Z(n3348) );
  MUX2_X1 U1987 ( .A(n3724), .B(DATAIN[14]), .S(n234), .Z(n3349) );
  MUX2_X1 U1988 ( .A(n3725), .B(DATAIN[15]), .S(n234), .Z(n3350) );
  MUX2_X1 U1989 ( .A(n3726), .B(DATAIN[16]), .S(n234), .Z(n3351) );
  MUX2_X1 U1990 ( .A(n3727), .B(DATAIN[17]), .S(n234), .Z(n3352) );
  MUX2_X1 U1991 ( .A(n3728), .B(DATAIN[18]), .S(n234), .Z(n3353) );
  MUX2_X1 U1992 ( .A(n3729), .B(DATAIN[19]), .S(n234), .Z(n3354) );
  MUX2_X1 U1993 ( .A(n3730), .B(DATAIN[20]), .S(n234), .Z(n3355) );
  MUX2_X1 U1994 ( .A(n3731), .B(DATAIN[21]), .S(n234), .Z(n3356) );
  MUX2_X1 U1995 ( .A(n3732), .B(DATAIN[22]), .S(n234), .Z(n3357) );
  MUX2_X1 U1996 ( .A(n3733), .B(DATAIN[23]), .S(n234), .Z(n3358) );
  MUX2_X1 U1997 ( .A(n3734), .B(DATAIN[24]), .S(n235), .Z(n3359) );
  MUX2_X1 U1998 ( .A(n3735), .B(DATAIN[25]), .S(n235), .Z(n3360) );
  MUX2_X1 U1999 ( .A(n3736), .B(DATAIN[26]), .S(n235), .Z(n3361) );
  MUX2_X1 U2000 ( .A(n3737), .B(DATAIN[27]), .S(n235), .Z(n3362) );
  MUX2_X1 U2001 ( .A(n3738), .B(DATAIN[28]), .S(n235), .Z(n3363) );
  MUX2_X1 U2002 ( .A(n3739), .B(DATAIN[29]), .S(n235), .Z(n3364) );
  MUX2_X1 U2003 ( .A(n3740), .B(DATAIN[30]), .S(n235), .Z(n3365) );
  MUX2_X1 U2004 ( .A(n3741), .B(DATAIN[31]), .S(n235), .Z(n3366) );
  MUX2_X1 U2005 ( .A(n1681), .B(DATAIN[0]), .S(n236), .Z(n4222) );
  MUX2_X1 U2006 ( .A(n1682), .B(DATAIN[1]), .S(n236), .Z(n4223) );
  MUX2_X1 U2007 ( .A(n1683), .B(DATAIN[2]), .S(n236), .Z(n4224) );
  MUX2_X1 U2008 ( .A(n1684), .B(DATAIN[3]), .S(n236), .Z(n4225) );
  MUX2_X1 U2009 ( .A(n1685), .B(DATAIN[4]), .S(n236), .Z(n4226) );
  MUX2_X1 U2010 ( .A(n1686), .B(DATAIN[5]), .S(n236), .Z(n4227) );
  MUX2_X1 U2011 ( .A(n1687), .B(DATAIN[6]), .S(n236), .Z(n4228) );
  MUX2_X1 U2012 ( .A(n1688), .B(DATAIN[7]), .S(n236), .Z(n4229) );
  MUX2_X1 U2013 ( .A(n1689), .B(DATAIN[8]), .S(n236), .Z(n4230) );
  MUX2_X1 U2014 ( .A(n1690), .B(DATAIN[9]), .S(n236), .Z(n4231) );
  MUX2_X1 U2015 ( .A(n1691), .B(DATAIN[10]), .S(n236), .Z(n4232) );
  MUX2_X1 U2016 ( .A(n1692), .B(DATAIN[11]), .S(n236), .Z(n4233) );
  MUX2_X1 U2017 ( .A(n1693), .B(DATAIN[12]), .S(n237), .Z(n4234) );
  MUX2_X1 U2018 ( .A(n1694), .B(DATAIN[13]), .S(n237), .Z(n4235) );
  MUX2_X1 U2019 ( .A(n1695), .B(DATAIN[14]), .S(n237), .Z(n4236) );
  MUX2_X1 U2020 ( .A(n1696), .B(DATAIN[15]), .S(n237), .Z(n4237) );
  MUX2_X1 U2021 ( .A(n1697), .B(DATAIN[16]), .S(n237), .Z(n4238) );
  MUX2_X1 U2022 ( .A(n1698), .B(DATAIN[17]), .S(n237), .Z(n4239) );
  MUX2_X1 U2023 ( .A(n1699), .B(DATAIN[18]), .S(n237), .Z(n4240) );
  MUX2_X1 U2024 ( .A(n1700), .B(DATAIN[19]), .S(n237), .Z(n4241) );
  MUX2_X1 U2025 ( .A(n1701), .B(DATAIN[20]), .S(n237), .Z(n4242) );
  MUX2_X1 U2026 ( .A(n1702), .B(DATAIN[21]), .S(n237), .Z(n4243) );
  MUX2_X1 U2027 ( .A(n1703), .B(DATAIN[22]), .S(n237), .Z(n4244) );
  MUX2_X1 U2028 ( .A(n1704), .B(DATAIN[23]), .S(n237), .Z(n4245) );
  MUX2_X1 U2029 ( .A(n1705), .B(DATAIN[24]), .S(n238), .Z(n4246) );
  MUX2_X1 U2030 ( .A(n1706), .B(DATAIN[25]), .S(n238), .Z(n4247) );
  MUX2_X1 U2031 ( .A(n1707), .B(DATAIN[26]), .S(n238), .Z(n4248) );
  MUX2_X1 U2032 ( .A(n1708), .B(DATAIN[27]), .S(n238), .Z(n4249) );
  MUX2_X1 U2033 ( .A(n1709), .B(DATAIN[28]), .S(n238), .Z(n4250) );
  MUX2_X1 U2034 ( .A(n1710), .B(DATAIN[29]), .S(n238), .Z(n4251) );
  MUX2_X1 U2035 ( .A(n1711), .B(DATAIN[30]), .S(n238), .Z(n4252) );
  MUX2_X1 U2036 ( .A(n1712), .B(DATAIN[31]), .S(n238), .Z(n4253) );
  MUX2_X1 U2037 ( .A(n1713), .B(DATAIN[0]), .S(n239), .Z(n4190) );
  MUX2_X1 U2038 ( .A(n1714), .B(DATAIN[1]), .S(n239), .Z(n4191) );
  MUX2_X1 U2039 ( .A(n1715), .B(DATAIN[2]), .S(n239), .Z(n4192) );
  MUX2_X1 U2040 ( .A(n1716), .B(DATAIN[3]), .S(n239), .Z(n4193) );
  MUX2_X1 U2041 ( .A(n1717), .B(DATAIN[4]), .S(n239), .Z(n4194) );
  MUX2_X1 U2042 ( .A(n1718), .B(DATAIN[5]), .S(n239), .Z(n4195) );
  MUX2_X1 U2043 ( .A(n1719), .B(DATAIN[6]), .S(n239), .Z(n4196) );
  MUX2_X1 U2044 ( .A(n1720), .B(DATAIN[7]), .S(n239), .Z(n4197) );
  MUX2_X1 U2045 ( .A(n1721), .B(DATAIN[8]), .S(n239), .Z(n4198) );
  MUX2_X1 U2046 ( .A(n1722), .B(DATAIN[9]), .S(n239), .Z(n4199) );
  MUX2_X1 U2047 ( .A(n1723), .B(DATAIN[10]), .S(n239), .Z(n4200) );
  MUX2_X1 U2048 ( .A(n1724), .B(DATAIN[11]), .S(n239), .Z(n4201) );
  MUX2_X1 U2049 ( .A(n1725), .B(DATAIN[12]), .S(n240), .Z(n4202) );
  MUX2_X1 U2050 ( .A(n1726), .B(DATAIN[13]), .S(n240), .Z(n4203) );
  MUX2_X1 U2051 ( .A(n1727), .B(DATAIN[14]), .S(n240), .Z(n4204) );
  MUX2_X1 U2052 ( .A(n1728), .B(DATAIN[15]), .S(n240), .Z(n4205) );
  MUX2_X1 U2053 ( .A(n1729), .B(DATAIN[16]), .S(n240), .Z(n4206) );
  MUX2_X1 U2054 ( .A(n1730), .B(DATAIN[17]), .S(n240), .Z(n4207) );
  MUX2_X1 U2055 ( .A(n1731), .B(DATAIN[18]), .S(n240), .Z(n4208) );
  MUX2_X1 U2056 ( .A(n1732), .B(DATAIN[19]), .S(n240), .Z(n4209) );
  MUX2_X1 U2057 ( .A(n1733), .B(DATAIN[20]), .S(n240), .Z(n4210) );
  MUX2_X1 U2058 ( .A(n1734), .B(DATAIN[21]), .S(n240), .Z(n4211) );
  MUX2_X1 U2059 ( .A(n1735), .B(DATAIN[22]), .S(n240), .Z(n4212) );
  MUX2_X1 U2060 ( .A(n1736), .B(DATAIN[23]), .S(n240), .Z(n4213) );
  MUX2_X1 U2061 ( .A(n1737), .B(DATAIN[24]), .S(n241), .Z(n4214) );
  MUX2_X1 U2062 ( .A(n1738), .B(DATAIN[25]), .S(n241), .Z(n4215) );
  MUX2_X1 U2063 ( .A(n1739), .B(DATAIN[26]), .S(n241), .Z(n4216) );
  MUX2_X1 U2064 ( .A(n1740), .B(DATAIN[27]), .S(n241), .Z(n4217) );
  MUX2_X1 U2065 ( .A(n1741), .B(DATAIN[28]), .S(n241), .Z(n4218) );
  MUX2_X1 U2066 ( .A(n1742), .B(DATAIN[29]), .S(n241), .Z(n4219) );
  MUX2_X1 U2067 ( .A(n1743), .B(DATAIN[30]), .S(n241), .Z(n4220) );
  MUX2_X1 U2068 ( .A(n1744), .B(DATAIN[31]), .S(n241), .Z(n4221) );
  MUX2_X1 U2069 ( .A(n3806), .B(DATAIN[0]), .S(n242), .Z(n3367) );
  MUX2_X1 U2070 ( .A(n3807), .B(DATAIN[1]), .S(n242), .Z(n3368) );
  MUX2_X1 U2071 ( .A(n3808), .B(DATAIN[2]), .S(n242), .Z(n3369) );
  MUX2_X1 U2072 ( .A(n3809), .B(DATAIN[3]), .S(n242), .Z(n3370) );
  MUX2_X1 U2073 ( .A(n3810), .B(DATAIN[4]), .S(n242), .Z(n3371) );
  MUX2_X1 U2074 ( .A(n3811), .B(DATAIN[5]), .S(n242), .Z(n3372) );
  MUX2_X1 U2075 ( .A(n3812), .B(DATAIN[6]), .S(n242), .Z(n3373) );
  MUX2_X1 U2076 ( .A(n3813), .B(DATAIN[7]), .S(n242), .Z(n3374) );
  MUX2_X1 U2077 ( .A(n3814), .B(DATAIN[8]), .S(n242), .Z(n3375) );
  MUX2_X1 U2078 ( .A(n3815), .B(DATAIN[9]), .S(n242), .Z(n3376) );
  MUX2_X1 U2079 ( .A(n3816), .B(DATAIN[10]), .S(n242), .Z(n3377) );
  MUX2_X1 U2080 ( .A(n3817), .B(DATAIN[11]), .S(n242), .Z(n3378) );
  MUX2_X1 U2081 ( .A(n3818), .B(DATAIN[12]), .S(n243), .Z(n3379) );
  MUX2_X1 U2082 ( .A(n3819), .B(DATAIN[13]), .S(n243), .Z(n3380) );
  MUX2_X1 U2083 ( .A(n3820), .B(DATAIN[14]), .S(n243), .Z(n3381) );
  MUX2_X1 U2084 ( .A(n3821), .B(DATAIN[15]), .S(n243), .Z(n3382) );
  MUX2_X1 U2085 ( .A(n3822), .B(DATAIN[16]), .S(n243), .Z(n3383) );
  MUX2_X1 U2086 ( .A(n3823), .B(DATAIN[17]), .S(n243), .Z(n3384) );
  MUX2_X1 U2087 ( .A(n3824), .B(DATAIN[18]), .S(n243), .Z(n3385) );
  MUX2_X1 U2088 ( .A(n3825), .B(DATAIN[19]), .S(n243), .Z(n3386) );
  MUX2_X1 U2089 ( .A(n3826), .B(DATAIN[20]), .S(n243), .Z(n3387) );
  MUX2_X1 U2090 ( .A(n3827), .B(DATAIN[21]), .S(n243), .Z(n3388) );
  MUX2_X1 U2091 ( .A(n3828), .B(DATAIN[22]), .S(n243), .Z(n3389) );
  MUX2_X1 U2092 ( .A(n3829), .B(DATAIN[23]), .S(n243), .Z(n3390) );
  MUX2_X1 U2093 ( .A(n3830), .B(DATAIN[24]), .S(n244), .Z(n3391) );
  MUX2_X1 U2094 ( .A(n3831), .B(DATAIN[25]), .S(n244), .Z(n3392) );
  MUX2_X1 U2095 ( .A(n3832), .B(DATAIN[26]), .S(n244), .Z(n3393) );
  MUX2_X1 U2096 ( .A(n3833), .B(DATAIN[27]), .S(n244), .Z(n3394) );
  MUX2_X1 U2097 ( .A(n3834), .B(DATAIN[28]), .S(n244), .Z(n3395) );
  MUX2_X1 U2098 ( .A(n3835), .B(DATAIN[29]), .S(n244), .Z(n3396) );
  MUX2_X1 U2099 ( .A(n3836), .B(DATAIN[30]), .S(n244), .Z(n3397) );
  MUX2_X1 U2100 ( .A(n3837), .B(DATAIN[31]), .S(n244), .Z(n3398) );
  MUX2_X1 U2101 ( .A(n3838), .B(DATAIN[0]), .S(n245), .Z(n3399) );
  MUX2_X1 U2102 ( .A(n3839), .B(DATAIN[1]), .S(n245), .Z(n3400) );
  MUX2_X1 U2103 ( .A(n3840), .B(DATAIN[2]), .S(n245), .Z(n3401) );
  MUX2_X1 U2104 ( .A(n3841), .B(DATAIN[3]), .S(n245), .Z(n3402) );
  MUX2_X1 U2105 ( .A(n3842), .B(DATAIN[4]), .S(n245), .Z(n3403) );
  MUX2_X1 U2106 ( .A(n3843), .B(DATAIN[5]), .S(n245), .Z(n3404) );
  MUX2_X1 U2107 ( .A(n3844), .B(DATAIN[6]), .S(n245), .Z(n3405) );
  MUX2_X1 U2108 ( .A(n3845), .B(DATAIN[7]), .S(n245), .Z(n3406) );
  MUX2_X1 U2109 ( .A(n3846), .B(DATAIN[8]), .S(n245), .Z(n3407) );
  MUX2_X1 U2110 ( .A(n3847), .B(DATAIN[9]), .S(n245), .Z(n3408) );
  MUX2_X1 U2111 ( .A(n3848), .B(DATAIN[10]), .S(n245), .Z(n3409) );
  MUX2_X1 U2112 ( .A(n3849), .B(DATAIN[11]), .S(n245), .Z(n3410) );
  MUX2_X1 U2113 ( .A(n3850), .B(DATAIN[12]), .S(n246), .Z(n3411) );
  MUX2_X1 U2114 ( .A(n3851), .B(DATAIN[13]), .S(n246), .Z(n3412) );
  MUX2_X1 U2115 ( .A(n3852), .B(DATAIN[14]), .S(n246), .Z(n3413) );
  MUX2_X1 U2116 ( .A(n3853), .B(DATAIN[15]), .S(n246), .Z(n3414) );
  MUX2_X1 U2117 ( .A(n3854), .B(DATAIN[16]), .S(n246), .Z(n3415) );
  MUX2_X1 U2118 ( .A(n3855), .B(DATAIN[17]), .S(n246), .Z(n3416) );
  MUX2_X1 U2119 ( .A(n3856), .B(DATAIN[18]), .S(n246), .Z(n3417) );
  MUX2_X1 U2120 ( .A(n3857), .B(DATAIN[19]), .S(n246), .Z(n3418) );
  MUX2_X1 U2121 ( .A(n3858), .B(DATAIN[20]), .S(n246), .Z(n3419) );
  MUX2_X1 U2122 ( .A(n3859), .B(DATAIN[21]), .S(n246), .Z(n3420) );
  MUX2_X1 U2123 ( .A(n3860), .B(DATAIN[22]), .S(n246), .Z(n3421) );
  MUX2_X1 U2124 ( .A(n3861), .B(DATAIN[23]), .S(n246), .Z(n3422) );
  MUX2_X1 U2125 ( .A(n3862), .B(DATAIN[24]), .S(n247), .Z(n3423) );
  MUX2_X1 U2126 ( .A(n3863), .B(DATAIN[25]), .S(n247), .Z(n3424) );
  MUX2_X1 U2127 ( .A(n3864), .B(DATAIN[26]), .S(n247), .Z(n3425) );
  MUX2_X1 U2128 ( .A(n3865), .B(DATAIN[27]), .S(n247), .Z(n3426) );
  MUX2_X1 U2129 ( .A(n3866), .B(DATAIN[28]), .S(n247), .Z(n3427) );
  MUX2_X1 U2130 ( .A(n3867), .B(DATAIN[29]), .S(n247), .Z(n3428) );
  MUX2_X1 U2131 ( .A(n3868), .B(DATAIN[30]), .S(n247), .Z(n3429) );
  MUX2_X1 U2132 ( .A(n3869), .B(DATAIN[31]), .S(n247), .Z(n3430) );
  MUX2_X1 U2133 ( .A(n1745), .B(DATAIN[0]), .S(n248), .Z(n4158) );
  MUX2_X1 U2134 ( .A(n1746), .B(DATAIN[1]), .S(n248), .Z(n4159) );
  MUX2_X1 U2135 ( .A(n1747), .B(DATAIN[2]), .S(n248), .Z(n4160) );
  MUX2_X1 U2136 ( .A(n1748), .B(DATAIN[3]), .S(n248), .Z(n4161) );
  MUX2_X1 U2137 ( .A(n1749), .B(DATAIN[4]), .S(n248), .Z(n4162) );
  MUX2_X1 U2138 ( .A(n1750), .B(DATAIN[5]), .S(n248), .Z(n4163) );
  MUX2_X1 U2139 ( .A(n1751), .B(DATAIN[6]), .S(n248), .Z(n4164) );
  MUX2_X1 U2140 ( .A(n1752), .B(DATAIN[7]), .S(n248), .Z(n4165) );
  MUX2_X1 U2141 ( .A(n1753), .B(DATAIN[8]), .S(n248), .Z(n4166) );
  MUX2_X1 U2142 ( .A(n1754), .B(DATAIN[9]), .S(n248), .Z(n4167) );
  MUX2_X1 U2143 ( .A(n1755), .B(DATAIN[10]), .S(n248), .Z(n4168) );
  MUX2_X1 U2144 ( .A(n1756), .B(DATAIN[11]), .S(n248), .Z(n4169) );
  MUX2_X1 U2145 ( .A(n1757), .B(DATAIN[12]), .S(n249), .Z(n4170) );
  MUX2_X1 U2146 ( .A(n1758), .B(DATAIN[13]), .S(n249), .Z(n4171) );
  MUX2_X1 U2147 ( .A(n1759), .B(DATAIN[14]), .S(n249), .Z(n4172) );
  MUX2_X1 U2148 ( .A(n1760), .B(DATAIN[15]), .S(n249), .Z(n4173) );
  MUX2_X1 U2149 ( .A(n1761), .B(DATAIN[16]), .S(n249), .Z(n4174) );
  MUX2_X1 U2150 ( .A(n1762), .B(DATAIN[17]), .S(n249), .Z(n4175) );
  MUX2_X1 U2151 ( .A(n1763), .B(DATAIN[18]), .S(n249), .Z(n4176) );
  MUX2_X1 U2152 ( .A(n1764), .B(DATAIN[19]), .S(n249), .Z(n4177) );
  MUX2_X1 U2153 ( .A(n1765), .B(DATAIN[20]), .S(n249), .Z(n4178) );
  MUX2_X1 U2154 ( .A(n1766), .B(DATAIN[21]), .S(n249), .Z(n4179) );
  MUX2_X1 U2155 ( .A(n1767), .B(DATAIN[22]), .S(n249), .Z(n4180) );
  MUX2_X1 U2156 ( .A(n1768), .B(DATAIN[23]), .S(n249), .Z(n4181) );
  MUX2_X1 U2157 ( .A(n1769), .B(DATAIN[24]), .S(n250), .Z(n4182) );
  MUX2_X1 U2158 ( .A(n1770), .B(DATAIN[25]), .S(n250), .Z(n4183) );
  MUX2_X1 U2159 ( .A(n1771), .B(DATAIN[26]), .S(n250), .Z(n4184) );
  MUX2_X1 U2160 ( .A(n1772), .B(DATAIN[27]), .S(n250), .Z(n4185) );
  MUX2_X1 U2161 ( .A(n1773), .B(DATAIN[28]), .S(n250), .Z(n4186) );
  MUX2_X1 U2162 ( .A(n1774), .B(DATAIN[29]), .S(n250), .Z(n4187) );
  MUX2_X1 U2163 ( .A(n1775), .B(DATAIN[30]), .S(n250), .Z(n4188) );
  MUX2_X1 U2164 ( .A(n1776), .B(DATAIN[31]), .S(n250), .Z(n4189) );
  MUX2_X1 U2165 ( .A(n1777), .B(DATAIN[0]), .S(n251), .Z(n4126) );
  MUX2_X1 U2166 ( .A(n1778), .B(DATAIN[1]), .S(n251), .Z(n4127) );
  MUX2_X1 U2167 ( .A(n1779), .B(DATAIN[2]), .S(n251), .Z(n4128) );
  MUX2_X1 U2168 ( .A(n1780), .B(DATAIN[3]), .S(n251), .Z(n4129) );
  MUX2_X1 U2169 ( .A(n1781), .B(DATAIN[4]), .S(n251), .Z(n4130) );
  MUX2_X1 U2170 ( .A(n1782), .B(DATAIN[5]), .S(n251), .Z(n4131) );
  MUX2_X1 U2171 ( .A(n1783), .B(DATAIN[6]), .S(n251), .Z(n4132) );
  MUX2_X1 U2172 ( .A(n1784), .B(DATAIN[7]), .S(n251), .Z(n4133) );
  MUX2_X1 U2173 ( .A(n1785), .B(DATAIN[8]), .S(n251), .Z(n4134) );
  MUX2_X1 U2174 ( .A(n1786), .B(DATAIN[9]), .S(n251), .Z(n4135) );
  MUX2_X1 U2175 ( .A(n1787), .B(DATAIN[10]), .S(n251), .Z(n4136) );
  MUX2_X1 U2176 ( .A(n1788), .B(DATAIN[11]), .S(n251), .Z(n4137) );
  MUX2_X1 U2177 ( .A(n1789), .B(DATAIN[12]), .S(n252), .Z(n4138) );
  MUX2_X1 U2178 ( .A(n1790), .B(DATAIN[13]), .S(n252), .Z(n4139) );
  MUX2_X1 U2179 ( .A(n1791), .B(DATAIN[14]), .S(n252), .Z(n4140) );
  MUX2_X1 U2180 ( .A(n1792), .B(DATAIN[15]), .S(n252), .Z(n4141) );
  MUX2_X1 U2181 ( .A(n1793), .B(DATAIN[16]), .S(n252), .Z(n4142) );
  MUX2_X1 U2182 ( .A(n1794), .B(DATAIN[17]), .S(n252), .Z(n4143) );
  MUX2_X1 U2183 ( .A(n1795), .B(DATAIN[18]), .S(n252), .Z(n4144) );
  MUX2_X1 U2184 ( .A(n1796), .B(DATAIN[19]), .S(n252), .Z(n4145) );
  MUX2_X1 U2185 ( .A(n1797), .B(DATAIN[20]), .S(n252), .Z(n4146) );
  MUX2_X1 U2186 ( .A(n1798), .B(DATAIN[21]), .S(n252), .Z(n4147) );
  MUX2_X1 U2187 ( .A(n1799), .B(DATAIN[22]), .S(n252), .Z(n4148) );
  MUX2_X1 U2188 ( .A(n1800), .B(DATAIN[23]), .S(n252), .Z(n4149) );
  MUX2_X1 U2189 ( .A(n1801), .B(DATAIN[24]), .S(n253), .Z(n4150) );
  MUX2_X1 U2190 ( .A(n1802), .B(DATAIN[25]), .S(n253), .Z(n4151) );
  MUX2_X1 U2191 ( .A(n1803), .B(DATAIN[26]), .S(n253), .Z(n4152) );
  MUX2_X1 U2192 ( .A(n1804), .B(DATAIN[27]), .S(n253), .Z(n4153) );
  MUX2_X1 U2193 ( .A(n1805), .B(DATAIN[28]), .S(n253), .Z(n4154) );
  MUX2_X1 U2194 ( .A(n1806), .B(DATAIN[29]), .S(n253), .Z(n4155) );
  MUX2_X1 U2195 ( .A(n1807), .B(DATAIN[30]), .S(n253), .Z(n4156) );
  MUX2_X1 U2196 ( .A(n1808), .B(DATAIN[31]), .S(n253), .Z(n4157) );
  MUX2_X1 U2197 ( .A(n3934), .B(DATAIN[0]), .S(n254), .Z(n3431) );
  MUX2_X1 U2198 ( .A(n3935), .B(DATAIN[1]), .S(n254), .Z(n3432) );
  MUX2_X1 U2199 ( .A(n3936), .B(DATAIN[2]), .S(n254), .Z(n3433) );
  MUX2_X1 U2200 ( .A(n3937), .B(DATAIN[3]), .S(n254), .Z(n3434) );
  MUX2_X1 U2201 ( .A(n3938), .B(DATAIN[4]), .S(n254), .Z(n3435) );
  MUX2_X1 U2202 ( .A(n3939), .B(DATAIN[5]), .S(n254), .Z(n3436) );
  MUX2_X1 U2203 ( .A(n3940), .B(DATAIN[6]), .S(n254), .Z(n3437) );
  MUX2_X1 U2204 ( .A(n3941), .B(DATAIN[7]), .S(n254), .Z(n3438) );
  MUX2_X1 U2205 ( .A(n3942), .B(DATAIN[8]), .S(n254), .Z(n3439) );
  MUX2_X1 U2206 ( .A(n3943), .B(DATAIN[9]), .S(n254), .Z(n3440) );
  MUX2_X1 U2207 ( .A(n3944), .B(DATAIN[10]), .S(n254), .Z(n3441) );
  MUX2_X1 U2208 ( .A(n3945), .B(DATAIN[11]), .S(n254), .Z(n3442) );
  MUX2_X1 U2209 ( .A(n3946), .B(DATAIN[12]), .S(n255), .Z(n3443) );
  MUX2_X1 U2210 ( .A(n3947), .B(DATAIN[13]), .S(n255), .Z(n3444) );
  MUX2_X1 U2211 ( .A(n3948), .B(DATAIN[14]), .S(n255), .Z(n3445) );
  MUX2_X1 U2212 ( .A(n3949), .B(DATAIN[15]), .S(n255), .Z(n3446) );
  MUX2_X1 U2213 ( .A(n3950), .B(DATAIN[16]), .S(n255), .Z(n3447) );
  MUX2_X1 U2214 ( .A(n3951), .B(DATAIN[17]), .S(n255), .Z(n3448) );
  MUX2_X1 U2215 ( .A(n3952), .B(DATAIN[18]), .S(n255), .Z(n3449) );
  MUX2_X1 U2216 ( .A(n3953), .B(DATAIN[19]), .S(n255), .Z(n3450) );
  MUX2_X1 U2217 ( .A(n3954), .B(DATAIN[20]), .S(n255), .Z(n3451) );
  MUX2_X1 U2218 ( .A(n3955), .B(DATAIN[21]), .S(n255), .Z(n3452) );
  MUX2_X1 U2219 ( .A(n3956), .B(DATAIN[22]), .S(n255), .Z(n3453) );
  MUX2_X1 U2220 ( .A(n3957), .B(DATAIN[23]), .S(n255), .Z(n3454) );
  MUX2_X1 U2221 ( .A(n3958), .B(DATAIN[24]), .S(n256), .Z(n3455) );
  MUX2_X1 U2222 ( .A(n3959), .B(DATAIN[25]), .S(n256), .Z(n3456) );
  MUX2_X1 U2223 ( .A(n3960), .B(DATAIN[26]), .S(n256), .Z(n3457) );
  MUX2_X1 U2224 ( .A(n3961), .B(DATAIN[27]), .S(n256), .Z(n3458) );
  MUX2_X1 U2225 ( .A(n3962), .B(DATAIN[28]), .S(n256), .Z(n3459) );
  MUX2_X1 U2226 ( .A(n3963), .B(DATAIN[29]), .S(n256), .Z(n3460) );
  MUX2_X1 U2227 ( .A(n3964), .B(DATAIN[30]), .S(n256), .Z(n3461) );
  MUX2_X1 U2228 ( .A(n3965), .B(DATAIN[31]), .S(n256), .Z(n3462) );
  MUX2_X1 U2229 ( .A(n3966), .B(DATAIN[0]), .S(n257), .Z(n3463) );
  MUX2_X1 U2230 ( .A(n3967), .B(DATAIN[1]), .S(n257), .Z(n3464) );
  MUX2_X1 U2231 ( .A(n3968), .B(DATAIN[2]), .S(n257), .Z(n3465) );
  MUX2_X1 U2232 ( .A(n3969), .B(DATAIN[3]), .S(n257), .Z(n3466) );
  MUX2_X1 U2233 ( .A(n3970), .B(DATAIN[4]), .S(n257), .Z(n3467) );
  MUX2_X1 U2234 ( .A(n3971), .B(DATAIN[5]), .S(n257), .Z(n3468) );
  MUX2_X1 U2235 ( .A(n3972), .B(DATAIN[6]), .S(n257), .Z(n3469) );
  MUX2_X1 U2236 ( .A(n3973), .B(DATAIN[7]), .S(n257), .Z(n3470) );
  MUX2_X1 U2237 ( .A(n3974), .B(DATAIN[8]), .S(n257), .Z(n3471) );
  MUX2_X1 U2238 ( .A(n3975), .B(DATAIN[9]), .S(n257), .Z(n3472) );
  MUX2_X1 U2239 ( .A(n3976), .B(DATAIN[10]), .S(n257), .Z(n3473) );
  MUX2_X1 U2240 ( .A(n3977), .B(DATAIN[11]), .S(n257), .Z(n3474) );
  MUX2_X1 U2241 ( .A(n3978), .B(DATAIN[12]), .S(n258), .Z(n3475) );
  MUX2_X1 U2242 ( .A(n3979), .B(DATAIN[13]), .S(n258), .Z(n3476) );
  MUX2_X1 U2243 ( .A(n3980), .B(DATAIN[14]), .S(n258), .Z(n3477) );
  MUX2_X1 U2244 ( .A(n3981), .B(DATAIN[15]), .S(n258), .Z(n3478) );
  MUX2_X1 U2245 ( .A(n3982), .B(DATAIN[16]), .S(n258), .Z(n3479) );
  MUX2_X1 U2246 ( .A(n3983), .B(DATAIN[17]), .S(n258), .Z(n3480) );
  MUX2_X1 U2247 ( .A(n3984), .B(DATAIN[18]), .S(n258), .Z(n3481) );
  MUX2_X1 U2248 ( .A(n3985), .B(DATAIN[19]), .S(n258), .Z(n3482) );
  MUX2_X1 U2249 ( .A(n3986), .B(DATAIN[20]), .S(n258), .Z(n3483) );
  MUX2_X1 U2250 ( .A(n3987), .B(DATAIN[21]), .S(n258), .Z(n3484) );
  MUX2_X1 U2251 ( .A(n3988), .B(DATAIN[22]), .S(n258), .Z(n3485) );
  MUX2_X1 U2252 ( .A(n3989), .B(DATAIN[23]), .S(n258), .Z(n3486) );
  MUX2_X1 U2253 ( .A(n3990), .B(DATAIN[24]), .S(n259), .Z(n3487) );
  MUX2_X1 U2254 ( .A(n3991), .B(DATAIN[25]), .S(n259), .Z(n3488) );
  MUX2_X1 U2255 ( .A(n3992), .B(DATAIN[26]), .S(n259), .Z(n3489) );
  MUX2_X1 U2256 ( .A(n3993), .B(DATAIN[27]), .S(n259), .Z(n3490) );
  MUX2_X1 U2257 ( .A(n3994), .B(DATAIN[28]), .S(n259), .Z(n3491) );
  MUX2_X1 U2258 ( .A(n3995), .B(DATAIN[29]), .S(n259), .Z(n3492) );
  MUX2_X1 U2259 ( .A(n3996), .B(DATAIN[30]), .S(n259), .Z(n3493) );
  MUX2_X1 U2260 ( .A(n3997), .B(DATAIN[31]), .S(n259), .Z(n3494) );
  MUX2_X1 U2261 ( .A(n1811), .B(DATAIN[0]), .S(n260), .Z(n4318) );
  MUX2_X1 U2262 ( .A(n1812), .B(DATAIN[1]), .S(n260), .Z(n4319) );
  MUX2_X1 U2263 ( .A(n1813), .B(DATAIN[2]), .S(n260), .Z(n4320) );
  MUX2_X1 U2264 ( .A(n1814), .B(DATAIN[3]), .S(n260), .Z(n4321) );
  MUX2_X1 U2265 ( .A(n1815), .B(DATAIN[4]), .S(n260), .Z(n4322) );
  MUX2_X1 U2266 ( .A(n1816), .B(DATAIN[5]), .S(n260), .Z(n4323) );
  MUX2_X1 U2267 ( .A(n1817), .B(DATAIN[6]), .S(n260), .Z(n4324) );
  MUX2_X1 U2268 ( .A(n1818), .B(DATAIN[7]), .S(n260), .Z(n4325) );
  MUX2_X1 U2269 ( .A(n1819), .B(DATAIN[8]), .S(n260), .Z(n4326) );
  MUX2_X1 U2270 ( .A(n1820), .B(DATAIN[9]), .S(n260), .Z(n4327) );
  MUX2_X1 U2271 ( .A(n1821), .B(DATAIN[10]), .S(n260), .Z(n4328) );
  MUX2_X1 U2272 ( .A(n1822), .B(DATAIN[11]), .S(n260), .Z(n4329) );
  MUX2_X1 U2273 ( .A(n1823), .B(DATAIN[12]), .S(n261), .Z(n4330) );
  MUX2_X1 U2274 ( .A(n1824), .B(DATAIN[13]), .S(n261), .Z(n4331) );
  MUX2_X1 U2275 ( .A(n1825), .B(DATAIN[14]), .S(n261), .Z(n4332) );
  MUX2_X1 U2276 ( .A(n1826), .B(DATAIN[15]), .S(n261), .Z(n4333) );
  MUX2_X1 U2277 ( .A(n1827), .B(DATAIN[16]), .S(n261), .Z(n4334) );
  MUX2_X1 U2278 ( .A(n1828), .B(DATAIN[17]), .S(n261), .Z(n4335) );
  MUX2_X1 U2279 ( .A(n1829), .B(DATAIN[18]), .S(n261), .Z(n4336) );
  MUX2_X1 U2280 ( .A(n1830), .B(DATAIN[19]), .S(n261), .Z(n4337) );
  MUX2_X1 U2281 ( .A(n1831), .B(DATAIN[20]), .S(n261), .Z(n4338) );
  MUX2_X1 U2282 ( .A(n1832), .B(DATAIN[21]), .S(n261), .Z(n4339) );
  MUX2_X1 U2283 ( .A(n1833), .B(DATAIN[22]), .S(n261), .Z(n4340) );
  MUX2_X1 U2284 ( .A(n1834), .B(DATAIN[23]), .S(n261), .Z(n4341) );
  MUX2_X1 U2285 ( .A(n1835), .B(DATAIN[24]), .S(n262), .Z(n4342) );
  MUX2_X1 U2286 ( .A(n1836), .B(DATAIN[25]), .S(n262), .Z(n4343) );
  MUX2_X1 U2287 ( .A(n1837), .B(DATAIN[26]), .S(n262), .Z(n4344) );
  MUX2_X1 U2288 ( .A(n1838), .B(DATAIN[27]), .S(n262), .Z(n4345) );
  MUX2_X1 U2289 ( .A(n1839), .B(DATAIN[28]), .S(n262), .Z(n4346) );
  MUX2_X1 U2290 ( .A(n1840), .B(DATAIN[29]), .S(n262), .Z(n4347) );
  MUX2_X1 U2291 ( .A(n1841), .B(DATAIN[30]), .S(n262), .Z(n4348) );
  MUX2_X1 U2292 ( .A(n1842), .B(DATAIN[31]), .S(n262), .Z(n4349) );
  MUX2_X1 U2293 ( .A(n1843), .B(DATAIN[0]), .S(n263), .Z(n4286) );
  MUX2_X1 U2294 ( .A(n1844), .B(DATAIN[1]), .S(n263), .Z(n4287) );
  MUX2_X1 U2295 ( .A(n1845), .B(DATAIN[2]), .S(n263), .Z(n4288) );
  MUX2_X1 U2296 ( .A(n1846), .B(DATAIN[3]), .S(n263), .Z(n4289) );
  MUX2_X1 U2297 ( .A(n1847), .B(DATAIN[4]), .S(n263), .Z(n4290) );
  MUX2_X1 U2298 ( .A(n1848), .B(DATAIN[5]), .S(n263), .Z(n4291) );
  MUX2_X1 U2299 ( .A(n1849), .B(DATAIN[6]), .S(n263), .Z(n4292) );
  MUX2_X1 U2300 ( .A(n1850), .B(DATAIN[7]), .S(n263), .Z(n4293) );
  MUX2_X1 U2301 ( .A(n1851), .B(DATAIN[8]), .S(n263), .Z(n4294) );
  MUX2_X1 U2302 ( .A(n1852), .B(DATAIN[9]), .S(n263), .Z(n4295) );
  MUX2_X1 U2303 ( .A(n1853), .B(DATAIN[10]), .S(n263), .Z(n4296) );
  MUX2_X1 U2304 ( .A(n1854), .B(DATAIN[11]), .S(n263), .Z(n4297) );
  MUX2_X1 U2305 ( .A(n1855), .B(DATAIN[12]), .S(n264), .Z(n4298) );
  MUX2_X1 U2306 ( .A(n1856), .B(DATAIN[13]), .S(n264), .Z(n4299) );
  MUX2_X1 U2307 ( .A(n1857), .B(DATAIN[14]), .S(n264), .Z(n4300) );
  MUX2_X1 U2308 ( .A(n1858), .B(DATAIN[15]), .S(n264), .Z(n4301) );
  MUX2_X1 U2309 ( .A(n1859), .B(DATAIN[16]), .S(n264), .Z(n4302) );
  MUX2_X1 U2310 ( .A(n1860), .B(DATAIN[17]), .S(n264), .Z(n4303) );
  MUX2_X1 U2311 ( .A(n1861), .B(DATAIN[18]), .S(n264), .Z(n4304) );
  MUX2_X1 U2312 ( .A(n1862), .B(DATAIN[19]), .S(n264), .Z(n4305) );
  MUX2_X1 U2313 ( .A(n1863), .B(DATAIN[20]), .S(n264), .Z(n4306) );
  MUX2_X1 U2314 ( .A(n1864), .B(DATAIN[21]), .S(n264), .Z(n4307) );
  MUX2_X1 U2315 ( .A(n1865), .B(DATAIN[22]), .S(n264), .Z(n4308) );
  MUX2_X1 U2316 ( .A(n1866), .B(DATAIN[23]), .S(n264), .Z(n4309) );
  MUX2_X1 U2317 ( .A(n1867), .B(DATAIN[24]), .S(n265), .Z(n4310) );
  MUX2_X1 U2318 ( .A(n1868), .B(DATAIN[25]), .S(n265), .Z(n4311) );
  MUX2_X1 U2319 ( .A(n1869), .B(DATAIN[26]), .S(n265), .Z(n4312) );
  MUX2_X1 U2320 ( .A(n1870), .B(DATAIN[27]), .S(n265), .Z(n4313) );
  MUX2_X1 U2321 ( .A(n1871), .B(DATAIN[28]), .S(n265), .Z(n4314) );
  MUX2_X1 U2322 ( .A(n1872), .B(DATAIN[29]), .S(n265), .Z(n4315) );
  MUX2_X1 U2323 ( .A(n1873), .B(DATAIN[30]), .S(n265), .Z(n4316) );
  MUX2_X1 U2324 ( .A(n1874), .B(DATAIN[31]), .S(n265), .Z(n4317) );
  MUX2_X1 U2325 ( .A(n4030), .B(DATAIN[0]), .S(n266), .Z(n3495) );
  MUX2_X1 U2326 ( .A(n4031), .B(DATAIN[1]), .S(n266), .Z(n3496) );
  MUX2_X1 U2327 ( .A(n4032), .B(DATAIN[2]), .S(n266), .Z(n3497) );
  MUX2_X1 U2328 ( .A(n4033), .B(DATAIN[3]), .S(n266), .Z(n3498) );
  MUX2_X1 U2329 ( .A(n4034), .B(DATAIN[4]), .S(n266), .Z(n3499) );
  MUX2_X1 U2330 ( .A(n4035), .B(DATAIN[5]), .S(n266), .Z(n3500) );
  MUX2_X1 U2331 ( .A(n4036), .B(DATAIN[6]), .S(n266), .Z(n3501) );
  MUX2_X1 U2332 ( .A(n4037), .B(DATAIN[7]), .S(n266), .Z(n3502) );
  MUX2_X1 U2333 ( .A(n4038), .B(DATAIN[8]), .S(n266), .Z(n3503) );
  MUX2_X1 U2334 ( .A(n4039), .B(DATAIN[9]), .S(n266), .Z(n3504) );
  MUX2_X1 U2335 ( .A(n4040), .B(DATAIN[10]), .S(n266), .Z(n3505) );
  MUX2_X1 U2336 ( .A(n4041), .B(DATAIN[11]), .S(n266), .Z(n3506) );
  MUX2_X1 U2337 ( .A(n4042), .B(DATAIN[12]), .S(n267), .Z(n3507) );
  MUX2_X1 U2338 ( .A(n4043), .B(DATAIN[13]), .S(n267), .Z(n3508) );
  MUX2_X1 U2339 ( .A(n4044), .B(DATAIN[14]), .S(n267), .Z(n3509) );
  MUX2_X1 U2340 ( .A(n4045), .B(DATAIN[15]), .S(n267), .Z(n3510) );
  MUX2_X1 U2341 ( .A(n4046), .B(DATAIN[16]), .S(n267), .Z(n3511) );
  MUX2_X1 U2342 ( .A(n4047), .B(DATAIN[17]), .S(n267), .Z(n3512) );
  MUX2_X1 U2343 ( .A(n4048), .B(DATAIN[18]), .S(n267), .Z(n3513) );
  MUX2_X1 U2344 ( .A(n4049), .B(DATAIN[19]), .S(n267), .Z(n3514) );
  MUX2_X1 U2345 ( .A(n4050), .B(DATAIN[20]), .S(n267), .Z(n3515) );
  MUX2_X1 U2346 ( .A(n4051), .B(DATAIN[21]), .S(n267), .Z(n3516) );
  MUX2_X1 U2347 ( .A(n4052), .B(DATAIN[22]), .S(n267), .Z(n3517) );
  MUX2_X1 U2348 ( .A(n4053), .B(DATAIN[23]), .S(n267), .Z(n3518) );
  MUX2_X1 U2349 ( .A(n4054), .B(DATAIN[24]), .S(n268), .Z(n3519) );
  MUX2_X1 U2350 ( .A(n4055), .B(DATAIN[25]), .S(n268), .Z(n3520) );
  MUX2_X1 U2351 ( .A(n4056), .B(DATAIN[26]), .S(n268), .Z(n3521) );
  MUX2_X1 U2352 ( .A(n4057), .B(DATAIN[27]), .S(n268), .Z(n3522) );
  MUX2_X1 U2353 ( .A(n4058), .B(DATAIN[28]), .S(n268), .Z(n3523) );
  MUX2_X1 U2354 ( .A(n4059), .B(DATAIN[29]), .S(n268), .Z(n3524) );
  MUX2_X1 U2355 ( .A(n4060), .B(DATAIN[30]), .S(n268), .Z(n3525) );
  MUX2_X1 U2356 ( .A(n4061), .B(DATAIN[31]), .S(n268), .Z(n3526) );
  MUX2_X1 U2357 ( .A(n4062), .B(DATAIN[0]), .S(n269), .Z(n3527) );
  MUX2_X1 U2358 ( .A(n4063), .B(DATAIN[1]), .S(n269), .Z(n3528) );
  MUX2_X1 U2359 ( .A(n4064), .B(DATAIN[2]), .S(n269), .Z(n3529) );
  MUX2_X1 U2360 ( .A(n4065), .B(DATAIN[3]), .S(n269), .Z(n3530) );
  MUX2_X1 U2361 ( .A(n4066), .B(DATAIN[4]), .S(n269), .Z(n3531) );
  MUX2_X1 U2362 ( .A(n4067), .B(DATAIN[5]), .S(n269), .Z(n3532) );
  MUX2_X1 U2363 ( .A(n4068), .B(DATAIN[6]), .S(n269), .Z(n3533) );
  MUX2_X1 U2364 ( .A(n4069), .B(DATAIN[7]), .S(n269), .Z(n3534) );
  MUX2_X1 U2365 ( .A(n4070), .B(DATAIN[8]), .S(n269), .Z(n3535) );
  MUX2_X1 U2366 ( .A(n4071), .B(DATAIN[9]), .S(n269), .Z(n3536) );
  MUX2_X1 U2367 ( .A(n4072), .B(DATAIN[10]), .S(n269), .Z(n3537) );
  MUX2_X1 U2368 ( .A(n4073), .B(DATAIN[11]), .S(n269), .Z(n3538) );
  MUX2_X1 U2369 ( .A(n4074), .B(DATAIN[12]), .S(n270), .Z(n3539) );
  MUX2_X1 U2370 ( .A(n4075), .B(DATAIN[13]), .S(n270), .Z(n3540) );
  MUX2_X1 U2371 ( .A(n4076), .B(DATAIN[14]), .S(n270), .Z(n3541) );
  MUX2_X1 U2372 ( .A(n4077), .B(DATAIN[15]), .S(n270), .Z(n3542) );
  MUX2_X1 U2373 ( .A(n4078), .B(DATAIN[16]), .S(n270), .Z(n3543) );
  MUX2_X1 U2374 ( .A(n4079), .B(DATAIN[17]), .S(n270), .Z(n3544) );
  MUX2_X1 U2375 ( .A(n4080), .B(DATAIN[18]), .S(n270), .Z(n3545) );
  MUX2_X1 U2376 ( .A(n4081), .B(DATAIN[19]), .S(n270), .Z(n3546) );
  MUX2_X1 U2377 ( .A(n4082), .B(DATAIN[20]), .S(n270), .Z(n3547) );
  MUX2_X1 U2378 ( .A(n4083), .B(DATAIN[21]), .S(n270), .Z(n3548) );
  MUX2_X1 U2379 ( .A(n4084), .B(DATAIN[22]), .S(n270), .Z(n3549) );
  MUX2_X1 U2380 ( .A(n4085), .B(DATAIN[23]), .S(n270), .Z(n3550) );
  MUX2_X1 U2381 ( .A(n4086), .B(DATAIN[24]), .S(n271), .Z(n3551) );
  MUX2_X1 U2382 ( .A(n4087), .B(DATAIN[25]), .S(n271), .Z(n3552) );
  MUX2_X1 U2383 ( .A(n4088), .B(DATAIN[26]), .S(n271), .Z(n3553) );
  MUX2_X1 U2384 ( .A(n4089), .B(DATAIN[27]), .S(n271), .Z(n3554) );
  MUX2_X1 U2385 ( .A(n4090), .B(DATAIN[28]), .S(n271), .Z(n3555) );
  MUX2_X1 U2386 ( .A(n4091), .B(DATAIN[29]), .S(n271), .Z(n3556) );
  MUX2_X1 U2387 ( .A(n4092), .B(DATAIN[30]), .S(n271), .Z(n3557) );
  MUX2_X1 U2388 ( .A(n4093), .B(DATAIN[31]), .S(n271), .Z(n3558) );
  MUX2_X1 U2389 ( .A(n1875), .B(DATAIN[0]), .S(n272), .Z(n4254) );
  MUX2_X1 U2390 ( .A(n1876), .B(DATAIN[1]), .S(n272), .Z(n4255) );
  MUX2_X1 U2391 ( .A(n1877), .B(DATAIN[2]), .S(n272), .Z(n4256) );
  MUX2_X1 U2392 ( .A(n1878), .B(DATAIN[3]), .S(n272), .Z(n4257) );
  MUX2_X1 U2393 ( .A(n1879), .B(DATAIN[4]), .S(n272), .Z(n4258) );
  MUX2_X1 U2394 ( .A(n1880), .B(DATAIN[5]), .S(n272), .Z(n4259) );
  MUX2_X1 U2395 ( .A(n1881), .B(DATAIN[6]), .S(n272), .Z(n4260) );
  MUX2_X1 U2396 ( .A(n1882), .B(DATAIN[7]), .S(n272), .Z(n4261) );
  MUX2_X1 U2397 ( .A(n1883), .B(DATAIN[8]), .S(n272), .Z(n4262) );
  MUX2_X1 U2398 ( .A(n1884), .B(DATAIN[9]), .S(n272), .Z(n4263) );
  MUX2_X1 U2399 ( .A(n1885), .B(DATAIN[10]), .S(n272), .Z(n4264) );
  MUX2_X1 U2400 ( .A(n1886), .B(DATAIN[11]), .S(n272), .Z(n4265) );
  MUX2_X1 U2401 ( .A(n1887), .B(DATAIN[12]), .S(n273), .Z(n4266) );
  MUX2_X1 U2402 ( .A(n1888), .B(DATAIN[13]), .S(n273), .Z(n4267) );
  MUX2_X1 U2403 ( .A(n1889), .B(DATAIN[14]), .S(n273), .Z(n4268) );
  MUX2_X1 U2404 ( .A(n1890), .B(DATAIN[15]), .S(n273), .Z(n4269) );
  MUX2_X1 U2405 ( .A(n1891), .B(DATAIN[16]), .S(n273), .Z(n4270) );
  MUX2_X1 U2406 ( .A(n1892), .B(DATAIN[17]), .S(n273), .Z(n4271) );
  MUX2_X1 U2407 ( .A(n1893), .B(DATAIN[18]), .S(n273), .Z(n4272) );
  MUX2_X1 U2408 ( .A(n1894), .B(DATAIN[19]), .S(n273), .Z(n4273) );
  MUX2_X1 U2409 ( .A(n1895), .B(DATAIN[20]), .S(n273), .Z(n4274) );
  MUX2_X1 U2410 ( .A(n1896), .B(DATAIN[21]), .S(n273), .Z(n4275) );
  MUX2_X1 U2411 ( .A(n1897), .B(DATAIN[22]), .S(n273), .Z(n4276) );
  MUX2_X1 U2412 ( .A(n1898), .B(DATAIN[23]), .S(n273), .Z(n4277) );
  MUX2_X1 U2413 ( .A(n1899), .B(DATAIN[24]), .S(n274), .Z(n4278) );
  MUX2_X1 U2414 ( .A(n1900), .B(DATAIN[25]), .S(n274), .Z(n4279) );
  MUX2_X1 U2415 ( .A(n1901), .B(DATAIN[26]), .S(n274), .Z(n4280) );
  MUX2_X1 U2416 ( .A(n1902), .B(DATAIN[27]), .S(n274), .Z(n4281) );
  MUX2_X1 U2417 ( .A(n1903), .B(DATAIN[28]), .S(n274), .Z(n4282) );
  MUX2_X1 U2418 ( .A(n1904), .B(DATAIN[29]), .S(n274), .Z(n4283) );
  MUX2_X1 U2419 ( .A(n1905), .B(DATAIN[30]), .S(n274), .Z(n4284) );
  MUX2_X1 U2420 ( .A(n1906), .B(DATAIN[31]), .S(n274), .Z(n4285) );
  AND2_X1 U2421 ( .A1(WR), .A2(ENABLE), .ZN(n1908) );
  OAI22_X1 U2422 ( .A1(n2974), .A2(n277), .B1(n1922), .B2(n280), .ZN(n1920) );
  AOI221_X1 U2423 ( .B1(n283), .B2(n3678), .C1(n286), .C2(n3710), .A(n1930), 
        .ZN(n1927) );
  OAI22_X1 U2424 ( .A1(n3742), .A2(n289), .B1(n3774), .B2(n292), .ZN(n1930) );
  AOI221_X1 U2425 ( .B1(n295), .B2(n3806), .C1(n298), .C2(n3838), .A(n1935), 
        .ZN(n1926) );
  OAI22_X1 U2426 ( .A1(n3870), .A2(n301), .B1(n3902), .B2(n304), .ZN(n1935) );
  OAI22_X1 U2427 ( .A1(n1940), .A2(n310), .B1(n1942), .B2(n313), .ZN(n1939) );
  OAI22_X1 U2428 ( .A1(n1946), .A2(n319), .B1(n1948), .B2(n322), .ZN(n1945) );
  OAI22_X1 U2429 ( .A1(n2975), .A2(n277), .B1(n1951), .B2(n280), .ZN(n1950) );
  AOI221_X1 U2430 ( .B1(n283), .B2(n3679), .C1(n286), .C2(n3711), .A(n1954), 
        .ZN(n1953) );
  OAI22_X1 U2431 ( .A1(n3743), .A2(n289), .B1(n3775), .B2(n292), .ZN(n1954) );
  AOI221_X1 U2432 ( .B1(n295), .B2(n3807), .C1(n298), .C2(n3839), .A(n1955), 
        .ZN(n1952) );
  OAI22_X1 U2433 ( .A1(n3871), .A2(n301), .B1(n3903), .B2(n304), .ZN(n1955) );
  OAI22_X1 U2434 ( .A1(n1957), .A2(n310), .B1(n1958), .B2(n313), .ZN(n1956) );
  OAI22_X1 U2435 ( .A1(n1960), .A2(n319), .B1(n1961), .B2(n322), .ZN(n1959) );
  OAI22_X1 U2436 ( .A1(n2976), .A2(n277), .B1(n1963), .B2(n280), .ZN(n1962) );
  AOI221_X1 U2437 ( .B1(n283), .B2(n3680), .C1(n286), .C2(n3712), .A(n1966), 
        .ZN(n1965) );
  OAI22_X1 U2438 ( .A1(n3744), .A2(n289), .B1(n3776), .B2(n292), .ZN(n1966) );
  AOI221_X1 U2439 ( .B1(n295), .B2(n3808), .C1(n298), .C2(n3840), .A(n1967), 
        .ZN(n1964) );
  OAI22_X1 U2440 ( .A1(n3872), .A2(n301), .B1(n3904), .B2(n304), .ZN(n1967) );
  OAI22_X1 U2441 ( .A1(n1969), .A2(n310), .B1(n1970), .B2(n313), .ZN(n1968) );
  OAI22_X1 U2442 ( .A1(n1972), .A2(n319), .B1(n1973), .B2(n322), .ZN(n1971) );
  OAI22_X1 U2443 ( .A1(n2977), .A2(n277), .B1(n1975), .B2(n280), .ZN(n1974) );
  AOI221_X1 U2444 ( .B1(n283), .B2(n3681), .C1(n286), .C2(n3713), .A(n1978), 
        .ZN(n1977) );
  OAI22_X1 U2445 ( .A1(n3745), .A2(n289), .B1(n3777), .B2(n292), .ZN(n1978) );
  AOI221_X1 U2446 ( .B1(n295), .B2(n3809), .C1(n298), .C2(n3841), .A(n1979), 
        .ZN(n1976) );
  OAI22_X1 U2447 ( .A1(n3873), .A2(n301), .B1(n3905), .B2(n304), .ZN(n1979) );
  OAI22_X1 U2448 ( .A1(n1981), .A2(n310), .B1(n1982), .B2(n313), .ZN(n1980) );
  OAI22_X1 U2449 ( .A1(n1984), .A2(n319), .B1(n1985), .B2(n322), .ZN(n1983) );
  OAI22_X1 U2450 ( .A1(n2978), .A2(n277), .B1(n1987), .B2(n280), .ZN(n1986) );
  AOI221_X1 U2451 ( .B1(n283), .B2(n3682), .C1(n286), .C2(n3714), .A(n1990), 
        .ZN(n1989) );
  OAI22_X1 U2452 ( .A1(n3746), .A2(n289), .B1(n3778), .B2(n292), .ZN(n1990) );
  AOI221_X1 U2453 ( .B1(n295), .B2(n3810), .C1(n298), .C2(n3842), .A(n1991), 
        .ZN(n1988) );
  OAI22_X1 U2454 ( .A1(n3874), .A2(n301), .B1(n3906), .B2(n304), .ZN(n1991) );
  OAI22_X1 U2455 ( .A1(n1993), .A2(n310), .B1(n1994), .B2(n313), .ZN(n1992) );
  OAI22_X1 U2456 ( .A1(n1996), .A2(n319), .B1(n1997), .B2(n322), .ZN(n1995) );
  OAI22_X1 U2457 ( .A1(n2979), .A2(n277), .B1(n1999), .B2(n280), .ZN(n1998) );
  AOI221_X1 U2458 ( .B1(n283), .B2(n3683), .C1(n286), .C2(n3715), .A(n2002), 
        .ZN(n2001) );
  OAI22_X1 U2459 ( .A1(n3747), .A2(n289), .B1(n3779), .B2(n292), .ZN(n2002) );
  AOI221_X1 U2460 ( .B1(n295), .B2(n3811), .C1(n298), .C2(n3843), .A(n2003), 
        .ZN(n2000) );
  OAI22_X1 U2461 ( .A1(n3875), .A2(n301), .B1(n3907), .B2(n304), .ZN(n2003) );
  OAI22_X1 U2462 ( .A1(n2005), .A2(n310), .B1(n2006), .B2(n313), .ZN(n2004) );
  OAI22_X1 U2463 ( .A1(n2008), .A2(n319), .B1(n2009), .B2(n322), .ZN(n2007) );
  OAI22_X1 U2464 ( .A1(n2980), .A2(n277), .B1(n2011), .B2(n280), .ZN(n2010) );
  AOI221_X1 U2465 ( .B1(n283), .B2(n3684), .C1(n286), .C2(n3716), .A(n2014), 
        .ZN(n2013) );
  OAI22_X1 U2466 ( .A1(n3748), .A2(n289), .B1(n3780), .B2(n292), .ZN(n2014) );
  AOI221_X1 U2467 ( .B1(n295), .B2(n3812), .C1(n298), .C2(n3844), .A(n2015), 
        .ZN(n2012) );
  OAI22_X1 U2468 ( .A1(n3876), .A2(n301), .B1(n3908), .B2(n304), .ZN(n2015) );
  OAI22_X1 U2469 ( .A1(n2017), .A2(n310), .B1(n2018), .B2(n313), .ZN(n2016) );
  OAI22_X1 U2470 ( .A1(n2020), .A2(n319), .B1(n2021), .B2(n322), .ZN(n2019) );
  OAI22_X1 U2471 ( .A1(n2981), .A2(n277), .B1(n2023), .B2(n280), .ZN(n2022) );
  AOI221_X1 U2472 ( .B1(n283), .B2(n3685), .C1(n286), .C2(n3717), .A(n2026), 
        .ZN(n2025) );
  OAI22_X1 U2473 ( .A1(n3749), .A2(n289), .B1(n3781), .B2(n292), .ZN(n2026) );
  AOI221_X1 U2474 ( .B1(n295), .B2(n3813), .C1(n298), .C2(n3845), .A(n2027), 
        .ZN(n2024) );
  OAI22_X1 U2475 ( .A1(n3877), .A2(n301), .B1(n3909), .B2(n304), .ZN(n2027) );
  OAI22_X1 U2476 ( .A1(n2029), .A2(n310), .B1(n2030), .B2(n313), .ZN(n2028) );
  OAI22_X1 U2477 ( .A1(n2032), .A2(n319), .B1(n2033), .B2(n322), .ZN(n2031) );
  OAI22_X1 U2478 ( .A1(n2982), .A2(n276), .B1(n2035), .B2(n279), .ZN(n2034) );
  AOI221_X1 U2479 ( .B1(n282), .B2(n3686), .C1(n285), .C2(n3718), .A(n2038), 
        .ZN(n2037) );
  OAI22_X1 U2480 ( .A1(n3750), .A2(n288), .B1(n3782), .B2(n291), .ZN(n2038) );
  AOI221_X1 U2481 ( .B1(n294), .B2(n3814), .C1(n297), .C2(n3846), .A(n2039), 
        .ZN(n2036) );
  OAI22_X1 U2482 ( .A1(n3878), .A2(n300), .B1(n3910), .B2(n303), .ZN(n2039) );
  OAI22_X1 U2483 ( .A1(n2041), .A2(n309), .B1(n2042), .B2(n312), .ZN(n2040) );
  OAI22_X1 U2484 ( .A1(n2044), .A2(n318), .B1(n2045), .B2(n321), .ZN(n2043) );
  OAI22_X1 U2485 ( .A1(n3559), .A2(n276), .B1(n2047), .B2(n279), .ZN(n2046) );
  AOI221_X1 U2486 ( .B1(n282), .B2(n3687), .C1(n285), .C2(n3719), .A(n2050), 
        .ZN(n2049) );
  OAI22_X1 U2487 ( .A1(n3751), .A2(n288), .B1(n3783), .B2(n291), .ZN(n2050) );
  AOI221_X1 U2488 ( .B1(n294), .B2(n3815), .C1(n297), .C2(n3847), .A(n2051), 
        .ZN(n2048) );
  OAI22_X1 U2489 ( .A1(n3879), .A2(n300), .B1(n3911), .B2(n303), .ZN(n2051) );
  OAI22_X1 U2490 ( .A1(n2053), .A2(n309), .B1(n2054), .B2(n312), .ZN(n2052) );
  OAI22_X1 U2491 ( .A1(n2056), .A2(n318), .B1(n2057), .B2(n321), .ZN(n2055) );
  OAI22_X1 U2492 ( .A1(n3560), .A2(n276), .B1(n2059), .B2(n279), .ZN(n2058) );
  AOI221_X1 U2493 ( .B1(n282), .B2(n3688), .C1(n285), .C2(n3720), .A(n2062), 
        .ZN(n2061) );
  OAI22_X1 U2494 ( .A1(n3752), .A2(n288), .B1(n3784), .B2(n291), .ZN(n2062) );
  AOI221_X1 U2495 ( .B1(n294), .B2(n3816), .C1(n297), .C2(n3848), .A(n2063), 
        .ZN(n2060) );
  OAI22_X1 U2496 ( .A1(n3880), .A2(n300), .B1(n3912), .B2(n303), .ZN(n2063) );
  OAI22_X1 U2497 ( .A1(n2065), .A2(n309), .B1(n2066), .B2(n312), .ZN(n2064) );
  OAI22_X1 U2498 ( .A1(n2068), .A2(n318), .B1(n2069), .B2(n321), .ZN(n2067) );
  OAI22_X1 U2499 ( .A1(n3561), .A2(n276), .B1(n2071), .B2(n279), .ZN(n2070) );
  AOI221_X1 U2500 ( .B1(n282), .B2(n3689), .C1(n285), .C2(n3721), .A(n2074), 
        .ZN(n2073) );
  OAI22_X1 U2501 ( .A1(n3753), .A2(n288), .B1(n3785), .B2(n291), .ZN(n2074) );
  AOI221_X1 U2502 ( .B1(n294), .B2(n3817), .C1(n297), .C2(n3849), .A(n2075), 
        .ZN(n2072) );
  OAI22_X1 U2503 ( .A1(n3881), .A2(n300), .B1(n3913), .B2(n303), .ZN(n2075) );
  OAI22_X1 U2504 ( .A1(n2077), .A2(n309), .B1(n2078), .B2(n312), .ZN(n2076) );
  OAI22_X1 U2505 ( .A1(n2080), .A2(n318), .B1(n2081), .B2(n321), .ZN(n2079) );
  OAI22_X1 U2506 ( .A1(n3562), .A2(n276), .B1(n2083), .B2(n279), .ZN(n2082) );
  AOI221_X1 U2507 ( .B1(n282), .B2(n3690), .C1(n285), .C2(n3722), .A(n2086), 
        .ZN(n2085) );
  OAI22_X1 U2508 ( .A1(n3754), .A2(n288), .B1(n3786), .B2(n291), .ZN(n2086) );
  AOI221_X1 U2509 ( .B1(n294), .B2(n3818), .C1(n297), .C2(n3850), .A(n2087), 
        .ZN(n2084) );
  OAI22_X1 U2510 ( .A1(n3882), .A2(n300), .B1(n3914), .B2(n303), .ZN(n2087) );
  OAI22_X1 U2511 ( .A1(n2089), .A2(n309), .B1(n2090), .B2(n312), .ZN(n2088) );
  OAI22_X1 U2512 ( .A1(n2092), .A2(n318), .B1(n2093), .B2(n321), .ZN(n2091) );
  OAI22_X1 U2513 ( .A1(n3563), .A2(n276), .B1(n2095), .B2(n279), .ZN(n2094) );
  AOI221_X1 U2514 ( .B1(n282), .B2(n3691), .C1(n285), .C2(n3723), .A(n2098), 
        .ZN(n2097) );
  OAI22_X1 U2515 ( .A1(n3755), .A2(n288), .B1(n3787), .B2(n291), .ZN(n2098) );
  AOI221_X1 U2516 ( .B1(n294), .B2(n3819), .C1(n297), .C2(n3851), .A(n2099), 
        .ZN(n2096) );
  OAI22_X1 U2517 ( .A1(n3883), .A2(n300), .B1(n3915), .B2(n303), .ZN(n2099) );
  OAI22_X1 U2518 ( .A1(n2101), .A2(n309), .B1(n2102), .B2(n312), .ZN(n2100) );
  OAI22_X1 U2519 ( .A1(n2104), .A2(n318), .B1(n2105), .B2(n321), .ZN(n2103) );
  OAI22_X1 U2520 ( .A1(n3564), .A2(n276), .B1(n2107), .B2(n279), .ZN(n2106) );
  AOI221_X1 U2521 ( .B1(n282), .B2(n3692), .C1(n285), .C2(n3724), .A(n2110), 
        .ZN(n2109) );
  OAI22_X1 U2522 ( .A1(n3756), .A2(n288), .B1(n3788), .B2(n291), .ZN(n2110) );
  AOI221_X1 U2523 ( .B1(n294), .B2(n3820), .C1(n297), .C2(n3852), .A(n2111), 
        .ZN(n2108) );
  OAI22_X1 U2524 ( .A1(n3884), .A2(n300), .B1(n3916), .B2(n303), .ZN(n2111) );
  OAI22_X1 U2525 ( .A1(n2113), .A2(n309), .B1(n2114), .B2(n312), .ZN(n2112) );
  OAI22_X1 U2526 ( .A1(n2116), .A2(n318), .B1(n2117), .B2(n321), .ZN(n2115) );
  OAI22_X1 U2527 ( .A1(n3565), .A2(n276), .B1(n2119), .B2(n279), .ZN(n2118) );
  AOI221_X1 U2528 ( .B1(n282), .B2(n3693), .C1(n285), .C2(n3725), .A(n2122), 
        .ZN(n2121) );
  OAI22_X1 U2529 ( .A1(n3757), .A2(n288), .B1(n3789), .B2(n291), .ZN(n2122) );
  AOI221_X1 U2530 ( .B1(n294), .B2(n3821), .C1(n297), .C2(n3853), .A(n2123), 
        .ZN(n2120) );
  OAI22_X1 U2531 ( .A1(n3885), .A2(n300), .B1(n3917), .B2(n303), .ZN(n2123) );
  OAI22_X1 U2532 ( .A1(n2125), .A2(n309), .B1(n2126), .B2(n312), .ZN(n2124) );
  OAI22_X1 U2533 ( .A1(n2128), .A2(n318), .B1(n2129), .B2(n321), .ZN(n2127) );
  OAI22_X1 U2534 ( .A1(n3566), .A2(n276), .B1(n2131), .B2(n279), .ZN(n2130) );
  AOI221_X1 U2535 ( .B1(n282), .B2(n3694), .C1(n285), .C2(n3726), .A(n2134), 
        .ZN(n2133) );
  OAI22_X1 U2536 ( .A1(n3758), .A2(n288), .B1(n3790), .B2(n291), .ZN(n2134) );
  AOI221_X1 U2537 ( .B1(n294), .B2(n3822), .C1(n297), .C2(n3854), .A(n2135), 
        .ZN(n2132) );
  OAI22_X1 U2538 ( .A1(n3886), .A2(n300), .B1(n3918), .B2(n303), .ZN(n2135) );
  OAI22_X1 U2539 ( .A1(n2137), .A2(n309), .B1(n2138), .B2(n312), .ZN(n2136) );
  OAI22_X1 U2540 ( .A1(n2140), .A2(n318), .B1(n2141), .B2(n321), .ZN(n2139) );
  OAI22_X1 U2541 ( .A1(n3567), .A2(n276), .B1(n2143), .B2(n279), .ZN(n2142) );
  AOI221_X1 U2542 ( .B1(n282), .B2(n3695), .C1(n285), .C2(n3727), .A(n2146), 
        .ZN(n2145) );
  OAI22_X1 U2543 ( .A1(n3759), .A2(n288), .B1(n3791), .B2(n291), .ZN(n2146) );
  AOI221_X1 U2544 ( .B1(n294), .B2(n3823), .C1(n297), .C2(n3855), .A(n2147), 
        .ZN(n2144) );
  OAI22_X1 U2545 ( .A1(n3887), .A2(n300), .B1(n3919), .B2(n303), .ZN(n2147) );
  OAI22_X1 U2546 ( .A1(n2149), .A2(n309), .B1(n2150), .B2(n312), .ZN(n2148) );
  OAI22_X1 U2547 ( .A1(n2152), .A2(n318), .B1(n2153), .B2(n321), .ZN(n2151) );
  OAI22_X1 U2548 ( .A1(n3568), .A2(n276), .B1(n2155), .B2(n279), .ZN(n2154) );
  AOI221_X1 U2549 ( .B1(n282), .B2(n3696), .C1(n285), .C2(n3728), .A(n2158), 
        .ZN(n2157) );
  OAI22_X1 U2550 ( .A1(n3760), .A2(n288), .B1(n3792), .B2(n291), .ZN(n2158) );
  AOI221_X1 U2551 ( .B1(n294), .B2(n3824), .C1(n297), .C2(n3856), .A(n2159), 
        .ZN(n2156) );
  OAI22_X1 U2552 ( .A1(n3888), .A2(n300), .B1(n3920), .B2(n303), .ZN(n2159) );
  OAI22_X1 U2553 ( .A1(n2161), .A2(n309), .B1(n2162), .B2(n312), .ZN(n2160) );
  OAI22_X1 U2554 ( .A1(n2164), .A2(n318), .B1(n2165), .B2(n321), .ZN(n2163) );
  OAI22_X1 U2555 ( .A1(n3569), .A2(n276), .B1(n2167), .B2(n279), .ZN(n2166) );
  AOI221_X1 U2556 ( .B1(n282), .B2(n3697), .C1(n285), .C2(n3729), .A(n2170), 
        .ZN(n2169) );
  OAI22_X1 U2557 ( .A1(n3761), .A2(n288), .B1(n3793), .B2(n291), .ZN(n2170) );
  AOI221_X1 U2558 ( .B1(n294), .B2(n3825), .C1(n297), .C2(n3857), .A(n2171), 
        .ZN(n2168) );
  OAI22_X1 U2559 ( .A1(n3889), .A2(n300), .B1(n3921), .B2(n303), .ZN(n2171) );
  OAI22_X1 U2560 ( .A1(n2173), .A2(n309), .B1(n2174), .B2(n312), .ZN(n2172) );
  OAI22_X1 U2561 ( .A1(n2176), .A2(n318), .B1(n2177), .B2(n321), .ZN(n2175) );
  OAI22_X1 U2562 ( .A1(n3570), .A2(n275), .B1(n2179), .B2(n278), .ZN(n2178) );
  AOI221_X1 U2563 ( .B1(n281), .B2(n3698), .C1(n284), .C2(n3730), .A(n2182), 
        .ZN(n2181) );
  OAI22_X1 U2564 ( .A1(n3762), .A2(n287), .B1(n3794), .B2(n290), .ZN(n2182) );
  AOI221_X1 U2565 ( .B1(n293), .B2(n3826), .C1(n296), .C2(n3858), .A(n2183), 
        .ZN(n2180) );
  OAI22_X1 U2566 ( .A1(n3890), .A2(n299), .B1(n3922), .B2(n302), .ZN(n2183) );
  OAI22_X1 U2567 ( .A1(n2185), .A2(n308), .B1(n2186), .B2(n311), .ZN(n2184) );
  OAI22_X1 U2568 ( .A1(n2188), .A2(n317), .B1(n2189), .B2(n320), .ZN(n2187) );
  OAI22_X1 U2569 ( .A1(n3571), .A2(n275), .B1(n2191), .B2(n278), .ZN(n2190) );
  AOI221_X1 U2570 ( .B1(n281), .B2(n3699), .C1(n284), .C2(n3731), .A(n2194), 
        .ZN(n2193) );
  OAI22_X1 U2571 ( .A1(n3763), .A2(n287), .B1(n3795), .B2(n290), .ZN(n2194) );
  AOI221_X1 U2572 ( .B1(n293), .B2(n3827), .C1(n296), .C2(n3859), .A(n2195), 
        .ZN(n2192) );
  OAI22_X1 U2573 ( .A1(n3891), .A2(n299), .B1(n3923), .B2(n302), .ZN(n2195) );
  OAI22_X1 U2574 ( .A1(n2197), .A2(n308), .B1(n2198), .B2(n311), .ZN(n2196) );
  OAI22_X1 U2575 ( .A1(n2200), .A2(n317), .B1(n2201), .B2(n320), .ZN(n2199) );
  OAI22_X1 U2576 ( .A1(n3572), .A2(n275), .B1(n2203), .B2(n278), .ZN(n2202) );
  AOI221_X1 U2577 ( .B1(n281), .B2(n3700), .C1(n284), .C2(n3732), .A(n2206), 
        .ZN(n2205) );
  OAI22_X1 U2578 ( .A1(n3764), .A2(n287), .B1(n3796), .B2(n290), .ZN(n2206) );
  AOI221_X1 U2579 ( .B1(n293), .B2(n3828), .C1(n296), .C2(n3860), .A(n2207), 
        .ZN(n2204) );
  OAI22_X1 U2580 ( .A1(n3892), .A2(n299), .B1(n3924), .B2(n302), .ZN(n2207) );
  OAI22_X1 U2581 ( .A1(n2209), .A2(n308), .B1(n2210), .B2(n311), .ZN(n2208) );
  OAI22_X1 U2582 ( .A1(n2212), .A2(n317), .B1(n2213), .B2(n320), .ZN(n2211) );
  OAI22_X1 U2583 ( .A1(n3573), .A2(n275), .B1(n2215), .B2(n278), .ZN(n2214) );
  AOI221_X1 U2584 ( .B1(n281), .B2(n3701), .C1(n284), .C2(n3733), .A(n2218), 
        .ZN(n2217) );
  OAI22_X1 U2585 ( .A1(n3765), .A2(n287), .B1(n3797), .B2(n290), .ZN(n2218) );
  AOI221_X1 U2586 ( .B1(n293), .B2(n3829), .C1(n296), .C2(n3861), .A(n2219), 
        .ZN(n2216) );
  OAI22_X1 U2587 ( .A1(n3893), .A2(n299), .B1(n3925), .B2(n302), .ZN(n2219) );
  OAI22_X1 U2588 ( .A1(n2221), .A2(n308), .B1(n2222), .B2(n311), .ZN(n2220) );
  OAI22_X1 U2589 ( .A1(n2224), .A2(n317), .B1(n2225), .B2(n320), .ZN(n2223) );
  OAI22_X1 U2590 ( .A1(n3574), .A2(n275), .B1(n2227), .B2(n278), .ZN(n2226) );
  AOI221_X1 U2591 ( .B1(n281), .B2(n3702), .C1(n284), .C2(n3734), .A(n2230), 
        .ZN(n2229) );
  OAI22_X1 U2592 ( .A1(n3766), .A2(n287), .B1(n3798), .B2(n290), .ZN(n2230) );
  AOI221_X1 U2593 ( .B1(n293), .B2(n3830), .C1(n296), .C2(n3862), .A(n2231), 
        .ZN(n2228) );
  OAI22_X1 U2594 ( .A1(n3894), .A2(n299), .B1(n3926), .B2(n302), .ZN(n2231) );
  OAI22_X1 U2595 ( .A1(n2233), .A2(n308), .B1(n2234), .B2(n311), .ZN(n2232) );
  OAI22_X1 U2596 ( .A1(n2236), .A2(n317), .B1(n2237), .B2(n320), .ZN(n2235) );
  OAI22_X1 U2597 ( .A1(n3575), .A2(n275), .B1(n2239), .B2(n278), .ZN(n2238) );
  AOI221_X1 U2598 ( .B1(n281), .B2(n3703), .C1(n284), .C2(n3735), .A(n2242), 
        .ZN(n2241) );
  OAI22_X1 U2599 ( .A1(n3767), .A2(n287), .B1(n3799), .B2(n290), .ZN(n2242) );
  AOI221_X1 U2600 ( .B1(n293), .B2(n3831), .C1(n296), .C2(n3863), .A(n2243), 
        .ZN(n2240) );
  OAI22_X1 U2601 ( .A1(n3895), .A2(n299), .B1(n3927), .B2(n302), .ZN(n2243) );
  OAI22_X1 U2602 ( .A1(n2245), .A2(n308), .B1(n2246), .B2(n311), .ZN(n2244) );
  OAI22_X1 U2603 ( .A1(n2248), .A2(n317), .B1(n2249), .B2(n320), .ZN(n2247) );
  OAI22_X1 U2604 ( .A1(n3576), .A2(n275), .B1(n2251), .B2(n278), .ZN(n2250) );
  AOI221_X1 U2605 ( .B1(n281), .B2(n3704), .C1(n284), .C2(n3736), .A(n2254), 
        .ZN(n2253) );
  OAI22_X1 U2606 ( .A1(n3768), .A2(n287), .B1(n3800), .B2(n290), .ZN(n2254) );
  AOI221_X1 U2607 ( .B1(n293), .B2(n3832), .C1(n296), .C2(n3864), .A(n2255), 
        .ZN(n2252) );
  OAI22_X1 U2608 ( .A1(n3896), .A2(n299), .B1(n3928), .B2(n302), .ZN(n2255) );
  OAI22_X1 U2609 ( .A1(n2257), .A2(n308), .B1(n2258), .B2(n311), .ZN(n2256) );
  OAI22_X1 U2610 ( .A1(n2260), .A2(n317), .B1(n2261), .B2(n320), .ZN(n2259) );
  OAI22_X1 U2611 ( .A1(n3577), .A2(n275), .B1(n2263), .B2(n278), .ZN(n2262) );
  AOI221_X1 U2612 ( .B1(n281), .B2(n3705), .C1(n284), .C2(n3737), .A(n2266), 
        .ZN(n2265) );
  OAI22_X1 U2613 ( .A1(n3769), .A2(n287), .B1(n3801), .B2(n290), .ZN(n2266) );
  AOI221_X1 U2614 ( .B1(n293), .B2(n3833), .C1(n296), .C2(n3865), .A(n2267), 
        .ZN(n2264) );
  OAI22_X1 U2615 ( .A1(n3897), .A2(n299), .B1(n3929), .B2(n302), .ZN(n2267) );
  OAI22_X1 U2616 ( .A1(n2269), .A2(n308), .B1(n2270), .B2(n311), .ZN(n2268) );
  OAI22_X1 U2617 ( .A1(n2272), .A2(n317), .B1(n2273), .B2(n320), .ZN(n2271) );
  OAI22_X1 U2618 ( .A1(n3578), .A2(n275), .B1(n2275), .B2(n278), .ZN(n2274) );
  AOI221_X1 U2619 ( .B1(n281), .B2(n3706), .C1(n284), .C2(n3738), .A(n2278), 
        .ZN(n2277) );
  OAI22_X1 U2620 ( .A1(n3770), .A2(n287), .B1(n3802), .B2(n290), .ZN(n2278) );
  AOI221_X1 U2621 ( .B1(n293), .B2(n3834), .C1(n296), .C2(n3866), .A(n2279), 
        .ZN(n2276) );
  OAI22_X1 U2622 ( .A1(n3898), .A2(n299), .B1(n3930), .B2(n302), .ZN(n2279) );
  OAI22_X1 U2623 ( .A1(n2281), .A2(n308), .B1(n2282), .B2(n311), .ZN(n2280) );
  OAI22_X1 U2624 ( .A1(n2284), .A2(n317), .B1(n2285), .B2(n320), .ZN(n2283) );
  OAI22_X1 U2625 ( .A1(n3579), .A2(n275), .B1(n2287), .B2(n278), .ZN(n2286) );
  AOI221_X1 U2626 ( .B1(n281), .B2(n3707), .C1(n284), .C2(n3739), .A(n2290), 
        .ZN(n2289) );
  OAI22_X1 U2627 ( .A1(n3771), .A2(n287), .B1(n3803), .B2(n290), .ZN(n2290) );
  AOI221_X1 U2628 ( .B1(n293), .B2(n3835), .C1(n296), .C2(n3867), .A(n2291), 
        .ZN(n2288) );
  OAI22_X1 U2629 ( .A1(n3899), .A2(n299), .B1(n3931), .B2(n302), .ZN(n2291) );
  OAI22_X1 U2630 ( .A1(n2293), .A2(n308), .B1(n2294), .B2(n311), .ZN(n2292) );
  OAI22_X1 U2631 ( .A1(n2296), .A2(n317), .B1(n2297), .B2(n320), .ZN(n2295) );
  OAI22_X1 U2632 ( .A1(n3580), .A2(n275), .B1(n2299), .B2(n278), .ZN(n2298) );
  AOI221_X1 U2633 ( .B1(n281), .B2(n3708), .C1(n284), .C2(n3740), .A(n2302), 
        .ZN(n2301) );
  OAI22_X1 U2634 ( .A1(n3772), .A2(n287), .B1(n3804), .B2(n290), .ZN(n2302) );
  AOI221_X1 U2635 ( .B1(n293), .B2(n3836), .C1(n296), .C2(n3868), .A(n2303), 
        .ZN(n2300) );
  OAI22_X1 U2636 ( .A1(n3900), .A2(n299), .B1(n3932), .B2(n302), .ZN(n2303) );
  OAI22_X1 U2637 ( .A1(n2305), .A2(n308), .B1(n2306), .B2(n311), .ZN(n2304) );
  OAI22_X1 U2638 ( .A1(n2308), .A2(n317), .B1(n2309), .B2(n320), .ZN(n2307) );
  AND2_X1 U2639 ( .A1(n2310), .A2(n2311), .ZN(n1912) );
  AND2_X1 U2640 ( .A1(n2310), .A2(n2312), .ZN(n1911) );
  NAND2_X1 U2641 ( .A1(n2313), .A2(n2314), .ZN(n1910) );
  NAND2_X1 U2642 ( .A1(n2315), .A2(n2311), .ZN(n1909) );
  AND2_X1 U2643 ( .A1(n2315), .A2(n2312), .ZN(n1916) );
  AND2_X1 U2644 ( .A1(n2315), .A2(n2314), .ZN(n1915) );
  NAND2_X1 U2645 ( .A1(n2310), .A2(n2314), .ZN(n1914) );
  NAND2_X1 U2646 ( .A1(n2310), .A2(n2316), .ZN(n1913) );
  NOR3_X1 U2647 ( .A1(n2317), .A2(ADD_RS2[0]), .A3(n2318), .ZN(n2310) );
  OAI22_X1 U2648 ( .A1(n3581), .A2(n275), .B1(n2320), .B2(n278), .ZN(n2319) );
  NAND2_X1 U2649 ( .A1(n2321), .A2(n2314), .ZN(n1923) );
  NAND2_X1 U2650 ( .A1(n2321), .A2(n2316), .ZN(n1921) );
  AND2_X1 U2651 ( .A1(n2313), .A2(n2311), .ZN(n1919) );
  AND2_X1 U2652 ( .A1(n2313), .A2(n2316), .ZN(n1918) );
  AND2_X1 U2653 ( .A1(n2321), .A2(n2312), .ZN(n1925) );
  AND2_X1 U2654 ( .A1(n2321), .A2(n2311), .ZN(n1924) );
  NOR3_X1 U2655 ( .A1(ADD_RS2[0]), .A2(ADD_RS2[3]), .A3(n2317), .ZN(n2321) );
  NAND2_X1 U2656 ( .A1(n2313), .A2(n2312), .ZN(n1917) );
  NOR3_X1 U2657 ( .A1(n2322), .A2(ADD_RS2[3]), .A3(n2317), .ZN(n2313) );
  AOI221_X1 U2658 ( .B1(n281), .B2(n3709), .C1(n284), .C2(n3741), .A(n2325), 
        .ZN(n2324) );
  OAI22_X1 U2659 ( .A1(n3773), .A2(n287), .B1(n3805), .B2(n290), .ZN(n2325) );
  NAND2_X1 U2660 ( .A1(n2316), .A2(n2326), .ZN(n1932) );
  NAND2_X1 U2661 ( .A1(n2316), .A2(n2327), .ZN(n1931) );
  AND2_X1 U2662 ( .A1(n2326), .A2(n2314), .ZN(n1929) );
  AND2_X1 U2663 ( .A1(n2314), .A2(n2327), .ZN(n1928) );
  AOI221_X1 U2664 ( .B1(n293), .B2(n3837), .C1(n296), .C2(n3869), .A(n2328), 
        .ZN(n2323) );
  OAI22_X1 U2665 ( .A1(n3901), .A2(n299), .B1(n3933), .B2(n302), .ZN(n2328) );
  NAND2_X1 U2666 ( .A1(n2312), .A2(n2326), .ZN(n1937) );
  NAND2_X1 U2667 ( .A1(n2312), .A2(n2327), .ZN(n1936) );
  AND2_X1 U2668 ( .A1(n2311), .A2(n2326), .ZN(n1934) );
  NOR3_X1 U2669 ( .A1(ADD_RS2[0]), .A2(ADD_RS2[4]), .A3(n2318), .ZN(n2326) );
  AND2_X1 U2670 ( .A1(n2311), .A2(n2327), .ZN(n1933) );
  NOR3_X1 U2671 ( .A1(n2322), .A2(ADD_RS2[4]), .A3(n2318), .ZN(n2327) );
  OAI22_X1 U2672 ( .A1(n2330), .A2(n308), .B1(n2331), .B2(n311), .ZN(n2329) );
  NAND2_X1 U2673 ( .A1(n2332), .A2(n2314), .ZN(n1943) );
  NAND2_X1 U2674 ( .A1(n2333), .A2(n2314), .ZN(n1941) );
  NOR2_X1 U2675 ( .A1(n2334), .A2(n2335), .ZN(n2314) );
  AND2_X1 U2676 ( .A1(n2333), .A2(n2316), .ZN(n1938) );
  OAI22_X1 U2677 ( .A1(n2337), .A2(n317), .B1(n2338), .B2(n320), .ZN(n2336) );
  NAND2_X1 U2678 ( .A1(n2332), .A2(n2311), .ZN(n1949) );
  NAND2_X1 U2679 ( .A1(n2333), .A2(n2311), .ZN(n1947) );
  NOR2_X1 U2680 ( .A1(n2335), .A2(ADD_RS2[2]), .ZN(n2311) );
  NOR3_X1 U2681 ( .A1(ADD_RS2[3]), .A2(ADD_RS2[4]), .A3(ADD_RS2[0]), .ZN(n2333) );
  AND2_X1 U2682 ( .A1(n2315), .A2(n2316), .ZN(n1944) );
  NOR2_X1 U2683 ( .A1(n2334), .A2(ADD_RS2[1]), .ZN(n2316) );
  INV_X1 U2684 ( .A(ADD_RS2[2]), .ZN(n2334) );
  NOR3_X1 U2685 ( .A1(n2317), .A2(n2322), .A3(n2318), .ZN(n2315) );
  INV_X1 U2686 ( .A(ADD_RS2[3]), .ZN(n2318) );
  INV_X1 U2687 ( .A(ADD_RS2[4]), .ZN(n2317) );
  NOR2_X1 U2688 ( .A1(ADD_RS2[1]), .A2(ADD_RS2[2]), .ZN(n2312) );
  NOR3_X1 U2689 ( .A1(ADD_RS2[3]), .A2(ADD_RS2[4]), .A3(n2322), .ZN(n2332) );
  INV_X1 U2690 ( .A(ADD_RS2[0]), .ZN(n2322) );
  NOR3_X1 U2691 ( .A1(n2343), .A2(n2344), .A3(n2345), .ZN(n2342) );
  XNOR2_X1 U2692 ( .A(ADD_WR[1]), .B(n2335), .ZN(n2345) );
  INV_X1 U2693 ( .A(ADD_RS2[1]), .ZN(n2335) );
  XNOR2_X1 U2694 ( .A(n1907), .B(ADD_RS2[0]), .ZN(n2343) );
  XNOR2_X1 U2695 ( .A(ADD_WR[3]), .B(ADD_RS2[3]), .ZN(n2341) );
  XNOR2_X1 U2696 ( .A(ADD_WR[4]), .B(ADD_RS2[4]), .ZN(n2340) );
  XNOR2_X1 U2697 ( .A(ADD_RS2[2]), .B(ADD_WR[2]), .ZN(n2339) );
  OAI22_X1 U2698 ( .A1(n3581), .A2(n325), .B1(n2320), .B2(n328), .ZN(n2357) );
  AOI221_X1 U2699 ( .B1(n331), .B2(n3709), .C1(n334), .C2(n3741), .A(n2366), 
        .ZN(n2363) );
  OAI22_X1 U2700 ( .A1(n3773), .A2(n337), .B1(n3805), .B2(n340), .ZN(n2366) );
  AOI221_X1 U2701 ( .B1(n343), .B2(n3837), .C1(n346), .C2(n3869), .A(n2371), 
        .ZN(n2362) );
  OAI22_X1 U2702 ( .A1(n3901), .A2(n349), .B1(n3933), .B2(n352), .ZN(n2371) );
  OAI22_X1 U2703 ( .A1(n2330), .A2(n358), .B1(n2331), .B2(n361), .ZN(n2375) );
  OAI22_X1 U2704 ( .A1(n2337), .A2(n367), .B1(n2338), .B2(n370), .ZN(n2379) );
  OAI22_X1 U2705 ( .A1(n3580), .A2(n325), .B1(n2299), .B2(n328), .ZN(n2382) );
  AOI221_X1 U2706 ( .B1(n331), .B2(n3708), .C1(n334), .C2(n3740), .A(n2385), 
        .ZN(n2384) );
  OAI22_X1 U2707 ( .A1(n3772), .A2(n337), .B1(n3804), .B2(n340), .ZN(n2385) );
  AOI221_X1 U2708 ( .B1(n343), .B2(n3836), .C1(n346), .C2(n3868), .A(n2386), 
        .ZN(n2383) );
  OAI22_X1 U2709 ( .A1(n3900), .A2(n349), .B1(n3932), .B2(n352), .ZN(n2386) );
  OAI22_X1 U2710 ( .A1(n2305), .A2(n358), .B1(n2306), .B2(n361), .ZN(n2387) );
  OAI22_X1 U2711 ( .A1(n2308), .A2(n367), .B1(n2309), .B2(n370), .ZN(n2388) );
  OAI22_X1 U2712 ( .A1(n3579), .A2(n325), .B1(n2287), .B2(n328), .ZN(n2389) );
  AOI221_X1 U2713 ( .B1(n331), .B2(n3707), .C1(n334), .C2(n3739), .A(n2392), 
        .ZN(n2391) );
  OAI22_X1 U2714 ( .A1(n3771), .A2(n337), .B1(n3803), .B2(n340), .ZN(n2392) );
  AOI221_X1 U2715 ( .B1(n343), .B2(n3835), .C1(n346), .C2(n3867), .A(n2393), 
        .ZN(n2390) );
  OAI22_X1 U2716 ( .A1(n3899), .A2(n349), .B1(n3931), .B2(n352), .ZN(n2393) );
  OAI22_X1 U2717 ( .A1(n2293), .A2(n358), .B1(n2294), .B2(n361), .ZN(n2394) );
  OAI22_X1 U2718 ( .A1(n2296), .A2(n367), .B1(n2297), .B2(n370), .ZN(n2395) );
  OAI22_X1 U2719 ( .A1(n3578), .A2(n325), .B1(n2275), .B2(n328), .ZN(n2396) );
  AOI221_X1 U2720 ( .B1(n331), .B2(n3706), .C1(n334), .C2(n3738), .A(n2399), 
        .ZN(n2398) );
  OAI22_X1 U2721 ( .A1(n3770), .A2(n337), .B1(n3802), .B2(n340), .ZN(n2399) );
  AOI221_X1 U2722 ( .B1(n343), .B2(n3834), .C1(n346), .C2(n3866), .A(n2400), 
        .ZN(n2397) );
  OAI22_X1 U2723 ( .A1(n3898), .A2(n349), .B1(n3930), .B2(n352), .ZN(n2400) );
  OAI22_X1 U2724 ( .A1(n2281), .A2(n358), .B1(n2282), .B2(n361), .ZN(n2401) );
  OAI22_X1 U2725 ( .A1(n2284), .A2(n367), .B1(n2285), .B2(n370), .ZN(n2402) );
  OAI22_X1 U2726 ( .A1(n3577), .A2(n325), .B1(n2263), .B2(n328), .ZN(n2403) );
  AOI221_X1 U2727 ( .B1(n331), .B2(n3705), .C1(n334), .C2(n3737), .A(n2406), 
        .ZN(n2405) );
  OAI22_X1 U2728 ( .A1(n3769), .A2(n337), .B1(n3801), .B2(n340), .ZN(n2406) );
  AOI221_X1 U2729 ( .B1(n343), .B2(n3833), .C1(n346), .C2(n3865), .A(n2407), 
        .ZN(n2404) );
  OAI22_X1 U2730 ( .A1(n3897), .A2(n349), .B1(n3929), .B2(n352), .ZN(n2407) );
  OAI22_X1 U2731 ( .A1(n2269), .A2(n358), .B1(n2270), .B2(n361), .ZN(n2408) );
  OAI22_X1 U2732 ( .A1(n2272), .A2(n367), .B1(n2273), .B2(n370), .ZN(n2409) );
  OAI22_X1 U2733 ( .A1(n3576), .A2(n325), .B1(n2251), .B2(n328), .ZN(n2410) );
  AOI221_X1 U2734 ( .B1(n331), .B2(n3704), .C1(n334), .C2(n3736), .A(n2413), 
        .ZN(n2412) );
  OAI22_X1 U2735 ( .A1(n3768), .A2(n337), .B1(n3800), .B2(n340), .ZN(n2413) );
  AOI221_X1 U2736 ( .B1(n343), .B2(n3832), .C1(n346), .C2(n3864), .A(n2414), 
        .ZN(n2411) );
  OAI22_X1 U2737 ( .A1(n3896), .A2(n349), .B1(n3928), .B2(n352), .ZN(n2414) );
  OAI22_X1 U2738 ( .A1(n2257), .A2(n358), .B1(n2258), .B2(n361), .ZN(n2415) );
  OAI22_X1 U2739 ( .A1(n2260), .A2(n367), .B1(n2261), .B2(n370), .ZN(n2416) );
  OAI22_X1 U2740 ( .A1(n3575), .A2(n325), .B1(n2239), .B2(n328), .ZN(n2417) );
  AOI221_X1 U2741 ( .B1(n331), .B2(n3703), .C1(n334), .C2(n3735), .A(n2420), 
        .ZN(n2419) );
  OAI22_X1 U2742 ( .A1(n3767), .A2(n337), .B1(n3799), .B2(n340), .ZN(n2420) );
  AOI221_X1 U2743 ( .B1(n343), .B2(n3831), .C1(n346), .C2(n3863), .A(n2421), 
        .ZN(n2418) );
  OAI22_X1 U2744 ( .A1(n3895), .A2(n349), .B1(n3927), .B2(n352), .ZN(n2421) );
  OAI22_X1 U2745 ( .A1(n2245), .A2(n358), .B1(n2246), .B2(n361), .ZN(n2422) );
  OAI22_X1 U2746 ( .A1(n2248), .A2(n367), .B1(n2249), .B2(n370), .ZN(n2423) );
  OAI22_X1 U2747 ( .A1(n3574), .A2(n325), .B1(n2227), .B2(n328), .ZN(n2424) );
  AOI221_X1 U2748 ( .B1(n331), .B2(n3702), .C1(n334), .C2(n3734), .A(n2427), 
        .ZN(n2426) );
  OAI22_X1 U2749 ( .A1(n3766), .A2(n337), .B1(n3798), .B2(n340), .ZN(n2427) );
  AOI221_X1 U2750 ( .B1(n343), .B2(n3830), .C1(n346), .C2(n3862), .A(n2428), 
        .ZN(n2425) );
  OAI22_X1 U2751 ( .A1(n3894), .A2(n349), .B1(n3926), .B2(n352), .ZN(n2428) );
  OAI22_X1 U2752 ( .A1(n2233), .A2(n358), .B1(n2234), .B2(n361), .ZN(n2429) );
  OAI22_X1 U2753 ( .A1(n2236), .A2(n367), .B1(n2237), .B2(n370), .ZN(n2430) );
  OAI22_X1 U2754 ( .A1(n3573), .A2(n324), .B1(n2215), .B2(n327), .ZN(n2431) );
  AOI221_X1 U2755 ( .B1(n330), .B2(n3701), .C1(n333), .C2(n3733), .A(n2434), 
        .ZN(n2433) );
  OAI22_X1 U2756 ( .A1(n3765), .A2(n336), .B1(n3797), .B2(n339), .ZN(n2434) );
  AOI221_X1 U2757 ( .B1(n342), .B2(n3829), .C1(n345), .C2(n3861), .A(n2435), 
        .ZN(n2432) );
  OAI22_X1 U2758 ( .A1(n3893), .A2(n348), .B1(n3925), .B2(n351), .ZN(n2435) );
  OAI22_X1 U2759 ( .A1(n2221), .A2(n357), .B1(n2222), .B2(n360), .ZN(n2436) );
  OAI22_X1 U2760 ( .A1(n2224), .A2(n366), .B1(n2225), .B2(n369), .ZN(n2437) );
  OAI22_X1 U2761 ( .A1(n3572), .A2(n324), .B1(n2203), .B2(n327), .ZN(n2438) );
  AOI221_X1 U2762 ( .B1(n330), .B2(n3700), .C1(n333), .C2(n3732), .A(n2441), 
        .ZN(n2440) );
  OAI22_X1 U2763 ( .A1(n3764), .A2(n336), .B1(n3796), .B2(n339), .ZN(n2441) );
  AOI221_X1 U2764 ( .B1(n342), .B2(n3828), .C1(n345), .C2(n3860), .A(n2442), 
        .ZN(n2439) );
  OAI22_X1 U2765 ( .A1(n3892), .A2(n348), .B1(n3924), .B2(n351), .ZN(n2442) );
  OAI22_X1 U2766 ( .A1(n2209), .A2(n357), .B1(n2210), .B2(n360), .ZN(n2443) );
  OAI22_X1 U2767 ( .A1(n2212), .A2(n366), .B1(n2213), .B2(n369), .ZN(n2444) );
  OAI22_X1 U2768 ( .A1(n3571), .A2(n324), .B1(n2191), .B2(n327), .ZN(n2445) );
  AOI221_X1 U2769 ( .B1(n330), .B2(n3699), .C1(n333), .C2(n3731), .A(n2448), 
        .ZN(n2447) );
  OAI22_X1 U2770 ( .A1(n3763), .A2(n336), .B1(n3795), .B2(n339), .ZN(n2448) );
  AOI221_X1 U2771 ( .B1(n342), .B2(n3827), .C1(n345), .C2(n3859), .A(n2449), 
        .ZN(n2446) );
  OAI22_X1 U2772 ( .A1(n3891), .A2(n348), .B1(n3923), .B2(n351), .ZN(n2449) );
  OAI22_X1 U2773 ( .A1(n2197), .A2(n357), .B1(n2198), .B2(n360), .ZN(n2450) );
  OAI22_X1 U2774 ( .A1(n2200), .A2(n366), .B1(n2201), .B2(n369), .ZN(n2451) );
  OAI22_X1 U2775 ( .A1(n3570), .A2(n324), .B1(n2179), .B2(n327), .ZN(n2452) );
  AOI221_X1 U2776 ( .B1(n330), .B2(n3698), .C1(n333), .C2(n3730), .A(n2455), 
        .ZN(n2454) );
  OAI22_X1 U2777 ( .A1(n3762), .A2(n336), .B1(n3794), .B2(n339), .ZN(n2455) );
  AOI221_X1 U2778 ( .B1(n342), .B2(n3826), .C1(n345), .C2(n3858), .A(n2456), 
        .ZN(n2453) );
  OAI22_X1 U2779 ( .A1(n3890), .A2(n348), .B1(n3922), .B2(n351), .ZN(n2456) );
  OAI22_X1 U2780 ( .A1(n2185), .A2(n357), .B1(n2186), .B2(n360), .ZN(n2457) );
  OAI22_X1 U2781 ( .A1(n2188), .A2(n366), .B1(n2189), .B2(n369), .ZN(n2458) );
  OAI22_X1 U2782 ( .A1(n3569), .A2(n324), .B1(n2167), .B2(n327), .ZN(n2459) );
  AOI221_X1 U2783 ( .B1(n330), .B2(n3697), .C1(n333), .C2(n3729), .A(n2462), 
        .ZN(n2461) );
  OAI22_X1 U2784 ( .A1(n3761), .A2(n336), .B1(n3793), .B2(n339), .ZN(n2462) );
  AOI221_X1 U2785 ( .B1(n342), .B2(n3825), .C1(n345), .C2(n3857), .A(n2463), 
        .ZN(n2460) );
  OAI22_X1 U2786 ( .A1(n3889), .A2(n348), .B1(n3921), .B2(n351), .ZN(n2463) );
  OAI22_X1 U2787 ( .A1(n2173), .A2(n357), .B1(n2174), .B2(n360), .ZN(n2464) );
  OAI22_X1 U2788 ( .A1(n2176), .A2(n366), .B1(n2177), .B2(n369), .ZN(n2465) );
  OAI22_X1 U2789 ( .A1(n3568), .A2(n324), .B1(n2155), .B2(n327), .ZN(n2466) );
  AOI221_X1 U2790 ( .B1(n330), .B2(n3696), .C1(n333), .C2(n3728), .A(n2469), 
        .ZN(n2468) );
  OAI22_X1 U2791 ( .A1(n3760), .A2(n336), .B1(n3792), .B2(n339), .ZN(n2469) );
  AOI221_X1 U2792 ( .B1(n342), .B2(n3824), .C1(n345), .C2(n3856), .A(n2470), 
        .ZN(n2467) );
  OAI22_X1 U2793 ( .A1(n3888), .A2(n348), .B1(n3920), .B2(n351), .ZN(n2470) );
  OAI22_X1 U2794 ( .A1(n2161), .A2(n357), .B1(n2162), .B2(n360), .ZN(n2471) );
  OAI22_X1 U2795 ( .A1(n2164), .A2(n366), .B1(n2165), .B2(n369), .ZN(n2472) );
  OAI22_X1 U2796 ( .A1(n3567), .A2(n324), .B1(n2143), .B2(n327), .ZN(n2473) );
  AOI221_X1 U2797 ( .B1(n330), .B2(n3695), .C1(n333), .C2(n3727), .A(n2476), 
        .ZN(n2475) );
  OAI22_X1 U2798 ( .A1(n3759), .A2(n336), .B1(n3791), .B2(n339), .ZN(n2476) );
  AOI221_X1 U2799 ( .B1(n342), .B2(n3823), .C1(n345), .C2(n3855), .A(n2477), 
        .ZN(n2474) );
  OAI22_X1 U2800 ( .A1(n3887), .A2(n348), .B1(n3919), .B2(n351), .ZN(n2477) );
  OAI22_X1 U2801 ( .A1(n2149), .A2(n357), .B1(n2150), .B2(n360), .ZN(n2478) );
  OAI22_X1 U2802 ( .A1(n2152), .A2(n366), .B1(n2153), .B2(n369), .ZN(n2479) );
  OAI22_X1 U2803 ( .A1(n3566), .A2(n324), .B1(n2131), .B2(n327), .ZN(n2480) );
  AOI221_X1 U2804 ( .B1(n330), .B2(n3694), .C1(n333), .C2(n3726), .A(n2483), 
        .ZN(n2482) );
  OAI22_X1 U2805 ( .A1(n3758), .A2(n336), .B1(n3790), .B2(n339), .ZN(n2483) );
  AOI221_X1 U2806 ( .B1(n342), .B2(n3822), .C1(n345), .C2(n3854), .A(n2484), 
        .ZN(n2481) );
  OAI22_X1 U2807 ( .A1(n3886), .A2(n348), .B1(n3918), .B2(n351), .ZN(n2484) );
  OAI22_X1 U2808 ( .A1(n2137), .A2(n357), .B1(n2138), .B2(n360), .ZN(n2485) );
  OAI22_X1 U2809 ( .A1(n2140), .A2(n366), .B1(n2141), .B2(n369), .ZN(n2486) );
  OAI22_X1 U2810 ( .A1(n3565), .A2(n324), .B1(n2119), .B2(n327), .ZN(n2487) );
  AOI221_X1 U2811 ( .B1(n330), .B2(n3693), .C1(n333), .C2(n3725), .A(n2490), 
        .ZN(n2489) );
  OAI22_X1 U2812 ( .A1(n3757), .A2(n336), .B1(n3789), .B2(n339), .ZN(n2490) );
  AOI221_X1 U2813 ( .B1(n342), .B2(n3821), .C1(n345), .C2(n3853), .A(n2491), 
        .ZN(n2488) );
  OAI22_X1 U2814 ( .A1(n3885), .A2(n348), .B1(n3917), .B2(n351), .ZN(n2491) );
  OAI22_X1 U2815 ( .A1(n2125), .A2(n357), .B1(n2126), .B2(n360), .ZN(n2492) );
  OAI22_X1 U2816 ( .A1(n2128), .A2(n366), .B1(n2129), .B2(n369), .ZN(n2493) );
  OAI22_X1 U2817 ( .A1(n3564), .A2(n324), .B1(n2107), .B2(n327), .ZN(n2494) );
  AOI221_X1 U2818 ( .B1(n330), .B2(n3692), .C1(n333), .C2(n3724), .A(n2497), 
        .ZN(n2496) );
  OAI22_X1 U2819 ( .A1(n3756), .A2(n336), .B1(n3788), .B2(n339), .ZN(n2497) );
  AOI221_X1 U2820 ( .B1(n342), .B2(n3820), .C1(n345), .C2(n3852), .A(n2498), 
        .ZN(n2495) );
  OAI22_X1 U2821 ( .A1(n3884), .A2(n348), .B1(n3916), .B2(n351), .ZN(n2498) );
  OAI22_X1 U2822 ( .A1(n2113), .A2(n357), .B1(n2114), .B2(n360), .ZN(n2499) );
  OAI22_X1 U2823 ( .A1(n2116), .A2(n366), .B1(n2117), .B2(n369), .ZN(n2500) );
  OAI22_X1 U2824 ( .A1(n3563), .A2(n324), .B1(n2095), .B2(n327), .ZN(n2501) );
  AOI221_X1 U2825 ( .B1(n330), .B2(n3691), .C1(n333), .C2(n3723), .A(n2504), 
        .ZN(n2503) );
  OAI22_X1 U2826 ( .A1(n3755), .A2(n336), .B1(n3787), .B2(n339), .ZN(n2504) );
  AOI221_X1 U2827 ( .B1(n342), .B2(n3819), .C1(n345), .C2(n3851), .A(n2505), 
        .ZN(n2502) );
  OAI22_X1 U2828 ( .A1(n3883), .A2(n348), .B1(n3915), .B2(n351), .ZN(n2505) );
  OAI22_X1 U2829 ( .A1(n2101), .A2(n357), .B1(n2102), .B2(n360), .ZN(n2506) );
  OAI22_X1 U2830 ( .A1(n2104), .A2(n366), .B1(n2105), .B2(n369), .ZN(n2507) );
  OAI22_X1 U2831 ( .A1(n3562), .A2(n324), .B1(n2083), .B2(n327), .ZN(n2508) );
  AOI221_X1 U2832 ( .B1(n330), .B2(n3690), .C1(n333), .C2(n3722), .A(n2511), 
        .ZN(n2510) );
  OAI22_X1 U2833 ( .A1(n3754), .A2(n336), .B1(n3786), .B2(n339), .ZN(n2511) );
  AOI221_X1 U2834 ( .B1(n342), .B2(n3818), .C1(n345), .C2(n3850), .A(n2512), 
        .ZN(n2509) );
  OAI22_X1 U2835 ( .A1(n3882), .A2(n348), .B1(n3914), .B2(n351), .ZN(n2512) );
  OAI22_X1 U2836 ( .A1(n2089), .A2(n357), .B1(n2090), .B2(n360), .ZN(n2513) );
  OAI22_X1 U2837 ( .A1(n2092), .A2(n366), .B1(n2093), .B2(n369), .ZN(n2514) );
  OAI22_X1 U2838 ( .A1(n3561), .A2(n323), .B1(n2071), .B2(n326), .ZN(n2515) );
  AOI221_X1 U2839 ( .B1(n329), .B2(n3689), .C1(n332), .C2(n3721), .A(n2518), 
        .ZN(n2517) );
  OAI22_X1 U2840 ( .A1(n3753), .A2(n335), .B1(n3785), .B2(n338), .ZN(n2518) );
  AOI221_X1 U2841 ( .B1(n341), .B2(n3817), .C1(n344), .C2(n3849), .A(n2519), 
        .ZN(n2516) );
  OAI22_X1 U2842 ( .A1(n3881), .A2(n347), .B1(n3913), .B2(n350), .ZN(n2519) );
  OAI22_X1 U2843 ( .A1(n2077), .A2(n356), .B1(n2078), .B2(n359), .ZN(n2520) );
  OAI22_X1 U2844 ( .A1(n2080), .A2(n365), .B1(n2081), .B2(n368), .ZN(n2521) );
  OAI22_X1 U2845 ( .A1(n3560), .A2(n323), .B1(n2059), .B2(n326), .ZN(n2522) );
  AOI221_X1 U2846 ( .B1(n329), .B2(n3688), .C1(n332), .C2(n3720), .A(n2525), 
        .ZN(n2524) );
  OAI22_X1 U2847 ( .A1(n3752), .A2(n335), .B1(n3784), .B2(n338), .ZN(n2525) );
  AOI221_X1 U2848 ( .B1(n341), .B2(n3816), .C1(n344), .C2(n3848), .A(n2526), 
        .ZN(n2523) );
  OAI22_X1 U2849 ( .A1(n3880), .A2(n347), .B1(n3912), .B2(n350), .ZN(n2526) );
  OAI22_X1 U2850 ( .A1(n2065), .A2(n356), .B1(n2066), .B2(n359), .ZN(n2527) );
  OAI22_X1 U2851 ( .A1(n2068), .A2(n365), .B1(n2069), .B2(n368), .ZN(n2528) );
  OAI22_X1 U2852 ( .A1(n3559), .A2(n323), .B1(n2047), .B2(n326), .ZN(n2529) );
  AOI221_X1 U2853 ( .B1(n329), .B2(n3687), .C1(n332), .C2(n3719), .A(n2532), 
        .ZN(n2531) );
  OAI22_X1 U2854 ( .A1(n3751), .A2(n335), .B1(n3783), .B2(n338), .ZN(n2532) );
  AOI221_X1 U2855 ( .B1(n341), .B2(n3815), .C1(n344), .C2(n3847), .A(n2533), 
        .ZN(n2530) );
  OAI22_X1 U2856 ( .A1(n3879), .A2(n347), .B1(n3911), .B2(n350), .ZN(n2533) );
  OAI22_X1 U2857 ( .A1(n2053), .A2(n356), .B1(n2054), .B2(n359), .ZN(n2534) );
  OAI22_X1 U2858 ( .A1(n2056), .A2(n365), .B1(n2057), .B2(n368), .ZN(n2535) );
  OAI22_X1 U2859 ( .A1(n2982), .A2(n323), .B1(n2035), .B2(n326), .ZN(n2536) );
  AOI221_X1 U2860 ( .B1(n329), .B2(n3686), .C1(n332), .C2(n3718), .A(n2539), 
        .ZN(n2538) );
  OAI22_X1 U2861 ( .A1(n3750), .A2(n335), .B1(n3782), .B2(n338), .ZN(n2539) );
  AOI221_X1 U2862 ( .B1(n341), .B2(n3814), .C1(n344), .C2(n3846), .A(n2540), 
        .ZN(n2537) );
  OAI22_X1 U2863 ( .A1(n3878), .A2(n347), .B1(n3910), .B2(n350), .ZN(n2540) );
  OAI22_X1 U2864 ( .A1(n2041), .A2(n356), .B1(n2042), .B2(n359), .ZN(n2541) );
  OAI22_X1 U2865 ( .A1(n2044), .A2(n365), .B1(n2045), .B2(n368), .ZN(n2542) );
  OAI22_X1 U2866 ( .A1(n2981), .A2(n323), .B1(n2023), .B2(n326), .ZN(n2543) );
  AOI221_X1 U2867 ( .B1(n329), .B2(n3685), .C1(n332), .C2(n3717), .A(n2546), 
        .ZN(n2545) );
  OAI22_X1 U2868 ( .A1(n3749), .A2(n335), .B1(n3781), .B2(n338), .ZN(n2546) );
  AOI221_X1 U2869 ( .B1(n341), .B2(n3813), .C1(n344), .C2(n3845), .A(n2547), 
        .ZN(n2544) );
  OAI22_X1 U2870 ( .A1(n3877), .A2(n347), .B1(n3909), .B2(n350), .ZN(n2547) );
  OAI22_X1 U2871 ( .A1(n2029), .A2(n356), .B1(n2030), .B2(n359), .ZN(n2548) );
  OAI22_X1 U2872 ( .A1(n2032), .A2(n365), .B1(n2033), .B2(n368), .ZN(n2549) );
  OAI22_X1 U2873 ( .A1(n2980), .A2(n323), .B1(n2011), .B2(n326), .ZN(n2550) );
  AOI221_X1 U2874 ( .B1(n329), .B2(n3684), .C1(n332), .C2(n3716), .A(n2553), 
        .ZN(n2552) );
  OAI22_X1 U2875 ( .A1(n3748), .A2(n335), .B1(n3780), .B2(n338), .ZN(n2553) );
  AOI221_X1 U2876 ( .B1(n341), .B2(n3812), .C1(n344), .C2(n3844), .A(n2554), 
        .ZN(n2551) );
  OAI22_X1 U2877 ( .A1(n3876), .A2(n347), .B1(n3908), .B2(n350), .ZN(n2554) );
  OAI22_X1 U2878 ( .A1(n2017), .A2(n356), .B1(n2018), .B2(n359), .ZN(n2555) );
  OAI22_X1 U2879 ( .A1(n2020), .A2(n365), .B1(n2021), .B2(n368), .ZN(n2556) );
  OAI22_X1 U2880 ( .A1(n2979), .A2(n323), .B1(n1999), .B2(n326), .ZN(n2557) );
  AOI221_X1 U2881 ( .B1(n329), .B2(n3683), .C1(n332), .C2(n3715), .A(n2560), 
        .ZN(n2559) );
  OAI22_X1 U2882 ( .A1(n3747), .A2(n335), .B1(n3779), .B2(n338), .ZN(n2560) );
  AOI221_X1 U2883 ( .B1(n341), .B2(n3811), .C1(n344), .C2(n3843), .A(n2561), 
        .ZN(n2558) );
  OAI22_X1 U2884 ( .A1(n3875), .A2(n347), .B1(n3907), .B2(n350), .ZN(n2561) );
  OAI22_X1 U2885 ( .A1(n2005), .A2(n356), .B1(n2006), .B2(n359), .ZN(n2562) );
  OAI22_X1 U2886 ( .A1(n2008), .A2(n365), .B1(n2009), .B2(n368), .ZN(n2563) );
  OAI22_X1 U2887 ( .A1(n2978), .A2(n323), .B1(n1987), .B2(n326), .ZN(n2564) );
  AOI221_X1 U2888 ( .B1(n329), .B2(n3682), .C1(n332), .C2(n3714), .A(n2567), 
        .ZN(n2566) );
  OAI22_X1 U2889 ( .A1(n3746), .A2(n335), .B1(n3778), .B2(n338), .ZN(n2567) );
  AOI221_X1 U2890 ( .B1(n341), .B2(n3810), .C1(n344), .C2(n3842), .A(n2568), 
        .ZN(n2565) );
  OAI22_X1 U2891 ( .A1(n3874), .A2(n347), .B1(n3906), .B2(n350), .ZN(n2568) );
  OAI22_X1 U2892 ( .A1(n1993), .A2(n356), .B1(n1994), .B2(n359), .ZN(n2569) );
  OAI22_X1 U2893 ( .A1(n1996), .A2(n365), .B1(n1997), .B2(n368), .ZN(n2570) );
  OAI22_X1 U2894 ( .A1(n2977), .A2(n323), .B1(n1975), .B2(n326), .ZN(n2571) );
  AOI221_X1 U2895 ( .B1(n329), .B2(n3681), .C1(n332), .C2(n3713), .A(n2574), 
        .ZN(n2573) );
  OAI22_X1 U2896 ( .A1(n3745), .A2(n335), .B1(n3777), .B2(n338), .ZN(n2574) );
  AOI221_X1 U2897 ( .B1(n341), .B2(n3809), .C1(n344), .C2(n3841), .A(n2575), 
        .ZN(n2572) );
  OAI22_X1 U2898 ( .A1(n3873), .A2(n347), .B1(n3905), .B2(n350), .ZN(n2575) );
  OAI22_X1 U2899 ( .A1(n1981), .A2(n356), .B1(n1982), .B2(n359), .ZN(n2576) );
  OAI22_X1 U2900 ( .A1(n1984), .A2(n365), .B1(n1985), .B2(n368), .ZN(n2577) );
  OAI22_X1 U2901 ( .A1(n2976), .A2(n323), .B1(n1963), .B2(n326), .ZN(n2578) );
  AOI221_X1 U2902 ( .B1(n329), .B2(n3680), .C1(n332), .C2(n3712), .A(n2581), 
        .ZN(n2580) );
  OAI22_X1 U2903 ( .A1(n3744), .A2(n335), .B1(n3776), .B2(n338), .ZN(n2581) );
  AOI221_X1 U2904 ( .B1(n341), .B2(n3808), .C1(n344), .C2(n3840), .A(n2582), 
        .ZN(n2579) );
  OAI22_X1 U2905 ( .A1(n3872), .A2(n347), .B1(n3904), .B2(n350), .ZN(n2582) );
  OAI22_X1 U2906 ( .A1(n1969), .A2(n356), .B1(n1970), .B2(n359), .ZN(n2583) );
  OAI22_X1 U2907 ( .A1(n1972), .A2(n365), .B1(n1973), .B2(n368), .ZN(n2584) );
  OAI22_X1 U2908 ( .A1(n2975), .A2(n323), .B1(n1951), .B2(n326), .ZN(n2585) );
  AOI221_X1 U2909 ( .B1(n329), .B2(n3679), .C1(n332), .C2(n3711), .A(n2588), 
        .ZN(n2587) );
  OAI22_X1 U2910 ( .A1(n3743), .A2(n335), .B1(n3775), .B2(n338), .ZN(n2588) );
  AOI221_X1 U2911 ( .B1(n341), .B2(n3807), .C1(n344), .C2(n3839), .A(n2589), 
        .ZN(n2586) );
  OAI22_X1 U2912 ( .A1(n3871), .A2(n347), .B1(n3903), .B2(n350), .ZN(n2589) );
  OAI22_X1 U2913 ( .A1(n1957), .A2(n356), .B1(n1958), .B2(n359), .ZN(n2590) );
  OAI22_X1 U2914 ( .A1(n1960), .A2(n365), .B1(n1961), .B2(n368), .ZN(n2591) );
  AND2_X1 U2915 ( .A1(n2592), .A2(n2593), .ZN(n2349) );
  AND2_X1 U2916 ( .A1(n2592), .A2(n2594), .ZN(n2348) );
  NAND2_X1 U2917 ( .A1(n2595), .A2(n2596), .ZN(n2347) );
  NAND2_X1 U2918 ( .A1(n2597), .A2(n2593), .ZN(n2346) );
  AND2_X1 U2919 ( .A1(n2597), .A2(n2594), .ZN(n2353) );
  AND2_X1 U2920 ( .A1(n2597), .A2(n2596), .ZN(n2352) );
  NAND2_X1 U2921 ( .A1(n2592), .A2(n2596), .ZN(n2351) );
  NAND2_X1 U2922 ( .A1(n2592), .A2(n2598), .ZN(n2350) );
  NOR3_X1 U2923 ( .A1(n2599), .A2(ADD_RS1[0]), .A3(n2600), .ZN(n2592) );
  OAI22_X1 U2924 ( .A1(n2974), .A2(n323), .B1(n1922), .B2(n326), .ZN(n2601) );
  NAND2_X1 U2925 ( .A1(n2602), .A2(n2596), .ZN(n2359) );
  NAND2_X1 U2926 ( .A1(n2602), .A2(n2598), .ZN(n2358) );
  AND2_X1 U2927 ( .A1(n2595), .A2(n2593), .ZN(n2356) );
  AND2_X1 U2928 ( .A1(n2595), .A2(n2598), .ZN(n2355) );
  AND2_X1 U2929 ( .A1(n2602), .A2(n2594), .ZN(n2361) );
  AND2_X1 U2930 ( .A1(n2602), .A2(n2593), .ZN(n2360) );
  NOR3_X1 U2931 ( .A1(ADD_RS1[0]), .A2(ADD_RS1[3]), .A3(n2599), .ZN(n2602) );
  NAND2_X1 U2932 ( .A1(n2595), .A2(n2594), .ZN(n2354) );
  NOR3_X1 U2933 ( .A1(n2603), .A2(ADD_RS1[3]), .A3(n2599), .ZN(n2595) );
  AOI221_X1 U2934 ( .B1(n329), .B2(n3678), .C1(n332), .C2(n3710), .A(n2606), 
        .ZN(n2605) );
  OAI22_X1 U2935 ( .A1(n3742), .A2(n335), .B1(n3774), .B2(n338), .ZN(n2606) );
  NAND2_X1 U2936 ( .A1(n2598), .A2(n2607), .ZN(n2368) );
  NAND2_X1 U2937 ( .A1(n2598), .A2(n2608), .ZN(n2367) );
  AND2_X1 U2938 ( .A1(n2607), .A2(n2596), .ZN(n2365) );
  AND2_X1 U2939 ( .A1(n2596), .A2(n2608), .ZN(n2364) );
  AOI221_X1 U2940 ( .B1(n341), .B2(n3806), .C1(n344), .C2(n3838), .A(n2609), 
        .ZN(n2604) );
  OAI22_X1 U2941 ( .A1(n3870), .A2(n347), .B1(n3902), .B2(n350), .ZN(n2609) );
  NAND2_X1 U2942 ( .A1(n2594), .A2(n2607), .ZN(n2373) );
  NAND2_X1 U2943 ( .A1(n2594), .A2(n2608), .ZN(n2372) );
  AND2_X1 U2944 ( .A1(n2593), .A2(n2607), .ZN(n2370) );
  NOR3_X1 U2945 ( .A1(ADD_RS1[0]), .A2(ADD_RS1[4]), .A3(n2600), .ZN(n2607) );
  AND2_X1 U2946 ( .A1(n2593), .A2(n2608), .ZN(n2369) );
  NOR3_X1 U2947 ( .A1(n2603), .A2(ADD_RS1[4]), .A3(n2600), .ZN(n2608) );
  OAI22_X1 U2948 ( .A1(n1940), .A2(n356), .B1(n1942), .B2(n359), .ZN(n2610) );
  NAND2_X1 U2949 ( .A1(n2611), .A2(n2596), .ZN(n2377) );
  NAND2_X1 U2950 ( .A1(n2612), .A2(n2596), .ZN(n2376) );
  NOR2_X1 U2951 ( .A1(n2613), .A2(n2614), .ZN(n2596) );
  AND2_X1 U2952 ( .A1(n2612), .A2(n2598), .ZN(n2374) );
  OAI22_X1 U2953 ( .A1(n1946), .A2(n365), .B1(n1948), .B2(n368), .ZN(n2615) );
  NAND2_X1 U2954 ( .A1(n2611), .A2(n2593), .ZN(n2381) );
  NAND2_X1 U2955 ( .A1(n2612), .A2(n2593), .ZN(n2380) );
  NOR2_X1 U2956 ( .A1(n2614), .A2(ADD_RS1[2]), .ZN(n2593) );
  NOR3_X1 U2957 ( .A1(ADD_RS1[3]), .A2(ADD_RS1[4]), .A3(ADD_RS1[0]), .ZN(n2612) );
  AND2_X1 U2958 ( .A1(n2597), .A2(n2598), .ZN(n2378) );
  NOR2_X1 U2959 ( .A1(n2613), .A2(ADD_RS1[1]), .ZN(n2598) );
  INV_X1 U2960 ( .A(ADD_RS1[2]), .ZN(n2613) );
  NOR3_X1 U2961 ( .A1(n2599), .A2(n2603), .A3(n2600), .ZN(n2597) );
  INV_X1 U2962 ( .A(ADD_RS1[3]), .ZN(n2600) );
  INV_X1 U2963 ( .A(ADD_RS1[4]), .ZN(n2599) );
  NOR2_X1 U2964 ( .A1(ADD_RS1[1]), .A2(ADD_RS1[2]), .ZN(n2594) );
  NOR3_X1 U2965 ( .A1(ADD_RS1[3]), .A2(ADD_RS1[4]), .A3(n2603), .ZN(n2611) );
  INV_X1 U2966 ( .A(ADD_RS1[0]), .ZN(n2603) );
  NOR3_X1 U2967 ( .A1(n2620), .A2(n2344), .A3(n2621), .ZN(n2619) );
  XNOR2_X1 U2968 ( .A(ADD_WR[1]), .B(n2614), .ZN(n2621) );
  INV_X1 U2969 ( .A(ADD_RS1[1]), .ZN(n2614) );
  INV_X1 U2970 ( .A(WR), .ZN(n2344) );
  XNOR2_X1 U2971 ( .A(n1907), .B(ADD_RS1[0]), .ZN(n2620) );
  XNOR2_X1 U2972 ( .A(ADD_WR[3]), .B(ADD_RS1[3]), .ZN(n2618) );
  XNOR2_X1 U2973 ( .A(ADD_WR[4]), .B(ADD_RS1[4]), .ZN(n2617) );
  XNOR2_X1 U2974 ( .A(ADD_RS1[2]), .B(ADD_WR[2]), .ZN(n2616) );
endmodule


module Decode ( CLK, RST, REG_LATCH_EN, RD1, RD2, RF_WE, ZERO_FLAG, PC_IN, 
        INS_IN, ADD_WR, DATA_WR_IN, PC_OUT, A_OUT, B_OUT, IMM_OUT, ADD_RS1_HDU, 
        ADD_RS2_HDU, ADD_WR_OUT, ADD_RS1_OUT, ADD_RS2_OUT );
  input [31:0] PC_IN;
  input [31:0] INS_IN;
  input [4:0] ADD_WR;
  input [31:0] DATA_WR_IN;
  output [31:0] PC_OUT;
  output [31:0] A_OUT;
  output [31:0] B_OUT;
  output [31:0] IMM_OUT;
  output [4:0] ADD_RS1_HDU;
  output [4:0] ADD_RS2_HDU;
  output [4:0] ADD_WR_OUT;
  output [4:0] ADD_RS1_OUT;
  output [4:0] ADD_RS2_OUT;
  input CLK, RST, REG_LATCH_EN, RD1, RD2, RF_WE, ZERO_FLAG;
  wire   sig_RST, sig_Rtype, sig_Itype, sig_Jtype, n1;
  wire   [4:0] sig_ADD_WR;
  wire   [31:0] sig_IMM;

  NOR2_X2 U2 ( .A1(ZERO_FLAG), .A2(n1), .ZN(sig_RST) );
  instruction_type ins_type ( .INST_IN(INS_IN), .Rtype(sig_Rtype), .Itype(
        sig_Itype), .Jtype(sig_Jtype) );
  instruction_decomposition ins_dec ( .INST_IN(INS_IN), .Rtype(sig_Rtype), 
        .Itype(sig_Itype), .Jtype(sig_Jtype), .ADD_RS1(ADD_RS1_HDU), .ADD_RS2(
        ADD_RS2_HDU), .ADD_WR(sig_ADD_WR), .IMM(sig_IMM) );
  regn_N32_8 regPC ( .DIN(PC_IN), .CLK(CLK), .EN(1'b1), .RST(sig_RST), .DOUT(
        PC_OUT) );
  regn_N32_7 regIMM ( .DIN(sig_IMM), .CLK(CLK), .EN(REG_LATCH_EN), .RST(
        sig_RST), .DOUT(IMM_OUT) );
  regn_N5_0 regWR ( .DIN(sig_ADD_WR), .CLK(CLK), .EN(REG_LATCH_EN), .RST(
        sig_RST), .DOUT(ADD_WR_OUT) );
  regn_N5_4 regRS1 ( .DIN(ADD_RS1_HDU), .CLK(CLK), .EN(REG_LATCH_EN), .RST(
        sig_RST), .DOUT(ADD_RS1_OUT) );
  regn_N5_3 regRS2 ( .DIN(ADD_RS2_HDU), .CLK(CLK), .EN(REG_LATCH_EN), .RST(
        sig_RST), .DOUT(ADD_RS2_OUT) );
  register_file_NBIT_ADD5_NBIT_DATA32 rf ( .CLK(CLK), .RST(RST), .ENABLE(
        REG_LATCH_EN), .RD1(RD1), .RD2(RD2), .WR(RF_WE), .ADD_WR(ADD_WR), 
        .ADD_RS1(ADD_RS1_HDU), .ADD_RS2(ADD_RS2_HDU), .DATAIN(DATA_WR_IN), 
        .OUT1(A_OUT), .OUT2(B_OUT) );
  INV_X1 U3 ( .A(RST), .ZN(n1) );
endmodule


module Branch_Cond_Unit_NBIT32 ( RST, A, .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , 
        \ALU_OPC[1] , \ALU_OPC[0] }), JUMP_TYPE, PC_SEL, ZERO );
  input [31:0] A;
  input [1:0] JUMP_TYPE;
  output [1:0] PC_SEL;
  input RST, \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] ;
  output ZERO;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n1, n2;
  wire   [3:0] ALU_OPC;

  NOR4_X1 U3 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n15) );
  NOR4_X1 U4 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n19) );
  NAND4_X1 U5 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .ZN(n11) );
  NOR4_X1 U6 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n12) );
  NOR4_X1 U7 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n13) );
  NOR4_X1 U8 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n14) );
  NAND4_X1 U9 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .ZN(n10) );
  NOR4_X1 U10 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n16) );
  NOR4_X1 U11 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n17) );
  NOR4_X1 U12 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n18) );
  NOR4_X1 U13 ( .A1(ALU_OPC[0]), .A2(n1), .A3(ALU_OPC[2]), .A4(ALU_OPC[1]), 
        .ZN(n7) );
  OAI211_X1 U14 ( .C1(n5), .C2(n6), .A(JUMP_TYPE[0]), .B(RST), .ZN(n4) );
  AND2_X1 U15 ( .A1(n7), .A2(n8), .ZN(n6) );
  NOR4_X1 U16 ( .A1(n8), .A2(n9), .A3(n7), .A4(n1), .ZN(n5) );
  NOR2_X1 U17 ( .A1(n10), .A2(n11), .ZN(n8) );
  NAND2_X1 U18 ( .A1(JUMP_TYPE[1]), .A2(RST), .ZN(n3) );
  INV_X1 U19 ( .A(ALU_OPC[3]), .ZN(n1) );
  NAND2_X1 U20 ( .A1(n3), .A2(n4), .ZN(ZERO) );
  OAI22_X1 U21 ( .A1(JUMP_TYPE[0]), .A2(n3), .B1(JUMP_TYPE[1]), .B2(n4), .ZN(
        PC_SEL[0]) );
  NOR2_X1 U22 ( .A1(n2), .A2(n3), .ZN(PC_SEL[1]) );
  INV_X1 U23 ( .A(JUMP_TYPE[0]), .ZN(n2) );
  OR2_X1 U24 ( .A1(ALU_OPC[1]), .A2(ALU_OPC[2]), .ZN(n9) );
endmodule


module ff_1 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n4, n5, n6;

  DFFR_X1 Q_reg ( .D(n4), .CK(CLK), .RN(RST), .Q(Q), .QN(n5) );
  OAI21_X1 U2 ( .B1(n5), .B2(EN), .A(n6), .ZN(n4) );
  NAND2_X1 U3 ( .A1(EN), .A2(D), .ZN(n6) );
endmodule


module regn_N2 ( DIN, CLK, EN, RST, DOUT );
  input [1:0] DIN;
  output [1:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n4, n5, n6;

  DFFR_X1 \DOUT_reg[1]  ( .D(n6), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n4) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n5), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n3) );
  OAI21_X1 U2 ( .B1(n3), .B2(EN), .A(n1), .ZN(n5) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n1) );
  OAI21_X1 U4 ( .B1(n4), .B2(EN), .A(n2), .ZN(n6) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n2) );
endmodule


module FWD_Unit ( RST, ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB, RF_WE_MEM, 
        RF_WE_WB, FWDA, FWDB );
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [4:0] ADD_WR_MEM;
  input [4:0] ADD_WR_WB;
  output [1:0] FWDA;
  output [1:0] FWDB;
  input RST, RF_WE_MEM, RF_WE_WB;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42;

  NOR2_X1 U3 ( .A1(n1), .A2(n2), .ZN(FWDB[1]) );
  AOI21_X1 U4 ( .B1(n3), .B2(n4), .A(n5), .ZN(n1) );
  INV_X1 U5 ( .A(n6), .ZN(n3) );
  NOR2_X1 U6 ( .A1(n2), .A2(n7), .ZN(FWDB[0]) );
  MUX2_X1 U7 ( .A(n6), .B(n8), .S(n5), .Z(n7) );
  AND4_X1 U8 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n5) );
  NOR2_X1 U9 ( .A1(n13), .A2(n14), .ZN(n12) );
  XOR2_X1 U10 ( .A(ADD_WR_MEM[4]), .B(ADD_RS2[4]), .Z(n14) );
  XOR2_X1 U11 ( .A(ADD_WR_MEM[3]), .B(ADD_RS2[3]), .Z(n13) );
  XNOR2_X1 U12 ( .A(ADD_RS2[1]), .B(ADD_WR_MEM[1]), .ZN(n11) );
  XNOR2_X1 U13 ( .A(ADD_RS2[2]), .B(ADD_WR_MEM[2]), .ZN(n10) );
  XNOR2_X1 U14 ( .A(ADD_RS2[0]), .B(ADD_WR_MEM[0]), .ZN(n9) );
  NAND4_X1 U15 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(n6) );
  NOR2_X1 U16 ( .A1(n19), .A2(n20), .ZN(n18) );
  XOR2_X1 U17 ( .A(ADD_WR_WB[3]), .B(ADD_RS2[3]), .Z(n20) );
  XOR2_X1 U18 ( .A(ADD_WR_WB[2]), .B(ADD_RS2[2]), .Z(n19) );
  XNOR2_X1 U19 ( .A(ADD_RS2[4]), .B(ADD_WR_WB[4]), .ZN(n17) );
  XNOR2_X1 U20 ( .A(ADD_RS2[1]), .B(ADD_WR_WB[1]), .ZN(n16) );
  XNOR2_X1 U21 ( .A(ADD_RS2[0]), .B(ADD_WR_WB[0]), .ZN(n15) );
  NOR2_X1 U22 ( .A1(n21), .A2(n2), .ZN(FWDA[1]) );
  AOI21_X1 U23 ( .B1(n22), .B2(n4), .A(n23), .ZN(n21) );
  OAI21_X1 U24 ( .B1(n24), .B2(n25), .A(RF_WE_WB), .ZN(n4) );
  OR2_X1 U25 ( .A1(ADD_WR_WB[0]), .A2(ADD_WR_WB[1]), .ZN(n25) );
  OR3_X1 U26 ( .A1(ADD_WR_WB[3]), .A2(ADD_WR_WB[4]), .A3(ADD_WR_WB[2]), .ZN(
        n24) );
  INV_X1 U27 ( .A(n26), .ZN(n22) );
  NOR2_X1 U28 ( .A1(n2), .A2(n27), .ZN(FWDA[0]) );
  MUX2_X1 U29 ( .A(n26), .B(n8), .S(n23), .Z(n27) );
  AND4_X1 U30 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n23) );
  NOR2_X1 U31 ( .A1(n32), .A2(n33), .ZN(n31) );
  XOR2_X1 U32 ( .A(ADD_WR_MEM[4]), .B(ADD_RS1[4]), .Z(n33) );
  XOR2_X1 U33 ( .A(ADD_WR_MEM[3]), .B(ADD_RS1[3]), .Z(n32) );
  XNOR2_X1 U34 ( .A(ADD_RS1[1]), .B(ADD_WR_MEM[1]), .ZN(n30) );
  XNOR2_X1 U35 ( .A(ADD_RS1[2]), .B(ADD_WR_MEM[2]), .ZN(n29) );
  XNOR2_X1 U36 ( .A(ADD_RS1[0]), .B(ADD_WR_MEM[0]), .ZN(n28) );
  INV_X1 U37 ( .A(n34), .ZN(n8) );
  OAI21_X1 U38 ( .B1(n35), .B2(n36), .A(RF_WE_MEM), .ZN(n34) );
  OR2_X1 U39 ( .A1(ADD_WR_MEM[0]), .A2(ADD_WR_MEM[1]), .ZN(n36) );
  OR3_X1 U40 ( .A1(ADD_WR_MEM[3]), .A2(ADD_WR_MEM[4]), .A3(ADD_WR_MEM[2]), 
        .ZN(n35) );
  NAND4_X1 U41 ( .A1(n37), .A2(n38), .A3(n39), .A4(n40), .ZN(n26) );
  NOR2_X1 U42 ( .A1(n41), .A2(n42), .ZN(n40) );
  XOR2_X1 U43 ( .A(ADD_WR_WB[3]), .B(ADD_RS1[3]), .Z(n42) );
  XOR2_X1 U44 ( .A(ADD_WR_WB[2]), .B(ADD_RS1[2]), .Z(n41) );
  XNOR2_X1 U45 ( .A(ADD_RS1[4]), .B(ADD_WR_WB[4]), .ZN(n39) );
  XNOR2_X1 U46 ( .A(ADD_RS1[1]), .B(ADD_WR_WB[1]), .ZN(n38) );
  XNOR2_X1 U47 ( .A(ADD_RS1[0]), .B(ADD_WR_WB[0]), .ZN(n37) );
  INV_X1 U48 ( .A(RST), .ZN(n2) );
endmodule


module mux41_NBIT32_0 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n1, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  BUF_X1 U1 ( .A(n6), .Z(n72) );
  BUF_X1 U2 ( .A(n6), .Z(n73) );
  BUF_X1 U3 ( .A(n4), .Z(n78) );
  BUF_X1 U4 ( .A(n4), .Z(n79) );
  BUF_X1 U5 ( .A(n7), .Z(n1) );
  BUF_X1 U6 ( .A(n7), .Z(n70) );
  BUF_X1 U7 ( .A(n5), .Z(n75) );
  BUF_X1 U8 ( .A(n5), .Z(n76) );
  BUF_X1 U9 ( .A(n6), .Z(n74) );
  BUF_X1 U10 ( .A(n4), .Z(n80) );
  BUF_X1 U11 ( .A(n7), .Z(n71) );
  BUF_X1 U12 ( .A(n5), .Z(n77) );
  NOR2_X1 U13 ( .A1(n81), .A2(S[1]), .ZN(n6) );
  NOR2_X1 U14 ( .A1(S[0]), .A2(S[1]), .ZN(n7) );
  AND2_X1 U15 ( .A1(S[1]), .A2(S[0]), .ZN(n4) );
  AND2_X1 U16 ( .A1(S[1]), .A2(n81), .ZN(n5) );
  INV_X1 U17 ( .A(S[0]), .ZN(n81) );
  NAND2_X1 U18 ( .A1(n44), .A2(n45), .ZN(Z[20]) );
  AOI22_X1 U19 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n45) );
  AOI22_X1 U20 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n44) );
  NAND2_X1 U21 ( .A1(n52), .A2(n53), .ZN(Z[17]) );
  AOI22_X1 U22 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n53) );
  AOI22_X1 U23 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n52) );
  NAND2_X1 U24 ( .A1(n60), .A2(n61), .ZN(Z[13]) );
  AOI22_X1 U25 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n61) );
  AOI22_X1 U26 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n60) );
  NAND2_X1 U27 ( .A1(n68), .A2(n69), .ZN(Z[0]) );
  AOI22_X1 U28 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n69) );
  AOI22_X1 U29 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n68) );
  NAND2_X1 U30 ( .A1(n12), .A2(n13), .ZN(Z[6]) );
  AOI22_X1 U31 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n13) );
  AOI22_X1 U32 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n12) );
  NAND2_X1 U33 ( .A1(n20), .A2(n21), .ZN(Z[31]) );
  AOI22_X1 U34 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n21) );
  AOI22_X1 U35 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n20) );
  NAND2_X1 U36 ( .A1(n28), .A2(n29), .ZN(Z[28]) );
  AOI22_X1 U37 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n29) );
  AOI22_X1 U38 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n28) );
  NAND2_X1 U39 ( .A1(n36), .A2(n37), .ZN(Z[24]) );
  AOI22_X1 U40 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n37) );
  AOI22_X1 U41 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n36) );
  NAND2_X1 U42 ( .A1(n42), .A2(n43), .ZN(Z[21]) );
  AOI22_X1 U43 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n43) );
  AOI22_X1 U44 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n42) );
  NAND2_X1 U45 ( .A1(n50), .A2(n51), .ZN(Z[18]) );
  AOI22_X1 U46 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n51) );
  AOI22_X1 U47 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n50) );
  NAND2_X1 U48 ( .A1(n58), .A2(n59), .ZN(Z[14]) );
  AOI22_X1 U49 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n59) );
  AOI22_X1 U50 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n58) );
  NAND2_X1 U51 ( .A1(n66), .A2(n67), .ZN(Z[10]) );
  AOI22_X1 U52 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n67) );
  AOI22_X1 U53 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n66) );
  NAND2_X1 U54 ( .A1(n10), .A2(n11), .ZN(Z[7]) );
  AOI22_X1 U55 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n11) );
  AOI22_X1 U56 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n10) );
  NAND2_X1 U57 ( .A1(n18), .A2(n19), .ZN(Z[3]) );
  AOI22_X1 U58 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n19) );
  AOI22_X1 U59 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n18) );
  NAND2_X1 U60 ( .A1(n26), .A2(n27), .ZN(Z[29]) );
  AOI22_X1 U61 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n27) );
  AOI22_X1 U62 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n26) );
  NAND2_X1 U63 ( .A1(n34), .A2(n35), .ZN(Z[25]) );
  AOI22_X1 U64 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n35) );
  AOI22_X1 U65 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n34) );
  NAND2_X1 U66 ( .A1(n40), .A2(n41), .ZN(Z[22]) );
  AOI22_X1 U67 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n41) );
  AOI22_X1 U68 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n40) );
  NAND2_X1 U69 ( .A1(n48), .A2(n49), .ZN(Z[19]) );
  AOI22_X1 U70 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n49) );
  AOI22_X1 U71 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n48) );
  NAND2_X1 U72 ( .A1(n56), .A2(n57), .ZN(Z[15]) );
  AOI22_X1 U73 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n57) );
  AOI22_X1 U74 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n56) );
  NAND2_X1 U75 ( .A1(n64), .A2(n65), .ZN(Z[11]) );
  AOI22_X1 U76 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n65) );
  AOI22_X1 U77 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n64) );
  NAND2_X1 U78 ( .A1(n8), .A2(n9), .ZN(Z[8]) );
  AOI22_X1 U79 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n9) );
  AOI22_X1 U80 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n8) );
  NAND2_X1 U81 ( .A1(n16), .A2(n17), .ZN(Z[4]) );
  AOI22_X1 U82 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n17) );
  AOI22_X1 U83 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n16) );
  NAND2_X1 U84 ( .A1(n24), .A2(n25), .ZN(Z[2]) );
  AOI22_X1 U85 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n25) );
  AOI22_X1 U86 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n24) );
  NAND2_X1 U87 ( .A1(n32), .A2(n33), .ZN(Z[26]) );
  AOI22_X1 U88 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n33) );
  AOI22_X1 U89 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n32) );
  NAND2_X1 U90 ( .A1(n38), .A2(n39), .ZN(Z[23]) );
  AOI22_X1 U91 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n39) );
  AOI22_X1 U92 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n38) );
  NAND2_X1 U93 ( .A1(n46), .A2(n47), .ZN(Z[1]) );
  AOI22_X1 U94 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n47) );
  AOI22_X1 U95 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n46) );
  NAND2_X1 U96 ( .A1(n54), .A2(n55), .ZN(Z[16]) );
  AOI22_X1 U97 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n55) );
  AOI22_X1 U98 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n54) );
  NAND2_X1 U99 ( .A1(n62), .A2(n63), .ZN(Z[12]) );
  AOI22_X1 U100 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n63) );
  AOI22_X1 U101 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n62) );
  NAND2_X1 U102 ( .A1(n2), .A2(n3), .ZN(Z[9]) );
  AOI22_X1 U103 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n3) );
  AOI22_X1 U104 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n2) );
  NAND2_X1 U105 ( .A1(n14), .A2(n15), .ZN(Z[5]) );
  AOI22_X1 U106 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n15) );
  AOI22_X1 U107 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n14) );
  NAND2_X1 U108 ( .A1(n22), .A2(n23), .ZN(Z[30]) );
  AOI22_X1 U109 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n23) );
  AOI22_X1 U110 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n22) );
  NAND2_X1 U111 ( .A1(n30), .A2(n31), .ZN(Z[27]) );
  AOI22_X1 U112 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n31) );
  AOI22_X1 U113 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n30) );
endmodule


module mux41_NBIT32_4 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149;

  BUF_X1 U1 ( .A(n145), .Z(n72) );
  BUF_X1 U2 ( .A(n145), .Z(n73) );
  BUF_X1 U3 ( .A(n147), .Z(n78) );
  BUF_X1 U4 ( .A(n147), .Z(n79) );
  BUF_X1 U5 ( .A(n144), .Z(n1) );
  BUF_X1 U6 ( .A(n144), .Z(n70) );
  BUF_X1 U7 ( .A(n146), .Z(n75) );
  BUF_X1 U8 ( .A(n146), .Z(n76) );
  BUF_X1 U9 ( .A(n145), .Z(n74) );
  BUF_X1 U10 ( .A(n147), .Z(n80) );
  BUF_X1 U11 ( .A(n144), .Z(n71) );
  BUF_X1 U12 ( .A(n146), .Z(n77) );
  NOR2_X1 U13 ( .A1(n81), .A2(S[1]), .ZN(n145) );
  NOR2_X1 U14 ( .A1(S[0]), .A2(S[1]), .ZN(n144) );
  AND2_X1 U15 ( .A1(S[1]), .A2(S[0]), .ZN(n147) );
  AND2_X1 U16 ( .A1(S[1]), .A2(n81), .ZN(n146) );
  INV_X1 U17 ( .A(S[0]), .ZN(n81) );
  NAND2_X1 U18 ( .A1(n135), .A2(n134), .ZN(Z[4]) );
  AOI22_X1 U19 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n134) );
  AOI22_X1 U20 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n135) );
  NAND2_X1 U21 ( .A1(n83), .A2(n82), .ZN(Z[0]) );
  AOI22_X1 U22 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n82) );
  AOI22_X1 U23 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n83) );
  NAND2_X1 U24 ( .A1(n143), .A2(n142), .ZN(Z[8]) );
  AOI22_X1 U25 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n142) );
  AOI22_X1 U26 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n143) );
  NAND2_X1 U27 ( .A1(n97), .A2(n96), .ZN(Z[16]) );
  AOI22_X1 U28 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n96) );
  AOI22_X1 U29 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n97) );
  NAND2_X1 U30 ( .A1(n89), .A2(n88), .ZN(Z[12]) );
  AOI22_X1 U31 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n88) );
  AOI22_X1 U32 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n89) );
  NAND2_X1 U33 ( .A1(n115), .A2(n114), .ZN(Z[24]) );
  AOI22_X1 U34 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n114) );
  AOI22_X1 U35 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n115) );
  NAND2_X1 U36 ( .A1(n105), .A2(n104), .ZN(Z[1]) );
  AOI22_X1 U37 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n104) );
  AOI22_X1 U38 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n105) );
  NAND2_X1 U39 ( .A1(n137), .A2(n136), .ZN(Z[5]) );
  AOI22_X1 U40 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n136) );
  AOI22_X1 U41 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n137) );
  NAND2_X1 U42 ( .A1(n149), .A2(n148), .ZN(Z[9]) );
  AOI22_X1 U43 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n148) );
  AOI22_X1 U44 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n149) );
  NAND2_X1 U45 ( .A1(n91), .A2(n90), .ZN(Z[13]) );
  AOI22_X1 U46 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n90) );
  AOI22_X1 U47 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n91) );
  NAND2_X1 U48 ( .A1(n99), .A2(n98), .ZN(Z[17]) );
  AOI22_X1 U49 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n98) );
  AOI22_X1 U50 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n99) );
  NAND2_X1 U51 ( .A1(n117), .A2(n116), .ZN(Z[25]) );
  AOI22_X1 U52 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n116) );
  AOI22_X1 U53 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n117) );
  NAND2_X1 U54 ( .A1(n109), .A2(n108), .ZN(Z[21]) );
  AOI22_X1 U55 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n108) );
  AOI22_X1 U56 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n109) );
  NAND2_X1 U57 ( .A1(n107), .A2(n106), .ZN(Z[20]) );
  AOI22_X1 U58 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n106) );
  AOI22_X1 U59 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n107) );
  NAND2_X1 U60 ( .A1(n125), .A2(n124), .ZN(Z[29]) );
  AOI22_X1 U61 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n124) );
  AOI22_X1 U62 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n125) );
  NAND2_X1 U63 ( .A1(n123), .A2(n122), .ZN(Z[28]) );
  AOI22_X1 U64 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n122) );
  AOI22_X1 U65 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n123) );
  NAND2_X1 U66 ( .A1(n127), .A2(n126), .ZN(Z[2]) );
  AOI22_X1 U67 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n126) );
  AOI22_X1 U68 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n127) );
  NAND2_X1 U69 ( .A1(n139), .A2(n138), .ZN(Z[6]) );
  AOI22_X1 U70 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n138) );
  AOI22_X1 U71 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n139) );
  NAND2_X1 U72 ( .A1(n85), .A2(n84), .ZN(Z[10]) );
  AOI22_X1 U73 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n84) );
  AOI22_X1 U74 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n85) );
  NAND2_X1 U75 ( .A1(n93), .A2(n92), .ZN(Z[14]) );
  AOI22_X1 U76 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n92) );
  AOI22_X1 U77 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n93) );
  NAND2_X1 U78 ( .A1(n101), .A2(n100), .ZN(Z[18]) );
  AOI22_X1 U79 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n100) );
  AOI22_X1 U80 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n101) );
  NAND2_X1 U81 ( .A1(n111), .A2(n110), .ZN(Z[22]) );
  AOI22_X1 U82 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n110) );
  AOI22_X1 U83 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n111) );
  NAND2_X1 U84 ( .A1(n119), .A2(n118), .ZN(Z[26]) );
  AOI22_X1 U85 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n118) );
  AOI22_X1 U86 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n119) );
  NAND2_X1 U87 ( .A1(n129), .A2(n128), .ZN(Z[30]) );
  AOI22_X1 U88 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n128) );
  AOI22_X1 U89 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n129) );
  NAND2_X1 U90 ( .A1(n133), .A2(n132), .ZN(Z[3]) );
  AOI22_X1 U91 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n132) );
  AOI22_X1 U92 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n133) );
  NAND2_X1 U93 ( .A1(n141), .A2(n140), .ZN(Z[7]) );
  AOI22_X1 U94 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n140) );
  AOI22_X1 U95 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n141) );
  NAND2_X1 U96 ( .A1(n87), .A2(n86), .ZN(Z[11]) );
  AOI22_X1 U97 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n86) );
  AOI22_X1 U98 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n87) );
  NAND2_X1 U99 ( .A1(n95), .A2(n94), .ZN(Z[15]) );
  AOI22_X1 U100 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n94) );
  AOI22_X1 U101 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n95) );
  NAND2_X1 U102 ( .A1(n103), .A2(n102), .ZN(Z[19]) );
  AOI22_X1 U103 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n102) );
  AOI22_X1 U104 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n103) );
  NAND2_X1 U105 ( .A1(n113), .A2(n112), .ZN(Z[23]) );
  AOI22_X1 U106 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n112) );
  AOI22_X1 U107 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n113) );
  NAND2_X1 U108 ( .A1(n121), .A2(n120), .ZN(Z[27]) );
  AOI22_X1 U109 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n120) );
  AOI22_X1 U110 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n121) );
  NAND2_X1 U111 ( .A1(n131), .A2(n130), .ZN(Z[31]) );
  AOI22_X1 U112 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n130) );
  AOI22_X1 U113 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n131) );
endmodule


module mux21_NBIT32_3 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100;

  BUF_X1 U1 ( .A(n68), .Z(n1) );
  BUF_X1 U2 ( .A(n68), .Z(n2) );
  BUF_X1 U3 ( .A(n68), .Z(n3) );
  INV_X1 U4 ( .A(n69), .ZN(Z[0]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n1), .B1(B[0]), .B2(S), .ZN(n69) );
  INV_X1 U6 ( .A(n85), .ZN(Z[24]) );
  AOI22_X1 U7 ( .A1(A[24]), .A2(n2), .B1(B[24]), .B2(S), .ZN(n85) );
  INV_X1 U8 ( .A(n73), .ZN(Z[13]) );
  AOI22_X1 U9 ( .A1(A[13]), .A2(n1), .B1(B[13]), .B2(S), .ZN(n73) );
  INV_X1 U10 ( .A(n77), .ZN(Z[17]) );
  AOI22_X1 U11 ( .A1(A[17]), .A2(n1), .B1(B[17]), .B2(S), .ZN(n77) );
  INV_X1 U12 ( .A(n81), .ZN(Z[20]) );
  AOI22_X1 U13 ( .A1(A[20]), .A2(n2), .B1(B[20]), .B2(S), .ZN(n81) );
  INV_X1 U14 ( .A(n89), .ZN(Z[28]) );
  AOI22_X1 U15 ( .A1(A[28]), .A2(n2), .B1(B[28]), .B2(S), .ZN(n89) );
  INV_X1 U16 ( .A(n97), .ZN(Z[6]) );
  AOI22_X1 U17 ( .A1(A[6]), .A2(n3), .B1(B[6]), .B2(S), .ZN(n97) );
  INV_X1 U18 ( .A(n93), .ZN(Z[31]) );
  AOI22_X1 U19 ( .A1(A[31]), .A2(n3), .B1(B[31]), .B2(S), .ZN(n93) );
  INV_X1 U20 ( .A(n86), .ZN(Z[25]) );
  AOI22_X1 U21 ( .A1(A[25]), .A2(n2), .B1(B[25]), .B2(S), .ZN(n86) );
  INV_X1 U22 ( .A(n82), .ZN(Z[21]) );
  AOI22_X1 U23 ( .A1(A[21]), .A2(n2), .B1(B[21]), .B2(S), .ZN(n82) );
  INV_X1 U24 ( .A(n90), .ZN(Z[29]) );
  AOI22_X1 U25 ( .A1(A[29]), .A2(n2), .B1(B[29]), .B2(S), .ZN(n90) );
  INV_X1 U26 ( .A(n70), .ZN(Z[10]) );
  AOI22_X1 U27 ( .A1(A[10]), .A2(n1), .B1(B[10]), .B2(S), .ZN(n70) );
  INV_X1 U28 ( .A(n74), .ZN(Z[14]) );
  AOI22_X1 U29 ( .A1(A[14]), .A2(n1), .B1(B[14]), .B2(S), .ZN(n74) );
  INV_X1 U30 ( .A(n78), .ZN(Z[18]) );
  AOI22_X1 U31 ( .A1(A[18]), .A2(n1), .B1(B[18]), .B2(S), .ZN(n78) );
  INV_X1 U32 ( .A(n94), .ZN(Z[3]) );
  AOI22_X1 U33 ( .A1(A[3]), .A2(n3), .B1(B[3]), .B2(S), .ZN(n94) );
  INV_X1 U34 ( .A(n98), .ZN(Z[7]) );
  AOI22_X1 U35 ( .A1(A[7]), .A2(n3), .B1(B[7]), .B2(S), .ZN(n98) );
  INV_X1 U36 ( .A(n95), .ZN(Z[4]) );
  AOI22_X1 U37 ( .A1(A[4]), .A2(n3), .B1(B[4]), .B2(S), .ZN(n95) );
  INV_X1 U38 ( .A(n99), .ZN(Z[8]) );
  AOI22_X1 U39 ( .A1(A[8]), .A2(n3), .B1(B[8]), .B2(S), .ZN(n99) );
  INV_X1 U40 ( .A(n91), .ZN(Z[2]) );
  AOI22_X1 U41 ( .A1(A[2]), .A2(n2), .B1(B[2]), .B2(S), .ZN(n91) );
  INV_X1 U42 ( .A(n83), .ZN(Z[22]) );
  AOI22_X1 U43 ( .A1(A[22]), .A2(n2), .B1(B[22]), .B2(S), .ZN(n83) );
  INV_X1 U44 ( .A(n87), .ZN(Z[26]) );
  AOI22_X1 U45 ( .A1(A[26]), .A2(n2), .B1(B[26]), .B2(S), .ZN(n87) );
  INV_X1 U46 ( .A(n71), .ZN(Z[11]) );
  AOI22_X1 U47 ( .A1(A[11]), .A2(n1), .B1(B[11]), .B2(S), .ZN(n71) );
  INV_X1 U48 ( .A(n75), .ZN(Z[15]) );
  AOI22_X1 U49 ( .A1(A[15]), .A2(n1), .B1(B[15]), .B2(S), .ZN(n75) );
  INV_X1 U50 ( .A(n79), .ZN(Z[19]) );
  AOI22_X1 U51 ( .A1(A[19]), .A2(n1), .B1(B[19]), .B2(S), .ZN(n79) );
  INV_X1 U52 ( .A(n76), .ZN(Z[16]) );
  AOI22_X1 U53 ( .A1(A[16]), .A2(n1), .B1(B[16]), .B2(S), .ZN(n76) );
  INV_X1 U54 ( .A(n72), .ZN(Z[12]) );
  AOI22_X1 U55 ( .A1(A[12]), .A2(n1), .B1(B[12]), .B2(S), .ZN(n72) );
  INV_X1 U56 ( .A(n80), .ZN(Z[1]) );
  AOI22_X1 U57 ( .A1(A[1]), .A2(n1), .B1(B[1]), .B2(S), .ZN(n80) );
  INV_X1 U58 ( .A(n96), .ZN(Z[5]) );
  AOI22_X1 U59 ( .A1(A[5]), .A2(n3), .B1(B[5]), .B2(S), .ZN(n96) );
  INV_X1 U60 ( .A(n92), .ZN(Z[30]) );
  AOI22_X1 U61 ( .A1(A[30]), .A2(n2), .B1(B[30]), .B2(S), .ZN(n92) );
  INV_X1 U62 ( .A(n84), .ZN(Z[23]) );
  AOI22_X1 U63 ( .A1(A[23]), .A2(n2), .B1(B[23]), .B2(S), .ZN(n84) );
  INV_X1 U64 ( .A(n88), .ZN(Z[27]) );
  AOI22_X1 U65 ( .A1(A[27]), .A2(n2), .B1(B[27]), .B2(S), .ZN(n88) );
  INV_X1 U66 ( .A(n100), .ZN(Z[9]) );
  AOI22_X1 U67 ( .A1(A[9]), .A2(n3), .B1(S), .B2(B[9]), .ZN(n100) );
  INV_X1 U68 ( .A(S), .ZN(n68) );
endmodule


module mux41_NBIT32_3 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149;

  BUF_X1 U1 ( .A(n145), .Z(n72) );
  BUF_X1 U2 ( .A(n147), .Z(n78) );
  BUF_X1 U3 ( .A(n145), .Z(n73) );
  BUF_X1 U4 ( .A(n147), .Z(n79) );
  BUF_X1 U5 ( .A(n144), .Z(n1) );
  BUF_X1 U6 ( .A(n146), .Z(n75) );
  BUF_X1 U7 ( .A(n144), .Z(n70) );
  BUF_X1 U8 ( .A(n146), .Z(n76) );
  BUF_X1 U9 ( .A(n145), .Z(n74) );
  BUF_X1 U10 ( .A(n147), .Z(n80) );
  BUF_X1 U11 ( .A(n144), .Z(n71) );
  BUF_X1 U12 ( .A(n146), .Z(n77) );
  NAND2_X1 U13 ( .A1(n135), .A2(n134), .ZN(Z[4]) );
  AOI22_X1 U14 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n134) );
  AOI22_X1 U15 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n135) );
  NAND2_X1 U16 ( .A1(n83), .A2(n82), .ZN(Z[0]) );
  AOI22_X1 U17 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n82) );
  AOI22_X1 U18 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n83) );
  NAND2_X1 U19 ( .A1(n143), .A2(n142), .ZN(Z[8]) );
  AOI22_X1 U20 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n142) );
  AOI22_X1 U21 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n143) );
  NAND2_X1 U22 ( .A1(n97), .A2(n96), .ZN(Z[16]) );
  AOI22_X1 U23 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n96) );
  AOI22_X1 U24 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n97) );
  NAND2_X1 U25 ( .A1(n89), .A2(n88), .ZN(Z[12]) );
  AOI22_X1 U26 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n88) );
  AOI22_X1 U27 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n89) );
  NAND2_X1 U28 ( .A1(n115), .A2(n114), .ZN(Z[24]) );
  AOI22_X1 U29 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n114) );
  AOI22_X1 U30 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n115) );
  NAND2_X1 U31 ( .A1(n105), .A2(n104), .ZN(Z[1]) );
  AOI22_X1 U32 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n104) );
  AOI22_X1 U33 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n105) );
  NAND2_X1 U34 ( .A1(n137), .A2(n136), .ZN(Z[5]) );
  AOI22_X1 U35 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n136) );
  AOI22_X1 U36 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n137) );
  NAND2_X1 U37 ( .A1(n149), .A2(n148), .ZN(Z[9]) );
  AOI22_X1 U38 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n148) );
  AOI22_X1 U39 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n149) );
  NAND2_X1 U40 ( .A1(n91), .A2(n90), .ZN(Z[13]) );
  AOI22_X1 U41 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n90) );
  AOI22_X1 U42 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n91) );
  NAND2_X1 U43 ( .A1(n99), .A2(n98), .ZN(Z[17]) );
  AOI22_X1 U44 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n98) );
  AOI22_X1 U45 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n99) );
  NAND2_X1 U46 ( .A1(n117), .A2(n116), .ZN(Z[25]) );
  AOI22_X1 U47 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n116) );
  AOI22_X1 U48 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n117) );
  NAND2_X1 U49 ( .A1(n109), .A2(n108), .ZN(Z[21]) );
  AOI22_X1 U50 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n108) );
  AOI22_X1 U51 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n109) );
  NAND2_X1 U52 ( .A1(n107), .A2(n106), .ZN(Z[20]) );
  AOI22_X1 U53 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n106) );
  AOI22_X1 U54 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n107) );
  NAND2_X1 U55 ( .A1(n125), .A2(n124), .ZN(Z[29]) );
  AOI22_X1 U56 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n124) );
  AOI22_X1 U57 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n125) );
  NAND2_X1 U58 ( .A1(n123), .A2(n122), .ZN(Z[28]) );
  AOI22_X1 U59 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n122) );
  AOI22_X1 U60 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n123) );
  NAND2_X1 U61 ( .A1(n127), .A2(n126), .ZN(Z[2]) );
  AOI22_X1 U62 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n126) );
  AOI22_X1 U63 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n127) );
  NAND2_X1 U64 ( .A1(n139), .A2(n138), .ZN(Z[6]) );
  AOI22_X1 U65 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n138) );
  AOI22_X1 U66 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n139) );
  NAND2_X1 U67 ( .A1(n85), .A2(n84), .ZN(Z[10]) );
  AOI22_X1 U68 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n84) );
  AOI22_X1 U69 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n85) );
  NAND2_X1 U70 ( .A1(n93), .A2(n92), .ZN(Z[14]) );
  AOI22_X1 U71 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n92) );
  AOI22_X1 U72 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n93) );
  NAND2_X1 U73 ( .A1(n101), .A2(n100), .ZN(Z[18]) );
  AOI22_X1 U74 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n100) );
  AOI22_X1 U75 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n101) );
  NAND2_X1 U76 ( .A1(n111), .A2(n110), .ZN(Z[22]) );
  AOI22_X1 U77 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n110) );
  AOI22_X1 U78 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n111) );
  NAND2_X1 U79 ( .A1(n119), .A2(n118), .ZN(Z[26]) );
  AOI22_X1 U80 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n118) );
  AOI22_X1 U81 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n119) );
  NAND2_X1 U82 ( .A1(n129), .A2(n128), .ZN(Z[30]) );
  AOI22_X1 U83 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n128) );
  AOI22_X1 U84 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n129) );
  NAND2_X1 U85 ( .A1(n133), .A2(n132), .ZN(Z[3]) );
  AOI22_X1 U86 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n132) );
  AOI22_X1 U87 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n133) );
  NAND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(Z[7]) );
  AOI22_X1 U89 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n140) );
  AOI22_X1 U90 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n141) );
  NAND2_X1 U91 ( .A1(n87), .A2(n86), .ZN(Z[11]) );
  AOI22_X1 U92 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n86) );
  AOI22_X1 U93 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n87) );
  NAND2_X1 U94 ( .A1(n95), .A2(n94), .ZN(Z[15]) );
  AOI22_X1 U95 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n94) );
  AOI22_X1 U96 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n95) );
  NAND2_X1 U97 ( .A1(n103), .A2(n102), .ZN(Z[19]) );
  AOI22_X1 U98 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n102) );
  AOI22_X1 U99 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n103) );
  NAND2_X1 U100 ( .A1(n113), .A2(n112), .ZN(Z[23]) );
  AOI22_X1 U101 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n112) );
  AOI22_X1 U102 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n113) );
  NAND2_X1 U103 ( .A1(n121), .A2(n120), .ZN(Z[27]) );
  AOI22_X1 U104 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n120) );
  AOI22_X1 U105 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n121) );
  NAND2_X1 U106 ( .A1(n131), .A2(n130), .ZN(Z[31]) );
  AOI22_X1 U107 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n130) );
  AOI22_X1 U108 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n131) );
  NOR2_X1 U109 ( .A1(n81), .A2(S[1]), .ZN(n145) );
  NOR2_X1 U110 ( .A1(S[0]), .A2(S[1]), .ZN(n144) );
  AND2_X1 U111 ( .A1(S[1]), .A2(S[0]), .ZN(n147) );
  AND2_X1 U112 ( .A1(S[1]), .A2(n81), .ZN(n146) );
  INV_X1 U113 ( .A(S[0]), .ZN(n81) );
endmodule


module comparator_NBIT32_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202;

  INV_X1 U1 ( .A(n142), .ZN(n10) );
  INV_X1 U2 ( .A(n130), .ZN(n14) );
  INV_X1 U3 ( .A(n118), .ZN(n18) );
  INV_X1 U4 ( .A(n106), .ZN(n22) );
  INV_X1 U5 ( .A(n94), .ZN(n26) );
  INV_X1 U6 ( .A(n82), .ZN(n30) );
  INV_X1 U7 ( .A(GE), .ZN(LT) );
  INV_X1 U8 ( .A(NE), .ZN(EQ) );
  INV_X1 U9 ( .A(n139), .ZN(n12) );
  INV_X1 U10 ( .A(n127), .ZN(n16) );
  INV_X1 U11 ( .A(n115), .ZN(n20) );
  INV_X1 U12 ( .A(n103), .ZN(n24) );
  INV_X1 U13 ( .A(n91), .ZN(n28) );
  INV_X1 U14 ( .A(n79), .ZN(n32) );
  INV_X1 U15 ( .A(GT), .ZN(LE) );
  INV_X1 U16 ( .A(n144), .ZN(n9) );
  INV_X1 U17 ( .A(n132), .ZN(n13) );
  INV_X1 U18 ( .A(n120), .ZN(n17) );
  INV_X1 U19 ( .A(n108), .ZN(n21) );
  INV_X1 U20 ( .A(n96), .ZN(n25) );
  INV_X1 U21 ( .A(n84), .ZN(n29) );
  INV_X1 U22 ( .A(n154), .ZN(n7) );
  INV_X1 U23 ( .A(n141), .ZN(n11) );
  INV_X1 U24 ( .A(n129), .ZN(n15) );
  INV_X1 U25 ( .A(n117), .ZN(n19) );
  INV_X1 U26 ( .A(n105), .ZN(n23) );
  INV_X1 U27 ( .A(n93), .ZN(n27) );
  INV_X1 U28 ( .A(n81), .ZN(n31) );
  INV_X1 U29 ( .A(n68), .ZN(n3) );
  INV_X1 U30 ( .A(A[30]), .ZN(n65) );
  INV_X1 U31 ( .A(n72), .ZN(n33) );
  INV_X1 U32 ( .A(n151), .ZN(n8) );
  INV_X1 U33 ( .A(n202), .ZN(n5) );
  INV_X1 U34 ( .A(B[30]), .ZN(n34) );
  INV_X1 U35 ( .A(A[0]), .ZN(n36) );
  INV_X1 U36 ( .A(A[3]), .ZN(n38) );
  INV_X1 U37 ( .A(A[5]), .ZN(n40) );
  INV_X1 U38 ( .A(A[7]), .ZN(n42) );
  INV_X1 U39 ( .A(A[9]), .ZN(n44) );
  INV_X1 U40 ( .A(A[11]), .ZN(n46) );
  INV_X1 U41 ( .A(A[13]), .ZN(n48) );
  INV_X1 U42 ( .A(A[15]), .ZN(n50) );
  INV_X1 U43 ( .A(A[17]), .ZN(n52) );
  INV_X1 U44 ( .A(A[19]), .ZN(n54) );
  INV_X1 U45 ( .A(A[21]), .ZN(n56) );
  INV_X1 U46 ( .A(A[23]), .ZN(n58) );
  INV_X1 U47 ( .A(A[25]), .ZN(n60) );
  INV_X1 U48 ( .A(A[27]), .ZN(n62) );
  INV_X1 U49 ( .A(A[29]), .ZN(n64) );
  INV_X1 U50 ( .A(B[31]), .ZN(n35) );
  INV_X1 U51 ( .A(B[1]), .ZN(n6) );
  INV_X1 U52 ( .A(A[4]), .ZN(n39) );
  INV_X1 U53 ( .A(A[8]), .ZN(n43) );
  INV_X1 U54 ( .A(A[12]), .ZN(n47) );
  INV_X1 U55 ( .A(A[16]), .ZN(n51) );
  INV_X1 U56 ( .A(A[20]), .ZN(n55) );
  INV_X1 U57 ( .A(A[24]), .ZN(n59) );
  INV_X1 U58 ( .A(A[28]), .ZN(n63) );
  INV_X1 U59 ( .A(A[2]), .ZN(n37) );
  INV_X1 U60 ( .A(A[6]), .ZN(n41) );
  INV_X1 U61 ( .A(A[10]), .ZN(n45) );
  INV_X1 U62 ( .A(A[14]), .ZN(n49) );
  INV_X1 U63 ( .A(A[18]), .ZN(n53) );
  INV_X1 U64 ( .A(A[22]), .ZN(n57) );
  INV_X1 U65 ( .A(A[26]), .ZN(n61) );
  NAND2_X1 U66 ( .A1(LE), .A2(GE), .ZN(NE) );
  AOI21_X1 U67 ( .B1(n66), .B2(n3), .A(n67), .ZN(GE) );
  AOI22_X1 U68 ( .A1(B[30]), .A2(n65), .B1(n69), .B2(n70), .ZN(n68) );
  AOI21_X1 U69 ( .B1(n71), .B2(n72), .A(n73), .ZN(n69) );
  AOI21_X1 U70 ( .B1(n74), .B2(n75), .A(n76), .ZN(n71) );
  AOI21_X1 U71 ( .B1(n77), .B2(n78), .A(n79), .ZN(n74) );
  AOI21_X1 U72 ( .B1(n80), .B2(n30), .A(n31), .ZN(n77) );
  AOI21_X1 U73 ( .B1(n83), .B2(n84), .A(n85), .ZN(n80) );
  AOI21_X1 U74 ( .B1(n86), .B2(n87), .A(n88), .ZN(n83) );
  AOI21_X1 U75 ( .B1(n89), .B2(n90), .A(n91), .ZN(n86) );
  AOI21_X1 U76 ( .B1(n92), .B2(n26), .A(n27), .ZN(n89) );
  AOI21_X1 U77 ( .B1(n95), .B2(n96), .A(n97), .ZN(n92) );
  AOI21_X1 U78 ( .B1(n98), .B2(n99), .A(n100), .ZN(n95) );
  AOI21_X1 U79 ( .B1(n101), .B2(n102), .A(n103), .ZN(n98) );
  AOI21_X1 U80 ( .B1(n104), .B2(n22), .A(n23), .ZN(n101) );
  AOI21_X1 U81 ( .B1(n107), .B2(n108), .A(n109), .ZN(n104) );
  AOI21_X1 U82 ( .B1(n110), .B2(n111), .A(n112), .ZN(n107) );
  AOI21_X1 U83 ( .B1(n113), .B2(n114), .A(n115), .ZN(n110) );
  AOI21_X1 U84 ( .B1(n116), .B2(n18), .A(n19), .ZN(n113) );
  AOI21_X1 U85 ( .B1(n119), .B2(n120), .A(n121), .ZN(n116) );
  AOI21_X1 U86 ( .B1(n122), .B2(n123), .A(n124), .ZN(n119) );
  AOI21_X1 U87 ( .B1(n125), .B2(n126), .A(n127), .ZN(n122) );
  AOI21_X1 U88 ( .B1(n128), .B2(n14), .A(n15), .ZN(n125) );
  AOI21_X1 U89 ( .B1(n131), .B2(n132), .A(n133), .ZN(n128) );
  AOI21_X1 U90 ( .B1(n134), .B2(n135), .A(n136), .ZN(n131) );
  AOI21_X1 U91 ( .B1(n137), .B2(n138), .A(n139), .ZN(n134) );
  AOI21_X1 U92 ( .B1(n140), .B2(n10), .A(n11), .ZN(n137) );
  AOI21_X1 U93 ( .B1(n143), .B2(n144), .A(n145), .ZN(n140) );
  AOI21_X1 U94 ( .B1(n146), .B2(n147), .A(n148), .ZN(n143) );
  AOI21_X1 U95 ( .B1(n149), .B2(n150), .A(n151), .ZN(n146) );
  AOI21_X1 U96 ( .B1(n152), .B2(n153), .A(n7), .ZN(n149) );
  AOI22_X1 U97 ( .A1(n155), .A2(n6), .B1(A[1]), .B2(n156), .ZN(n152) );
  OR2_X1 U98 ( .A1(n156), .A2(A[1]), .ZN(n155) );
  NAND2_X1 U99 ( .A1(B[0]), .A2(n36), .ZN(n156) );
  OAI21_X1 U100 ( .B1(n67), .B2(n157), .A(n66), .ZN(GT) );
  NAND2_X1 U101 ( .A1(A[31]), .A2(n35), .ZN(n66) );
  AOI22_X1 U102 ( .A1(A[30]), .A2(n34), .B1(n158), .B2(n70), .ZN(n157) );
  XOR2_X1 U103 ( .A(A[30]), .B(n34), .Z(n70) );
  AOI21_X1 U104 ( .B1(n159), .B2(n160), .A(n33), .ZN(n158) );
  NAND2_X1 U105 ( .A1(B[29]), .A2(n64), .ZN(n72) );
  OAI211_X1 U106 ( .C1(n161), .C2(n162), .A(n78), .B(n75), .ZN(n160) );
  NOR2_X1 U107 ( .A1(n163), .A2(n76), .ZN(n75) );
  AND2_X1 U108 ( .A1(B[28]), .A2(n63), .ZN(n76) );
  NAND2_X1 U109 ( .A1(B[27]), .A2(n62), .ZN(n78) );
  NAND2_X1 U110 ( .A1(n32), .A2(n164), .ZN(n162) );
  NOR2_X1 U111 ( .A1(n62), .A2(B[27]), .ZN(n79) );
  AOI211_X1 U112 ( .C1(n165), .C2(n166), .A(n82), .B(n29), .ZN(n161) );
  NAND2_X1 U113 ( .A1(B[25]), .A2(n60), .ZN(n84) );
  NAND2_X1 U114 ( .A1(n164), .A2(n81), .ZN(n82) );
  NAND2_X1 U115 ( .A1(B[26]), .A2(n61), .ZN(n81) );
  OR2_X1 U116 ( .A1(n61), .A2(B[26]), .ZN(n164) );
  OAI211_X1 U117 ( .C1(n167), .C2(n168), .A(n90), .B(n87), .ZN(n166) );
  NOR2_X1 U118 ( .A1(n169), .A2(n88), .ZN(n87) );
  AND2_X1 U119 ( .A1(B[24]), .A2(n59), .ZN(n88) );
  NAND2_X1 U120 ( .A1(B[23]), .A2(n58), .ZN(n90) );
  NAND2_X1 U121 ( .A1(n28), .A2(n170), .ZN(n168) );
  NOR2_X1 U122 ( .A1(n58), .A2(B[23]), .ZN(n91) );
  AOI211_X1 U123 ( .C1(n171), .C2(n172), .A(n94), .B(n25), .ZN(n167) );
  NAND2_X1 U124 ( .A1(B[21]), .A2(n56), .ZN(n96) );
  NAND2_X1 U125 ( .A1(n170), .A2(n93), .ZN(n94) );
  NAND2_X1 U126 ( .A1(B[22]), .A2(n57), .ZN(n93) );
  OR2_X1 U127 ( .A1(n57), .A2(B[22]), .ZN(n170) );
  OAI211_X1 U128 ( .C1(n173), .C2(n174), .A(n102), .B(n99), .ZN(n172) );
  NOR2_X1 U129 ( .A1(n175), .A2(n100), .ZN(n99) );
  AND2_X1 U130 ( .A1(B[20]), .A2(n55), .ZN(n100) );
  NAND2_X1 U131 ( .A1(B[19]), .A2(n54), .ZN(n102) );
  NAND2_X1 U132 ( .A1(n24), .A2(n176), .ZN(n174) );
  NOR2_X1 U133 ( .A1(n54), .A2(B[19]), .ZN(n103) );
  AOI211_X1 U134 ( .C1(n177), .C2(n178), .A(n106), .B(n21), .ZN(n173) );
  NAND2_X1 U135 ( .A1(B[17]), .A2(n52), .ZN(n108) );
  NAND2_X1 U136 ( .A1(n176), .A2(n105), .ZN(n106) );
  NAND2_X1 U137 ( .A1(B[18]), .A2(n53), .ZN(n105) );
  OR2_X1 U138 ( .A1(n53), .A2(B[18]), .ZN(n176) );
  OAI211_X1 U139 ( .C1(n179), .C2(n180), .A(n114), .B(n111), .ZN(n178) );
  NOR2_X1 U140 ( .A1(n181), .A2(n112), .ZN(n111) );
  AND2_X1 U141 ( .A1(B[16]), .A2(n51), .ZN(n112) );
  NAND2_X1 U142 ( .A1(B[15]), .A2(n50), .ZN(n114) );
  NAND2_X1 U143 ( .A1(n20), .A2(n182), .ZN(n180) );
  NOR2_X1 U144 ( .A1(n50), .A2(B[15]), .ZN(n115) );
  AOI211_X1 U145 ( .C1(n183), .C2(n184), .A(n118), .B(n17), .ZN(n179) );
  NAND2_X1 U146 ( .A1(B[13]), .A2(n48), .ZN(n120) );
  NAND2_X1 U147 ( .A1(n182), .A2(n117), .ZN(n118) );
  NAND2_X1 U148 ( .A1(B[14]), .A2(n49), .ZN(n117) );
  OR2_X1 U149 ( .A1(n49), .A2(B[14]), .ZN(n182) );
  OAI211_X1 U150 ( .C1(n185), .C2(n186), .A(n126), .B(n123), .ZN(n184) );
  NOR2_X1 U151 ( .A1(n187), .A2(n124), .ZN(n123) );
  AND2_X1 U152 ( .A1(B[12]), .A2(n47), .ZN(n124) );
  NAND2_X1 U153 ( .A1(B[11]), .A2(n46), .ZN(n126) );
  NAND2_X1 U154 ( .A1(n16), .A2(n188), .ZN(n186) );
  NOR2_X1 U155 ( .A1(n46), .A2(B[11]), .ZN(n127) );
  AOI211_X1 U156 ( .C1(n189), .C2(n190), .A(n130), .B(n13), .ZN(n185) );
  NAND2_X1 U157 ( .A1(B[9]), .A2(n44), .ZN(n132) );
  NAND2_X1 U158 ( .A1(n188), .A2(n129), .ZN(n130) );
  NAND2_X1 U159 ( .A1(B[10]), .A2(n45), .ZN(n129) );
  OR2_X1 U160 ( .A1(n45), .A2(B[10]), .ZN(n188) );
  OAI211_X1 U161 ( .C1(n191), .C2(n192), .A(n138), .B(n135), .ZN(n190) );
  NOR2_X1 U162 ( .A1(n193), .A2(n136), .ZN(n135) );
  AND2_X1 U163 ( .A1(B[8]), .A2(n43), .ZN(n136) );
  NAND2_X1 U164 ( .A1(B[7]), .A2(n42), .ZN(n138) );
  NAND2_X1 U165 ( .A1(n12), .A2(n194), .ZN(n192) );
  NOR2_X1 U166 ( .A1(n42), .A2(B[7]), .ZN(n139) );
  AOI211_X1 U167 ( .C1(n195), .C2(n196), .A(n142), .B(n9), .ZN(n191) );
  NAND2_X1 U168 ( .A1(B[5]), .A2(n40), .ZN(n144) );
  NAND2_X1 U169 ( .A1(n194), .A2(n141), .ZN(n142) );
  NAND2_X1 U170 ( .A1(B[6]), .A2(n41), .ZN(n141) );
  OR2_X1 U171 ( .A1(n41), .A2(B[6]), .ZN(n194) );
  NAND3_X1 U172 ( .A1(n197), .A2(n150), .A3(n147), .ZN(n196) );
  NOR2_X1 U173 ( .A1(n198), .A2(n148), .ZN(n147) );
  AND2_X1 U174 ( .A1(B[4]), .A2(n39), .ZN(n148) );
  NAND2_X1 U175 ( .A1(B[3]), .A2(n38), .ZN(n150) );
  NAND3_X1 U176 ( .A1(n8), .A2(n199), .A3(n200), .ZN(n197) );
  OAI211_X1 U177 ( .C1(A[1]), .C2(n201), .A(n5), .B(n153), .ZN(n200) );
  AND2_X1 U178 ( .A1(n199), .A2(n154), .ZN(n153) );
  NAND2_X1 U179 ( .A1(B[2]), .A2(n37), .ZN(n154) );
  AOI21_X1 U180 ( .B1(A[1]), .B2(n201), .A(n6), .ZN(n202) );
  NOR2_X1 U181 ( .A1(n36), .A2(B[0]), .ZN(n201) );
  OR2_X1 U182 ( .A1(n37), .A2(B[2]), .ZN(n199) );
  NOR2_X1 U183 ( .A1(n38), .A2(B[3]), .ZN(n151) );
  NOR2_X1 U184 ( .A1(n198), .A2(n145), .ZN(n195) );
  NOR2_X1 U185 ( .A1(n40), .A2(B[5]), .ZN(n145) );
  NOR2_X1 U186 ( .A1(n39), .A2(B[4]), .ZN(n198) );
  NOR2_X1 U187 ( .A1(n193), .A2(n133), .ZN(n189) );
  NOR2_X1 U188 ( .A1(n44), .A2(B[9]), .ZN(n133) );
  NOR2_X1 U189 ( .A1(n43), .A2(B[8]), .ZN(n193) );
  NOR2_X1 U190 ( .A1(n187), .A2(n121), .ZN(n183) );
  NOR2_X1 U191 ( .A1(n48), .A2(B[13]), .ZN(n121) );
  NOR2_X1 U192 ( .A1(n47), .A2(B[12]), .ZN(n187) );
  NOR2_X1 U193 ( .A1(n181), .A2(n109), .ZN(n177) );
  NOR2_X1 U194 ( .A1(n52), .A2(B[17]), .ZN(n109) );
  NOR2_X1 U195 ( .A1(n51), .A2(B[16]), .ZN(n181) );
  NOR2_X1 U196 ( .A1(n175), .A2(n97), .ZN(n171) );
  NOR2_X1 U197 ( .A1(n56), .A2(B[21]), .ZN(n97) );
  NOR2_X1 U198 ( .A1(n55), .A2(B[20]), .ZN(n175) );
  NOR2_X1 U199 ( .A1(n169), .A2(n85), .ZN(n165) );
  NOR2_X1 U200 ( .A1(n60), .A2(B[25]), .ZN(n85) );
  NOR2_X1 U201 ( .A1(n59), .A2(B[24]), .ZN(n169) );
  NOR2_X1 U202 ( .A1(n163), .A2(n73), .ZN(n159) );
  NOR2_X1 U203 ( .A1(n64), .A2(B[29]), .ZN(n73) );
  NOR2_X1 U204 ( .A1(n63), .A2(B[28]), .ZN(n163) );
  NOR2_X1 U205 ( .A1(n35), .A2(A[31]), .ZN(n67) );
endmodule


module comparator_NBIT32 ( A, B, .OPSel({\OPSel[2] , \OPSel[1] , \OPSel[0] }), 
        RES );
  input [31:0] A;
  input [31:0] B;
  output [31:0] RES;
  input \OPSel[2] , \OPSel[1] , \OPSel[0] ;
  wire   N26, N27, N28, N29, N30, N31, n15, n16, n17, n18, n19, n20, n2, n3,
         n4;
  wire   [2:0] OPSel;
  assign RES[1] = 1'b0;
  assign RES[2] = 1'b0;
  assign RES[3] = 1'b0;
  assign RES[4] = 1'b0;
  assign RES[5] = 1'b0;
  assign RES[6] = 1'b0;
  assign RES[7] = 1'b0;
  assign RES[8] = 1'b0;
  assign RES[9] = 1'b0;
  assign RES[10] = 1'b0;
  assign RES[11] = 1'b0;
  assign RES[12] = 1'b0;
  assign RES[13] = 1'b0;
  assign RES[14] = 1'b0;
  assign RES[15] = 1'b0;
  assign RES[16] = 1'b0;
  assign RES[17] = 1'b0;
  assign RES[18] = 1'b0;
  assign RES[19] = 1'b0;
  assign RES[20] = 1'b0;
  assign RES[21] = 1'b0;
  assign RES[22] = 1'b0;
  assign RES[23] = 1'b0;
  assign RES[24] = 1'b0;
  assign RES[25] = 1'b0;
  assign RES[26] = 1'b0;
  assign RES[27] = 1'b0;
  assign RES[28] = 1'b0;
  assign RES[29] = 1'b0;
  assign RES[30] = 1'b0;
  assign RES[31] = 1'b0;

  comparator_NBIT32_DW01_cmp6_0 r57 ( .A(A), .B(B), .TC(1'b0), .LT(N30), .GT(
        N28), .EQ(N26), .LE(N31), .GE(N29), .NE(N27) );
  INV_X1 U3 ( .A(n15), .ZN(RES[0]) );
  AOI21_X1 U4 ( .B1(n16), .B2(n4), .A(n17), .ZN(n15) );
  NOR3_X1 U5 ( .A1(n4), .A2(OPSel[1]), .A3(n18), .ZN(n17) );
  OAI22_X1 U6 ( .A1(n19), .A2(n3), .B1(OPSel[1]), .B2(n20), .ZN(n16) );
  INV_X1 U7 ( .A(OPSel[1]), .ZN(n3) );
  AOI22_X1 U8 ( .A1(N28), .A2(n2), .B1(N29), .B2(OPSel[0]), .ZN(n19) );
  INV_X1 U9 ( .A(OPSel[0]), .ZN(n2) );
  AOI22_X1 U10 ( .A1(N30), .A2(n2), .B1(OPSel[0]), .B2(N31), .ZN(n18) );
  AOI22_X1 U11 ( .A1(N26), .A2(n2), .B1(N27), .B2(OPSel[0]), .ZN(n20) );
  INV_X1 U12 ( .A(OPSel[2]), .ZN(n4) );
endmodule


module PG_net_0 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_30 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_29 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_28 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_27 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_26 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_25 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_24 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_23 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_22 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_21 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_20 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_19 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_18 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_17 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_16 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_15 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_14 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_13 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_12 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_11 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_10 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_9 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_8 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_7 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_6 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_5 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_4 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_3 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_2 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_1 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module Gblock_0 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n2) );
endmodule


module Gblock_8 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_7 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_6 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_5 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_4 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_3 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_2 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_1 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module PGblock_0 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n2) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_26 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_25 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_24 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_23 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_22 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_21 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_20 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_19 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_18 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_17 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_16 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_15 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_14 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_13 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_12 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_11 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_10 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_9 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_8 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_7 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_6 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_5 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_4 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_3 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_2 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_1 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module carry_generator_NBIT32_NBIT_PER_BLOCK4 ( A, B, Cin, Co );
  input [32:1] A;
  input [32:1] B;
  output [7:0] Co;
  input Cin;
  wire   \G[16][16] , \G[16][15] , \G[16][13] , \G[16][9] , \G[15][15] ,
         \G[14][14] , \G[14][13] , \G[13][13] , \G[12][12] , \G[12][11] ,
         \G[12][9] , \G[11][11] , \G[10][10] , \G[10][9] , \G[9][9] ,
         \G[8][8] , \G[8][7] , \G[8][5] , \G[7][7] , \G[6][6] , \G[6][5] ,
         \G[5][5] , \G[4][4] , \G[4][3] , \G[3][3] , \G[2][2] , \G[2][1] ,
         \G[1][1] , \P[16][16] , \P[16][15] , \P[16][13] , \P[16][9] ,
         \P[15][15] , \P[14][14] , \P[14][13] , \P[13][13] , \P[12][12] ,
         \P[12][11] , \P[12][9] , \P[11][11] , \P[10][10] , \P[10][9] ,
         \P[9][9] , \P[8][8] , \P[8][7] , \P[8][5] , \P[7][7] , \P[6][6] ,
         \P[6][5] , \P[5][5] , \P[4][4] , \P[4][3] , \P[3][3] , \P[2][2] ,
         \G[32][32] , \G[32][31] , \G[32][29] , \G[32][25] , \G[32][17] ,
         \G[31][31] , \G[30][30] , \G[30][29] , \G[29][29] , \G[28][28] ,
         \G[28][27] , \G[28][25] , \G[28][17] , \G[27][27] , \G[26][26] ,
         \G[26][25] , \G[25][25] , \G[24][24] , \G[24][23] , \G[24][21] ,
         \G[24][17] , \G[23][23] , \G[22][22] , \G[22][21] , \G[21][21] ,
         \G[20][20] , \G[20][19] , \G[20][17] , \G[19][19] , \G[18][18] ,
         \G[18][17] , \G[17][17] , \P[32][32] , \P[32][31] , \P[32][29] ,
         \P[32][25] , \P[32][17] , \P[31][31] , \P[30][30] , \P[30][29] ,
         \P[29][29] , \P[28][28] , \P[28][27] , \P[28][25] , \P[28][17] ,
         \P[27][27] , \P[26][26] , \P[26][25] , \P[25][25] , \P[24][24] ,
         \P[24][23] , \P[24][21] , \P[24][17] , \P[23][23] , \P[22][22] ,
         \P[22][21] , \P[21][21] , \P[20][20] , \P[20][19] , \P[20][17] ,
         \P[19][19] , \P[18][18] , \P[18][17] , \P[17][17] , n3, n1, n2;

  PG_net_0 PGnetblock_2 ( .a(A[2]), .b(B[2]), .p(\P[2][2] ), .g(\G[2][2] ) );
  PG_net_30 PGnetblock_3 ( .a(A[3]), .b(B[3]), .p(\P[3][3] ), .g(\G[3][3] ) );
  PG_net_29 PGnetblock_4 ( .a(A[4]), .b(B[4]), .p(\P[4][4] ), .g(\G[4][4] ) );
  PG_net_28 PGnetblock_5 ( .a(A[5]), .b(B[5]), .p(\P[5][5] ), .g(\G[5][5] ) );
  PG_net_27 PGnetblock_6 ( .a(A[6]), .b(B[6]), .p(\P[6][6] ), .g(\G[6][6] ) );
  PG_net_26 PGnetblock_7 ( .a(A[7]), .b(B[7]), .p(\P[7][7] ), .g(\G[7][7] ) );
  PG_net_25 PGnetblock_8 ( .a(A[8]), .b(B[8]), .p(\P[8][8] ), .g(\G[8][8] ) );
  PG_net_24 PGnetblock_9 ( .a(A[9]), .b(B[9]), .p(\P[9][9] ), .g(\G[9][9] ) );
  PG_net_23 PGnetblock_10 ( .a(A[10]), .b(B[10]), .p(\P[10][10] ), .g(
        \G[10][10] ) );
  PG_net_22 PGnetblock_11 ( .a(A[11]), .b(B[11]), .p(\P[11][11] ), .g(
        \G[11][11] ) );
  PG_net_21 PGnetblock_12 ( .a(A[12]), .b(B[12]), .p(\P[12][12] ), .g(
        \G[12][12] ) );
  PG_net_20 PGnetblock_13 ( .a(A[13]), .b(B[13]), .p(\P[13][13] ), .g(
        \G[13][13] ) );
  PG_net_19 PGnetblock_14 ( .a(A[14]), .b(B[14]), .p(\P[14][14] ), .g(
        \G[14][14] ) );
  PG_net_18 PGnetblock_15 ( .a(A[15]), .b(B[15]), .p(\P[15][15] ), .g(
        \G[15][15] ) );
  PG_net_17 PGnetblock_16 ( .a(A[16]), .b(B[16]), .p(\P[16][16] ), .g(
        \G[16][16] ) );
  PG_net_16 PGnetblock_17 ( .a(A[17]), .b(B[17]), .p(\P[17][17] ), .g(
        \G[17][17] ) );
  PG_net_15 PGnetblock_18 ( .a(A[18]), .b(B[18]), .p(\P[18][18] ), .g(
        \G[18][18] ) );
  PG_net_14 PGnetblock_19 ( .a(A[19]), .b(B[19]), .p(\P[19][19] ), .g(
        \G[19][19] ) );
  PG_net_13 PGnetblock_20 ( .a(A[20]), .b(B[20]), .p(\P[20][20] ), .g(
        \G[20][20] ) );
  PG_net_12 PGnetblock_21 ( .a(A[21]), .b(B[21]), .p(\P[21][21] ), .g(
        \G[21][21] ) );
  PG_net_11 PGnetblock_22 ( .a(A[22]), .b(B[22]), .p(\P[22][22] ), .g(
        \G[22][22] ) );
  PG_net_10 PGnetblock_23 ( .a(A[23]), .b(B[23]), .p(\P[23][23] ), .g(
        \G[23][23] ) );
  PG_net_9 PGnetblock_24 ( .a(A[24]), .b(B[24]), .p(\P[24][24] ), .g(
        \G[24][24] ) );
  PG_net_8 PGnetblock_25 ( .a(A[25]), .b(B[25]), .p(\P[25][25] ), .g(
        \G[25][25] ) );
  PG_net_7 PGnetblock_26 ( .a(A[26]), .b(B[26]), .p(\P[26][26] ), .g(
        \G[26][26] ) );
  PG_net_6 PGnetblock_27 ( .a(A[27]), .b(B[27]), .p(\P[27][27] ), .g(
        \G[27][27] ) );
  PG_net_5 PGnetblock_28 ( .a(A[28]), .b(B[28]), .p(\P[28][28] ), .g(
        \G[28][28] ) );
  PG_net_4 PGnetblock_29 ( .a(A[29]), .b(B[29]), .p(\P[29][29] ), .g(
        \G[29][29] ) );
  PG_net_3 PGnetblock_30 ( .a(A[30]), .b(B[30]), .p(\P[30][30] ), .g(
        \G[30][30] ) );
  PG_net_2 PGnetblock_31 ( .a(A[31]), .b(B[31]), .p(\P[31][31] ), .g(
        \G[31][31] ) );
  PG_net_1 PGnetblock_32 ( .a(A[32]), .b(B[32]), .p(\P[32][32] ), .g(
        \G[32][32] ) );
  Gblock_0 GB_low_1_2 ( .Pik(\P[2][2] ), .Gik(\G[2][2] ), .Gk_1j(\G[1][1] ), 
        .Gij(\G[2][1] ) );
  Gblock_8 GB_low_2_4 ( .Pik(\P[4][3] ), .Gik(\G[4][3] ), .Gk_1j(\G[2][1] ), 
        .Gij(Co[0]) );
  Gblock_7 GB_low_3_8 ( .Pik(\P[8][5] ), .Gik(\G[8][5] ), .Gk_1j(Co[0]), .Gij(
        Co[1]) );
  Gblock_6 GB_high_4_16_0 ( .Pik(\P[16][9] ), .Gik(\G[16][9] ), .Gk_1j(Co[1]), 
        .Gij(Co[3]) );
  Gblock_5 GB_high_4_16_1 ( .Pik(\P[12][9] ), .Gik(\G[12][9] ), .Gk_1j(Co[1]), 
        .Gij(Co[2]) );
  Gblock_4 GB_high_5_32_0 ( .Pik(\P[32][17] ), .Gik(\G[32][17] ), .Gk_1j(Co[3]), .Gij(Co[7]) );
  Gblock_3 GB_high_5_32_1 ( .Pik(\P[28][17] ), .Gik(\G[28][17] ), .Gk_1j(Co[3]), .Gij(Co[6]) );
  Gblock_2 GB_high_5_32_2 ( .Pik(\P[24][17] ), .Gik(\G[24][17] ), .Gk_1j(Co[3]), .Gij(Co[5]) );
  Gblock_1 GB_high_5_32_3 ( .Pik(\P[20][17] ), .Gik(\G[20][17] ), .Gk_1j(Co[3]), .Gij(Co[4]) );
  PGblock_0 PGB_low_1_4 ( .Pik(\P[4][4] ), .Gik(\G[4][4] ), .Pk_1j(\P[3][3] ), 
        .Gk_1j(\G[3][3] ), .Pij(\P[4][3] ), .Gij(\G[4][3] ) );
  PGblock_26 PGB_low_1_6 ( .Pik(\P[6][6] ), .Gik(\G[6][6] ), .Pk_1j(\P[5][5] ), 
        .Gk_1j(\G[5][5] ), .Pij(\P[6][5] ), .Gij(\G[6][5] ) );
  PGblock_25 PGB_low_1_8 ( .Pik(\P[8][8] ), .Gik(\G[8][8] ), .Pk_1j(\P[7][7] ), 
        .Gk_1j(\G[7][7] ), .Pij(\P[8][7] ), .Gij(\G[8][7] ) );
  PGblock_24 PGB_low_1_10 ( .Pik(\P[10][10] ), .Gik(\G[10][10] ), .Pk_1j(
        \P[9][9] ), .Gk_1j(\G[9][9] ), .Pij(\P[10][9] ), .Gij(\G[10][9] ) );
  PGblock_23 PGB_low_1_12 ( .Pik(\P[12][12] ), .Gik(\G[12][12] ), .Pk_1j(
        \P[11][11] ), .Gk_1j(\G[11][11] ), .Pij(\P[12][11] ), .Gij(\G[12][11] ) );
  PGblock_22 PGB_low_1_14 ( .Pik(\P[14][14] ), .Gik(\G[14][14] ), .Pk_1j(
        \P[13][13] ), .Gk_1j(\G[13][13] ), .Pij(\P[14][13] ), .Gij(\G[14][13] ) );
  PGblock_21 PGB_low_1_16 ( .Pik(\P[16][16] ), .Gik(\G[16][16] ), .Pk_1j(
        \P[15][15] ), .Gk_1j(\G[15][15] ), .Pij(\P[16][15] ), .Gij(\G[16][15] ) );
  PGblock_20 PGB_low_1_18 ( .Pik(\P[18][18] ), .Gik(\G[18][18] ), .Pk_1j(
        \P[17][17] ), .Gk_1j(\G[17][17] ), .Pij(\P[18][17] ), .Gij(\G[18][17] ) );
  PGblock_19 PGB_low_1_20 ( .Pik(\P[20][20] ), .Gik(\G[20][20] ), .Pk_1j(
        \P[19][19] ), .Gk_1j(\G[19][19] ), .Pij(\P[20][19] ), .Gij(\G[20][19] ) );
  PGblock_18 PGB_low_1_22 ( .Pik(\P[22][22] ), .Gik(\G[22][22] ), .Pk_1j(
        \P[21][21] ), .Gk_1j(\G[21][21] ), .Pij(\P[22][21] ), .Gij(\G[22][21] ) );
  PGblock_17 PGB_low_1_24 ( .Pik(\P[24][24] ), .Gik(\G[24][24] ), .Pk_1j(
        \P[23][23] ), .Gk_1j(\G[23][23] ), .Pij(\P[24][23] ), .Gij(\G[24][23] ) );
  PGblock_16 PGB_low_1_26 ( .Pik(\P[26][26] ), .Gik(\G[26][26] ), .Pk_1j(
        \P[25][25] ), .Gk_1j(\G[25][25] ), .Pij(\P[26][25] ), .Gij(\G[26][25] ) );
  PGblock_15 PGB_low_1_28 ( .Pik(\P[28][28] ), .Gik(\G[28][28] ), .Pk_1j(
        \P[27][27] ), .Gk_1j(\G[27][27] ), .Pij(\P[28][27] ), .Gij(\G[28][27] ) );
  PGblock_14 PGB_low_1_30 ( .Pik(\P[30][30] ), .Gik(\G[30][30] ), .Pk_1j(
        \P[29][29] ), .Gk_1j(\G[29][29] ), .Pij(\P[30][29] ), .Gij(\G[30][29] ) );
  PGblock_13 PGB_low_1_32 ( .Pik(\P[32][32] ), .Gik(\G[32][32] ), .Pk_1j(
        \P[31][31] ), .Gk_1j(\G[31][31] ), .Pij(\P[32][31] ), .Gij(\G[32][31] ) );
  PGblock_12 PGB_low_2_8 ( .Pik(\P[8][7] ), .Gik(\G[8][7] ), .Pk_1j(\P[6][5] ), 
        .Gk_1j(\G[6][5] ), .Pij(\P[8][5] ), .Gij(\G[8][5] ) );
  PGblock_11 PGB_low_2_12 ( .Pik(\P[12][11] ), .Gik(\G[12][11] ), .Pk_1j(
        \P[10][9] ), .Gk_1j(\G[10][9] ), .Pij(\P[12][9] ), .Gij(\G[12][9] ) );
  PGblock_10 PGB_low_2_16 ( .Pik(\P[16][15] ), .Gik(\G[16][15] ), .Pk_1j(
        \P[14][13] ), .Gk_1j(\G[14][13] ), .Pij(\P[16][13] ), .Gij(\G[16][13] ) );
  PGblock_9 PGB_low_2_20 ( .Pik(\P[20][19] ), .Gik(\G[20][19] ), .Pk_1j(
        \P[18][17] ), .Gk_1j(\G[18][17] ), .Pij(\P[20][17] ), .Gij(\G[20][17] ) );
  PGblock_8 PGB_low_2_24 ( .Pik(\P[24][23] ), .Gik(\G[24][23] ), .Pk_1j(
        \P[22][21] ), .Gk_1j(\G[22][21] ), .Pij(\P[24][21] ), .Gij(\G[24][21] ) );
  PGblock_7 PGB_low_2_28 ( .Pik(\P[28][27] ), .Gik(\G[28][27] ), .Pk_1j(
        \P[26][25] ), .Gk_1j(\G[26][25] ), .Pij(\P[28][25] ), .Gij(\G[28][25] ) );
  PGblock_6 PGB_low_2_32 ( .Pik(\P[32][31] ), .Gik(\G[32][31] ), .Pk_1j(
        \P[30][29] ), .Gk_1j(\G[30][29] ), .Pij(\P[32][29] ), .Gij(\G[32][29] ) );
  PGblock_5 PGB_low_3_16 ( .Pik(\P[16][13] ), .Gik(\G[16][13] ), .Pk_1j(
        \P[12][9] ), .Gk_1j(\G[12][9] ), .Pij(\P[16][9] ), .Gij(\G[16][9] ) );
  PGblock_4 PGB_low_3_24 ( .Pik(\P[24][21] ), .Gik(\G[24][21] ), .Pk_1j(
        \P[20][17] ), .Gk_1j(\G[20][17] ), .Pij(\P[24][17] ), .Gij(\G[24][17] ) );
  PGblock_3 PGB_low_3_32 ( .Pik(\P[32][29] ), .Gik(\G[32][29] ), .Pk_1j(
        \P[28][25] ), .Gk_1j(\G[28][25] ), .Pij(\P[32][25] ), .Gij(\G[32][25] ) );
  PGblock_2 PGB_high_4_32_0 ( .Pik(\P[32][25] ), .Gik(\G[32][25] ), .Pk_1j(
        \P[24][17] ), .Gk_1j(\G[24][17] ), .Pij(\P[32][17] ), .Gij(\G[32][17] ) );
  PGblock_1 PGB_high_4_32_1 ( .Pik(\P[28][25] ), .Gik(\G[28][25] ), .Pk_1j(
        \P[24][17] ), .Gk_1j(\G[24][17] ), .Pij(\P[28][17] ), .Gij(\G[28][17] ) );
  INV_X1 U1 ( .A(A[1]), .ZN(n1) );
  OAI21_X1 U2 ( .B1(n1), .B2(n2), .A(n3), .ZN(\G[1][1] ) );
  OAI21_X1 U3 ( .B1(A[1]), .B2(B[1]), .A(Cin), .ZN(n3) );
  INV_X1 U4 ( .A(B[1]), .ZN(n2) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_0 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n6, n7, n8, n9, n1;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_0 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_15 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  AOI22_X1 U3 ( .A1(Y1[2]), .A2(n1), .B1(Y2[2]), .B2(C_i), .ZN(n7) );
  AOI22_X1 U4 ( .A1(Y1[3]), .A2(n1), .B1(Y2[3]), .B2(C_i), .ZN(n6) );
  AOI22_X1 U5 ( .A1(Y1[1]), .A2(n1), .B1(Y2[1]), .B2(C_i), .ZN(n8) );
  AOI22_X1 U6 ( .A1(Y1[0]), .A2(n1), .B1(Y2[0]), .B2(C_i), .ZN(n9) );
  INV_X1 U7 ( .A(n6), .ZN(S[3]) );
  INV_X1 U8 ( .A(n9), .ZN(S[0]) );
  INV_X1 U9 ( .A(n8), .ZN(S[1]) );
  INV_X1 U10 ( .A(n7), .ZN(S[2]) );
  INV_X1 U11 ( .A(C_i), .ZN(n1) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_7 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_14 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_13 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  AOI22_X1 U4 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  AOI22_X1 U5 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  AOI22_X1 U6 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  AOI22_X1 U7 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
  INV_X1 U8 ( .A(n10), .ZN(S[0]) );
  INV_X1 U9 ( .A(n11), .ZN(S[1]) );
  INV_X1 U10 ( .A(n12), .ZN(S[2]) );
  INV_X1 U11 ( .A(n13), .ZN(S[3]) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_6 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_12 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_11 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  AOI22_X1 U4 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  AOI22_X1 U5 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  AOI22_X1 U6 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  AOI22_X1 U7 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
  INV_X1 U8 ( .A(n10), .ZN(S[0]) );
  INV_X1 U9 ( .A(n11), .ZN(S[1]) );
  INV_X1 U10 ( .A(n12), .ZN(S[2]) );
  INV_X1 U11 ( .A(n13), .ZN(S[3]) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_5 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_10 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_9 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  AOI22_X1 U4 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  AOI22_X1 U5 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  AOI22_X1 U6 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  AOI22_X1 U7 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
  INV_X1 U8 ( .A(n10), .ZN(S[0]) );
  INV_X1 U9 ( .A(n11), .ZN(S[1]) );
  INV_X1 U10 ( .A(n12), .ZN(S[2]) );
  INV_X1 U11 ( .A(n13), .ZN(S[3]) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_4 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_8 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_7 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  AOI22_X1 U4 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  AOI22_X1 U5 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  AOI22_X1 U6 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  AOI22_X1 U7 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
  INV_X1 U8 ( .A(n10), .ZN(S[0]) );
  INV_X1 U9 ( .A(n11), .ZN(S[1]) );
  INV_X1 U10 ( .A(n12), .ZN(S[2]) );
  INV_X1 U11 ( .A(n13), .ZN(S[3]) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_3 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_6 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_5 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  AOI22_X1 U4 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  AOI22_X1 U5 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  AOI22_X1 U6 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  AOI22_X1 U7 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
  INV_X1 U8 ( .A(n10), .ZN(S[0]) );
  INV_X1 U9 ( .A(n11), .ZN(S[1]) );
  INV_X1 U10 ( .A(n12), .ZN(S[2]) );
  INV_X1 U11 ( .A(n13), .ZN(S[3]) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_2 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_4 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_3 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  AOI22_X1 U4 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  AOI22_X1 U5 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  AOI22_X1 U6 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  AOI22_X1 U7 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
  INV_X1 U8 ( .A(n10), .ZN(S[0]) );
  INV_X1 U9 ( .A(n11), .ZN(S[1]) );
  INV_X1 U10 ( .A(n12), .ZN(S[2]) );
  INV_X1 U11 ( .A(n13), .ZN(S[3]) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_1 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_2 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_1 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  AOI22_X1 U4 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  AOI22_X1 U5 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  AOI22_X1 U6 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  AOI22_X1 U7 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
  INV_X1 U8 ( .A(n13), .ZN(S[3]) );
  INV_X1 U9 ( .A(n10), .ZN(S[0]) );
  INV_X1 U10 ( .A(n11), .ZN(S[1]) );
  INV_X1 U11 ( .A(n12), .ZN(S[2]) );
endmodule


module SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_select_basic_N4_0 CSBI_1 ( .A(A[3:0]), .B(B[3:0]), .C_i(Ci[0]), .S(
        S[3:0]) );
  carry_select_basic_N4_7 CSBI_2 ( .A(A[7:4]), .B(B[7:4]), .C_i(Ci[1]), .S(
        S[7:4]) );
  carry_select_basic_N4_6 CSBI_3 ( .A(A[11:8]), .B(B[11:8]), .C_i(Ci[2]), .S(
        S[11:8]) );
  carry_select_basic_N4_5 CSBI_4 ( .A(A[15:12]), .B(B[15:12]), .C_i(Ci[3]), 
        .S(S[15:12]) );
  carry_select_basic_N4_4 CSBI_5 ( .A(A[19:16]), .B(B[19:16]), .C_i(Ci[4]), 
        .S(S[19:16]) );
  carry_select_basic_N4_3 CSBI_6 ( .A(A[23:20]), .B(B[23:20]), .C_i(Ci[5]), 
        .S(S[23:20]) );
  carry_select_basic_N4_2 CSBI_7 ( .A(A[27:24]), .B(B[27:24]), .C_i(Ci[6]), 
        .S(S[27:24]) );
  carry_select_basic_N4_1 CSBI_8 ( .A(A[31:28]), .B(B[31:28]), .C_i(Ci[7]), 
        .S(S[31:28]) );
endmodule


module P4Adder_NBIT32 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;

  wire   [7:1] Csum;

  carry_generator_NBIT32_NBIT_PER_BLOCK4 Carrygen0 ( .A(A), .B(B), .Cin(Cin), 
        .Co({Cout, Csum}) );
  SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 Sumgen0 ( .A(A), .B(B), .Ci({Csum, 
        Cin}), .S(S) );
endmodule


module mux41_NBIT32_1 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149;

  BUF_X1 U1 ( .A(n145), .Z(n72) );
  BUF_X1 U2 ( .A(n145), .Z(n73) );
  BUF_X1 U3 ( .A(n147), .Z(n78) );
  BUF_X1 U4 ( .A(n147), .Z(n79) );
  BUF_X1 U5 ( .A(n144), .Z(n1) );
  BUF_X1 U6 ( .A(n144), .Z(n70) );
  BUF_X1 U7 ( .A(n146), .Z(n75) );
  BUF_X1 U8 ( .A(n146), .Z(n76) );
  BUF_X1 U9 ( .A(n145), .Z(n74) );
  BUF_X1 U10 ( .A(n147), .Z(n80) );
  BUF_X1 U11 ( .A(n144), .Z(n71) );
  BUF_X1 U12 ( .A(n146), .Z(n77) );
  NOR2_X1 U13 ( .A1(S[0]), .A2(S[1]), .ZN(n144) );
  NOR2_X1 U14 ( .A1(n81), .A2(S[1]), .ZN(n145) );
  AND2_X1 U15 ( .A1(S[1]), .A2(S[0]), .ZN(n147) );
  AND2_X1 U16 ( .A1(S[1]), .A2(n81), .ZN(n146) );
  INV_X1 U17 ( .A(S[0]), .ZN(n81) );
  NAND2_X1 U18 ( .A1(n133), .A2(n132), .ZN(Z[3]) );
  AOI22_X1 U19 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n132) );
  AOI22_X1 U20 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n133) );
  NAND2_X1 U21 ( .A1(n135), .A2(n134), .ZN(Z[4]) );
  AOI22_X1 U22 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n134) );
  AOI22_X1 U23 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n135) );
  NAND2_X1 U24 ( .A1(n137), .A2(n136), .ZN(Z[5]) );
  AOI22_X1 U25 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n136) );
  AOI22_X1 U26 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n137) );
  NAND2_X1 U27 ( .A1(n139), .A2(n138), .ZN(Z[6]) );
  AOI22_X1 U28 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n138) );
  AOI22_X1 U29 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n139) );
  NAND2_X1 U30 ( .A1(n141), .A2(n140), .ZN(Z[7]) );
  AOI22_X1 U31 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n140) );
  AOI22_X1 U32 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n141) );
  NAND2_X1 U33 ( .A1(n143), .A2(n142), .ZN(Z[8]) );
  AOI22_X1 U34 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n142) );
  AOI22_X1 U35 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n143) );
  NAND2_X1 U36 ( .A1(n149), .A2(n148), .ZN(Z[9]) );
  AOI22_X1 U37 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n148) );
  AOI22_X1 U38 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n149) );
  NAND2_X1 U39 ( .A1(n131), .A2(n130), .ZN(Z[31]) );
  AOI22_X1 U40 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n130) );
  AOI22_X1 U41 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n131) );
  NAND2_X1 U42 ( .A1(n83), .A2(n82), .ZN(Z[0]) );
  AOI22_X1 U43 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n83) );
  AOI22_X1 U44 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n82) );
  NAND2_X1 U45 ( .A1(n105), .A2(n104), .ZN(Z[1]) );
  AOI22_X1 U46 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n104) );
  AOI22_X1 U47 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n105) );
  NAND2_X1 U48 ( .A1(n127), .A2(n126), .ZN(Z[2]) );
  AOI22_X1 U49 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n126) );
  AOI22_X1 U50 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n127) );
  NAND2_X1 U51 ( .A1(n85), .A2(n84), .ZN(Z[10]) );
  AOI22_X1 U52 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n84) );
  AOI22_X1 U53 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n85) );
  NAND2_X1 U54 ( .A1(n87), .A2(n86), .ZN(Z[11]) );
  AOI22_X1 U55 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n86) );
  AOI22_X1 U56 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n87) );
  NAND2_X1 U57 ( .A1(n89), .A2(n88), .ZN(Z[12]) );
  AOI22_X1 U58 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n88) );
  AOI22_X1 U59 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n89) );
  NAND2_X1 U60 ( .A1(n91), .A2(n90), .ZN(Z[13]) );
  AOI22_X1 U61 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n90) );
  AOI22_X1 U62 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n91) );
  NAND2_X1 U63 ( .A1(n93), .A2(n92), .ZN(Z[14]) );
  AOI22_X1 U64 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n92) );
  AOI22_X1 U65 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n93) );
  NAND2_X1 U66 ( .A1(n95), .A2(n94), .ZN(Z[15]) );
  AOI22_X1 U67 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n94) );
  AOI22_X1 U68 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n95) );
  NAND2_X1 U69 ( .A1(n97), .A2(n96), .ZN(Z[16]) );
  AOI22_X1 U70 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n96) );
  AOI22_X1 U71 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n97) );
  NAND2_X1 U72 ( .A1(n99), .A2(n98), .ZN(Z[17]) );
  AOI22_X1 U73 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n98) );
  AOI22_X1 U74 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n99) );
  NAND2_X1 U75 ( .A1(n101), .A2(n100), .ZN(Z[18]) );
  AOI22_X1 U76 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n100) );
  AOI22_X1 U77 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n101) );
  NAND2_X1 U78 ( .A1(n103), .A2(n102), .ZN(Z[19]) );
  AOI22_X1 U79 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n102) );
  AOI22_X1 U80 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n103) );
  NAND2_X1 U81 ( .A1(n107), .A2(n106), .ZN(Z[20]) );
  AOI22_X1 U82 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n106) );
  AOI22_X1 U83 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n107) );
  NAND2_X1 U84 ( .A1(n109), .A2(n108), .ZN(Z[21]) );
  AOI22_X1 U85 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n108) );
  AOI22_X1 U86 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n109) );
  NAND2_X1 U87 ( .A1(n111), .A2(n110), .ZN(Z[22]) );
  AOI22_X1 U88 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n110) );
  AOI22_X1 U89 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n111) );
  NAND2_X1 U90 ( .A1(n113), .A2(n112), .ZN(Z[23]) );
  AOI22_X1 U91 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n112) );
  AOI22_X1 U92 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n113) );
  NAND2_X1 U93 ( .A1(n115), .A2(n114), .ZN(Z[24]) );
  AOI22_X1 U94 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n114) );
  AOI22_X1 U95 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n115) );
  NAND2_X1 U96 ( .A1(n117), .A2(n116), .ZN(Z[25]) );
  AOI22_X1 U97 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n116) );
  AOI22_X1 U98 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n117) );
  NAND2_X1 U99 ( .A1(n119), .A2(n118), .ZN(Z[26]) );
  AOI22_X1 U100 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n118) );
  AOI22_X1 U101 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n119) );
  NAND2_X1 U102 ( .A1(n121), .A2(n120), .ZN(Z[27]) );
  AOI22_X1 U103 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n120) );
  AOI22_X1 U104 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n121) );
  NAND2_X1 U105 ( .A1(n123), .A2(n122), .ZN(Z[28]) );
  AOI22_X1 U106 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n122) );
  AOI22_X1 U107 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n123) );
  NAND2_X1 U108 ( .A1(n125), .A2(n124), .ZN(Z[29]) );
  AOI22_X1 U109 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n124) );
  AOI22_X1 U110 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n125) );
  NAND2_X1 U111 ( .A1(n129), .A2(n128), .ZN(Z[30]) );
  AOI22_X1 U112 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n128) );
  AOI22_X1 U113 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n129) );
endmodule


module mux21_NBIT32_1 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n11) );
  BUF_X1 U6 ( .A(n2), .Z(n9) );
  BUF_X1 U7 ( .A(n1), .Z(n8) );
  BUF_X1 U8 ( .A(n2), .Z(n10) );
  BUF_X1 U9 ( .A(n1), .Z(n7) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(S), .Z(n3) );
  BUF_X1 U13 ( .A(S), .Z(n2) );
  BUF_X1 U14 ( .A(S), .Z(n1) );
  INV_X1 U15 ( .A(n79), .ZN(Z[0]) );
  AOI22_X1 U16 ( .A1(A[0]), .A2(n4), .B1(B[0]), .B2(n13), .ZN(n79) );
  INV_X1 U17 ( .A(n90), .ZN(Z[1]) );
  AOI22_X1 U18 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(n10), .ZN(n90) );
  INV_X1 U19 ( .A(n101), .ZN(Z[2]) );
  AOI22_X1 U20 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n7), .ZN(n101) );
  INV_X1 U21 ( .A(n104), .ZN(Z[3]) );
  AOI22_X1 U22 ( .A1(A[3]), .A2(n4), .B1(B[3]), .B2(n7), .ZN(n104) );
  INV_X1 U23 ( .A(n105), .ZN(Z[4]) );
  AOI22_X1 U24 ( .A1(A[4]), .A2(n5), .B1(B[4]), .B2(n7), .ZN(n105) );
  INV_X1 U25 ( .A(n106), .ZN(Z[5]) );
  AOI22_X1 U26 ( .A1(A[5]), .A2(n4), .B1(B[5]), .B2(n6), .ZN(n106) );
  INV_X1 U27 ( .A(n107), .ZN(Z[6]) );
  AOI22_X1 U28 ( .A1(A[6]), .A2(n5), .B1(B[6]), .B2(n6), .ZN(n107) );
  INV_X1 U29 ( .A(n108), .ZN(Z[7]) );
  AOI22_X1 U30 ( .A1(A[7]), .A2(n4), .B1(B[7]), .B2(n6), .ZN(n108) );
  INV_X1 U31 ( .A(n109), .ZN(Z[8]) );
  AOI22_X1 U32 ( .A1(A[8]), .A2(n5), .B1(B[8]), .B2(n6), .ZN(n109) );
  INV_X1 U33 ( .A(n110), .ZN(Z[9]) );
  AOI22_X1 U34 ( .A1(A[9]), .A2(n4), .B1(n13), .B2(B[9]), .ZN(n110) );
  INV_X1 U35 ( .A(n80), .ZN(Z[10]) );
  AOI22_X1 U36 ( .A1(A[10]), .A2(n4), .B1(B[10]), .B2(n13), .ZN(n80) );
  INV_X1 U37 ( .A(n81), .ZN(Z[11]) );
  AOI22_X1 U38 ( .A1(A[11]), .A2(n4), .B1(B[11]), .B2(n13), .ZN(n81) );
  INV_X1 U39 ( .A(n82), .ZN(Z[12]) );
  AOI22_X1 U40 ( .A1(A[12]), .A2(n4), .B1(B[12]), .B2(n12), .ZN(n82) );
  INV_X1 U41 ( .A(n83), .ZN(Z[13]) );
  AOI22_X1 U42 ( .A1(A[13]), .A2(n4), .B1(B[13]), .B2(n12), .ZN(n83) );
  INV_X1 U43 ( .A(n84), .ZN(Z[14]) );
  AOI22_X1 U44 ( .A1(A[14]), .A2(n4), .B1(B[14]), .B2(n12), .ZN(n84) );
  INV_X1 U45 ( .A(n85), .ZN(Z[15]) );
  AOI22_X1 U46 ( .A1(A[15]), .A2(n4), .B1(B[15]), .B2(n12), .ZN(n85) );
  INV_X1 U47 ( .A(n86), .ZN(Z[16]) );
  AOI22_X1 U48 ( .A1(A[16]), .A2(n4), .B1(B[16]), .B2(n11), .ZN(n86) );
  INV_X1 U49 ( .A(n87), .ZN(Z[17]) );
  AOI22_X1 U50 ( .A1(A[17]), .A2(n4), .B1(B[17]), .B2(n11), .ZN(n87) );
  INV_X1 U51 ( .A(n88), .ZN(Z[18]) );
  AOI22_X1 U52 ( .A1(A[18]), .A2(n4), .B1(B[18]), .B2(n11), .ZN(n88) );
  INV_X1 U53 ( .A(n89), .ZN(Z[19]) );
  AOI22_X1 U54 ( .A1(A[19]), .A2(n4), .B1(B[19]), .B2(n11), .ZN(n89) );
  INV_X1 U55 ( .A(n91), .ZN(Z[20]) );
  AOI22_X1 U56 ( .A1(A[20]), .A2(n5), .B1(B[20]), .B2(n10), .ZN(n91) );
  INV_X1 U57 ( .A(n92), .ZN(Z[21]) );
  AOI22_X1 U58 ( .A1(A[21]), .A2(n5), .B1(B[21]), .B2(n10), .ZN(n92) );
  INV_X1 U59 ( .A(n93), .ZN(Z[22]) );
  AOI22_X1 U60 ( .A1(A[22]), .A2(n5), .B1(B[22]), .B2(n9), .ZN(n93) );
  INV_X1 U61 ( .A(n94), .ZN(Z[23]) );
  AOI22_X1 U62 ( .A1(A[23]), .A2(n5), .B1(B[23]), .B2(n9), .ZN(n94) );
  INV_X1 U63 ( .A(n95), .ZN(Z[24]) );
  AOI22_X1 U64 ( .A1(A[24]), .A2(n5), .B1(B[24]), .B2(n9), .ZN(n95) );
  INV_X1 U65 ( .A(n96), .ZN(Z[25]) );
  AOI22_X1 U66 ( .A1(A[25]), .A2(n5), .B1(B[25]), .B2(n9), .ZN(n96) );
  INV_X1 U67 ( .A(n97), .ZN(Z[26]) );
  AOI22_X1 U68 ( .A1(A[26]), .A2(n5), .B1(B[26]), .B2(n8), .ZN(n97) );
  INV_X1 U69 ( .A(n98), .ZN(Z[27]) );
  AOI22_X1 U70 ( .A1(A[27]), .A2(n5), .B1(B[27]), .B2(n8), .ZN(n98) );
  INV_X1 U71 ( .A(n99), .ZN(Z[28]) );
  AOI22_X1 U72 ( .A1(A[28]), .A2(n5), .B1(B[28]), .B2(n8), .ZN(n99) );
  INV_X1 U73 ( .A(n100), .ZN(Z[29]) );
  AOI22_X1 U74 ( .A1(A[29]), .A2(n5), .B1(B[29]), .B2(n8), .ZN(n100) );
  INV_X1 U75 ( .A(n102), .ZN(Z[30]) );
  AOI22_X1 U76 ( .A1(A[30]), .A2(n5), .B1(B[30]), .B2(n10), .ZN(n102) );
  INV_X1 U77 ( .A(n103), .ZN(Z[31]) );
  AOI22_X1 U78 ( .A1(A[31]), .A2(n5), .B1(B[31]), .B2(n7), .ZN(n103) );
endmodule


module ALU_NBIT32 ( OP1, OP2, .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , 
        \ALU_OPC[1] , \ALU_OPC[0] }), ALU_RES );
  input [31:0] OP1;
  input [31:0] OP2;
  output [31:0] ALU_RES;
  input \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] ;
  wire   select_zero_sig, LOGIC_ARITH, \OPSel[0] , n78, n79, n80, n81, n82,
         n83, n84, n85, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n86, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186;
  wire   [3:0] ALU_OPC;
  wire   [1:0] select_type_sig;
  wire   [31:0] A_SHF;
  wire   [31:0] B_SHF;
  wire   [31:0] A_ADD;
  wire   [31:0] B_ADD;
  wire   [31:0] LOGIC_RES;
  wire   [31:0] COMP_RES;
  wire   [31:0] SHIFT_RES;
  wire   [31:0] ADD_SUB_RES;
  wire   [31:0] sig_intraMux;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  NAND3_X1 U317 ( .A1(n185), .A2(n184), .A3(n186), .ZN(n79) );
  NAND3_X1 U318 ( .A1(n84), .A2(n83), .A3(n87), .ZN(\OPSel[0] ) );
  NAND3_X1 U319 ( .A1(ALU_OPC[3]), .A2(n186), .A3(n88), .ZN(n87) );
  NAND3_X1 U320 ( .A1(ALU_OPC[3]), .A2(n186), .A3(n89), .ZN(n83) );
  NAND3_X1 U321 ( .A1(ALU_OPC[3]), .A2(ALU_OPC[0]), .A3(n89), .ZN(n84) );
  NAND3_X1 U322 ( .A1(ALU_OPC[2]), .A2(ALU_OPC[1]), .A3(n155), .ZN(n157) );
  NAND3_X1 U323 ( .A1(ALU_OPC[2]), .A2(ALU_OPC[1]), .A3(n154), .ZN(n85) );
  NAND3_X1 U324 ( .A1(n185), .A2(n184), .A3(n155), .ZN(n156) );
  comparator_NBIT32 Comp ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .OPSel({n183, n182, 
        \OPSel[0] }), .RES({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, COMP_RES[0]}) );
  shifter Shift ( .A(A_SHF), .B(B_SHF), .LOGIC_ARITH(LOGIC_ARITH), 
        .LEFT_RIGHT(n180), .RES(SHIFT_RES) );
  P4Adder_NBIT32 Add_Sub_unit ( .A(A_ADD), .B(B_ADD), .Cin(n1), .S(ADD_SUB_RES) );
  mux41_NBIT32_1 Res_mux ( .A(ADD_SUB_RES), .B(LOGIC_RES), .C(SHIFT_RES), .D({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, COMP_RES[0]}), .S(
        select_type_sig), .Z(sig_intraMux) );
  mux21_NBIT32_1 Zeros_mux ( .A(sig_intraMux), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .S(select_zero_sig), .Z(ALU_RES) );
  BUF_X1 U2 ( .A(n158), .Z(n23) );
  BUF_X1 U3 ( .A(n158), .Z(n24) );
  BUF_X1 U4 ( .A(n158), .Z(n25) );
  BUF_X1 U5 ( .A(n177), .Z(n5) );
  BUF_X1 U6 ( .A(n177), .Z(n6) );
  BUF_X1 U7 ( .A(n177), .Z(n7) );
  BUF_X1 U8 ( .A(n177), .Z(n9) );
  BUF_X1 U9 ( .A(n177), .Z(n8) );
  BUF_X1 U10 ( .A(n179), .Z(n17) );
  BUF_X1 U11 ( .A(n179), .Z(n18) );
  BUF_X1 U12 ( .A(n179), .Z(n21) );
  BUF_X1 U13 ( .A(n179), .Z(n20) );
  BUF_X1 U14 ( .A(n179), .Z(n19) );
  BUF_X1 U15 ( .A(n176), .Z(n2) );
  BUF_X1 U16 ( .A(n176), .Z(n3) );
  BUF_X1 U17 ( .A(n176), .Z(n4) );
  AND2_X1 U18 ( .A1(n28), .A2(n29), .ZN(n158) );
  NOR2_X1 U19 ( .A1(n23), .A2(n31), .ZN(A_ADD[0]) );
  NOR2_X1 U20 ( .A1(n25), .A2(n57), .ZN(A_ADD[4]) );
  NOR2_X1 U21 ( .A1(n25), .A2(n61), .ZN(A_ADD[8]) );
  NOR2_X1 U22 ( .A1(n25), .A2(n58), .ZN(A_ADD[5]) );
  NOR2_X1 U23 ( .A1(n25), .A2(n62), .ZN(A_ADD[9]) );
  NOR2_X1 U24 ( .A1(n25), .A2(n59), .ZN(A_ADD[6]) );
  NOR2_X1 U25 ( .A1(n25), .A2(n56), .ZN(A_ADD[3]) );
  NOR2_X1 U26 ( .A1(n25), .A2(n60), .ZN(A_ADD[7]) );
  NOR2_X1 U27 ( .A1(n25), .A2(n55), .ZN(A_ADD[31]) );
  NOR2_X1 U28 ( .A1(n23), .A2(n38), .ZN(A_ADD[16]) );
  NOR2_X1 U29 ( .A1(n23), .A2(n34), .ZN(A_ADD[12]) );
  NOR2_X1 U30 ( .A1(n24), .A2(n47), .ZN(A_ADD[24]) );
  NOR2_X1 U31 ( .A1(n23), .A2(n42), .ZN(A_ADD[1]) );
  NOR2_X1 U32 ( .A1(n23), .A2(n35), .ZN(A_ADD[13]) );
  NOR2_X1 U33 ( .A1(n23), .A2(n39), .ZN(A_ADD[17]) );
  NOR2_X1 U34 ( .A1(n24), .A2(n48), .ZN(A_ADD[25]) );
  NOR2_X1 U35 ( .A1(n24), .A2(n44), .ZN(A_ADD[21]) );
  NOR2_X1 U36 ( .A1(n24), .A2(n43), .ZN(A_ADD[20]) );
  NOR2_X1 U37 ( .A1(n24), .A2(n52), .ZN(A_ADD[29]) );
  NOR2_X1 U38 ( .A1(n24), .A2(n51), .ZN(A_ADD[28]) );
  NOR2_X1 U39 ( .A1(n24), .A2(n53), .ZN(A_ADD[2]) );
  NOR2_X1 U40 ( .A1(n23), .A2(n32), .ZN(A_ADD[10]) );
  NOR2_X1 U41 ( .A1(n23), .A2(n36), .ZN(A_ADD[14]) );
  NOR2_X1 U42 ( .A1(n23), .A2(n40), .ZN(A_ADD[18]) );
  NOR2_X1 U43 ( .A1(n24), .A2(n45), .ZN(A_ADD[22]) );
  NOR2_X1 U44 ( .A1(n24), .A2(n49), .ZN(A_ADD[26]) );
  NOR2_X1 U45 ( .A1(n24), .A2(n54), .ZN(A_ADD[30]) );
  NOR2_X1 U46 ( .A1(n23), .A2(n33), .ZN(A_ADD[11]) );
  NOR2_X1 U47 ( .A1(n23), .A2(n37), .ZN(A_ADD[15]) );
  NOR2_X1 U48 ( .A1(n23), .A2(n41), .ZN(A_ADD[19]) );
  NOR2_X1 U49 ( .A1(n24), .A2(n46), .ZN(A_ADD[23]) );
  NOR2_X1 U50 ( .A1(n24), .A2(n50), .ZN(A_ADD[27]) );
  BUF_X1 U51 ( .A(n178), .Z(n14) );
  BUF_X1 U52 ( .A(n178), .Z(n15) );
  BUF_X1 U53 ( .A(n178), .Z(n11) );
  BUF_X1 U54 ( .A(n178), .Z(n12) );
  BUF_X1 U55 ( .A(n178), .Z(n13) );
  BUF_X1 U56 ( .A(n156), .Z(n27) );
  BUF_X1 U57 ( .A(n156), .Z(n26) );
  NAND4_X1 U58 ( .A1(n80), .A2(n81), .A3(n82), .A4(n181), .ZN(
        select_type_sig[0]) );
  INV_X1 U59 ( .A(n81), .ZN(n179) );
  NAND2_X1 U60 ( .A1(n16), .A2(n181), .ZN(select_type_sig[1]) );
  BUF_X1 U61 ( .A(n156), .Z(n28) );
  INV_X1 U62 ( .A(n80), .ZN(n177) );
  NOR2_X1 U63 ( .A1(n16), .A2(n171), .ZN(B_SHF[6]) );
  NOR2_X1 U64 ( .A1(n16), .A2(n172), .ZN(B_SHF[7]) );
  NOR2_X1 U65 ( .A1(n16), .A2(n173), .ZN(B_SHF[8]) );
  NOR2_X1 U66 ( .A1(n16), .A2(n174), .ZN(B_SHF[9]) );
  INV_X1 U67 ( .A(n82), .ZN(n176) );
  NOR2_X1 U68 ( .A1(n13), .A2(n63), .ZN(B_SHF[0]) );
  NOR2_X1 U69 ( .A1(n14), .A2(n74), .ZN(B_SHF[1]) );
  NOR2_X1 U70 ( .A1(n15), .A2(n165), .ZN(B_SHF[2]) );
  NOR2_X1 U71 ( .A1(n15), .A2(n168), .ZN(B_SHF[3]) );
  NOR2_X1 U72 ( .A1(n15), .A2(n169), .ZN(B_SHF[4]) );
  NOR2_X1 U73 ( .A1(n15), .A2(n170), .ZN(B_SHF[5]) );
  NOR2_X1 U74 ( .A1(n13), .A2(n64), .ZN(B_SHF[10]) );
  NOR2_X1 U75 ( .A1(n13), .A2(n65), .ZN(B_SHF[11]) );
  NOR2_X1 U76 ( .A1(n13), .A2(n66), .ZN(B_SHF[12]) );
  NOR2_X1 U77 ( .A1(n14), .A2(n67), .ZN(B_SHF[13]) );
  NOR2_X1 U78 ( .A1(n14), .A2(n68), .ZN(B_SHF[14]) );
  NOR2_X1 U79 ( .A1(n14), .A2(n69), .ZN(B_SHF[15]) );
  NOR2_X1 U80 ( .A1(n14), .A2(n70), .ZN(B_SHF[16]) );
  NOR2_X1 U81 ( .A1(n14), .A2(n71), .ZN(B_SHF[17]) );
  NOR2_X1 U82 ( .A1(n14), .A2(n72), .ZN(B_SHF[18]) );
  NOR2_X1 U83 ( .A1(n14), .A2(n73), .ZN(B_SHF[19]) );
  NOR2_X1 U84 ( .A1(n14), .A2(n75), .ZN(B_SHF[20]) );
  NOR2_X1 U85 ( .A1(n14), .A2(n76), .ZN(B_SHF[21]) );
  NOR2_X1 U86 ( .A1(n14), .A2(n77), .ZN(B_SHF[22]) );
  NOR2_X1 U87 ( .A1(n14), .A2(n86), .ZN(B_SHF[23]) );
  NOR2_X1 U88 ( .A1(n15), .A2(n159), .ZN(B_SHF[24]) );
  NOR2_X1 U89 ( .A1(n15), .A2(n160), .ZN(B_SHF[25]) );
  NOR2_X1 U90 ( .A1(n15), .A2(n161), .ZN(B_SHF[26]) );
  NOR2_X1 U91 ( .A1(n15), .A2(n162), .ZN(B_SHF[27]) );
  NOR2_X1 U92 ( .A1(n15), .A2(n163), .ZN(B_SHF[28]) );
  NOR2_X1 U93 ( .A1(n15), .A2(n164), .ZN(B_SHF[29]) );
  NOR2_X1 U94 ( .A1(n15), .A2(n166), .ZN(B_SHF[30]) );
  NOR2_X1 U95 ( .A1(n15), .A2(n167), .ZN(B_SHF[31]) );
  NOR2_X1 U96 ( .A1(n11), .A2(n31), .ZN(A_SHF[0]) );
  NOR2_X1 U97 ( .A1(n11), .A2(n42), .ZN(A_SHF[1]) );
  NOR2_X1 U98 ( .A1(n12), .A2(n53), .ZN(A_SHF[2]) );
  NOR2_X1 U99 ( .A1(n13), .A2(n56), .ZN(A_SHF[3]) );
  NOR2_X1 U100 ( .A1(n13), .A2(n57), .ZN(A_SHF[4]) );
  NOR2_X1 U101 ( .A1(n13), .A2(n58), .ZN(A_SHF[5]) );
  NOR2_X1 U102 ( .A1(n13), .A2(n59), .ZN(A_SHF[6]) );
  NOR2_X1 U103 ( .A1(n13), .A2(n60), .ZN(A_SHF[7]) );
  NOR2_X1 U104 ( .A1(n13), .A2(n61), .ZN(A_SHF[8]) );
  NOR2_X1 U105 ( .A1(n13), .A2(n62), .ZN(A_SHF[9]) );
  NOR2_X1 U106 ( .A1(n11), .A2(n32), .ZN(A_SHF[10]) );
  NOR2_X1 U107 ( .A1(n11), .A2(n33), .ZN(A_SHF[11]) );
  NOR2_X1 U108 ( .A1(n11), .A2(n34), .ZN(A_SHF[12]) );
  NOR2_X1 U109 ( .A1(n11), .A2(n35), .ZN(A_SHF[13]) );
  NOR2_X1 U110 ( .A1(n11), .A2(n36), .ZN(A_SHF[14]) );
  NOR2_X1 U111 ( .A1(n11), .A2(n37), .ZN(A_SHF[15]) );
  NOR2_X1 U112 ( .A1(n11), .A2(n38), .ZN(A_SHF[16]) );
  NOR2_X1 U113 ( .A1(n11), .A2(n39), .ZN(A_SHF[17]) );
  NOR2_X1 U114 ( .A1(n11), .A2(n40), .ZN(A_SHF[18]) );
  NOR2_X1 U115 ( .A1(n11), .A2(n41), .ZN(A_SHF[19]) );
  NOR2_X1 U116 ( .A1(n12), .A2(n43), .ZN(A_SHF[20]) );
  NOR2_X1 U117 ( .A1(n12), .A2(n44), .ZN(A_SHF[21]) );
  NOR2_X1 U118 ( .A1(n12), .A2(n45), .ZN(A_SHF[22]) );
  NOR2_X1 U119 ( .A1(n12), .A2(n46), .ZN(A_SHF[23]) );
  NOR2_X1 U120 ( .A1(n12), .A2(n47), .ZN(A_SHF[24]) );
  NOR2_X1 U121 ( .A1(n12), .A2(n48), .ZN(A_SHF[25]) );
  NOR2_X1 U122 ( .A1(n12), .A2(n49), .ZN(A_SHF[26]) );
  NOR2_X1 U123 ( .A1(n12), .A2(n50), .ZN(A_SHF[27]) );
  NOR2_X1 U124 ( .A1(n12), .A2(n51), .ZN(A_SHF[28]) );
  NOR2_X1 U125 ( .A1(n12), .A2(n52), .ZN(A_SHF[29]) );
  NOR2_X1 U126 ( .A1(n12), .A2(n54), .ZN(A_SHF[30]) );
  NOR2_X1 U127 ( .A1(n13), .A2(n55), .ZN(A_SHF[31]) );
  OAI22_X1 U128 ( .A1(n63), .A2(n28), .B1(OP2[0]), .B2(n29), .ZN(B_ADD[0]) );
  OAI22_X1 U129 ( .A1(n169), .A2(n26), .B1(OP2[4]), .B2(n29), .ZN(B_ADD[4]) );
  OAI22_X1 U130 ( .A1(n173), .A2(n26), .B1(OP2[8]), .B2(n29), .ZN(B_ADD[8]) );
  OAI22_X1 U131 ( .A1(n159), .A2(n27), .B1(OP2[24]), .B2(n30), .ZN(B_ADD[24])
         );
  OAI22_X1 U132 ( .A1(n74), .A2(n27), .B1(OP2[1]), .B2(n30), .ZN(B_ADD[1]) );
  OAI22_X1 U133 ( .A1(n170), .A2(n26), .B1(OP2[5]), .B2(n29), .ZN(B_ADD[5]) );
  OAI22_X1 U134 ( .A1(n174), .A2(n26), .B1(OP2[9]), .B2(n29), .ZN(B_ADD[9]) );
  OAI22_X1 U135 ( .A1(n71), .A2(n27), .B1(OP2[17]), .B2(n30), .ZN(B_ADD[17])
         );
  OAI22_X1 U136 ( .A1(n160), .A2(n27), .B1(OP2[25]), .B2(n30), .ZN(B_ADD[25])
         );
  OAI22_X1 U137 ( .A1(n76), .A2(n27), .B1(OP2[21]), .B2(n30), .ZN(B_ADD[21])
         );
  OAI22_X1 U138 ( .A1(n75), .A2(n27), .B1(OP2[20]), .B2(n30), .ZN(B_ADD[20])
         );
  OAI22_X1 U139 ( .A1(n164), .A2(n26), .B1(OP2[29]), .B2(n29), .ZN(B_ADD[29])
         );
  OAI22_X1 U140 ( .A1(n163), .A2(n26), .B1(OP2[28]), .B2(n29), .ZN(B_ADD[28])
         );
  OAI22_X1 U141 ( .A1(n165), .A2(n26), .B1(OP2[2]), .B2(n29), .ZN(B_ADD[2]) );
  OAI22_X1 U142 ( .A1(n171), .A2(n26), .B1(OP2[6]), .B2(n29), .ZN(B_ADD[6]) );
  OAI22_X1 U143 ( .A1(n72), .A2(n27), .B1(OP2[18]), .B2(n30), .ZN(B_ADD[18])
         );
  OAI22_X1 U144 ( .A1(n77), .A2(n27), .B1(OP2[22]), .B2(n30), .ZN(B_ADD[22])
         );
  OAI22_X1 U145 ( .A1(n161), .A2(n27), .B1(OP2[26]), .B2(n30), .ZN(B_ADD[26])
         );
  OAI22_X1 U146 ( .A1(n166), .A2(n26), .B1(OP2[30]), .B2(n29), .ZN(B_ADD[30])
         );
  OAI22_X1 U147 ( .A1(n168), .A2(n26), .B1(OP2[3]), .B2(n29), .ZN(B_ADD[3]) );
  OAI22_X1 U148 ( .A1(n172), .A2(n26), .B1(OP2[7]), .B2(n29), .ZN(B_ADD[7]) );
  OAI22_X1 U149 ( .A1(n73), .A2(n27), .B1(OP2[19]), .B2(n30), .ZN(B_ADD[19])
         );
  OAI22_X1 U150 ( .A1(n86), .A2(n27), .B1(OP2[23]), .B2(n30), .ZN(B_ADD[23])
         );
  OAI22_X1 U151 ( .A1(n162), .A2(n27), .B1(OP2[27]), .B2(n30), .ZN(B_ADD[27])
         );
  OAI22_X1 U152 ( .A1(n167), .A2(n26), .B1(OP2[31]), .B2(n29), .ZN(B_ADD[31])
         );
  OAI22_X1 U153 ( .A1(n70), .A2(n28), .B1(OP2[16]), .B2(n30), .ZN(B_ADD[16])
         );
  OAI22_X1 U154 ( .A1(n66), .A2(n28), .B1(OP2[12]), .B2(n29), .ZN(B_ADD[12])
         );
  OAI22_X1 U155 ( .A1(n67), .A2(n28), .B1(OP2[13]), .B2(n30), .ZN(B_ADD[13])
         );
  OAI22_X1 U156 ( .A1(n64), .A2(n28), .B1(OP2[10]), .B2(n29), .ZN(B_ADD[10])
         );
  OAI22_X1 U157 ( .A1(n68), .A2(n28), .B1(OP2[14]), .B2(n30), .ZN(B_ADD[14])
         );
  OAI22_X1 U158 ( .A1(n65), .A2(n28), .B1(OP2[11]), .B2(n29), .ZN(B_ADD[11])
         );
  OAI22_X1 U159 ( .A1(n69), .A2(n28), .B1(OP2[15]), .B2(n30), .ZN(B_ADD[15])
         );
  OAI22_X1 U160 ( .A1(n152), .A2(n63), .B1(n153), .B2(n31), .ZN(LOGIC_RES[0])
         );
  AOI21_X1 U161 ( .B1(n7), .B2(n63), .A(n19), .ZN(n153) );
  AOI221_X1 U162 ( .B1(OP1[0]), .B2(n4), .C1(n5), .C2(n31), .A(n17), .ZN(n152)
         );
  OAI22_X1 U163 ( .A1(n130), .A2(n74), .B1(n131), .B2(n42), .ZN(LOGIC_RES[1])
         );
  AOI21_X1 U164 ( .B1(n9), .B2(n74), .A(n21), .ZN(n131) );
  AOI221_X1 U165 ( .B1(OP1[1]), .B2(n3), .C1(n6), .C2(n42), .A(n18), .ZN(n130)
         );
  OAI22_X1 U166 ( .A1(n108), .A2(n165), .B1(n109), .B2(n53), .ZN(LOGIC_RES[2])
         );
  AOI21_X1 U167 ( .B1(n8), .B2(n165), .A(n20), .ZN(n109) );
  AOI221_X1 U168 ( .B1(OP1[2]), .B2(n2), .C1(n7), .C2(n53), .A(n19), .ZN(n108)
         );
  OAI22_X1 U169 ( .A1(n102), .A2(n168), .B1(n103), .B2(n56), .ZN(LOGIC_RES[3])
         );
  AOI21_X1 U170 ( .B1(n8), .B2(n168), .A(n20), .ZN(n103) );
  AOI221_X1 U171 ( .B1(OP1[3]), .B2(n2), .C1(n6), .C2(n56), .A(n18), .ZN(n102)
         );
  OAI22_X1 U172 ( .A1(n100), .A2(n169), .B1(n101), .B2(n57), .ZN(LOGIC_RES[4])
         );
  AOI21_X1 U173 ( .B1(n8), .B2(n169), .A(n20), .ZN(n101) );
  AOI221_X1 U174 ( .B1(OP1[4]), .B2(n2), .C1(n6), .C2(n57), .A(n18), .ZN(n100)
         );
  OAI22_X1 U175 ( .A1(n98), .A2(n170), .B1(n99), .B2(n58), .ZN(LOGIC_RES[5])
         );
  AOI21_X1 U176 ( .B1(n7), .B2(n170), .A(n19), .ZN(n99) );
  AOI221_X1 U177 ( .B1(OP1[5]), .B2(n2), .C1(n6), .C2(n58), .A(n18), .ZN(n98)
         );
  OAI22_X1 U178 ( .A1(n96), .A2(n171), .B1(n97), .B2(n59), .ZN(LOGIC_RES[6])
         );
  AOI21_X1 U179 ( .B1(n7), .B2(n171), .A(n19), .ZN(n97) );
  AOI221_X1 U180 ( .B1(OP1[6]), .B2(n2), .C1(n5), .C2(n59), .A(n17), .ZN(n96)
         );
  OAI22_X1 U181 ( .A1(n94), .A2(n172), .B1(n95), .B2(n60), .ZN(LOGIC_RES[7])
         );
  AOI21_X1 U182 ( .B1(n8), .B2(n172), .A(n20), .ZN(n95) );
  AOI221_X1 U183 ( .B1(OP1[7]), .B2(n2), .C1(n5), .C2(n60), .A(n17), .ZN(n94)
         );
  OAI22_X1 U184 ( .A1(n92), .A2(n173), .B1(n93), .B2(n61), .ZN(LOGIC_RES[8])
         );
  AOI21_X1 U185 ( .B1(n7), .B2(n173), .A(n19), .ZN(n93) );
  AOI221_X1 U186 ( .B1(OP1[8]), .B2(n2), .C1(n5), .C2(n61), .A(n17), .ZN(n92)
         );
  OAI22_X1 U187 ( .A1(n90), .A2(n174), .B1(n91), .B2(n62), .ZN(LOGIC_RES[9])
         );
  AOI21_X1 U188 ( .B1(n8), .B2(n174), .A(n20), .ZN(n91) );
  AOI221_X1 U189 ( .B1(n2), .B2(OP1[9]), .C1(n5), .C2(n62), .A(n17), .ZN(n90)
         );
  OAI22_X1 U190 ( .A1(n150), .A2(n64), .B1(n151), .B2(n32), .ZN(LOGIC_RES[10])
         );
  AOI21_X1 U191 ( .B1(n10), .B2(n64), .A(n22), .ZN(n151) );
  AOI221_X1 U192 ( .B1(OP1[10]), .B2(n4), .C1(n5), .C2(n32), .A(n17), .ZN(n150) );
  OAI22_X1 U193 ( .A1(n148), .A2(n65), .B1(n149), .B2(n33), .ZN(LOGIC_RES[11])
         );
  AOI21_X1 U194 ( .B1(n10), .B2(n65), .A(n22), .ZN(n149) );
  AOI221_X1 U195 ( .B1(OP1[11]), .B2(n4), .C1(n5), .C2(n33), .A(n17), .ZN(n148) );
  OAI22_X1 U196 ( .A1(n146), .A2(n66), .B1(n147), .B2(n34), .ZN(LOGIC_RES[12])
         );
  AOI21_X1 U197 ( .B1(n10), .B2(n66), .A(n21), .ZN(n147) );
  AOI221_X1 U198 ( .B1(OP1[12]), .B2(n4), .C1(n5), .C2(n34), .A(n17), .ZN(n146) );
  OAI22_X1 U199 ( .A1(n144), .A2(n67), .B1(n145), .B2(n35), .ZN(LOGIC_RES[13])
         );
  AOI21_X1 U200 ( .B1(n10), .B2(n67), .A(n21), .ZN(n145) );
  AOI221_X1 U201 ( .B1(OP1[13]), .B2(n4), .C1(n5), .C2(n35), .A(n17), .ZN(n144) );
  OAI22_X1 U202 ( .A1(n142), .A2(n68), .B1(n143), .B2(n36), .ZN(LOGIC_RES[14])
         );
  AOI21_X1 U203 ( .B1(n9), .B2(n68), .A(n21), .ZN(n143) );
  AOI221_X1 U204 ( .B1(OP1[14]), .B2(n4), .C1(n5), .C2(n36), .A(n17), .ZN(n142) );
  OAI22_X1 U205 ( .A1(n140), .A2(n69), .B1(n141), .B2(n37), .ZN(LOGIC_RES[15])
         );
  AOI21_X1 U206 ( .B1(n9), .B2(n69), .A(n21), .ZN(n141) );
  AOI221_X1 U207 ( .B1(OP1[15]), .B2(n4), .C1(n5), .C2(n37), .A(n17), .ZN(n140) );
  OAI22_X1 U208 ( .A1(n138), .A2(n70), .B1(n139), .B2(n38), .ZN(LOGIC_RES[16])
         );
  AOI21_X1 U209 ( .B1(n9), .B2(n70), .A(n21), .ZN(n139) );
  AOI221_X1 U210 ( .B1(OP1[16]), .B2(n4), .C1(n5), .C2(n38), .A(n17), .ZN(n138) );
  OAI22_X1 U211 ( .A1(n136), .A2(n71), .B1(n137), .B2(n39), .ZN(LOGIC_RES[17])
         );
  AOI21_X1 U212 ( .B1(n9), .B2(n71), .A(n21), .ZN(n137) );
  AOI221_X1 U213 ( .B1(OP1[17]), .B2(n3), .C1(n6), .C2(n39), .A(n18), .ZN(n136) );
  OAI22_X1 U214 ( .A1(n134), .A2(n72), .B1(n135), .B2(n40), .ZN(LOGIC_RES[18])
         );
  AOI21_X1 U215 ( .B1(n9), .B2(n72), .A(n21), .ZN(n135) );
  AOI221_X1 U216 ( .B1(OP1[18]), .B2(n3), .C1(n6), .C2(n40), .A(n18), .ZN(n134) );
  OAI22_X1 U217 ( .A1(n132), .A2(n73), .B1(n133), .B2(n41), .ZN(LOGIC_RES[19])
         );
  AOI21_X1 U218 ( .B1(n9), .B2(n73), .A(n21), .ZN(n133) );
  AOI221_X1 U219 ( .B1(OP1[19]), .B2(n3), .C1(n6), .C2(n41), .A(n18), .ZN(n132) );
  OAI22_X1 U220 ( .A1(n128), .A2(n75), .B1(n129), .B2(n43), .ZN(LOGIC_RES[20])
         );
  AOI21_X1 U221 ( .B1(n9), .B2(n75), .A(n21), .ZN(n129) );
  AOI221_X1 U222 ( .B1(OP1[20]), .B2(n3), .C1(n6), .C2(n43), .A(n18), .ZN(n128) );
  OAI22_X1 U223 ( .A1(n126), .A2(n76), .B1(n127), .B2(n44), .ZN(LOGIC_RES[21])
         );
  AOI21_X1 U224 ( .B1(n9), .B2(n76), .A(n21), .ZN(n127) );
  AOI221_X1 U225 ( .B1(OP1[21]), .B2(n3), .C1(n6), .C2(n44), .A(n18), .ZN(n126) );
  OAI22_X1 U226 ( .A1(n124), .A2(n77), .B1(n125), .B2(n45), .ZN(LOGIC_RES[22])
         );
  AOI21_X1 U227 ( .B1(n9), .B2(n77), .A(n21), .ZN(n125) );
  AOI221_X1 U228 ( .B1(OP1[22]), .B2(n3), .C1(n6), .C2(n45), .A(n18), .ZN(n124) );
  OAI22_X1 U229 ( .A1(n122), .A2(n86), .B1(n123), .B2(n46), .ZN(LOGIC_RES[23])
         );
  AOI21_X1 U230 ( .B1(n9), .B2(n86), .A(n21), .ZN(n123) );
  AOI221_X1 U231 ( .B1(OP1[23]), .B2(n3), .C1(n6), .C2(n46), .A(n18), .ZN(n122) );
  OAI22_X1 U232 ( .A1(n120), .A2(n159), .B1(n121), .B2(n47), .ZN(LOGIC_RES[24]) );
  AOI21_X1 U233 ( .B1(n9), .B2(n159), .A(n20), .ZN(n121) );
  AOI221_X1 U234 ( .B1(OP1[24]), .B2(n3), .C1(n7), .C2(n47), .A(n19), .ZN(n120) );
  OAI22_X1 U235 ( .A1(n118), .A2(n160), .B1(n119), .B2(n48), .ZN(LOGIC_RES[25]) );
  AOI21_X1 U236 ( .B1(n8), .B2(n160), .A(n20), .ZN(n119) );
  AOI221_X1 U237 ( .B1(OP1[25]), .B2(n3), .C1(n7), .C2(n48), .A(n19), .ZN(n118) );
  OAI22_X1 U238 ( .A1(n116), .A2(n161), .B1(n117), .B2(n49), .ZN(LOGIC_RES[26]) );
  AOI21_X1 U239 ( .B1(n8), .B2(n161), .A(n20), .ZN(n117) );
  AOI221_X1 U240 ( .B1(OP1[26]), .B2(n3), .C1(n6), .C2(n49), .A(n18), .ZN(n116) );
  OAI22_X1 U241 ( .A1(n114), .A2(n162), .B1(n115), .B2(n50), .ZN(LOGIC_RES[27]) );
  AOI21_X1 U242 ( .B1(n8), .B2(n162), .A(n20), .ZN(n115) );
  AOI221_X1 U243 ( .B1(OP1[27]), .B2(n3), .C1(n7), .C2(n50), .A(n19), .ZN(n114) );
  OAI22_X1 U244 ( .A1(n112), .A2(n163), .B1(n113), .B2(n51), .ZN(LOGIC_RES[28]) );
  AOI21_X1 U245 ( .B1(n8), .B2(n163), .A(n20), .ZN(n113) );
  AOI221_X1 U246 ( .B1(OP1[28]), .B2(n2), .C1(n7), .C2(n51), .A(n19), .ZN(n112) );
  OAI22_X1 U247 ( .A1(n110), .A2(n164), .B1(n111), .B2(n52), .ZN(LOGIC_RES[29]) );
  AOI21_X1 U248 ( .B1(n8), .B2(n164), .A(n20), .ZN(n111) );
  AOI221_X1 U249 ( .B1(OP1[29]), .B2(n2), .C1(n7), .C2(n52), .A(n19), .ZN(n110) );
  OAI22_X1 U250 ( .A1(n106), .A2(n166), .B1(n107), .B2(n54), .ZN(LOGIC_RES[30]) );
  AOI21_X1 U251 ( .B1(n8), .B2(n166), .A(n20), .ZN(n107) );
  AOI221_X1 U252 ( .B1(OP1[30]), .B2(n2), .C1(n7), .C2(n54), .A(n19), .ZN(n106) );
  OAI22_X1 U253 ( .A1(n104), .A2(n167), .B1(n105), .B2(n55), .ZN(LOGIC_RES[31]) );
  AOI21_X1 U254 ( .B1(n8), .B2(n167), .A(n20), .ZN(n105) );
  AOI221_X1 U255 ( .B1(OP1[31]), .B2(n2), .C1(n7), .C2(n55), .A(n19), .ZN(n104) );
  INV_X1 U256 ( .A(\OPSel[0] ), .ZN(n181) );
  INV_X1 U257 ( .A(OP1[4]), .ZN(n57) );
  INV_X1 U258 ( .A(OP1[0]), .ZN(n31) );
  INV_X1 U259 ( .A(OP1[8]), .ZN(n61) );
  INV_X1 U260 ( .A(OP1[16]), .ZN(n38) );
  INV_X1 U261 ( .A(OP1[12]), .ZN(n34) );
  INV_X1 U262 ( .A(OP1[24]), .ZN(n47) );
  INV_X1 U263 ( .A(OP1[1]), .ZN(n42) );
  INV_X1 U264 ( .A(OP1[5]), .ZN(n58) );
  INV_X1 U265 ( .A(OP1[9]), .ZN(n62) );
  INV_X1 U266 ( .A(OP1[13]), .ZN(n35) );
  INV_X1 U267 ( .A(OP1[17]), .ZN(n39) );
  INV_X1 U268 ( .A(OP1[25]), .ZN(n48) );
  INV_X1 U269 ( .A(OP1[21]), .ZN(n44) );
  INV_X1 U270 ( .A(OP1[20]), .ZN(n43) );
  INV_X1 U271 ( .A(OP1[29]), .ZN(n52) );
  INV_X1 U272 ( .A(OP1[28]), .ZN(n51) );
  INV_X1 U273 ( .A(OP1[2]), .ZN(n53) );
  INV_X1 U274 ( .A(OP1[6]), .ZN(n59) );
  INV_X1 U275 ( .A(OP1[10]), .ZN(n32) );
  INV_X1 U276 ( .A(OP1[14]), .ZN(n36) );
  INV_X1 U277 ( .A(OP1[18]), .ZN(n40) );
  INV_X1 U278 ( .A(OP1[22]), .ZN(n45) );
  INV_X1 U279 ( .A(OP1[26]), .ZN(n49) );
  INV_X1 U280 ( .A(OP1[30]), .ZN(n54) );
  INV_X1 U281 ( .A(OP1[3]), .ZN(n56) );
  INV_X1 U282 ( .A(OP1[7]), .ZN(n60) );
  INV_X1 U283 ( .A(OP1[11]), .ZN(n33) );
  INV_X1 U284 ( .A(OP1[15]), .ZN(n37) );
  INV_X1 U285 ( .A(OP1[19]), .ZN(n41) );
  INV_X1 U286 ( .A(OP1[23]), .ZN(n46) );
  INV_X1 U287 ( .A(OP1[27]), .ZN(n50) );
  INV_X1 U288 ( .A(OP1[31]), .ZN(n55) );
  INV_X1 U289 ( .A(OP2[4]), .ZN(n169) );
  INV_X1 U290 ( .A(OP2[0]), .ZN(n63) );
  INV_X1 U291 ( .A(OP2[8]), .ZN(n173) );
  INV_X1 U292 ( .A(OP2[16]), .ZN(n70) );
  INV_X1 U293 ( .A(OP2[12]), .ZN(n66) );
  INV_X1 U294 ( .A(OP2[24]), .ZN(n159) );
  INV_X1 U295 ( .A(OP2[1]), .ZN(n74) );
  INV_X1 U296 ( .A(OP2[5]), .ZN(n170) );
  INV_X1 U297 ( .A(OP2[9]), .ZN(n174) );
  INV_X1 U298 ( .A(OP2[13]), .ZN(n67) );
  INV_X1 U299 ( .A(OP2[17]), .ZN(n71) );
  INV_X1 U300 ( .A(OP2[25]), .ZN(n160) );
  INV_X1 U301 ( .A(OP2[21]), .ZN(n76) );
  INV_X1 U302 ( .A(OP2[20]), .ZN(n75) );
  INV_X1 U303 ( .A(OP2[29]), .ZN(n164) );
  INV_X1 U304 ( .A(OP2[28]), .ZN(n163) );
  INV_X1 U305 ( .A(OP2[2]), .ZN(n165) );
  INV_X1 U306 ( .A(OP2[6]), .ZN(n171) );
  INV_X1 U307 ( .A(OP2[10]), .ZN(n64) );
  INV_X1 U308 ( .A(OP2[14]), .ZN(n68) );
  INV_X1 U309 ( .A(OP2[18]), .ZN(n72) );
  INV_X1 U310 ( .A(OP2[22]), .ZN(n77) );
  INV_X1 U311 ( .A(OP2[26]), .ZN(n161) );
  INV_X1 U312 ( .A(OP2[30]), .ZN(n166) );
  INV_X1 U313 ( .A(OP2[3]), .ZN(n168) );
  INV_X1 U314 ( .A(OP2[7]), .ZN(n172) );
  INV_X1 U315 ( .A(OP2[11]), .ZN(n65) );
  INV_X1 U316 ( .A(OP2[15]), .ZN(n69) );
  INV_X1 U325 ( .A(OP2[19]), .ZN(n73) );
  INV_X1 U326 ( .A(OP2[23]), .ZN(n86) );
  INV_X1 U327 ( .A(OP2[27]), .ZN(n162) );
  INV_X1 U328 ( .A(OP2[31]), .ZN(n167) );
  AND2_X1 U329 ( .A1(n154), .A2(n89), .ZN(n1) );
  INV_X1 U330 ( .A(n83), .ZN(n182) );
  NAND2_X1 U331 ( .A1(n155), .A2(n89), .ZN(n82) );
  INV_X1 U332 ( .A(LOGIC_ARITH), .ZN(n178) );
  NAND2_X1 U333 ( .A1(n155), .A2(n88), .ZN(n80) );
  NAND2_X1 U334 ( .A1(n154), .A2(n88), .ZN(n81) );
  INV_X1 U335 ( .A(n84), .ZN(n183) );
  INV_X1 U336 ( .A(n85), .ZN(n180) );
  NOR2_X1 U337 ( .A1(n185), .A2(ALU_OPC[2]), .ZN(n89) );
  NOR2_X1 U338 ( .A1(n186), .A2(ALU_OPC[3]), .ZN(n155) );
  NOR2_X1 U339 ( .A1(n184), .A2(ALU_OPC[1]), .ZN(n88) );
  NOR2_X1 U340 ( .A1(ALU_OPC[3]), .A2(ALU_OPC[0]), .ZN(n154) );
  OAI21_X1 U341 ( .B1(n78), .B2(n175), .A(n79), .ZN(select_zero_sig) );
  INV_X1 U342 ( .A(ALU_OPC[3]), .ZN(n175) );
  AOI22_X1 U343 ( .A1(ALU_OPC[0]), .A2(n185), .B1(ALU_OPC[2]), .B2(ALU_OPC[1]), 
        .ZN(n78) );
  INV_X1 U344 ( .A(ALU_OPC[1]), .ZN(n185) );
  INV_X1 U345 ( .A(ALU_OPC[0]), .ZN(n186) );
  INV_X1 U346 ( .A(ALU_OPC[2]), .ZN(n184) );
  NAND2_X1 U347 ( .A1(n85), .A2(n157), .ZN(LOGIC_ARITH) );
  CLKBUF_X1 U348 ( .A(n177), .Z(n10) );
  CLKBUF_X1 U349 ( .A(n178), .Z(n16) );
  CLKBUF_X1 U350 ( .A(n179), .Z(n22) );
  INV_X1 U351 ( .A(n1), .ZN(n29) );
  INV_X1 U352 ( .A(n1), .ZN(n30) );
endmodule


module regn_N32_6 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n68, n69, n70;

  DFFR_X1 \DOUT_reg[31]  ( .D(n36), .CK(CLK), .RN(n3), .Q(DOUT[31]) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n37), .CK(CLK), .RN(n3), .Q(DOUT[30]) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n38), .CK(CLK), .RN(n3), .Q(DOUT[29]) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n39), .CK(CLK), .RN(n3), .Q(DOUT[28]) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n40), .CK(CLK), .RN(n3), .Q(DOUT[27]) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n41), .CK(CLK), .RN(n3), .Q(DOUT[26]) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n42), .CK(CLK), .RN(n3), .Q(DOUT[25]) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n43), .CK(CLK), .RN(n3), .Q(DOUT[24]) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n44), .CK(CLK), .RN(n2), .Q(DOUT[23]) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n45), .CK(CLK), .RN(n2), .Q(DOUT[22]) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n46), .CK(CLK), .RN(n2), .Q(DOUT[21]) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n47), .CK(CLK), .RN(n2), .Q(DOUT[20]) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n48), .CK(CLK), .RN(n2), .Q(DOUT[19]) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n49), .CK(CLK), .RN(n2), .Q(DOUT[18]) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n50), .CK(CLK), .RN(n2), .Q(DOUT[17]) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n51), .CK(CLK), .RN(n2), .Q(DOUT[16]) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n52), .CK(CLK), .RN(n2), .Q(DOUT[15]) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n53), .CK(CLK), .RN(n2), .Q(DOUT[14]) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n54), .CK(CLK), .RN(n2), .Q(DOUT[13]) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n55), .CK(CLK), .RN(n2), .Q(DOUT[12]) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n56), .CK(CLK), .RN(n1), .Q(DOUT[11]) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n57), .CK(CLK), .RN(n1), .Q(DOUT[10]) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n58), .CK(CLK), .RN(n1), .Q(DOUT[9]) );
  DFFR_X1 \DOUT_reg[8]  ( .D(n59), .CK(CLK), .RN(n1), .Q(DOUT[8]) );
  DFFR_X1 \DOUT_reg[7]  ( .D(n60), .CK(CLK), .RN(n1), .Q(DOUT[7]) );
  DFFR_X1 \DOUT_reg[6]  ( .D(n61), .CK(CLK), .RN(n1), .Q(DOUT[6]) );
  DFFR_X1 \DOUT_reg[5]  ( .D(n62), .CK(CLK), .RN(n1), .Q(DOUT[5]) );
  DFFR_X1 \DOUT_reg[4]  ( .D(n63), .CK(CLK), .RN(n1), .Q(DOUT[4]) );
  DFFR_X1 \DOUT_reg[3]  ( .D(n64), .CK(CLK), .RN(n1), .Q(DOUT[3]) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n68), .CK(CLK), .RN(n1), .Q(DOUT[2]) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n69), .CK(CLK), .RN(n1), .Q(DOUT[1]) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n70), .CK(CLK), .RN(n1), .Q(DOUT[0]) );
  BUF_X1 U2 ( .A(RST), .Z(n1) );
  BUF_X1 U3 ( .A(RST), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n3) );
  MUX2_X1 U5 ( .A(DOUT[0]), .B(DIN[0]), .S(EN), .Z(n70) );
  MUX2_X1 U6 ( .A(DOUT[1]), .B(DIN[1]), .S(EN), .Z(n69) );
  MUX2_X1 U7 ( .A(DOUT[2]), .B(DIN[2]), .S(EN), .Z(n68) );
  MUX2_X1 U8 ( .A(DOUT[3]), .B(DIN[3]), .S(EN), .Z(n64) );
  MUX2_X1 U9 ( .A(DOUT[4]), .B(DIN[4]), .S(EN), .Z(n63) );
  MUX2_X1 U10 ( .A(DOUT[5]), .B(DIN[5]), .S(EN), .Z(n62) );
  MUX2_X1 U11 ( .A(DOUT[6]), .B(DIN[6]), .S(EN), .Z(n61) );
  MUX2_X1 U12 ( .A(DOUT[7]), .B(DIN[7]), .S(EN), .Z(n60) );
  MUX2_X1 U13 ( .A(DOUT[8]), .B(DIN[8]), .S(EN), .Z(n59) );
  MUX2_X1 U14 ( .A(DOUT[9]), .B(DIN[9]), .S(EN), .Z(n58) );
  MUX2_X1 U15 ( .A(DOUT[10]), .B(DIN[10]), .S(EN), .Z(n57) );
  MUX2_X1 U16 ( .A(DOUT[11]), .B(DIN[11]), .S(EN), .Z(n56) );
  MUX2_X1 U17 ( .A(DOUT[12]), .B(DIN[12]), .S(EN), .Z(n55) );
  MUX2_X1 U18 ( .A(DOUT[13]), .B(DIN[13]), .S(EN), .Z(n54) );
  MUX2_X1 U19 ( .A(DOUT[14]), .B(DIN[14]), .S(EN), .Z(n53) );
  MUX2_X1 U20 ( .A(DOUT[15]), .B(DIN[15]), .S(EN), .Z(n52) );
  MUX2_X1 U21 ( .A(DOUT[16]), .B(DIN[16]), .S(EN), .Z(n51) );
  MUX2_X1 U22 ( .A(DOUT[17]), .B(DIN[17]), .S(EN), .Z(n50) );
  MUX2_X1 U23 ( .A(DOUT[18]), .B(DIN[18]), .S(EN), .Z(n49) );
  MUX2_X1 U24 ( .A(DOUT[19]), .B(DIN[19]), .S(EN), .Z(n48) );
  MUX2_X1 U25 ( .A(DOUT[20]), .B(DIN[20]), .S(EN), .Z(n47) );
  MUX2_X1 U26 ( .A(DOUT[21]), .B(DIN[21]), .S(EN), .Z(n46) );
  MUX2_X1 U27 ( .A(DOUT[22]), .B(DIN[22]), .S(EN), .Z(n45) );
  MUX2_X1 U28 ( .A(DOUT[23]), .B(DIN[23]), .S(EN), .Z(n44) );
  MUX2_X1 U29 ( .A(DOUT[24]), .B(DIN[24]), .S(EN), .Z(n43) );
  MUX2_X1 U30 ( .A(DOUT[25]), .B(DIN[25]), .S(EN), .Z(n42) );
  MUX2_X1 U31 ( .A(DOUT[26]), .B(DIN[26]), .S(EN), .Z(n41) );
  MUX2_X1 U32 ( .A(DOUT[27]), .B(DIN[27]), .S(EN), .Z(n40) );
  MUX2_X1 U33 ( .A(DOUT[28]), .B(DIN[28]), .S(EN), .Z(n39) );
  MUX2_X1 U34 ( .A(DOUT[29]), .B(DIN[29]), .S(EN), .Z(n38) );
  MUX2_X1 U35 ( .A(DOUT[30]), .B(DIN[30]), .S(EN), .Z(n37) );
  MUX2_X1 U36 ( .A(DOUT[31]), .B(DIN[31]), .S(EN), .Z(n36) );
endmodule


module regn_N32_5 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n68, n69, n70;

  DFFR_X1 \DOUT_reg[31]  ( .D(n36), .CK(CLK), .RN(n3), .Q(DOUT[31]) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n37), .CK(CLK), .RN(n3), .Q(DOUT[30]) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n38), .CK(CLK), .RN(n3), .Q(DOUT[29]) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n39), .CK(CLK), .RN(n3), .Q(DOUT[28]) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n40), .CK(CLK), .RN(n3), .Q(DOUT[27]) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n41), .CK(CLK), .RN(n3), .Q(DOUT[26]) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n42), .CK(CLK), .RN(n3), .Q(DOUT[25]) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n43), .CK(CLK), .RN(n3), .Q(DOUT[24]) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n44), .CK(CLK), .RN(n2), .Q(DOUT[23]) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n45), .CK(CLK), .RN(n2), .Q(DOUT[22]) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n46), .CK(CLK), .RN(n2), .Q(DOUT[21]) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n47), .CK(CLK), .RN(n2), .Q(DOUT[20]) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n48), .CK(CLK), .RN(n2), .Q(DOUT[19]) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n49), .CK(CLK), .RN(n2), .Q(DOUT[18]) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n50), .CK(CLK), .RN(n2), .Q(DOUT[17]) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n51), .CK(CLK), .RN(n2), .Q(DOUT[16]) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n52), .CK(CLK), .RN(n2), .Q(DOUT[15]) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n53), .CK(CLK), .RN(n2), .Q(DOUT[14]) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n54), .CK(CLK), .RN(n2), .Q(DOUT[13]) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n55), .CK(CLK), .RN(n2), .Q(DOUT[12]) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n56), .CK(CLK), .RN(n1), .Q(DOUT[11]) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n57), .CK(CLK), .RN(n1), .Q(DOUT[10]) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n58), .CK(CLK), .RN(n1), .Q(DOUT[9]) );
  DFFR_X1 \DOUT_reg[8]  ( .D(n59), .CK(CLK), .RN(n1), .Q(DOUT[8]) );
  DFFR_X1 \DOUT_reg[7]  ( .D(n60), .CK(CLK), .RN(n1), .Q(DOUT[7]) );
  DFFR_X1 \DOUT_reg[6]  ( .D(n61), .CK(CLK), .RN(n1), .Q(DOUT[6]) );
  DFFR_X1 \DOUT_reg[5]  ( .D(n62), .CK(CLK), .RN(n1), .Q(DOUT[5]) );
  DFFR_X1 \DOUT_reg[4]  ( .D(n63), .CK(CLK), .RN(n1), .Q(DOUT[4]) );
  DFFR_X1 \DOUT_reg[3]  ( .D(n64), .CK(CLK), .RN(n1), .Q(DOUT[3]) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n68), .CK(CLK), .RN(n1), .Q(DOUT[2]) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n69), .CK(CLK), .RN(n1), .Q(DOUT[1]) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n70), .CK(CLK), .RN(n1), .Q(DOUT[0]) );
  BUF_X1 U2 ( .A(RST), .Z(n1) );
  BUF_X1 U3 ( .A(RST), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n3) );
  MUX2_X1 U5 ( .A(DOUT[0]), .B(DIN[0]), .S(EN), .Z(n70) );
  MUX2_X1 U6 ( .A(DOUT[1]), .B(DIN[1]), .S(EN), .Z(n69) );
  MUX2_X1 U7 ( .A(DOUT[2]), .B(DIN[2]), .S(EN), .Z(n68) );
  MUX2_X1 U8 ( .A(DOUT[3]), .B(DIN[3]), .S(EN), .Z(n64) );
  MUX2_X1 U9 ( .A(DOUT[4]), .B(DIN[4]), .S(EN), .Z(n63) );
  MUX2_X1 U10 ( .A(DOUT[5]), .B(DIN[5]), .S(EN), .Z(n62) );
  MUX2_X1 U11 ( .A(DOUT[6]), .B(DIN[6]), .S(EN), .Z(n61) );
  MUX2_X1 U12 ( .A(DOUT[7]), .B(DIN[7]), .S(EN), .Z(n60) );
  MUX2_X1 U13 ( .A(DOUT[8]), .B(DIN[8]), .S(EN), .Z(n59) );
  MUX2_X1 U14 ( .A(DOUT[9]), .B(DIN[9]), .S(EN), .Z(n58) );
  MUX2_X1 U15 ( .A(DOUT[10]), .B(DIN[10]), .S(EN), .Z(n57) );
  MUX2_X1 U16 ( .A(DOUT[11]), .B(DIN[11]), .S(EN), .Z(n56) );
  MUX2_X1 U17 ( .A(DOUT[12]), .B(DIN[12]), .S(EN), .Z(n55) );
  MUX2_X1 U18 ( .A(DOUT[13]), .B(DIN[13]), .S(EN), .Z(n54) );
  MUX2_X1 U19 ( .A(DOUT[14]), .B(DIN[14]), .S(EN), .Z(n53) );
  MUX2_X1 U20 ( .A(DOUT[15]), .B(DIN[15]), .S(EN), .Z(n52) );
  MUX2_X1 U21 ( .A(DOUT[16]), .B(DIN[16]), .S(EN), .Z(n51) );
  MUX2_X1 U22 ( .A(DOUT[17]), .B(DIN[17]), .S(EN), .Z(n50) );
  MUX2_X1 U23 ( .A(DOUT[18]), .B(DIN[18]), .S(EN), .Z(n49) );
  MUX2_X1 U24 ( .A(DOUT[19]), .B(DIN[19]), .S(EN), .Z(n48) );
  MUX2_X1 U25 ( .A(DOUT[20]), .B(DIN[20]), .S(EN), .Z(n47) );
  MUX2_X1 U26 ( .A(DOUT[21]), .B(DIN[21]), .S(EN), .Z(n46) );
  MUX2_X1 U27 ( .A(DOUT[22]), .B(DIN[22]), .S(EN), .Z(n45) );
  MUX2_X1 U28 ( .A(DOUT[23]), .B(DIN[23]), .S(EN), .Z(n44) );
  MUX2_X1 U29 ( .A(DOUT[24]), .B(DIN[24]), .S(EN), .Z(n43) );
  MUX2_X1 U30 ( .A(DOUT[25]), .B(DIN[25]), .S(EN), .Z(n42) );
  MUX2_X1 U31 ( .A(DOUT[26]), .B(DIN[26]), .S(EN), .Z(n41) );
  MUX2_X1 U32 ( .A(DOUT[27]), .B(DIN[27]), .S(EN), .Z(n40) );
  MUX2_X1 U33 ( .A(DOUT[28]), .B(DIN[28]), .S(EN), .Z(n39) );
  MUX2_X1 U34 ( .A(DOUT[29]), .B(DIN[29]), .S(EN), .Z(n38) );
  MUX2_X1 U35 ( .A(DOUT[30]), .B(DIN[30]), .S(EN), .Z(n37) );
  MUX2_X1 U36 ( .A(DOUT[31]), .B(DIN[31]), .S(EN), .Z(n36) );
endmodule


module regn_N5_2 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n6, n7, n8, n9, n10;

  DFFR_X1 \DOUT_reg[4]  ( .D(n6), .CK(CLK), .RN(RST), .Q(DOUT[4]) );
  DFFR_X1 \DOUT_reg[3]  ( .D(n7), .CK(CLK), .RN(RST), .Q(DOUT[3]) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n8), .CK(CLK), .RN(RST), .Q(DOUT[2]) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n9), .CK(CLK), .RN(RST), .Q(DOUT[1]) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n10), .CK(CLK), .RN(RST), .Q(DOUT[0]) );
  MUX2_X1 U2 ( .A(DOUT[0]), .B(DIN[0]), .S(EN), .Z(n10) );
  MUX2_X1 U3 ( .A(DOUT[1]), .B(DIN[1]), .S(EN), .Z(n9) );
  MUX2_X1 U4 ( .A(DOUT[2]), .B(DIN[2]), .S(EN), .Z(n8) );
  MUX2_X1 U5 ( .A(DOUT[3]), .B(DIN[3]), .S(EN), .Z(n7) );
  MUX2_X1 U6 ( .A(DOUT[4]), .B(DIN[4]), .S(EN), .Z(n6) );
endmodule


module regn_N32_4 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17, n18,
         n19, n20, n22, n23, n24, n25, n26, n28, n29, n30, n31, n32, n33, n34,
         n42, n50, n56, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151;

  DFFR_X1 \DOUT_reg[31]  ( .D(n50), .CK(CLK), .RN(n3), .Q(DOUT[31]), .QN(n125)
         );
  DFFR_X1 \DOUT_reg[30]  ( .D(n56), .CK(CLK), .RN(n3), .Q(DOUT[30]), .QN(n126)
         );
  DFFR_X1 \DOUT_reg[29]  ( .D(n95), .CK(CLK), .RN(n3), .Q(DOUT[29]), .QN(n127)
         );
  DFFR_X1 \DOUT_reg[28]  ( .D(n96), .CK(CLK), .RN(n3), .Q(DOUT[28]), .QN(n128)
         );
  DFFR_X1 \DOUT_reg[27]  ( .D(n97), .CK(CLK), .RN(n3), .Q(DOUT[27]), .QN(n129)
         );
  DFFR_X1 \DOUT_reg[26]  ( .D(n98), .CK(CLK), .RN(n3), .Q(DOUT[26]), .QN(n130)
         );
  DFFR_X1 \DOUT_reg[25]  ( .D(n99), .CK(CLK), .RN(n3), .Q(DOUT[25]), .QN(n131)
         );
  DFFR_X1 \DOUT_reg[24]  ( .D(n100), .CK(CLK), .RN(n3), .Q(DOUT[24]), .QN(n132) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n101), .CK(CLK), .RN(n2), .Q(DOUT[23]) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n102), .CK(CLK), .RN(n2), .Q(DOUT[22]), .QN(n133) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n103), .CK(CLK), .RN(n2), .Q(DOUT[21]), .QN(n134) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n104), .CK(CLK), .RN(n2), .Q(DOUT[20]), .QN(n135) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n105), .CK(CLK), .RN(n2), .Q(DOUT[19]), .QN(n136) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n106), .CK(CLK), .RN(n2), .Q(DOUT[18]), .QN(n137) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n107), .CK(CLK), .RN(n2), .Q(DOUT[17]) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n108), .CK(CLK), .RN(n2), .Q(DOUT[16]), .QN(n138) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n109), .CK(CLK), .RN(n2), .Q(DOUT[15]), .QN(n139) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n110), .CK(CLK), .RN(n2), .Q(DOUT[14]), .QN(n140) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n111), .CK(CLK), .RN(n2), .Q(DOUT[13]), .QN(n141) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n112), .CK(CLK), .RN(n2), .Q(DOUT[12]), .QN(n142) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n113), .CK(CLK), .RN(n1), .Q(DOUT[11]), .QN(n143) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n114), .CK(CLK), .RN(n1), .Q(DOUT[10]), .QN(n144) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n115), .CK(CLK), .RN(n1), .Q(DOUT[9]) );
  DFFR_X1 \DOUT_reg[8]  ( .D(n116), .CK(CLK), .RN(n1), .Q(DOUT[8]), .QN(n145)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n117), .CK(CLK), .RN(n1), .Q(DOUT[7]), .QN(n146)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n118), .CK(CLK), .RN(n1), .Q(DOUT[6]), .QN(n147)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n119), .CK(CLK), .RN(n1), .Q(DOUT[5]), .QN(n148)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n120), .CK(CLK), .RN(n1), .Q(DOUT[4]), .QN(n149)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n121), .CK(CLK), .RN(n1), .Q(DOUT[3]), .QN(n150)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n122), .CK(CLK), .RN(n1), .Q(DOUT[2]), .QN(n151)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n123), .CK(CLK), .RN(n1), .Q(DOUT[1]) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n124), .CK(CLK), .RN(n1), .Q(DOUT[0]) );
  BUF_X1 U2 ( .A(RST), .Z(n1) );
  BUF_X1 U3 ( .A(RST), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n3) );
  MUX2_X1 U5 ( .A(DOUT[0]), .B(DIN[0]), .S(EN), .Z(n124) );
  MUX2_X1 U6 ( .A(DOUT[1]), .B(DIN[1]), .S(EN), .Z(n123) );
  INV_X1 U7 ( .A(n151), .ZN(n6) );
  MUX2_X1 U8 ( .A(n6), .B(DIN[2]), .S(EN), .Z(n122) );
  INV_X1 U9 ( .A(n150), .ZN(n7) );
  MUX2_X1 U10 ( .A(n7), .B(DIN[3]), .S(EN), .Z(n121) );
  INV_X1 U11 ( .A(n149), .ZN(n8) );
  MUX2_X1 U12 ( .A(n8), .B(DIN[4]), .S(EN), .Z(n120) );
  INV_X1 U13 ( .A(n148), .ZN(n9) );
  MUX2_X1 U14 ( .A(n9), .B(DIN[5]), .S(EN), .Z(n119) );
  INV_X1 U15 ( .A(n147), .ZN(n10) );
  MUX2_X1 U16 ( .A(n10), .B(DIN[6]), .S(EN), .Z(n118) );
  INV_X1 U17 ( .A(n146), .ZN(n11) );
  MUX2_X1 U18 ( .A(n11), .B(DIN[7]), .S(EN), .Z(n117) );
  INV_X1 U19 ( .A(n145), .ZN(n12) );
  MUX2_X1 U20 ( .A(n12), .B(DIN[8]), .S(EN), .Z(n116) );
  MUX2_X1 U21 ( .A(DOUT[9]), .B(DIN[9]), .S(EN), .Z(n115) );
  INV_X1 U22 ( .A(n144), .ZN(n14) );
  MUX2_X1 U23 ( .A(n14), .B(DIN[10]), .S(EN), .Z(n114) );
  INV_X1 U24 ( .A(n143), .ZN(n15) );
  MUX2_X1 U25 ( .A(n15), .B(DIN[11]), .S(EN), .Z(n113) );
  INV_X1 U26 ( .A(n142), .ZN(n16) );
  MUX2_X1 U27 ( .A(n16), .B(DIN[12]), .S(EN), .Z(n112) );
  INV_X1 U28 ( .A(n141), .ZN(n17) );
  MUX2_X1 U29 ( .A(n17), .B(DIN[13]), .S(EN), .Z(n111) );
  INV_X1 U30 ( .A(n140), .ZN(n18) );
  MUX2_X1 U31 ( .A(n18), .B(DIN[14]), .S(EN), .Z(n110) );
  INV_X1 U32 ( .A(n139), .ZN(n19) );
  MUX2_X1 U33 ( .A(n19), .B(DIN[15]), .S(EN), .Z(n109) );
  INV_X1 U34 ( .A(n138), .ZN(n20) );
  MUX2_X1 U35 ( .A(n20), .B(DIN[16]), .S(EN), .Z(n108) );
  MUX2_X1 U36 ( .A(DOUT[17]), .B(DIN[17]), .S(EN), .Z(n107) );
  INV_X1 U37 ( .A(n137), .ZN(n22) );
  MUX2_X1 U38 ( .A(n22), .B(DIN[18]), .S(EN), .Z(n106) );
  INV_X1 U39 ( .A(n136), .ZN(n23) );
  MUX2_X1 U40 ( .A(n23), .B(DIN[19]), .S(EN), .Z(n105) );
  INV_X1 U41 ( .A(n135), .ZN(n24) );
  MUX2_X1 U42 ( .A(n24), .B(DIN[20]), .S(EN), .Z(n104) );
  INV_X1 U43 ( .A(n134), .ZN(n25) );
  MUX2_X1 U44 ( .A(n25), .B(DIN[21]), .S(EN), .Z(n103) );
  INV_X1 U45 ( .A(n133), .ZN(n26) );
  MUX2_X1 U46 ( .A(n26), .B(DIN[22]), .S(EN), .Z(n102) );
  MUX2_X1 U47 ( .A(DOUT[23]), .B(DIN[23]), .S(EN), .Z(n101) );
  INV_X1 U48 ( .A(n132), .ZN(n28) );
  MUX2_X1 U49 ( .A(n28), .B(DIN[24]), .S(EN), .Z(n100) );
  INV_X1 U50 ( .A(n131), .ZN(n29) );
  MUX2_X1 U51 ( .A(n29), .B(DIN[25]), .S(EN), .Z(n99) );
  INV_X1 U52 ( .A(n130), .ZN(n30) );
  MUX2_X1 U53 ( .A(n30), .B(DIN[26]), .S(EN), .Z(n98) );
  INV_X1 U54 ( .A(n129), .ZN(n31) );
  MUX2_X1 U55 ( .A(n31), .B(DIN[27]), .S(EN), .Z(n97) );
  INV_X1 U56 ( .A(n128), .ZN(n32) );
  MUX2_X1 U57 ( .A(n32), .B(DIN[28]), .S(EN), .Z(n96) );
  INV_X1 U58 ( .A(n127), .ZN(n33) );
  MUX2_X1 U59 ( .A(n33), .B(DIN[29]), .S(EN), .Z(n95) );
  INV_X1 U60 ( .A(n126), .ZN(n34) );
  MUX2_X1 U61 ( .A(n34), .B(DIN[30]), .S(EN), .Z(n56) );
  INV_X1 U62 ( .A(n125), .ZN(n42) );
  MUX2_X1 U63 ( .A(n42), .B(DIN[31]), .S(EN), .Z(n50) );
endmodule


module regn_N32_3 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \DOUT_reg[31]  ( .D(n100), .CK(CLK), .RN(n3), .Q(DOUT[31]), .QN(n132) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n101), .CK(CLK), .RN(n3), .Q(DOUT[30]), .QN(n133) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n102), .CK(CLK), .RN(n3), .Q(DOUT[29]), .QN(n134) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n103), .CK(CLK), .RN(n3), .Q(DOUT[28]), .QN(n135) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n104), .CK(CLK), .RN(n3), .Q(DOUT[27]), .QN(n136) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n105), .CK(CLK), .RN(n3), .Q(DOUT[26]), .QN(n137) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n106), .CK(CLK), .RN(n3), .Q(DOUT[25]), .QN(n138) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n107), .CK(CLK), .RN(n3), .Q(DOUT[24]), .QN(n139) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n108), .CK(CLK), .RN(n2), .Q(DOUT[23]), .QN(n140) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n109), .CK(CLK), .RN(n2), .Q(DOUT[22]), .QN(n141) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n110), .CK(CLK), .RN(n2), .Q(DOUT[21]), .QN(n142) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n111), .CK(CLK), .RN(n2), .Q(DOUT[20]), .QN(n143) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n112), .CK(CLK), .RN(n2), .Q(DOUT[19]), .QN(n144) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n113), .CK(CLK), .RN(n2), .Q(DOUT[18]), .QN(n145) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n114), .CK(CLK), .RN(n2), .Q(DOUT[17]), .QN(n146) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n115), .CK(CLK), .RN(n2), .Q(DOUT[16]), .QN(n147) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n116), .CK(CLK), .RN(n2), .Q(DOUT[15]), .QN(n148) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n117), .CK(CLK), .RN(n2), .Q(DOUT[14]), .QN(n149) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n118), .CK(CLK), .RN(n2), .Q(DOUT[13]), .QN(n150) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n119), .CK(CLK), .RN(n2), .Q(DOUT[12]), .QN(n151) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n120), .CK(CLK), .RN(n1), .Q(DOUT[11]), .QN(n152) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n121), .CK(CLK), .RN(n1), .Q(DOUT[10]), .QN(n153) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n122), .CK(CLK), .RN(n1), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 \DOUT_reg[8]  ( .D(n123), .CK(CLK), .RN(n1), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 \DOUT_reg[7]  ( .D(n124), .CK(CLK), .RN(n1), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 \DOUT_reg[6]  ( .D(n125), .CK(CLK), .RN(n1), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 \DOUT_reg[5]  ( .D(n126), .CK(CLK), .RN(n1), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 \DOUT_reg[4]  ( .D(n127), .CK(CLK), .RN(n1), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 \DOUT_reg[3]  ( .D(n128), .CK(CLK), .RN(n1), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 \DOUT_reg[2]  ( .D(n129), .CK(CLK), .RN(n1), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 \DOUT_reg[1]  ( .D(n130), .CK(CLK), .RN(n1), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 \DOUT_reg[0]  ( .D(n131), .CK(CLK), .RN(n1), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n1) );
  BUF_X1 U3 ( .A(RST), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n3) );
  INV_X1 U5 ( .A(n163), .ZN(n4) );
  MUX2_X1 U6 ( .A(n4), .B(DIN[0]), .S(EN), .Z(n131) );
  INV_X1 U7 ( .A(n162), .ZN(n5) );
  MUX2_X1 U8 ( .A(n5), .B(DIN[1]), .S(EN), .Z(n130) );
  INV_X1 U9 ( .A(n161), .ZN(n6) );
  MUX2_X1 U10 ( .A(n6), .B(DIN[2]), .S(EN), .Z(n129) );
  INV_X1 U11 ( .A(n160), .ZN(n7) );
  MUX2_X1 U12 ( .A(n7), .B(DIN[3]), .S(EN), .Z(n128) );
  INV_X1 U13 ( .A(n159), .ZN(n8) );
  MUX2_X1 U14 ( .A(n8), .B(DIN[4]), .S(EN), .Z(n127) );
  INV_X1 U15 ( .A(n158), .ZN(n9) );
  MUX2_X1 U16 ( .A(n9), .B(DIN[5]), .S(EN), .Z(n126) );
  INV_X1 U17 ( .A(n157), .ZN(n10) );
  MUX2_X1 U18 ( .A(n10), .B(DIN[6]), .S(EN), .Z(n125) );
  INV_X1 U19 ( .A(n156), .ZN(n11) );
  MUX2_X1 U20 ( .A(n11), .B(DIN[7]), .S(EN), .Z(n124) );
  INV_X1 U21 ( .A(n155), .ZN(n12) );
  MUX2_X1 U22 ( .A(n12), .B(DIN[8]), .S(EN), .Z(n123) );
  INV_X1 U23 ( .A(n154), .ZN(n13) );
  MUX2_X1 U24 ( .A(n13), .B(DIN[9]), .S(EN), .Z(n122) );
  INV_X1 U25 ( .A(n153), .ZN(n14) );
  MUX2_X1 U26 ( .A(n14), .B(DIN[10]), .S(EN), .Z(n121) );
  INV_X1 U27 ( .A(n152), .ZN(n15) );
  MUX2_X1 U28 ( .A(n15), .B(DIN[11]), .S(EN), .Z(n120) );
  INV_X1 U29 ( .A(n151), .ZN(n16) );
  MUX2_X1 U30 ( .A(n16), .B(DIN[12]), .S(EN), .Z(n119) );
  INV_X1 U31 ( .A(n150), .ZN(n17) );
  MUX2_X1 U32 ( .A(n17), .B(DIN[13]), .S(EN), .Z(n118) );
  INV_X1 U33 ( .A(n149), .ZN(n18) );
  MUX2_X1 U34 ( .A(n18), .B(DIN[14]), .S(EN), .Z(n117) );
  INV_X1 U35 ( .A(n148), .ZN(n19) );
  MUX2_X1 U36 ( .A(n19), .B(DIN[15]), .S(EN), .Z(n116) );
  INV_X1 U37 ( .A(n147), .ZN(n20) );
  MUX2_X1 U38 ( .A(n20), .B(DIN[16]), .S(EN), .Z(n115) );
  INV_X1 U39 ( .A(n146), .ZN(n21) );
  MUX2_X1 U40 ( .A(n21), .B(DIN[17]), .S(EN), .Z(n114) );
  INV_X1 U41 ( .A(n145), .ZN(n22) );
  MUX2_X1 U42 ( .A(n22), .B(DIN[18]), .S(EN), .Z(n113) );
  INV_X1 U43 ( .A(n144), .ZN(n23) );
  MUX2_X1 U44 ( .A(n23), .B(DIN[19]), .S(EN), .Z(n112) );
  INV_X1 U45 ( .A(n143), .ZN(n24) );
  MUX2_X1 U46 ( .A(n24), .B(DIN[20]), .S(EN), .Z(n111) );
  INV_X1 U47 ( .A(n142), .ZN(n25) );
  MUX2_X1 U48 ( .A(n25), .B(DIN[21]), .S(EN), .Z(n110) );
  INV_X1 U49 ( .A(n141), .ZN(n26) );
  MUX2_X1 U50 ( .A(n26), .B(DIN[22]), .S(EN), .Z(n109) );
  INV_X1 U51 ( .A(n140), .ZN(n27) );
  MUX2_X1 U52 ( .A(n27), .B(DIN[23]), .S(EN), .Z(n108) );
  INV_X1 U53 ( .A(n139), .ZN(n28) );
  MUX2_X1 U54 ( .A(n28), .B(DIN[24]), .S(EN), .Z(n107) );
  INV_X1 U55 ( .A(n138), .ZN(n29) );
  MUX2_X1 U56 ( .A(n29), .B(DIN[25]), .S(EN), .Z(n106) );
  INV_X1 U57 ( .A(n137), .ZN(n30) );
  MUX2_X1 U58 ( .A(n30), .B(DIN[26]), .S(EN), .Z(n105) );
  INV_X1 U59 ( .A(n136), .ZN(n31) );
  MUX2_X1 U60 ( .A(n31), .B(DIN[27]), .S(EN), .Z(n104) );
  INV_X1 U61 ( .A(n135), .ZN(n32) );
  MUX2_X1 U62 ( .A(n32), .B(DIN[28]), .S(EN), .Z(n103) );
  INV_X1 U63 ( .A(n134), .ZN(n97) );
  MUX2_X1 U64 ( .A(n97), .B(DIN[29]), .S(EN), .Z(n102) );
  INV_X1 U65 ( .A(n133), .ZN(n98) );
  MUX2_X1 U66 ( .A(n98), .B(DIN[30]), .S(EN), .Z(n101) );
  INV_X1 U67 ( .A(n132), .ZN(n99) );
  MUX2_X1 U68 ( .A(n99), .B(DIN[31]), .S(EN), .Z(n100) );
endmodule


module Execute_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \B[0] , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57;
  assign SUM[1] = B[1];
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR2_X1 U1 ( .A(B[31]), .B(n57), .ZN(SUM[31]) );
  NAND2_X1 U2 ( .A1(B[30]), .A2(n56), .ZN(n57) );
  INV_X1 U3 ( .A(B[2]), .ZN(SUM[2]) );
  XOR2_X1 U4 ( .A(B[3]), .B(B[2]), .Z(SUM[3]) );
  XOR2_X1 U5 ( .A(B[4]), .B(n30), .Z(SUM[4]) );
  XOR2_X1 U6 ( .A(B[5]), .B(n31), .Z(SUM[5]) );
  XOR2_X1 U7 ( .A(B[6]), .B(n32), .Z(SUM[6]) );
  XOR2_X1 U8 ( .A(B[7]), .B(n33), .Z(SUM[7]) );
  XOR2_X1 U9 ( .A(B[8]), .B(n34), .Z(SUM[8]) );
  XOR2_X1 U10 ( .A(B[9]), .B(n35), .Z(SUM[9]) );
  XOR2_X1 U11 ( .A(B[10]), .B(n36), .Z(SUM[10]) );
  XOR2_X1 U12 ( .A(B[11]), .B(n37), .Z(SUM[11]) );
  XOR2_X1 U13 ( .A(B[12]), .B(n38), .Z(SUM[12]) );
  XOR2_X1 U14 ( .A(B[13]), .B(n39), .Z(SUM[13]) );
  XOR2_X1 U15 ( .A(B[14]), .B(n40), .Z(SUM[14]) );
  XOR2_X1 U16 ( .A(B[15]), .B(n41), .Z(SUM[15]) );
  XOR2_X1 U17 ( .A(B[16]), .B(n42), .Z(SUM[16]) );
  XOR2_X1 U18 ( .A(B[17]), .B(n43), .Z(SUM[17]) );
  XOR2_X1 U19 ( .A(B[18]), .B(n44), .Z(SUM[18]) );
  XOR2_X1 U20 ( .A(B[19]), .B(n45), .Z(SUM[19]) );
  XOR2_X1 U21 ( .A(B[20]), .B(n46), .Z(SUM[20]) );
  XOR2_X1 U22 ( .A(B[21]), .B(n47), .Z(SUM[21]) );
  XOR2_X1 U23 ( .A(B[22]), .B(n48), .Z(SUM[22]) );
  XOR2_X1 U24 ( .A(B[23]), .B(n49), .Z(SUM[23]) );
  XOR2_X1 U25 ( .A(B[24]), .B(n50), .Z(SUM[24]) );
  XOR2_X1 U26 ( .A(B[25]), .B(n51), .Z(SUM[25]) );
  XOR2_X1 U27 ( .A(B[26]), .B(n52), .Z(SUM[26]) );
  XOR2_X1 U28 ( .A(B[27]), .B(n53), .Z(SUM[27]) );
  XOR2_X1 U29 ( .A(B[28]), .B(n54), .Z(SUM[28]) );
  XOR2_X1 U30 ( .A(B[29]), .B(n55), .Z(SUM[29]) );
  XOR2_X1 U31 ( .A(B[30]), .B(n56), .Z(SUM[30]) );
  AND2_X1 U32 ( .A1(B[3]), .A2(B[2]), .ZN(n30) );
  AND2_X1 U33 ( .A1(B[4]), .A2(n30), .ZN(n31) );
  AND2_X1 U34 ( .A1(B[5]), .A2(n31), .ZN(n32) );
  AND2_X1 U35 ( .A1(B[6]), .A2(n32), .ZN(n33) );
  AND2_X1 U36 ( .A1(B[7]), .A2(n33), .ZN(n34) );
  AND2_X1 U37 ( .A1(B[8]), .A2(n34), .ZN(n35) );
  AND2_X1 U38 ( .A1(B[9]), .A2(n35), .ZN(n36) );
  AND2_X1 U39 ( .A1(B[10]), .A2(n36), .ZN(n37) );
  AND2_X1 U40 ( .A1(B[11]), .A2(n37), .ZN(n38) );
  AND2_X1 U41 ( .A1(B[12]), .A2(n38), .ZN(n39) );
  AND2_X1 U42 ( .A1(B[13]), .A2(n39), .ZN(n40) );
  AND2_X1 U43 ( .A1(B[14]), .A2(n40), .ZN(n41) );
  AND2_X1 U44 ( .A1(B[15]), .A2(n41), .ZN(n42) );
  AND2_X1 U45 ( .A1(B[16]), .A2(n42), .ZN(n43) );
  AND2_X1 U46 ( .A1(B[17]), .A2(n43), .ZN(n44) );
  AND2_X1 U47 ( .A1(B[18]), .A2(n44), .ZN(n45) );
  AND2_X1 U48 ( .A1(B[19]), .A2(n45), .ZN(n46) );
  AND2_X1 U49 ( .A1(B[20]), .A2(n46), .ZN(n47) );
  AND2_X1 U50 ( .A1(B[21]), .A2(n47), .ZN(n48) );
  AND2_X1 U51 ( .A1(B[22]), .A2(n48), .ZN(n49) );
  AND2_X1 U52 ( .A1(B[23]), .A2(n49), .ZN(n50) );
  AND2_X1 U53 ( .A1(B[24]), .A2(n50), .ZN(n51) );
  AND2_X1 U54 ( .A1(B[25]), .A2(n51), .ZN(n52) );
  AND2_X1 U55 ( .A1(B[26]), .A2(n52), .ZN(n53) );
  AND2_X1 U56 ( .A1(B[27]), .A2(n53), .ZN(n54) );
  AND2_X1 U57 ( .A1(B[28]), .A2(n54), .ZN(n55) );
  AND2_X1 U58 ( .A1(B[29]), .A2(n55), .ZN(n56) );
endmodule


module Execute_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module Execute ( CLK, RST, MUX_A_SEL, MUX_B_SEL, .ALU_OPC({\ALU_OPC[3] , 
        \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), ALU_OUTREG_EN, JUMP_TYPE, 
        PC_IN, A_IN, B_IN, IMM_IN, ADD_WR_IN, ADD_RS1_IN, ADD_RS2_IN, 
        ADD_WR_MEM, ADD_WR_WB, RF_WE_MEM, RF_WE_WB, OP_MEM, OP_WB, PC_SEL, 
        ZERO_FLAG, NPC_ABS, NPC_REL, ALU_RES, B_OUT, ADD_WR_OUT );
  input [1:0] MUX_B_SEL;
  input [1:0] JUMP_TYPE;
  input [31:0] PC_IN;
  input [31:0] A_IN;
  input [31:0] B_IN;
  input [31:0] IMM_IN;
  input [4:0] ADD_WR_IN;
  input [4:0] ADD_RS1_IN;
  input [4:0] ADD_RS2_IN;
  input [4:0] ADD_WR_MEM;
  input [4:0] ADD_WR_WB;
  input [31:0] OP_MEM;
  input [31:0] OP_WB;
  output [1:0] PC_SEL;
  output [31:0] NPC_ABS;
  output [31:0] NPC_REL;
  output [31:0] ALU_RES;
  output [31:0] B_OUT;
  output [4:0] ADD_WR_OUT;
  input CLK, RST, MUX_A_SEL, \ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] ,
         \ALU_OPC[0] , ALU_OUTREG_EN, RF_WE_MEM, RF_WE_WB;
  output ZERO_FLAG;
  wire   sig_RST, sig_ZERO_FLAG, N9, N8, N7, N6, N5, N4, N31, N30, N3, N29,
         N28, N27, N26, N25, N24, N23, N22, N21, N20, N2, N19, N18, N17, N16,
         N15, N14, N13, N12, N11, N10, N1, N0, n1;
  wire   [3:0] ALU_OPC;
  wire   [31:0] sig_NPC_ABS;
  wire   [31:0] sig_NPC_REL;
  wire   [1:0] sig_PC_SEL;
  wire   [1:0] FWDA;
  wire   [1:0] FWDB;
  wire   [31:0] OP2_FW;
  wire   [31:0] sig_OP1;
  wire   [31:0] sig_OP2;
  wire   [31:0] sig_ALU_RES;

  Branch_Cond_Unit_NBIT32 Branch_Cond ( .RST(sig_RST), .A(sig_NPC_ABS), 
        .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), 
        .JUMP_TYPE(JUMP_TYPE), .PC_SEL(sig_PC_SEL), .ZERO(sig_ZERO_FLAG) );
  ff_1 ff0 ( .D(sig_ZERO_FLAG), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(ZERO_FLAG)
         );
  regn_N2 reg0 ( .DIN(sig_PC_SEL), .CLK(CLK), .EN(1'b1), .RST(RST), .DOUT(
        PC_SEL) );
  FWD_Unit FWD ( .RST(sig_RST), .ADD_RS1(ADD_RS1_IN), .ADD_RS2(ADD_RS2_IN), 
        .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_WB(ADD_WR_WB), .RF_WE_MEM(RF_WE_MEM), 
        .RF_WE_WB(RF_WE_WB), .FWDA(FWDA), .FWDB(FWDB) );
  mux41_NBIT32_0 FW1 ( .A(A_IN), .B(OP_WB), .C(OP_MEM), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(FWDA), .Z(sig_NPC_ABS) );
  mux41_NBIT32_4 FW2 ( .A(B_IN), .B(OP_WB), .C(OP_MEM), .D({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(FWDB), .Z(OP2_FW) );
  mux21_NBIT32_3 muxA ( .A(sig_NPC_ABS), .B(PC_IN), .S(MUX_A_SEL), .Z(sig_OP1)
         );
  mux41_NBIT32_3 muxB ( .A(OP2_FW), .B(IMM_IN), .C({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(MUX_B_SEL), .Z(sig_OP2) );
  ALU_NBIT32 alu0 ( .OP1(sig_OP1), .OP2(sig_OP2), .ALU_OPC({\ALU_OPC[3] , 
        \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), .ALU_RES(sig_ALU_RES) );
  regn_N32_6 alureg ( .DIN(sig_ALU_RES), .CLK(CLK), .EN(ALU_OUTREG_EN), .RST(
        RST), .DOUT(ALU_RES) );
  regn_N32_5 B_reg ( .DIN(OP2_FW), .CLK(CLK), .EN(ALU_OUTREG_EN), .RST(RST), 
        .DOUT(B_OUT) );
  regn_N5_2 ADD_WR_reg ( .DIN(ADD_WR_IN), .CLK(CLK), .EN(ALU_OUTREG_EN), .RST(
        RST), .DOUT(ADD_WR_OUT) );
  regn_N32_4 NPC_ABS_reg ( .DIN(sig_NPC_ABS), .CLK(CLK), .EN(ALU_OUTREG_EN), 
        .RST(RST), .DOUT(NPC_ABS) );
  regn_N32_3 NPC_REL_reg ( .DIN(sig_NPC_REL), .CLK(CLK), .EN(ALU_OUTREG_EN), 
        .RST(RST), .DOUT(NPC_REL) );
  Execute_DW01_add_1 add_1_root_add_0_root_add_118_2 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .B(IMM_IN), .CI(1'b0), .SUM({N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0})
         );
  Execute_DW01_add_0 add_0_root_add_0_root_add_118_2 ( .A(PC_IN), .B({N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}), 
        .CI(1'b0), .SUM(sig_NPC_REL) );
  NOR2_X1 U3 ( .A1(ZERO_FLAG), .A2(n1), .ZN(sig_RST) );
  INV_X1 U4 ( .A(RST), .ZN(n1) );
endmodule


module ff_0 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n2, n3;

  DFFR_X1 Q_reg ( .D(n3), .CK(CLK), .RN(RST), .Q(Q), .QN(n2) );
  OAI21_X1 U2 ( .B1(n2), .B2(EN), .A(n1), .ZN(n3) );
  NAND2_X1 U3 ( .A1(EN), .A2(D), .ZN(n1) );
endmodule


module regn_N32_2 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n68, n69, n70;

  DFFR_X1 \DOUT_reg[31]  ( .D(n36), .CK(CLK), .RN(n3), .Q(DOUT[31]) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n37), .CK(CLK), .RN(n3), .Q(DOUT[30]) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n38), .CK(CLK), .RN(n3), .Q(DOUT[29]) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n39), .CK(CLK), .RN(n3), .Q(DOUT[28]) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n40), .CK(CLK), .RN(n3), .Q(DOUT[27]) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n41), .CK(CLK), .RN(n3), .Q(DOUT[26]) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n42), .CK(CLK), .RN(n3), .Q(DOUT[25]) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n43), .CK(CLK), .RN(n3), .Q(DOUT[24]) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n44), .CK(CLK), .RN(n2), .Q(DOUT[23]) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n45), .CK(CLK), .RN(n2), .Q(DOUT[22]) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n46), .CK(CLK), .RN(n2), .Q(DOUT[21]) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n47), .CK(CLK), .RN(n2), .Q(DOUT[20]) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n48), .CK(CLK), .RN(n2), .Q(DOUT[19]) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n49), .CK(CLK), .RN(n2), .Q(DOUT[18]) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n50), .CK(CLK), .RN(n2), .Q(DOUT[17]) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n51), .CK(CLK), .RN(n2), .Q(DOUT[16]) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n52), .CK(CLK), .RN(n2), .Q(DOUT[15]) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n53), .CK(CLK), .RN(n2), .Q(DOUT[14]) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n54), .CK(CLK), .RN(n2), .Q(DOUT[13]) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n55), .CK(CLK), .RN(n2), .Q(DOUT[12]) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n56), .CK(CLK), .RN(n1), .Q(DOUT[11]) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n57), .CK(CLK), .RN(n1), .Q(DOUT[10]) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n58), .CK(CLK), .RN(n1), .Q(DOUT[9]) );
  DFFR_X1 \DOUT_reg[8]  ( .D(n59), .CK(CLK), .RN(n1), .Q(DOUT[8]) );
  DFFR_X1 \DOUT_reg[7]  ( .D(n60), .CK(CLK), .RN(n1), .Q(DOUT[7]) );
  DFFR_X1 \DOUT_reg[6]  ( .D(n61), .CK(CLK), .RN(n1), .Q(DOUT[6]) );
  DFFR_X1 \DOUT_reg[5]  ( .D(n62), .CK(CLK), .RN(n1), .Q(DOUT[5]) );
  DFFR_X1 \DOUT_reg[4]  ( .D(n63), .CK(CLK), .RN(n1), .Q(DOUT[4]) );
  DFFR_X1 \DOUT_reg[3]  ( .D(n64), .CK(CLK), .RN(n1), .Q(DOUT[3]) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n68), .CK(CLK), .RN(n1), .Q(DOUT[2]) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n69), .CK(CLK), .RN(n1), .Q(DOUT[1]) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n70), .CK(CLK), .RN(n1), .Q(DOUT[0]) );
  BUF_X1 U2 ( .A(RST), .Z(n1) );
  BUF_X1 U3 ( .A(RST), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n3) );
  MUX2_X1 U5 ( .A(DOUT[0]), .B(DIN[0]), .S(EN), .Z(n70) );
  MUX2_X1 U6 ( .A(DOUT[1]), .B(DIN[1]), .S(EN), .Z(n69) );
  MUX2_X1 U7 ( .A(DOUT[2]), .B(DIN[2]), .S(EN), .Z(n68) );
  MUX2_X1 U8 ( .A(DOUT[3]), .B(DIN[3]), .S(EN), .Z(n64) );
  MUX2_X1 U9 ( .A(DOUT[4]), .B(DIN[4]), .S(EN), .Z(n63) );
  MUX2_X1 U10 ( .A(DOUT[5]), .B(DIN[5]), .S(EN), .Z(n62) );
  MUX2_X1 U11 ( .A(DOUT[6]), .B(DIN[6]), .S(EN), .Z(n61) );
  MUX2_X1 U12 ( .A(DOUT[7]), .B(DIN[7]), .S(EN), .Z(n60) );
  MUX2_X1 U13 ( .A(DOUT[8]), .B(DIN[8]), .S(EN), .Z(n59) );
  MUX2_X1 U14 ( .A(DOUT[9]), .B(DIN[9]), .S(EN), .Z(n58) );
  MUX2_X1 U15 ( .A(DOUT[10]), .B(DIN[10]), .S(EN), .Z(n57) );
  MUX2_X1 U16 ( .A(DOUT[11]), .B(DIN[11]), .S(EN), .Z(n56) );
  MUX2_X1 U17 ( .A(DOUT[12]), .B(DIN[12]), .S(EN), .Z(n55) );
  MUX2_X1 U18 ( .A(DOUT[13]), .B(DIN[13]), .S(EN), .Z(n54) );
  MUX2_X1 U19 ( .A(DOUT[14]), .B(DIN[14]), .S(EN), .Z(n53) );
  MUX2_X1 U20 ( .A(DOUT[15]), .B(DIN[15]), .S(EN), .Z(n52) );
  MUX2_X1 U21 ( .A(DOUT[16]), .B(DIN[16]), .S(EN), .Z(n51) );
  MUX2_X1 U22 ( .A(DOUT[17]), .B(DIN[17]), .S(EN), .Z(n50) );
  MUX2_X1 U23 ( .A(DOUT[18]), .B(DIN[18]), .S(EN), .Z(n49) );
  MUX2_X1 U24 ( .A(DOUT[19]), .B(DIN[19]), .S(EN), .Z(n48) );
  MUX2_X1 U25 ( .A(DOUT[20]), .B(DIN[20]), .S(EN), .Z(n47) );
  MUX2_X1 U26 ( .A(DOUT[21]), .B(DIN[21]), .S(EN), .Z(n46) );
  MUX2_X1 U27 ( .A(DOUT[22]), .B(DIN[22]), .S(EN), .Z(n45) );
  MUX2_X1 U28 ( .A(DOUT[23]), .B(DIN[23]), .S(EN), .Z(n44) );
  MUX2_X1 U29 ( .A(DOUT[24]), .B(DIN[24]), .S(EN), .Z(n43) );
  MUX2_X1 U30 ( .A(DOUT[25]), .B(DIN[25]), .S(EN), .Z(n42) );
  MUX2_X1 U31 ( .A(DOUT[26]), .B(DIN[26]), .S(EN), .Z(n41) );
  MUX2_X1 U32 ( .A(DOUT[27]), .B(DIN[27]), .S(EN), .Z(n40) );
  MUX2_X1 U33 ( .A(DOUT[28]), .B(DIN[28]), .S(EN), .Z(n39) );
  MUX2_X1 U34 ( .A(DOUT[29]), .B(DIN[29]), .S(EN), .Z(n38) );
  MUX2_X1 U35 ( .A(DOUT[30]), .B(DIN[30]), .S(EN), .Z(n37) );
  MUX2_X1 U36 ( .A(DOUT[31]), .B(DIN[31]), .S(EN), .Z(n36) );
endmodule


module regn_N5_1 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n6, n7, n8, n9, n10;

  DFFR_X1 \DOUT_reg[4]  ( .D(n6), .CK(CLK), .RN(RST), .Q(DOUT[4]) );
  DFFR_X1 \DOUT_reg[3]  ( .D(n7), .CK(CLK), .RN(RST), .Q(DOUT[3]) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n8), .CK(CLK), .RN(RST), .Q(DOUT[2]) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n9), .CK(CLK), .RN(RST), .Q(DOUT[1]) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n10), .CK(CLK), .RN(RST), .Q(DOUT[0]) );
  MUX2_X1 U2 ( .A(DOUT[0]), .B(DIN[0]), .S(EN), .Z(n10) );
  MUX2_X1 U3 ( .A(DOUT[1]), .B(DIN[1]), .S(EN), .Z(n9) );
  MUX2_X1 U4 ( .A(DOUT[2]), .B(DIN[2]), .S(EN), .Z(n8) );
  MUX2_X1 U5 ( .A(DOUT[3]), .B(DIN[3]), .S(EN), .Z(n7) );
  MUX2_X1 U6 ( .A(DOUT[4]), .B(DIN[4]), .S(EN), .Z(n6) );
endmodule


module regn_N32_1 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n68, n69, n70;

  DFFR_X1 \DOUT_reg[31]  ( .D(n36), .CK(CLK), .RN(n3), .Q(DOUT[31]) );
  DFFR_X1 \DOUT_reg[30]  ( .D(n37), .CK(CLK), .RN(n3), .Q(DOUT[30]) );
  DFFR_X1 \DOUT_reg[29]  ( .D(n38), .CK(CLK), .RN(n3), .Q(DOUT[29]) );
  DFFR_X1 \DOUT_reg[28]  ( .D(n39), .CK(CLK), .RN(n3), .Q(DOUT[28]) );
  DFFR_X1 \DOUT_reg[27]  ( .D(n40), .CK(CLK), .RN(n3), .Q(DOUT[27]) );
  DFFR_X1 \DOUT_reg[26]  ( .D(n41), .CK(CLK), .RN(n3), .Q(DOUT[26]) );
  DFFR_X1 \DOUT_reg[25]  ( .D(n42), .CK(CLK), .RN(n3), .Q(DOUT[25]) );
  DFFR_X1 \DOUT_reg[24]  ( .D(n43), .CK(CLK), .RN(n3), .Q(DOUT[24]) );
  DFFR_X1 \DOUT_reg[23]  ( .D(n44), .CK(CLK), .RN(n2), .Q(DOUT[23]) );
  DFFR_X1 \DOUT_reg[22]  ( .D(n45), .CK(CLK), .RN(n2), .Q(DOUT[22]) );
  DFFR_X1 \DOUT_reg[21]  ( .D(n46), .CK(CLK), .RN(n2), .Q(DOUT[21]) );
  DFFR_X1 \DOUT_reg[20]  ( .D(n47), .CK(CLK), .RN(n2), .Q(DOUT[20]) );
  DFFR_X1 \DOUT_reg[19]  ( .D(n48), .CK(CLK), .RN(n2), .Q(DOUT[19]) );
  DFFR_X1 \DOUT_reg[18]  ( .D(n49), .CK(CLK), .RN(n2), .Q(DOUT[18]) );
  DFFR_X1 \DOUT_reg[17]  ( .D(n50), .CK(CLK), .RN(n2), .Q(DOUT[17]) );
  DFFR_X1 \DOUT_reg[16]  ( .D(n51), .CK(CLK), .RN(n2), .Q(DOUT[16]) );
  DFFR_X1 \DOUT_reg[15]  ( .D(n52), .CK(CLK), .RN(n2), .Q(DOUT[15]) );
  DFFR_X1 \DOUT_reg[14]  ( .D(n53), .CK(CLK), .RN(n2), .Q(DOUT[14]) );
  DFFR_X1 \DOUT_reg[13]  ( .D(n54), .CK(CLK), .RN(n2), .Q(DOUT[13]) );
  DFFR_X1 \DOUT_reg[12]  ( .D(n55), .CK(CLK), .RN(n2), .Q(DOUT[12]) );
  DFFR_X1 \DOUT_reg[11]  ( .D(n56), .CK(CLK), .RN(n1), .Q(DOUT[11]) );
  DFFR_X1 \DOUT_reg[10]  ( .D(n57), .CK(CLK), .RN(n1), .Q(DOUT[10]) );
  DFFR_X1 \DOUT_reg[9]  ( .D(n58), .CK(CLK), .RN(n1), .Q(DOUT[9]) );
  DFFR_X1 \DOUT_reg[8]  ( .D(n59), .CK(CLK), .RN(n1), .Q(DOUT[8]) );
  DFFR_X1 \DOUT_reg[7]  ( .D(n60), .CK(CLK), .RN(n1), .Q(DOUT[7]) );
  DFFR_X1 \DOUT_reg[6]  ( .D(n61), .CK(CLK), .RN(n1), .Q(DOUT[6]) );
  DFFR_X1 \DOUT_reg[5]  ( .D(n62), .CK(CLK), .RN(n1), .Q(DOUT[5]) );
  DFFR_X1 \DOUT_reg[4]  ( .D(n63), .CK(CLK), .RN(n1), .Q(DOUT[4]) );
  DFFR_X1 \DOUT_reg[3]  ( .D(n64), .CK(CLK), .RN(n1), .Q(DOUT[3]) );
  DFFR_X1 \DOUT_reg[2]  ( .D(n68), .CK(CLK), .RN(n1), .Q(DOUT[2]) );
  DFFR_X1 \DOUT_reg[1]  ( .D(n69), .CK(CLK), .RN(n1), .Q(DOUT[1]) );
  DFFR_X1 \DOUT_reg[0]  ( .D(n70), .CK(CLK), .RN(n1), .Q(DOUT[0]) );
  BUF_X1 U2 ( .A(RST), .Z(n1) );
  BUF_X1 U3 ( .A(RST), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n3) );
  MUX2_X1 U5 ( .A(DOUT[0]), .B(DIN[0]), .S(EN), .Z(n70) );
  MUX2_X1 U6 ( .A(DOUT[1]), .B(DIN[1]), .S(EN), .Z(n69) );
  MUX2_X1 U7 ( .A(DOUT[2]), .B(DIN[2]), .S(EN), .Z(n68) );
  MUX2_X1 U8 ( .A(DOUT[3]), .B(DIN[3]), .S(EN), .Z(n64) );
  MUX2_X1 U9 ( .A(DOUT[4]), .B(DIN[4]), .S(EN), .Z(n63) );
  MUX2_X1 U10 ( .A(DOUT[5]), .B(DIN[5]), .S(EN), .Z(n62) );
  MUX2_X1 U11 ( .A(DOUT[6]), .B(DIN[6]), .S(EN), .Z(n61) );
  MUX2_X1 U12 ( .A(DOUT[7]), .B(DIN[7]), .S(EN), .Z(n60) );
  MUX2_X1 U13 ( .A(DOUT[8]), .B(DIN[8]), .S(EN), .Z(n59) );
  MUX2_X1 U14 ( .A(DOUT[9]), .B(DIN[9]), .S(EN), .Z(n58) );
  MUX2_X1 U15 ( .A(DOUT[10]), .B(DIN[10]), .S(EN), .Z(n57) );
  MUX2_X1 U16 ( .A(DOUT[11]), .B(DIN[11]), .S(EN), .Z(n56) );
  MUX2_X1 U17 ( .A(DOUT[12]), .B(DIN[12]), .S(EN), .Z(n55) );
  MUX2_X1 U18 ( .A(DOUT[13]), .B(DIN[13]), .S(EN), .Z(n54) );
  MUX2_X1 U19 ( .A(DOUT[14]), .B(DIN[14]), .S(EN), .Z(n53) );
  MUX2_X1 U20 ( .A(DOUT[15]), .B(DIN[15]), .S(EN), .Z(n52) );
  MUX2_X1 U21 ( .A(DOUT[16]), .B(DIN[16]), .S(EN), .Z(n51) );
  MUX2_X1 U22 ( .A(DOUT[17]), .B(DIN[17]), .S(EN), .Z(n50) );
  MUX2_X1 U23 ( .A(DOUT[18]), .B(DIN[18]), .S(EN), .Z(n49) );
  MUX2_X1 U24 ( .A(DOUT[19]), .B(DIN[19]), .S(EN), .Z(n48) );
  MUX2_X1 U25 ( .A(DOUT[20]), .B(DIN[20]), .S(EN), .Z(n47) );
  MUX2_X1 U26 ( .A(DOUT[21]), .B(DIN[21]), .S(EN), .Z(n46) );
  MUX2_X1 U27 ( .A(DOUT[22]), .B(DIN[22]), .S(EN), .Z(n45) );
  MUX2_X1 U28 ( .A(DOUT[23]), .B(DIN[23]), .S(EN), .Z(n44) );
  MUX2_X1 U29 ( .A(DOUT[24]), .B(DIN[24]), .S(EN), .Z(n43) );
  MUX2_X1 U30 ( .A(DOUT[25]), .B(DIN[25]), .S(EN), .Z(n42) );
  MUX2_X1 U31 ( .A(DOUT[26]), .B(DIN[26]), .S(EN), .Z(n41) );
  MUX2_X1 U32 ( .A(DOUT[27]), .B(DIN[27]), .S(EN), .Z(n40) );
  MUX2_X1 U33 ( .A(DOUT[28]), .B(DIN[28]), .S(EN), .Z(n39) );
  MUX2_X1 U34 ( .A(DOUT[29]), .B(DIN[29]), .S(EN), .Z(n38) );
  MUX2_X1 U35 ( .A(DOUT[30]), .B(DIN[30]), .S(EN), .Z(n37) );
  MUX2_X1 U36 ( .A(DOUT[31]), .B(DIN[31]), .S(EN), .Z(n36) );
endmodule


module mux41_NBIT32_2 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103;

  BUF_X1 U1 ( .A(S[1]), .Z(n1) );
  BUF_X1 U2 ( .A(n30), .Z(n2) );
  BUF_X1 U3 ( .A(n30), .Z(n3) );
  BUF_X2 U4 ( .A(n28), .Z(n4) );
  BUF_X2 U5 ( .A(n28), .Z(n5) );
  BUF_X1 U6 ( .A(n30), .Z(n38) );
  BUF_X1 U7 ( .A(n30), .Z(n6) );
  BUF_X1 U8 ( .A(n30), .Z(n40) );
  BUF_X1 U9 ( .A(n30), .Z(n7) );
  AND2_X2 U10 ( .A1(n44), .A2(n45), .ZN(n28) );
  AND2_X2 U11 ( .A1(S[0]), .A2(n45), .ZN(n30) );
  AND2_X1 U12 ( .A1(n99), .A2(n26), .ZN(n8) );
  OAI221_X1 U13 ( .B1(n9), .B2(n10), .C1(n11), .C2(n12), .A(n72), .ZN(Z[14])
         );
  INV_X1 U14 ( .A(A[14]), .ZN(n9) );
  INV_X1 U15 ( .A(n28), .ZN(n10) );
  INV_X1 U16 ( .A(B[14]), .ZN(n11) );
  INV_X1 U17 ( .A(n30), .ZN(n12) );
  OAI211_X1 U18 ( .C1(n13), .C2(n15), .A(n27), .B(n101), .ZN(Z[30]) );
  INV_X1 U19 ( .A(A[30]), .ZN(n13) );
  AOI22_X1 U20 ( .A1(A[15]), .A2(n28), .B1(B[15]), .B2(n40), .ZN(n73) );
  OAI221_X1 U21 ( .B1(n14), .B2(n15), .C1(n16), .C2(n17), .A(n100), .ZN(Z[29])
         );
  INV_X1 U22 ( .A(A[29]), .ZN(n14) );
  INV_X1 U23 ( .A(n28), .ZN(n15) );
  INV_X1 U24 ( .A(B[29]), .ZN(n16) );
  INV_X1 U25 ( .A(n30), .ZN(n17) );
  OAI221_X1 U26 ( .B1(n18), .B2(n19), .C1(n20), .C2(n21), .A(n64), .ZN(Z[9])
         );
  INV_X1 U27 ( .A(A[9]), .ZN(n18) );
  INV_X1 U28 ( .A(n28), .ZN(n19) );
  INV_X1 U29 ( .A(B[9]), .ZN(n20) );
  INV_X1 U30 ( .A(n30), .ZN(n21) );
  OAI221_X1 U31 ( .B1(n22), .B2(n23), .C1(n24), .C2(n17), .A(n71), .ZN(Z[13])
         );
  INV_X1 U32 ( .A(A[13]), .ZN(n22) );
  INV_X1 U33 ( .A(n28), .ZN(n23) );
  INV_X1 U34 ( .A(B[13]), .ZN(n24) );
  NAND2_X1 U35 ( .A1(A[28]), .A2(n36), .ZN(n25) );
  NAND2_X1 U36 ( .A1(B[28]), .A2(n38), .ZN(n26) );
  BUF_X2 U37 ( .A(n28), .Z(n35) );
  NAND2_X1 U38 ( .A1(B[30]), .A2(n40), .ZN(n27) );
  BUF_X2 U39 ( .A(n29), .Z(n33) );
  BUF_X2 U40 ( .A(n29), .Z(n34) );
  BUF_X1 U41 ( .A(n28), .Z(n36) );
  BUF_X1 U42 ( .A(n28), .Z(n37) );
  BUF_X1 U43 ( .A(n29), .Z(n32) );
  BUF_X1 U44 ( .A(n30), .Z(n39) );
  BUF_X1 U45 ( .A(n31), .Z(n41) );
  BUF_X1 U46 ( .A(n31), .Z(n42) );
  BUF_X1 U47 ( .A(n31), .Z(n43) );
  AND2_X1 U48 ( .A1(n44), .A2(n1), .ZN(n29) );
  AND2_X1 U49 ( .A1(S[0]), .A2(n1), .ZN(n31) );
  INV_X1 U50 ( .A(S[0]), .ZN(n44) );
  AOI22_X1 U51 ( .A1(C[0]), .A2(n33), .B1(D[0]), .B2(n42), .ZN(n47) );
  INV_X1 U52 ( .A(S[1]), .ZN(n45) );
  AOI22_X1 U53 ( .A1(A[0]), .A2(n36), .B1(B[0]), .B2(n39), .ZN(n46) );
  NAND2_X1 U54 ( .A1(n46), .A2(n47), .ZN(Z[0]) );
  AOI22_X1 U55 ( .A1(C[1]), .A2(n34), .B1(D[1]), .B2(n41), .ZN(n49) );
  AOI22_X1 U56 ( .A1(A[1]), .A2(n35), .B1(B[1]), .B2(n2), .ZN(n48) );
  NAND2_X1 U57 ( .A1(n48), .A2(n49), .ZN(Z[1]) );
  AOI22_X1 U58 ( .A1(C[2]), .A2(n34), .B1(D[2]), .B2(n43), .ZN(n51) );
  AOI22_X1 U59 ( .A1(A[2]), .A2(n35), .B1(n6), .B2(B[2]), .ZN(n50) );
  NAND2_X1 U60 ( .A1(n50), .A2(n51), .ZN(Z[2]) );
  AOI22_X1 U61 ( .A1(C[3]), .A2(n34), .B1(D[3]), .B2(n43), .ZN(n53) );
  AOI22_X1 U62 ( .A1(A[3]), .A2(n35), .B1(n7), .B2(B[3]), .ZN(n52) );
  NAND2_X1 U63 ( .A1(n52), .A2(n53), .ZN(Z[3]) );
  AOI22_X1 U64 ( .A1(C[4]), .A2(n34), .B1(D[4]), .B2(n43), .ZN(n55) );
  AOI22_X1 U65 ( .A1(A[4]), .A2(n35), .B1(n30), .B2(B[4]), .ZN(n54) );
  NAND2_X1 U66 ( .A1(n54), .A2(n55), .ZN(Z[4]) );
  AOI22_X1 U67 ( .A1(C[5]), .A2(n33), .B1(D[5]), .B2(n43), .ZN(n57) );
  AOI22_X1 U68 ( .A1(A[5]), .A2(n35), .B1(B[5]), .B2(n6), .ZN(n56) );
  NAND2_X1 U69 ( .A1(n56), .A2(n57), .ZN(Z[5]) );
  AOI22_X1 U70 ( .A1(C[6]), .A2(n33), .B1(D[6]), .B2(n43), .ZN(n59) );
  AOI22_X1 U71 ( .A1(A[6]), .A2(n4), .B1(B[6]), .B2(n3), .ZN(n58) );
  NAND2_X1 U72 ( .A1(n58), .A2(n59), .ZN(Z[6]) );
  AOI22_X1 U73 ( .A1(C[7]), .A2(n33), .B1(D[7]), .B2(n43), .ZN(n61) );
  AOI22_X1 U74 ( .A1(A[7]), .A2(n36), .B1(B[7]), .B2(n3), .ZN(n60) );
  NAND2_X1 U75 ( .A1(n60), .A2(n61), .ZN(Z[7]) );
  AOI22_X1 U76 ( .A1(C[8]), .A2(n33), .B1(D[8]), .B2(n42), .ZN(n63) );
  AOI22_X1 U77 ( .A1(A[8]), .A2(n37), .B1(B[8]), .B2(n40), .ZN(n62) );
  NAND2_X1 U78 ( .A1(n62), .A2(n63), .ZN(Z[8]) );
  AOI22_X1 U79 ( .A1(C[9]), .A2(n33), .B1(D[9]), .B2(n43), .ZN(n64) );
  AOI22_X1 U80 ( .A1(C[10]), .A2(n33), .B1(D[10]), .B2(n42), .ZN(n66) );
  AOI22_X1 U81 ( .A1(A[10]), .A2(n5), .B1(B[10]), .B2(n7), .ZN(n65) );
  NAND2_X1 U82 ( .A1(n65), .A2(n66), .ZN(Z[10]) );
  AOI22_X1 U83 ( .A1(C[11]), .A2(n33), .B1(D[11]), .B2(n42), .ZN(n68) );
  AOI22_X1 U84 ( .A1(A[11]), .A2(n5), .B1(B[11]), .B2(n2), .ZN(n67) );
  NAND2_X1 U85 ( .A1(n67), .A2(n68), .ZN(Z[11]) );
  AOI22_X1 U86 ( .A1(C[12]), .A2(n33), .B1(D[12]), .B2(n42), .ZN(n70) );
  AOI22_X1 U87 ( .A1(A[12]), .A2(n5), .B1(B[12]), .B2(n38), .ZN(n69) );
  NAND2_X1 U88 ( .A1(n69), .A2(n70), .ZN(Z[12]) );
  AOI22_X1 U89 ( .A1(C[13]), .A2(n33), .B1(D[13]), .B2(n42), .ZN(n71) );
  AOI22_X1 U90 ( .A1(C[14]), .A2(n33), .B1(D[14]), .B2(n42), .ZN(n72) );
  AOI22_X1 U91 ( .A1(C[15]), .A2(n33), .B1(D[15]), .B2(n42), .ZN(n74) );
  NAND2_X1 U92 ( .A1(n73), .A2(n74), .ZN(Z[15]) );
  AOI22_X1 U93 ( .A1(C[16]), .A2(n32), .B1(D[16]), .B2(n42), .ZN(n76) );
  AOI22_X1 U94 ( .A1(A[16]), .A2(n37), .B1(B[16]), .B2(n38), .ZN(n75) );
  NAND2_X1 U95 ( .A1(n75), .A2(n76), .ZN(Z[16]) );
  AOI22_X1 U96 ( .A1(C[17]), .A2(n32), .B1(D[17]), .B2(n42), .ZN(n78) );
  AOI22_X1 U97 ( .A1(A[17]), .A2(n4), .B1(B[17]), .B2(n7), .ZN(n77) );
  NAND2_X1 U98 ( .A1(n77), .A2(n78), .ZN(Z[17]) );
  AOI22_X1 U99 ( .A1(C[18]), .A2(n32), .B1(D[18]), .B2(n42), .ZN(n80) );
  AOI22_X1 U100 ( .A1(A[18]), .A2(n5), .B1(B[18]), .B2(n3), .ZN(n79) );
  NAND2_X1 U101 ( .A1(n79), .A2(n80), .ZN(Z[18]) );
  AOI22_X1 U102 ( .A1(A[19]), .A2(n37), .B1(C[19]), .B2(n34), .ZN(n82) );
  AOI22_X1 U103 ( .A1(D[19]), .A2(n41), .B1(B[19]), .B2(n40), .ZN(n81) );
  NAND2_X1 U104 ( .A1(n82), .A2(n81), .ZN(Z[19]) );
  AOI22_X1 U105 ( .A1(C[20]), .A2(n32), .B1(D[20]), .B2(n42), .ZN(n84) );
  AOI22_X1 U106 ( .A1(A[20]), .A2(n36), .B1(B[20]), .B2(n2), .ZN(n83) );
  NAND2_X1 U107 ( .A1(n83), .A2(n84), .ZN(Z[20]) );
  AOI22_X1 U108 ( .A1(C[21]), .A2(n32), .B1(D[21]), .B2(n41), .ZN(n86) );
  AOI22_X1 U109 ( .A1(A[21]), .A2(n4), .B1(B[21]), .B2(n6), .ZN(n85) );
  NAND2_X1 U110 ( .A1(n85), .A2(n86), .ZN(Z[21]) );
  AOI22_X1 U111 ( .A1(C[22]), .A2(n32), .B1(D[22]), .B2(n41), .ZN(n88) );
  AOI22_X1 U112 ( .A1(A[22]), .A2(n4), .B1(B[22]), .B2(n38), .ZN(n87) );
  NAND2_X1 U113 ( .A1(n87), .A2(n88), .ZN(Z[22]) );
  NAND2_X1 U114 ( .A1(A[23]), .A2(n5), .ZN(n90) );
  AOI222_X1 U115 ( .A1(B[23]), .A2(n3), .B1(C[23]), .B2(n34), .C1(D[23]), .C2(
        n43), .ZN(n89) );
  NAND2_X1 U116 ( .A1(n90), .A2(n89), .ZN(Z[23]) );
  AOI22_X1 U117 ( .A1(C[24]), .A2(n32), .B1(D[24]), .B2(n41), .ZN(n92) );
  AOI22_X1 U118 ( .A1(A[24]), .A2(n36), .B1(B[24]), .B2(n39), .ZN(n91) );
  NAND2_X1 U119 ( .A1(n91), .A2(n92), .ZN(Z[24]) );
  AOI22_X1 U120 ( .A1(C[25]), .A2(n32), .B1(D[25]), .B2(n41), .ZN(n94) );
  AOI22_X1 U121 ( .A1(A[25]), .A2(n37), .B1(B[25]), .B2(n6), .ZN(n93) );
  NAND2_X1 U122 ( .A1(n93), .A2(n94), .ZN(Z[25]) );
  AOI22_X1 U123 ( .A1(C[26]), .A2(n32), .B1(D[26]), .B2(n41), .ZN(n96) );
  AOI22_X1 U124 ( .A1(A[26]), .A2(n37), .B1(B[26]), .B2(n39), .ZN(n95) );
  NAND2_X1 U125 ( .A1(n95), .A2(n96), .ZN(Z[26]) );
  AOI22_X1 U126 ( .A1(A[27]), .A2(n5), .B1(C[27]), .B2(n34), .ZN(n98) );
  AOI22_X1 U127 ( .A1(D[27]), .A2(n41), .B1(B[27]), .B2(n39), .ZN(n97) );
  NAND2_X1 U128 ( .A1(n98), .A2(n97), .ZN(Z[27]) );
  AOI22_X1 U129 ( .A1(C[28]), .A2(n32), .B1(D[28]), .B2(n41), .ZN(n99) );
  NAND2_X1 U130 ( .A1(n25), .A2(n8), .ZN(Z[28]) );
  AOI22_X1 U131 ( .A1(C[29]), .A2(n32), .B1(D[29]), .B2(n41), .ZN(n100) );
  AOI22_X1 U132 ( .A1(C[30]), .A2(n32), .B1(D[30]), .B2(n41), .ZN(n101) );
  AOI22_X1 U133 ( .A1(A[31]), .A2(n4), .B1(C[31]), .B2(n34), .ZN(n103) );
  AOI22_X1 U134 ( .A1(D[31]), .A2(n41), .B1(B[31]), .B2(n7), .ZN(n102) );
  NAND2_X1 U135 ( .A1(n103), .A2(n102), .ZN(Z[31]) );
endmodule


module Memory ( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, DRAM_EN_IN, PC_SEL, 
        NPC_IN, NPC_ABS, NPC_REL, ALU_RES_IN, B_IN, ADD_WR_IN, DRAM_DATA_IN, 
        PC_OUT, DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, DRAM_ADDR_OUT, 
        DRAM_DATA_OUT, DATA_OUT, ALU_RES_OUT, OP_MEM, ADD_WR_MEM, ADD_WR_OUT
 );
  input [1:0] PC_SEL;
  input [31:0] NPC_IN;
  input [31:0] NPC_ABS;
  input [31:0] NPC_REL;
  input [31:0] ALU_RES_IN;
  input [31:0] B_IN;
  input [4:0] ADD_WR_IN;
  input [31:0] DRAM_DATA_IN;
  output [31:0] PC_OUT;
  output [31:0] DRAM_ADDR_OUT;
  output [31:0] DRAM_DATA_OUT;
  output [31:0] DATA_OUT;
  output [31:0] ALU_RES_OUT;
  output [31:0] OP_MEM;
  output [4:0] ADD_WR_MEM;
  output [4:0] ADD_WR_OUT;
  input CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, DRAM_EN_IN;
  output DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT;
  wire   DRAM_EN_IN, DRAM_R_IN, DRAM_W_IN;
  assign DRAM_EN_OUT = DRAM_EN_IN;
  assign DRAM_R_OUT = DRAM_R_IN;
  assign DRAM_W_OUT = DRAM_W_IN;
  assign OP_MEM[31] = ALU_RES_IN[31];
  assign DRAM_ADDR_OUT[31] = ALU_RES_IN[31];
  assign OP_MEM[30] = ALU_RES_IN[30];
  assign DRAM_ADDR_OUT[30] = ALU_RES_IN[30];
  assign OP_MEM[29] = ALU_RES_IN[29];
  assign DRAM_ADDR_OUT[29] = ALU_RES_IN[29];
  assign OP_MEM[28] = ALU_RES_IN[28];
  assign DRAM_ADDR_OUT[28] = ALU_RES_IN[28];
  assign OP_MEM[27] = ALU_RES_IN[27];
  assign DRAM_ADDR_OUT[27] = ALU_RES_IN[27];
  assign OP_MEM[26] = ALU_RES_IN[26];
  assign DRAM_ADDR_OUT[26] = ALU_RES_IN[26];
  assign OP_MEM[25] = ALU_RES_IN[25];
  assign DRAM_ADDR_OUT[25] = ALU_RES_IN[25];
  assign OP_MEM[24] = ALU_RES_IN[24];
  assign DRAM_ADDR_OUT[24] = ALU_RES_IN[24];
  assign OP_MEM[23] = ALU_RES_IN[23];
  assign DRAM_ADDR_OUT[23] = ALU_RES_IN[23];
  assign OP_MEM[22] = ALU_RES_IN[22];
  assign DRAM_ADDR_OUT[22] = ALU_RES_IN[22];
  assign OP_MEM[21] = ALU_RES_IN[21];
  assign DRAM_ADDR_OUT[21] = ALU_RES_IN[21];
  assign OP_MEM[20] = ALU_RES_IN[20];
  assign DRAM_ADDR_OUT[20] = ALU_RES_IN[20];
  assign OP_MEM[19] = ALU_RES_IN[19];
  assign DRAM_ADDR_OUT[19] = ALU_RES_IN[19];
  assign OP_MEM[18] = ALU_RES_IN[18];
  assign DRAM_ADDR_OUT[18] = ALU_RES_IN[18];
  assign OP_MEM[17] = ALU_RES_IN[17];
  assign DRAM_ADDR_OUT[17] = ALU_RES_IN[17];
  assign OP_MEM[16] = ALU_RES_IN[16];
  assign DRAM_ADDR_OUT[16] = ALU_RES_IN[16];
  assign OP_MEM[15] = ALU_RES_IN[15];
  assign DRAM_ADDR_OUT[15] = ALU_RES_IN[15];
  assign OP_MEM[14] = ALU_RES_IN[14];
  assign DRAM_ADDR_OUT[14] = ALU_RES_IN[14];
  assign OP_MEM[13] = ALU_RES_IN[13];
  assign DRAM_ADDR_OUT[13] = ALU_RES_IN[13];
  assign OP_MEM[12] = ALU_RES_IN[12];
  assign DRAM_ADDR_OUT[12] = ALU_RES_IN[12];
  assign OP_MEM[11] = ALU_RES_IN[11];
  assign DRAM_ADDR_OUT[11] = ALU_RES_IN[11];
  assign OP_MEM[10] = ALU_RES_IN[10];
  assign DRAM_ADDR_OUT[10] = ALU_RES_IN[10];
  assign OP_MEM[9] = ALU_RES_IN[9];
  assign DRAM_ADDR_OUT[9] = ALU_RES_IN[9];
  assign OP_MEM[8] = ALU_RES_IN[8];
  assign DRAM_ADDR_OUT[8] = ALU_RES_IN[8];
  assign OP_MEM[7] = ALU_RES_IN[7];
  assign DRAM_ADDR_OUT[7] = ALU_RES_IN[7];
  assign OP_MEM[6] = ALU_RES_IN[6];
  assign DRAM_ADDR_OUT[6] = ALU_RES_IN[6];
  assign OP_MEM[5] = ALU_RES_IN[5];
  assign DRAM_ADDR_OUT[5] = ALU_RES_IN[5];
  assign OP_MEM[4] = ALU_RES_IN[4];
  assign DRAM_ADDR_OUT[4] = ALU_RES_IN[4];
  assign OP_MEM[3] = ALU_RES_IN[3];
  assign DRAM_ADDR_OUT[3] = ALU_RES_IN[3];
  assign OP_MEM[2] = ALU_RES_IN[2];
  assign DRAM_ADDR_OUT[2] = ALU_RES_IN[2];
  assign OP_MEM[1] = ALU_RES_IN[1];
  assign DRAM_ADDR_OUT[1] = ALU_RES_IN[1];
  assign OP_MEM[0] = ALU_RES_IN[0];
  assign DRAM_ADDR_OUT[0] = ALU_RES_IN[0];
  assign DRAM_DATA_OUT[31] = B_IN[31];
  assign DRAM_DATA_OUT[30] = B_IN[30];
  assign DRAM_DATA_OUT[29] = B_IN[29];
  assign DRAM_DATA_OUT[28] = B_IN[28];
  assign DRAM_DATA_OUT[27] = B_IN[27];
  assign DRAM_DATA_OUT[26] = B_IN[26];
  assign DRAM_DATA_OUT[25] = B_IN[25];
  assign DRAM_DATA_OUT[24] = B_IN[24];
  assign DRAM_DATA_OUT[23] = B_IN[23];
  assign DRAM_DATA_OUT[22] = B_IN[22];
  assign DRAM_DATA_OUT[21] = B_IN[21];
  assign DRAM_DATA_OUT[20] = B_IN[20];
  assign DRAM_DATA_OUT[19] = B_IN[19];
  assign DRAM_DATA_OUT[18] = B_IN[18];
  assign DRAM_DATA_OUT[17] = B_IN[17];
  assign DRAM_DATA_OUT[16] = B_IN[16];
  assign DRAM_DATA_OUT[15] = B_IN[15];
  assign DRAM_DATA_OUT[14] = B_IN[14];
  assign DRAM_DATA_OUT[13] = B_IN[13];
  assign DRAM_DATA_OUT[12] = B_IN[12];
  assign DRAM_DATA_OUT[11] = B_IN[11];
  assign DRAM_DATA_OUT[10] = B_IN[10];
  assign DRAM_DATA_OUT[9] = B_IN[9];
  assign DRAM_DATA_OUT[8] = B_IN[8];
  assign DRAM_DATA_OUT[7] = B_IN[7];
  assign DRAM_DATA_OUT[6] = B_IN[6];
  assign DRAM_DATA_OUT[5] = B_IN[5];
  assign DRAM_DATA_OUT[4] = B_IN[4];
  assign DRAM_DATA_OUT[3] = B_IN[3];
  assign DRAM_DATA_OUT[2] = B_IN[2];
  assign DRAM_DATA_OUT[1] = B_IN[1];
  assign DRAM_DATA_OUT[0] = B_IN[0];
  assign ADD_WR_MEM[4] = ADD_WR_IN[4];
  assign ADD_WR_MEM[3] = ADD_WR_IN[3];
  assign ADD_WR_MEM[2] = ADD_WR_IN[2];
  assign ADD_WR_MEM[1] = ADD_WR_IN[1];
  assign ADD_WR_MEM[0] = ADD_WR_IN[0];

  regn_N32_2 LMD ( .DIN(DRAM_DATA_IN), .CLK(CLK), .EN(MEM_EN_IN), .RST(RST), 
        .DOUT(DATA_OUT) );
  regn_N5_1 reg0 ( .DIN(ADD_WR_IN), .CLK(CLK), .EN(MEM_EN_IN), .RST(RST), 
        .DOUT(ADD_WR_OUT) );
  regn_N32_1 reg1 ( .DIN(ALU_RES_IN), .CLK(CLK), .EN(MEM_EN_IN), .RST(RST), 
        .DOUT(ALU_RES_OUT) );
  mux41_NBIT32_2 PCsel ( .A(NPC_IN), .B(NPC_REL), .C(NPC_ABS), .D({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(PC_SEL), .Z(PC_OUT) );
endmodule


module ff_2 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n4, n5, n6;

  DFFR_X1 Q_reg ( .D(n4), .CK(CLK), .RN(RST), .Q(Q), .QN(n5) );
  OAI21_X1 U2 ( .B1(n5), .B2(EN), .A(n6), .ZN(n4) );
  NAND2_X1 U3 ( .A1(EN), .A2(D), .ZN(n6) );
endmodule


module mux21_NBIT32_2 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100;

  BUF_X1 U1 ( .A(n68), .Z(n1) );
  BUF_X1 U2 ( .A(n68), .Z(n2) );
  BUF_X1 U3 ( .A(n68), .Z(n3) );
  INV_X1 U4 ( .A(n81), .ZN(Z[20]) );
  AOI22_X1 U5 ( .A1(A[20]), .A2(n2), .B1(B[20]), .B2(S), .ZN(n81) );
  INV_X1 U6 ( .A(n82), .ZN(Z[21]) );
  AOI22_X1 U7 ( .A1(A[21]), .A2(n2), .B1(B[21]), .B2(S), .ZN(n82) );
  INV_X1 U8 ( .A(n83), .ZN(Z[22]) );
  AOI22_X1 U9 ( .A1(A[22]), .A2(n2), .B1(B[22]), .B2(S), .ZN(n83) );
  INV_X1 U10 ( .A(n77), .ZN(Z[17]) );
  AOI22_X1 U11 ( .A1(A[17]), .A2(n1), .B1(B[17]), .B2(S), .ZN(n77) );
  INV_X1 U12 ( .A(n78), .ZN(Z[18]) );
  AOI22_X1 U13 ( .A1(A[18]), .A2(n1), .B1(B[18]), .B2(S), .ZN(n78) );
  INV_X1 U14 ( .A(n80), .ZN(Z[1]) );
  AOI22_X1 U15 ( .A1(A[1]), .A2(n1), .B1(B[1]), .B2(S), .ZN(n80) );
  INV_X1 U16 ( .A(n73), .ZN(Z[13]) );
  AOI22_X1 U17 ( .A1(A[13]), .A2(n1), .B1(B[13]), .B2(S), .ZN(n73) );
  INV_X1 U18 ( .A(n74), .ZN(Z[14]) );
  AOI22_X1 U19 ( .A1(A[14]), .A2(n1), .B1(B[14]), .B2(S), .ZN(n74) );
  INV_X1 U20 ( .A(n76), .ZN(Z[16]) );
  AOI22_X1 U21 ( .A1(A[16]), .A2(n1), .B1(B[16]), .B2(S), .ZN(n76) );
  INV_X1 U22 ( .A(n69), .ZN(Z[0]) );
  AOI22_X1 U23 ( .A1(A[0]), .A2(n1), .B1(B[0]), .B2(S), .ZN(n69) );
  INV_X1 U24 ( .A(n70), .ZN(Z[10]) );
  AOI22_X1 U25 ( .A1(A[10]), .A2(n1), .B1(B[10]), .B2(S), .ZN(n70) );
  INV_X1 U26 ( .A(n72), .ZN(Z[12]) );
  AOI22_X1 U27 ( .A1(A[12]), .A2(n1), .B1(B[12]), .B2(S), .ZN(n72) );
  INV_X1 U28 ( .A(n97), .ZN(Z[6]) );
  AOI22_X1 U29 ( .A1(A[6]), .A2(n3), .B1(B[6]), .B2(S), .ZN(n97) );
  INV_X1 U30 ( .A(n99), .ZN(Z[8]) );
  AOI22_X1 U31 ( .A1(A[8]), .A2(n3), .B1(B[8]), .B2(S), .ZN(n99) );
  INV_X1 U32 ( .A(n95), .ZN(Z[4]) );
  AOI22_X1 U33 ( .A1(A[4]), .A2(n3), .B1(B[4]), .B2(S), .ZN(n95) );
  INV_X1 U34 ( .A(n96), .ZN(Z[5]) );
  AOI22_X1 U35 ( .A1(A[5]), .A2(n3), .B1(B[5]), .B2(S), .ZN(n96) );
  INV_X1 U36 ( .A(n89), .ZN(Z[28]) );
  AOI22_X1 U37 ( .A1(A[28]), .A2(n2), .B1(B[28]), .B2(S), .ZN(n89) );
  INV_X1 U38 ( .A(n90), .ZN(Z[29]) );
  AOI22_X1 U39 ( .A1(A[29]), .A2(n2), .B1(B[29]), .B2(S), .ZN(n90) );
  INV_X1 U40 ( .A(n91), .ZN(Z[2]) );
  AOI22_X1 U41 ( .A1(A[2]), .A2(n2), .B1(B[2]), .B2(S), .ZN(n91) );
  INV_X1 U42 ( .A(n92), .ZN(Z[30]) );
  AOI22_X1 U43 ( .A1(A[30]), .A2(n2), .B1(B[30]), .B2(S), .ZN(n92) );
  INV_X1 U44 ( .A(n85), .ZN(Z[24]) );
  AOI22_X1 U45 ( .A1(A[24]), .A2(n2), .B1(B[24]), .B2(S), .ZN(n85) );
  INV_X1 U46 ( .A(n86), .ZN(Z[25]) );
  AOI22_X1 U47 ( .A1(A[25]), .A2(n2), .B1(B[25]), .B2(S), .ZN(n86) );
  INV_X1 U48 ( .A(n87), .ZN(Z[26]) );
  AOI22_X1 U49 ( .A1(A[26]), .A2(n2), .B1(B[26]), .B2(S), .ZN(n87) );
  INV_X1 U50 ( .A(n94), .ZN(Z[3]) );
  AOI22_X1 U51 ( .A1(A[3]), .A2(n3), .B1(B[3]), .B2(S), .ZN(n94) );
  INV_X1 U52 ( .A(n98), .ZN(Z[7]) );
  AOI22_X1 U53 ( .A1(A[7]), .A2(n3), .B1(B[7]), .B2(S), .ZN(n98) );
  INV_X1 U54 ( .A(n71), .ZN(Z[11]) );
  AOI22_X1 U55 ( .A1(A[11]), .A2(n1), .B1(B[11]), .B2(S), .ZN(n71) );
  INV_X1 U56 ( .A(n75), .ZN(Z[15]) );
  AOI22_X1 U57 ( .A1(A[15]), .A2(n1), .B1(B[15]), .B2(S), .ZN(n75) );
  INV_X1 U58 ( .A(n79), .ZN(Z[19]) );
  AOI22_X1 U59 ( .A1(A[19]), .A2(n1), .B1(B[19]), .B2(S), .ZN(n79) );
  INV_X1 U60 ( .A(n84), .ZN(Z[23]) );
  AOI22_X1 U61 ( .A1(A[23]), .A2(n2), .B1(B[23]), .B2(S), .ZN(n84) );
  INV_X1 U62 ( .A(n88), .ZN(Z[27]) );
  AOI22_X1 U63 ( .A1(A[27]), .A2(n2), .B1(B[27]), .B2(S), .ZN(n88) );
  INV_X1 U64 ( .A(n93), .ZN(Z[31]) );
  AOI22_X1 U65 ( .A1(A[31]), .A2(n3), .B1(B[31]), .B2(S), .ZN(n93) );
  INV_X1 U66 ( .A(n100), .ZN(Z[9]) );
  AOI22_X1 U67 ( .A1(A[9]), .A2(n3), .B1(S), .B2(B[9]), .ZN(n100) );
  INV_X1 U68 ( .A(S), .ZN(n68) );
endmodule


module Writeback ( WB_MUX_SEL, DATA_IN, ALU_RES_IN, ADD_WR_IN, DATA_OUT, 
        ADD_WR_OUT );
  input [31:0] DATA_IN;
  input [31:0] ALU_RES_IN;
  input [4:0] ADD_WR_IN;
  output [31:0] DATA_OUT;
  output [4:0] ADD_WR_OUT;
  input WB_MUX_SEL;

  assign ADD_WR_OUT[4] = ADD_WR_IN[4];
  assign ADD_WR_OUT[3] = ADD_WR_IN[3];
  assign ADD_WR_OUT[2] = ADD_WR_IN[2];
  assign ADD_WR_OUT[1] = ADD_WR_IN[1];
  assign ADD_WR_OUT[0] = ADD_WR_IN[0];

  mux21_NBIT32_2 WBmux ( .A(DATA_IN), .B(ALU_RES_IN), .S(WB_MUX_SEL), .Z(
        DATA_OUT) );
endmodule


module HazardDetection_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \A[0] ;
  wire   [32:0] carry;
  assign DIFF[1] = A[1];
  assign DIFF[0] = \A[0] ;
  assign \A[0]  = A[0];

  XNOR2_X1 U1 ( .A(A[5]), .B(carry[5]), .ZN(DIFF[5]) );
  XNOR2_X1 U2 ( .A(A[6]), .B(carry[6]), .ZN(DIFF[6]) );
  XNOR2_X1 U3 ( .A(A[10]), .B(carry[10]), .ZN(DIFF[10]) );
  XNOR2_X1 U4 ( .A(A[13]), .B(carry[13]), .ZN(DIFF[13]) );
  XNOR2_X1 U5 ( .A(A[11]), .B(carry[11]), .ZN(DIFF[11]) );
  XNOR2_X1 U6 ( .A(A[14]), .B(carry[14]), .ZN(DIFF[14]) );
  XNOR2_X1 U7 ( .A(A[15]), .B(carry[15]), .ZN(DIFF[15]) );
  XNOR2_X1 U8 ( .A(A[17]), .B(carry[17]), .ZN(DIFF[17]) );
  XNOR2_X1 U9 ( .A(A[4]), .B(carry[4]), .ZN(DIFF[4]) );
  XNOR2_X1 U10 ( .A(A[8]), .B(carry[8]), .ZN(DIFF[8]) );
  XNOR2_X1 U11 ( .A(A[9]), .B(carry[9]), .ZN(DIFF[9]) );
  INV_X1 U12 ( .A(A[2]), .ZN(DIFF[2]) );
  XNOR2_X1 U13 ( .A(A[20]), .B(carry[20]), .ZN(DIFF[20]) );
  XNOR2_X1 U14 ( .A(A[21]), .B(carry[21]), .ZN(DIFF[21]) );
  XNOR2_X1 U15 ( .A(A[22]), .B(carry[22]), .ZN(DIFF[22]) );
  XNOR2_X1 U16 ( .A(A[23]), .B(carry[23]), .ZN(DIFF[23]) );
  XNOR2_X1 U17 ( .A(A[24]), .B(carry[24]), .ZN(DIFF[24]) );
  XNOR2_X1 U18 ( .A(A[25]), .B(carry[25]), .ZN(DIFF[25]) );
  XNOR2_X1 U19 ( .A(A[26]), .B(carry[26]), .ZN(DIFF[26]) );
  XNOR2_X1 U20 ( .A(A[28]), .B(carry[28]), .ZN(DIFF[28]) );
  XNOR2_X1 U21 ( .A(A[29]), .B(carry[29]), .ZN(DIFF[29]) );
  XNOR2_X1 U22 ( .A(A[30]), .B(carry[30]), .ZN(DIFF[30]) );
  XNOR2_X1 U23 ( .A(A[31]), .B(carry[31]), .ZN(DIFF[31]) );
  XNOR2_X1 U24 ( .A(A[7]), .B(carry[7]), .ZN(DIFF[7]) );
  XNOR2_X1 U25 ( .A(A[12]), .B(carry[12]), .ZN(DIFF[12]) );
  XNOR2_X1 U26 ( .A(A[16]), .B(carry[16]), .ZN(DIFF[16]) );
  XNOR2_X1 U27 ( .A(A[3]), .B(A[2]), .ZN(DIFF[3]) );
  XNOR2_X1 U28 ( .A(A[18]), .B(carry[18]), .ZN(DIFF[18]) );
  XNOR2_X1 U29 ( .A(A[19]), .B(carry[19]), .ZN(DIFF[19]) );
  XNOR2_X1 U30 ( .A(A[27]), .B(carry[27]), .ZN(DIFF[27]) );
  OR2_X1 U31 ( .A1(A[3]), .A2(A[2]), .ZN(carry[4]) );
  OR2_X1 U32 ( .A1(A[4]), .A2(carry[4]), .ZN(carry[5]) );
  OR2_X1 U33 ( .A1(A[5]), .A2(carry[5]), .ZN(carry[6]) );
  OR2_X1 U34 ( .A1(A[6]), .A2(carry[6]), .ZN(carry[7]) );
  OR2_X1 U35 ( .A1(A[7]), .A2(carry[7]), .ZN(carry[8]) );
  OR2_X1 U36 ( .A1(A[8]), .A2(carry[8]), .ZN(carry[9]) );
  OR2_X1 U37 ( .A1(A[9]), .A2(carry[9]), .ZN(carry[10]) );
  OR2_X1 U38 ( .A1(A[10]), .A2(carry[10]), .ZN(carry[11]) );
  OR2_X1 U39 ( .A1(A[11]), .A2(carry[11]), .ZN(carry[12]) );
  OR2_X1 U40 ( .A1(A[12]), .A2(carry[12]), .ZN(carry[13]) );
  OR2_X1 U41 ( .A1(A[13]), .A2(carry[13]), .ZN(carry[14]) );
  OR2_X1 U42 ( .A1(A[14]), .A2(carry[14]), .ZN(carry[15]) );
  OR2_X1 U43 ( .A1(A[15]), .A2(carry[15]), .ZN(carry[16]) );
  OR2_X1 U44 ( .A1(A[16]), .A2(carry[16]), .ZN(carry[17]) );
  OR2_X1 U45 ( .A1(A[17]), .A2(carry[17]), .ZN(carry[18]) );
  OR2_X1 U46 ( .A1(A[18]), .A2(carry[18]), .ZN(carry[19]) );
  OR2_X1 U47 ( .A1(A[19]), .A2(carry[19]), .ZN(carry[20]) );
  OR2_X1 U48 ( .A1(A[20]), .A2(carry[20]), .ZN(carry[21]) );
  OR2_X1 U49 ( .A1(A[21]), .A2(carry[21]), .ZN(carry[22]) );
  OR2_X1 U50 ( .A1(A[22]), .A2(carry[22]), .ZN(carry[23]) );
  OR2_X1 U51 ( .A1(A[23]), .A2(carry[23]), .ZN(carry[24]) );
  OR2_X1 U52 ( .A1(A[24]), .A2(carry[24]), .ZN(carry[25]) );
  OR2_X1 U53 ( .A1(A[25]), .A2(carry[25]), .ZN(carry[26]) );
  OR2_X1 U54 ( .A1(A[26]), .A2(carry[26]), .ZN(carry[27]) );
  OR2_X1 U55 ( .A1(A[27]), .A2(carry[27]), .ZN(carry[28]) );
  OR2_X1 U56 ( .A1(A[28]), .A2(carry[28]), .ZN(carry[29]) );
  OR2_X1 U57 ( .A1(A[29]), .A2(carry[29]), .ZN(carry[30]) );
  OR2_X1 U58 ( .A1(A[30]), .A2(carry[30]), .ZN(carry[31]) );
endmodule


module HazardDetection ( RST, ADD_RS1, ADD_RS2, ADD_WR, DRAM_R, INS_IN, PC_IN, 
        Bubble, HDU_INS_OUT, HDU_PC_OUT, HDU_NPC_OUT );
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [4:0] ADD_WR;
  input [31:0] INS_IN;
  input [31:0] PC_IN;
  output [31:0] HDU_INS_OUT;
  output [31:0] HDU_PC_OUT;
  output [31:0] HDU_NPC_OUT;
  input RST, DRAM_R;
  output Bubble;
  wire   n1, n2, n3, n4, n5, n6, n9, n10, n12, n13, n14, n15, n16;
  assign HDU_INS_OUT[31] = INS_IN[31];
  assign HDU_INS_OUT[30] = INS_IN[30];
  assign HDU_INS_OUT[29] = INS_IN[29];
  assign HDU_INS_OUT[28] = INS_IN[28];
  assign HDU_INS_OUT[27] = INS_IN[27];
  assign HDU_INS_OUT[26] = INS_IN[26];
  assign HDU_INS_OUT[25] = INS_IN[25];
  assign HDU_INS_OUT[24] = INS_IN[24];
  assign HDU_INS_OUT[23] = INS_IN[23];
  assign HDU_INS_OUT[22] = INS_IN[22];
  assign HDU_INS_OUT[21] = INS_IN[21];
  assign HDU_INS_OUT[20] = INS_IN[20];
  assign HDU_INS_OUT[19] = INS_IN[19];
  assign HDU_INS_OUT[18] = INS_IN[18];
  assign HDU_INS_OUT[17] = INS_IN[17];
  assign HDU_INS_OUT[16] = INS_IN[16];
  assign HDU_INS_OUT[15] = INS_IN[15];
  assign HDU_INS_OUT[14] = INS_IN[14];
  assign HDU_INS_OUT[13] = INS_IN[13];
  assign HDU_INS_OUT[12] = INS_IN[12];
  assign HDU_INS_OUT[11] = INS_IN[11];
  assign HDU_INS_OUT[10] = INS_IN[10];
  assign HDU_INS_OUT[9] = INS_IN[9];
  assign HDU_INS_OUT[8] = INS_IN[8];
  assign HDU_INS_OUT[7] = INS_IN[7];
  assign HDU_INS_OUT[6] = INS_IN[6];
  assign HDU_INS_OUT[5] = INS_IN[5];
  assign HDU_INS_OUT[4] = INS_IN[4];
  assign HDU_INS_OUT[3] = INS_IN[3];
  assign HDU_INS_OUT[2] = INS_IN[2];
  assign HDU_INS_OUT[1] = INS_IN[1];
  assign HDU_INS_OUT[0] = INS_IN[0];
  assign HDU_NPC_OUT[31] = PC_IN[31];
  assign HDU_NPC_OUT[30] = PC_IN[30];
  assign HDU_NPC_OUT[29] = PC_IN[29];
  assign HDU_NPC_OUT[28] = PC_IN[28];
  assign HDU_NPC_OUT[27] = PC_IN[27];
  assign HDU_NPC_OUT[26] = PC_IN[26];
  assign HDU_NPC_OUT[25] = PC_IN[25];
  assign HDU_NPC_OUT[24] = PC_IN[24];
  assign HDU_NPC_OUT[23] = PC_IN[23];
  assign HDU_NPC_OUT[22] = PC_IN[22];
  assign HDU_NPC_OUT[21] = PC_IN[21];
  assign HDU_NPC_OUT[20] = PC_IN[20];
  assign HDU_NPC_OUT[19] = PC_IN[19];
  assign HDU_NPC_OUT[18] = PC_IN[18];
  assign HDU_NPC_OUT[17] = PC_IN[17];
  assign HDU_NPC_OUT[16] = PC_IN[16];
  assign HDU_NPC_OUT[15] = PC_IN[15];
  assign HDU_NPC_OUT[14] = PC_IN[14];
  assign HDU_NPC_OUT[13] = PC_IN[13];
  assign HDU_NPC_OUT[12] = PC_IN[12];
  assign HDU_NPC_OUT[11] = PC_IN[11];
  assign HDU_NPC_OUT[10] = PC_IN[10];
  assign HDU_NPC_OUT[9] = PC_IN[9];
  assign HDU_NPC_OUT[8] = PC_IN[8];
  assign HDU_NPC_OUT[7] = PC_IN[7];
  assign HDU_NPC_OUT[6] = PC_IN[6];
  assign HDU_NPC_OUT[5] = PC_IN[5];
  assign HDU_NPC_OUT[4] = PC_IN[4];
  assign HDU_NPC_OUT[3] = PC_IN[3];
  assign HDU_NPC_OUT[2] = PC_IN[2];
  assign HDU_NPC_OUT[1] = PC_IN[1];
  assign HDU_NPC_OUT[0] = PC_IN[0];

  HazardDetection_DW01_sub_0 sub_25 ( .A(PC_IN), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .DIFF(HDU_PC_OUT) );
  AND3_X1 U4 ( .A1(DRAM_R), .A2(n1), .A3(RST), .ZN(Bubble) );
  OAI33_X1 U5 ( .A1(n2), .A2(n3), .A3(n4), .B1(n5), .B2(n6), .B3(n9), .ZN(n1)
         );
  XOR2_X1 U6 ( .A(ADD_WR[4]), .B(ADD_RS2[4]), .Z(n9) );
  XOR2_X1 U8 ( .A(ADD_WR[2]), .B(ADD_RS2[2]), .Z(n6) );
  NAND3_X1 U9 ( .A1(n10), .A2(n12), .A3(n13), .ZN(n5) );
  XNOR2_X1 U11 ( .A(ADD_WR[0]), .B(ADD_RS2[0]), .ZN(n13) );
  XNOR2_X1 U12 ( .A(ADD_WR[1]), .B(ADD_RS2[1]), .ZN(n12) );
  XNOR2_X1 U13 ( .A(ADD_WR[3]), .B(ADD_RS2[3]), .ZN(n10) );
  XOR2_X1 U14 ( .A(ADD_WR[4]), .B(ADD_RS1[4]), .Z(n4) );
  XOR2_X1 U15 ( .A(ADD_WR[2]), .B(ADD_RS1[2]), .Z(n3) );
  NAND3_X1 U16 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n2) );
  XNOR2_X1 U17 ( .A(ADD_WR[0]), .B(ADD_RS1[0]), .ZN(n16) );
  XNOR2_X1 U18 ( .A(ADD_WR[1]), .B(ADD_RS1[1]), .ZN(n15) );
  XNOR2_X1 U19 ( .A(ADD_WR[3]), .B(ADD_RS1[3]), .ZN(n14) );
endmodule


module Datapath ( CLK, RST, INS_IN, DATA_IN, REG_LATCH_EN, RD1, RD2, MUX_A_SEL, 
        MUX_B_SEL, .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , 
        \ALU_OPC[0] }), ALU_OUTREG_EN, JUMP_TYPE, DRAM_R_IN, MEM_EN_IN, 
        DRAM_W_IN, RF_WE, DRAM_EN_IN, WB_MUX_SEL, INS_OUT, IRAM_ADDR_OUT, 
        DRAM_ADDR_OUT, DATA_OUT, DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, 
        Bubble_out );
  input [31:0] INS_IN;
  input [31:0] DATA_IN;
  input [1:0] MUX_B_SEL;
  input [1:0] JUMP_TYPE;
  output [31:0] INS_OUT;
  output [31:0] IRAM_ADDR_OUT;
  output [31:0] DRAM_ADDR_OUT;
  output [31:0] DATA_OUT;
  input CLK, RST, REG_LATCH_EN, RD1, RD2, MUX_A_SEL, \ALU_OPC[3] ,
         \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] , ALU_OUTREG_EN, DRAM_R_IN,
         MEM_EN_IN, DRAM_W_IN, RF_WE, DRAM_EN_IN, WB_MUX_SEL;
  output DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble_out;
  wire   ZERO_FLAG_EX, RF_WE_WB, DRAM_R_MEM;
  wire   [3:0] ALU_OPC;
  wire   [31:0] PC_MEM_OUT;
  wire   [31:0] sig_HDU_INS_OUT;
  wire   [31:0] sig_HDU_PC_OUT;
  wire   [31:0] sig_HDU_NPC_OUT;
  wire   [31:0] PC_FETCH_OUT;
  wire   [31:0] NPC_FETCH_OUT;
  wire   [4:0] ADD_WR_WB;
  wire   [31:0] OP_WB;
  wire   [31:0] PC_DECODE_OUT;
  wire   [31:0] A_DECODE_OUT;
  wire   [31:0] B_DECODE_OUT;
  wire   [31:0] IMM_DECODE_OUT;
  wire   [4:0] ADD_RS1_HDU;
  wire   [4:0] ADD_RS2_HDU;
  wire   [4:0] ADD_WR_DECODE_OUT;
  wire   [4:0] ADD_RS1_DECODE_OUT;
  wire   [4:0] ADD_RS2_DECODE_OUT;
  wire   [4:0] ADD_WR_MEM;
  wire   [31:0] OP_MEM;
  wire   [1:0] PC_SEL_EX;
  wire   [31:0] NPC_ABS_EX;
  wire   [31:0] NPC_REL_EX;
  wire   [31:0] ALU_RES_EX;
  wire   [31:0] B_EX_OUT;
  wire   [4:0] ADD_WR_EX_OUT;
  wire   [31:0] DATA_MEM_OUT;
  wire   [31:0] ALU_RES_MEM;
  wire   [4:0] ADD_WR_MEM_OUT;

  Fetch FetchStage ( .CLK(CLK), .RST(RST), .ZERO_FLAG(ZERO_FLAG_EX), .PC_EXT(
        PC_MEM_OUT), .INS_IN(INS_IN), .Bubble_in(Bubble_out), .HDU_INS_IN(
        sig_HDU_INS_OUT), .HDU_PC_IN(sig_HDU_PC_OUT), .HDU_NPC_IN(
        sig_HDU_NPC_OUT), .PC_OUT(PC_FETCH_OUT), .ADDR_OUT(IRAM_ADDR_OUT), 
        .NPC_OUT(NPC_FETCH_OUT), .INS_OUT(INS_OUT) );
  Decode DecodeStage ( .CLK(CLK), .RST(RST), .REG_LATCH_EN(REG_LATCH_EN), 
        .RD1(RD1), .RD2(RD2), .RF_WE(RF_WE_WB), .ZERO_FLAG(ZERO_FLAG_EX), 
        .PC_IN(PC_FETCH_OUT), .INS_IN(INS_OUT), .ADD_WR(ADD_WR_WB), 
        .DATA_WR_IN(OP_WB), .PC_OUT(PC_DECODE_OUT), .A_OUT(A_DECODE_OUT), 
        .B_OUT(B_DECODE_OUT), .IMM_OUT(IMM_DECODE_OUT), .ADD_RS1_HDU(
        ADD_RS1_HDU), .ADD_RS2_HDU(ADD_RS2_HDU), .ADD_WR_OUT(ADD_WR_DECODE_OUT), .ADD_RS1_OUT(ADD_RS1_DECODE_OUT), .ADD_RS2_OUT(ADD_RS2_DECODE_OUT) );
  Execute ExecuteStage ( .CLK(CLK), .RST(RST), .MUX_A_SEL(MUX_A_SEL), 
        .MUX_B_SEL(MUX_B_SEL), .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , 
        \ALU_OPC[1] , \ALU_OPC[0] }), .ALU_OUTREG_EN(ALU_OUTREG_EN), 
        .JUMP_TYPE(JUMP_TYPE), .PC_IN(PC_DECODE_OUT), .A_IN(A_DECODE_OUT), 
        .B_IN(B_DECODE_OUT), .IMM_IN(IMM_DECODE_OUT), .ADD_WR_IN(
        ADD_WR_DECODE_OUT), .ADD_RS1_IN(ADD_RS1_DECODE_OUT), .ADD_RS2_IN(
        ADD_RS2_DECODE_OUT), .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_WB(ADD_WR_WB), 
        .RF_WE_MEM(RF_WE), .RF_WE_WB(RF_WE_WB), .OP_MEM(OP_MEM), .OP_WB(OP_WB), 
        .PC_SEL(PC_SEL_EX), .ZERO_FLAG(ZERO_FLAG_EX), .NPC_ABS(NPC_ABS_EX), 
        .NPC_REL(NPC_REL_EX), .ALU_RES(ALU_RES_EX), .B_OUT(B_EX_OUT), 
        .ADD_WR_OUT(ADD_WR_EX_OUT) );
  ff_0 DRAM_R_ff ( .D(DRAM_R_IN), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(
        DRAM_R_MEM) );
  Memory MemoryStage ( .CLK(CLK), .RST(RST), .MEM_EN_IN(MEM_EN_IN), 
        .DRAM_R_IN(DRAM_R_MEM), .DRAM_W_IN(DRAM_W_IN), .DRAM_EN_IN(DRAM_EN_IN), 
        .PC_SEL(PC_SEL_EX), .NPC_IN(NPC_FETCH_OUT), .NPC_ABS(NPC_ABS_EX), 
        .NPC_REL(NPC_REL_EX), .ALU_RES_IN(ALU_RES_EX), .B_IN(B_EX_OUT), 
        .ADD_WR_IN(ADD_WR_EX_OUT), .DRAM_DATA_IN(DATA_IN), .PC_OUT(PC_MEM_OUT), 
        .DRAM_EN_OUT(DRAM_EN_OUT), .DRAM_R_OUT(DRAM_R_OUT), .DRAM_W_OUT(
        DRAM_W_OUT), .DRAM_ADDR_OUT(DRAM_ADDR_OUT), .DRAM_DATA_OUT(DATA_OUT), 
        .DATA_OUT(DATA_MEM_OUT), .ALU_RES_OUT(ALU_RES_MEM), .OP_MEM(OP_MEM), 
        .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_OUT(ADD_WR_MEM_OUT) );
  ff_2 RF_WE_ff ( .D(RF_WE), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(RF_WE_WB) );
  Writeback WritebackStage ( .WB_MUX_SEL(WB_MUX_SEL), .DATA_IN(DATA_MEM_OUT), 
        .ALU_RES_IN(ALU_RES_MEM), .ADD_WR_IN(ADD_WR_MEM_OUT), .DATA_OUT(OP_WB), 
        .ADD_WR_OUT(ADD_WR_WB) );
  HazardDetection HDU ( .RST(RST), .ADD_RS1(ADD_RS1_HDU), .ADD_RS2(ADD_RS2_HDU), .ADD_WR(ADD_WR_DECODE_OUT), .DRAM_R(DRAM_R_IN), .INS_IN(INS_OUT), .PC_IN(
        PC_FETCH_OUT), .Bubble(Bubble_out), .HDU_INS_OUT(sig_HDU_INS_OUT), 
        .HDU_PC_OUT(sig_HDU_PC_OUT), .HDU_NPC_OUT(sig_HDU_NPC_OUT) );
endmodule


module hardwired_cu_NBIT32 ( REG_LATCH_EN, RD1, RD2, MUX_A_SEL, MUX_B_SEL, 
    .ALU_OPC({\ALU_OPC[3] , \ALU_OPC[2] , \ALU_OPC[1] , \ALU_OPC[0] }), 
        ALU_OUTREG_EN, DRAM_R_IN, JUMP_TYPE, MEM_EN_IN, DRAM_W_IN, RF_WE, 
        DRAM_EN_IN, WB_MUX_SEL, INS_IN, Bubble, Clk, Rst );
  output [1:0] MUX_B_SEL;
  output [1:0] JUMP_TYPE;
  input [31:0] INS_IN;
  input Bubble, Clk, Rst;
  output REG_LATCH_EN, RD1, RD2, MUX_A_SEL, \ALU_OPC[3] , \ALU_OPC[2] ,
         \ALU_OPC[1] , \ALU_OPC[0] , ALU_OUTREG_EN, DRAM_R_IN, MEM_EN_IN,
         DRAM_W_IN, RF_WE, DRAM_EN_IN, WB_MUX_SEL;
  wire   INS_IN_31, INS_IN_30, INS_IN_29, INS_IN_28, INS_IN_27, INS_IN_26, N24,
         N25, N26, N27, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n58,
         n59, n60, n61, n62, n63, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18;
  wire   [3:0] ALU_OPC;
  wire   [3:0] AluOP_E;
  assign REG_LATCH_EN = 1'b0;
  assign RD1 = 1'b0;
  assign RD2 = 1'b0;
  assign MUX_A_SEL = 1'b0;
  assign MUX_B_SEL[1] = 1'b0;
  assign MUX_B_SEL[0] = 1'b0;
  assign ALU_OUTREG_EN = 1'b0;
  assign DRAM_R_IN = 1'b0;
  assign JUMP_TYPE[1] = 1'b0;
  assign JUMP_TYPE[0] = 1'b0;
  assign MEM_EN_IN = 1'b0;
  assign DRAM_W_IN = 1'b0;
  assign RF_WE = 1'b0;
  assign DRAM_EN_IN = 1'b0;
  assign WB_MUX_SEL = 1'b0;
  assign INS_IN_31 = INS_IN[31];
  assign INS_IN_30 = INS_IN[30];
  assign INS_IN_29 = INS_IN[29];
  assign INS_IN_28 = INS_IN[28];
  assign INS_IN_27 = INS_IN[27];
  assign INS_IN_26 = INS_IN[26];

  DFFR_X1 \AluOP_E_reg[3]  ( .D(N27), .CK(Clk), .RN(Rst), .Q(AluOP_E[3]) );
  DFFR_X1 \ALU_OPC_reg[3]  ( .D(AluOP_E[3]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[3]) );
  DFFR_X1 \AluOP_E_reg[2]  ( .D(N26), .CK(Clk), .RN(Rst), .Q(AluOP_E[2]) );
  DFFR_X1 \ALU_OPC_reg[2]  ( .D(AluOP_E[2]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[2]) );
  DFFR_X1 \AluOP_E_reg[1]  ( .D(N25), .CK(Clk), .RN(Rst), .Q(AluOP_E[1]) );
  DFFR_X1 \ALU_OPC_reg[1]  ( .D(AluOP_E[1]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[1]) );
  DFFR_X1 \AluOP_E_reg[0]  ( .D(N24), .CK(Clk), .RN(Rst), .Q(AluOP_E[0]) );
  DFFR_X1 \ALU_OPC_reg[0]  ( .D(AluOP_E[0]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[0]) );
  XOR2_X1 U74 ( .A(n2), .B(INS_IN[1]), .Z(n33) );
  NAND3_X1 U75 ( .A1(n16), .A2(n13), .A3(INS_IN_30), .ZN(n37) );
  OAI33_X1 U76 ( .A1(n26), .A2(n13), .A3(n17), .B1(n46), .B2(INS_IN_30), .B3(
        INS_IN_28), .ZN(n43) );
  OAI33_X1 U77 ( .A1(n24), .A2(n25), .A3(n17), .B1(n3), .B2(n8), .B3(n34), 
        .ZN(n50) );
  OAI33_X1 U78 ( .A1(n12), .A2(n56), .A3(n11), .B1(n27), .B2(INS_IN_30), .B3(
        n25), .ZN(n55) );
  NAND3_X1 U79 ( .A1(n51), .A2(n7), .A3(INS_IN[5]), .ZN(n35) );
  OAI33_X1 U80 ( .A1(n58), .A2(n13), .A3(n17), .B1(n59), .B2(n39), .B3(n6), 
        .ZN(n48) );
  NAND3_X1 U81 ( .A1(INS_IN[3]), .A2(n51), .A3(INS_IN[5]), .ZN(n39) );
  NAND3_X1 U82 ( .A1(n15), .A2(n18), .A3(INS_IN_28), .ZN(n24) );
  NAND3_X1 U83 ( .A1(n10), .A2(n13), .A3(n63), .ZN(n34) );
  NAND3_X1 U84 ( .A1(n16), .A2(n17), .A3(INS_IN_28), .ZN(n36) );
  INV_X1 U18 ( .A(n25), .ZN(n10) );
  NAND2_X1 U19 ( .A1(n12), .A2(n11), .ZN(n25) );
  AOI21_X1 U20 ( .B1(n40), .B2(n41), .A(Bubble), .ZN(N25) );
  AOI211_X1 U21 ( .C1(n14), .C2(n10), .A(n38), .B(n48), .ZN(n40) );
  AOI221_X1 U22 ( .B1(n42), .B2(n5), .C1(n16), .C2(n43), .A(n44), .ZN(n41) );
  INV_X1 U23 ( .A(n47), .ZN(n5) );
  AOI21_X1 U24 ( .B1(n28), .B2(n29), .A(Bubble), .ZN(N26) );
  AOI21_X1 U25 ( .B1(n20), .B2(n6), .A(n38), .ZN(n28) );
  NOR3_X1 U26 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n29) );
  AOI21_X1 U27 ( .B1(n36), .B2(n37), .A(n26), .ZN(n30) );
  INV_X1 U28 ( .A(n36), .ZN(n14) );
  INV_X1 U29 ( .A(n27), .ZN(n16) );
  OR2_X1 U30 ( .A1(n49), .A2(n50), .ZN(n38) );
  INV_X1 U31 ( .A(n52), .ZN(n3) );
  INV_X1 U32 ( .A(n51), .ZN(n8) );
  NAND2_X1 U33 ( .A1(n16), .A2(n10), .ZN(n58) );
  OR3_X1 U34 ( .A1(INS_IN[0]), .A2(INS_IN[1]), .A3(n34), .ZN(n59) );
  NOR4_X1 U35 ( .A1(INS_IN[6]), .A2(INS_IN[4]), .A3(INS_IN[10]), .A4(n62), 
        .ZN(n51) );
  OR3_X1 U36 ( .A1(INS_IN[9]), .A2(INS_IN[8]), .A3(INS_IN[7]), .ZN(n62) );
  NAND2_X1 U37 ( .A1(INS_IN_27), .A2(n11), .ZN(n46) );
  NOR3_X1 U38 ( .A1(INS_IN_29), .A2(INS_IN_31), .A3(INS_IN_30), .ZN(n63) );
  NOR4_X1 U39 ( .A1(n2), .A2(n39), .A3(n34), .A4(INS_IN[1]), .ZN(n20) );
  NOR4_X1 U40 ( .A1(n6), .A2(INS_IN[0]), .A3(INS_IN[3]), .A4(INS_IN[5]), .ZN(
        n52) );
  NOR4_X1 U41 ( .A1(n33), .A2(n34), .A3(n6), .A4(n35), .ZN(n32) );
  NOR4_X1 U42 ( .A1(INS_IN[1]), .A2(n4), .A3(n34), .A4(n6), .ZN(n44) );
  INV_X1 U43 ( .A(n45), .ZN(n4) );
  OAI21_X1 U44 ( .B1(n35), .B2(INS_IN[0]), .A(n39), .ZN(n45) );
  NOR3_X1 U45 ( .A1(n34), .A2(INS_IN[0]), .A3(n35), .ZN(n42) );
  INV_X1 U46 ( .A(INS_IN[3]), .ZN(n7) );
  NOR3_X1 U47 ( .A1(n36), .A2(INS_IN_26), .A3(n12), .ZN(n31) );
  INV_X1 U48 ( .A(INS_IN[2]), .ZN(n6) );
  INV_X1 U49 ( .A(INS_IN_30), .ZN(n17) );
  AOI22_X1 U50 ( .A1(n15), .A2(n18), .B1(INS_IN_31), .B2(n17), .ZN(n56) );
  NAND2_X1 U51 ( .A1(INS_IN_26), .A2(n12), .ZN(n26) );
  INV_X1 U52 ( .A(INS_IN_27), .ZN(n12) );
  AOI21_X1 U53 ( .B1(n53), .B2(n54), .A(Bubble), .ZN(N24) );
  AOI211_X1 U54 ( .C1(n14), .C2(n10), .A(n49), .B(n23), .ZN(n53) );
  AOI221_X1 U55 ( .B1(n42), .B2(n47), .C1(n55), .C2(n13), .A(n31), .ZN(n54) );
  INV_X1 U56 ( .A(INS_IN_28), .ZN(n13) );
  NAND2_X1 U57 ( .A1(INS_IN_29), .A2(n18), .ZN(n27) );
  OR2_X1 U58 ( .A1(n48), .A2(n1), .ZN(n23) );
  NOR3_X1 U59 ( .A1(n26), .A2(INS_IN_30), .A3(n24), .ZN(n1) );
  NAND2_X1 U60 ( .A1(INS_IN[1]), .A2(n6), .ZN(n47) );
  INV_X1 U61 ( .A(INS_IN_31), .ZN(n18) );
  INV_X1 U62 ( .A(INS_IN_26), .ZN(n11) );
  NAND2_X1 U63 ( .A1(n60), .A2(n61), .ZN(n49) );
  OR4_X1 U64 ( .A1(n12), .A2(n24), .A3(n17), .A4(INS_IN_26), .ZN(n61) );
  NAND4_X1 U65 ( .A1(INS_IN[1]), .A2(n52), .A3(n9), .A4(n51), .ZN(n60) );
  INV_X1 U66 ( .A(n34), .ZN(n9) );
  NOR2_X1 U67 ( .A1(Bubble), .A2(n19), .ZN(N27) );
  NOR4_X1 U68 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n19) );
  NOR3_X1 U69 ( .A1(n26), .A2(n27), .A3(n17), .ZN(n21) );
  NOR3_X1 U70 ( .A1(n24), .A2(INS_IN_30), .A3(n25), .ZN(n22) );
  INV_X1 U71 ( .A(INS_IN[0]), .ZN(n2) );
  INV_X1 U72 ( .A(INS_IN_29), .ZN(n15) );
endmodule


module DLX ( Clk, Rst );
  input Clk, Rst;
  wire   DRAM_EN_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble;
  wire   [31:0] INS_IN;
  wire   [31:0] DATA_IN;
  wire   [1:0] MUX_B_SEL;
  wire   [3:0] ALU_OPC;
  wire   [1:0] JUMP_TYPE;
  wire   [31:0] IRAM_ADDR_OUT;
  wire   [31:0] DRAM_ADDR_OUT;
  wire   [31:0] DATA_OUT;

  Datapath DP ( .CLK(Clk), .RST(Rst), .INS_IN(INS_IN), .DATA_IN(DATA_IN), 
        .REG_LATCH_EN(1'b0), .RD1(1'b0), .RD2(1'b0), .MUX_A_SEL(1'b0), 
        .MUX_B_SEL({1'b0, 1'b0}), .ALU_OPC(ALU_OPC), .ALU_OUTREG_EN(1'b0), 
        .JUMP_TYPE({1'b0, 1'b0}), .DRAM_R_IN(1'b0), .MEM_EN_IN(1'b0), 
        .DRAM_W_IN(1'b0), .RF_WE(1'b0), .DRAM_EN_IN(1'b0), .WB_MUX_SEL(1'b0), 
        .IRAM_ADDR_OUT(IRAM_ADDR_OUT), .DRAM_ADDR_OUT(DRAM_ADDR_OUT), 
        .DATA_OUT(DATA_OUT), .DRAM_EN_OUT(DRAM_EN_OUT), .DRAM_R_OUT(DRAM_R_OUT), .DRAM_W_OUT(DRAM_W_OUT), .Bubble_out(Bubble) );
  hardwired_cu_NBIT32 CU ( .ALU_OPC(ALU_OPC), .INS_IN(INS_IN), .Bubble(Bubble), 
        .Clk(Clk), .Rst(Rst) );
  IRAM IRAM_I ( .Rst(Rst), .Addr(IRAM_ADDR_OUT), .Iout(INS_IN) );
  DRAM DRAM_I ( .En(DRAM_EN_OUT), .Rst(Rst), .ADDR_IN(DRAM_ADDR_OUT), 
        .DATA_IN(DATA_OUT), .DRAM_W(DRAM_W_OUT), .DRAM_R(DRAM_R_OUT), 
        .DATA_OUT(DATA_IN) );
endmodule

